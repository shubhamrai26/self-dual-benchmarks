module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 , y9658 , y9659 , y9660 , y9661 , y9662 , y9663 , y9664 , y9665 , y9666 , y9667 , y9668 , y9669 , y9670 , y9671 , y9672 , y9673 , y9674 , y9675 , y9676 , y9677 , y9678 , y9679 , y9680 , y9681 , y9682 , y9683 , y9684 , y9685 , y9686 , y9687 , y9688 , y9689 , y9690 , y9691 , y9692 , y9693 , y9694 , y9695 , y9696 , y9697 , y9698 , y9699 , y9700 , y9701 , y9702 , y9703 , y9704 , y9705 , y9706 , y9707 , y9708 , y9709 , y9710 , y9711 , y9712 , y9713 , y9714 , y9715 , y9716 , y9717 , y9718 , y9719 , y9720 , y9721 , y9722 , y9723 , y9724 , y9725 , y9726 , y9727 , y9728 , y9729 , y9730 , y9731 , y9732 , y9733 , y9734 , y9735 , y9736 , y9737 , y9738 , y9739 , y9740 , y9741 , y9742 , y9743 , y9744 , y9745 , y9746 , y9747 , y9748 , y9749 , y9750 , y9751 , y9752 , y9753 , y9754 , y9755 , y9756 , y9757 , y9758 , y9759 , y9760 , y9761 , y9762 , y9763 , y9764 , y9765 , y9766 , y9767 , y9768 , y9769 , y9770 , y9771 , y9772 , y9773 , y9774 , y9775 , y9776 , y9777 , y9778 , y9779 , y9780 , y9781 , y9782 , y9783 , y9784 , y9785 , y9786 , y9787 , y9788 , y9789 , y9790 , y9791 , y9792 , y9793 , y9794 , y9795 , y9796 , y9797 , y9798 , y9799 , y9800 , y9801 , y9802 , y9803 , y9804 , y9805 , y9806 , y9807 , y9808 , y9809 , y9810 , y9811 , y9812 , y9813 , y9814 , y9815 , y9816 , y9817 , y9818 , y9819 , y9820 , y9821 , y9822 , y9823 , y9824 , y9825 , y9826 , y9827 , y9828 , y9829 , y9830 , y9831 , y9832 , y9833 , y9834 , y9835 , y9836 , y9837 , y9838 , y9839 , y9840 , y9841 , y9842 , y9843 , y9844 , y9845 , y9846 , y9847 , y9848 , y9849 , y9850 , y9851 , y9852 , y9853 , y9854 , y9855 , y9856 , y9857 , y9858 , y9859 , y9860 , y9861 , y9862 , y9863 , y9864 , y9865 , y9866 , y9867 , y9868 , y9869 , y9870 , y9871 , y9872 , y9873 , y9874 , y9875 , y9876 , y9877 , y9878 , y9879 , y9880 , y9881 , y9882 , y9883 , y9884 , y9885 , y9886 , y9887 , y9888 , y9889 , y9890 , y9891 , y9892 , y9893 , y9894 , y9895 , y9896 , y9897 , y9898 , y9899 , y9900 , y9901 , y9902 , y9903 , y9904 , y9905 , y9906 , y9907 , y9908 , y9909 , y9910 , y9911 , y9912 , y9913 , y9914 , y9915 , y9916 , y9917 , y9918 , y9919 , y9920 , y9921 , y9922 , y9923 , y9924 , y9925 , y9926 , y9927 , y9928 , y9929 , y9930 , y9931 , y9932 , y9933 , y9934 , y9935 , y9936 , y9937 , y9938 , y9939 , y9940 , y9941 , y9942 , y9943 , y9944 , y9945 , y9946 , y9947 , y9948 , y9949 , y9950 , y9951 , y9952 , y9953 , y9954 , y9955 , y9956 , y9957 , y9958 , y9959 , y9960 , y9961 , y9962 , y9963 , y9964 , y9965 , y9966 , y9967 , y9968 , y9969 , y9970 , y9971 , y9972 , y9973 , y9974 , y9975 , y9976 , y9977 , y9978 , y9979 , y9980 , y9981 , y9982 , y9983 , y9984 , y9985 , y9986 , y9987 , y9988 , y9989 , y9990 , y9991 , y9992 , y9993 , y9994 , y9995 , y9996 , y9997 , y9998 , y9999 , y10000 , y10001 , y10002 , y10003 , y10004 , y10005 , y10006 , y10007 , y10008 , y10009 , y10010 , y10011 , y10012 , y10013 , y10014 , y10015 , y10016 , y10017 , y10018 , y10019 , y10020 , y10021 , y10022 , y10023 , y10024 , y10025 , y10026 , y10027 , y10028 , y10029 , y10030 , y10031 , y10032 , y10033 , y10034 , y10035 , y10036 , y10037 , y10038 , y10039 , y10040 , y10041 , y10042 , y10043 , y10044 , y10045 , y10046 , y10047 , y10048 , y10049 , y10050 , y10051 , y10052 , y10053 , y10054 , y10055 , y10056 , y10057 , y10058 , y10059 , y10060 , y10061 , y10062 , y10063 , y10064 , y10065 , y10066 , y10067 , y10068 , y10069 , y10070 , y10071 , y10072 , y10073 , y10074 , y10075 , y10076 , y10077 , y10078 , y10079 , y10080 , y10081 , y10082 , y10083 , y10084 , y10085 , y10086 , y10087 , y10088 , y10089 , y10090 , y10091 , y10092 , y10093 , y10094 , y10095 , y10096 , y10097 , y10098 , y10099 , y10100 , y10101 , y10102 , y10103 , y10104 , y10105 , y10106 , y10107 , y10108 , y10109 , y10110 , y10111 , y10112 , y10113 , y10114 , y10115 , y10116 , y10117 , y10118 , y10119 , y10120 , y10121 , y10122 , y10123 , y10124 , y10125 , y10126 , y10127 , y10128 , y10129 , y10130 , y10131 , y10132 , y10133 , y10134 , y10135 , y10136 , y10137 , y10138 , y10139 , y10140 , y10141 , y10142 , y10143 , y10144 , y10145 , y10146 , y10147 , y10148 , y10149 , y10150 , y10151 , y10152 , y10153 , y10154 , y10155 , y10156 , y10157 , y10158 , y10159 , y10160 , y10161 , y10162 , y10163 , y10164 , y10165 , y10166 , y10167 , y10168 , y10169 , y10170 , y10171 , y10172 , y10173 , y10174 , y10175 , y10176 , y10177 , y10178 , y10179 , y10180 , y10181 , y10182 , y10183 , y10184 , y10185 , y10186 , y10187 , y10188 , y10189 , y10190 , y10191 , y10192 , y10193 , y10194 , y10195 , y10196 , y10197 , y10198 , y10199 , y10200 , y10201 , y10202 , y10203 , y10204 , y10205 , y10206 , y10207 , y10208 , y10209 , y10210 , y10211 , y10212 , y10213 , y10214 , y10215 , y10216 , y10217 , y10218 , y10219 , y10220 , y10221 , y10222 , y10223 , y10224 , y10225 , y10226 , y10227 , y10228 , y10229 , y10230 , y10231 , y10232 , y10233 , y10234 , y10235 , y10236 , y10237 , y10238 , y10239 , y10240 , y10241 , y10242 , y10243 , y10244 , y10245 , y10246 , y10247 , y10248 , y10249 , y10250 , y10251 , y10252 , y10253 , y10254 , y10255 , y10256 , y10257 , y10258 , y10259 , y10260 , y10261 , y10262 , y10263 , y10264 , y10265 , y10266 , y10267 , y10268 , y10269 , y10270 , y10271 , y10272 , y10273 , y10274 , y10275 , y10276 , y10277 , y10278 , y10279 , y10280 , y10281 , y10282 , y10283 , y10284 , y10285 , y10286 , y10287 , y10288 , y10289 , y10290 , y10291 , y10292 , y10293 , y10294 , y10295 , y10296 , y10297 , y10298 , y10299 , y10300 , y10301 , y10302 , y10303 , y10304 , y10305 , y10306 , y10307 , y10308 , y10309 , y10310 , y10311 , y10312 , y10313 , y10314 , y10315 , y10316 , y10317 , y10318 , y10319 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 ;
  assign n129 = ( ~x30 & x44 ) | ( ~x30 & x91 ) | ( x44 & x91 ) ;
  assign n130 = ( x6 & x108 ) | ( x6 & ~x116 ) | ( x108 & ~x116 ) ;
  assign n131 = ( x31 & x54 ) | ( x31 & ~x95 ) | ( x54 & ~x95 ) ;
  assign n132 = ( ~x102 & x107 ) | ( ~x102 & x111 ) | ( x107 & x111 ) ;
  assign n133 = n132 ^ x74 ^ x36 ;
  assign n134 = x80 ^ x24 ^ 1'b0 ;
  assign n135 = x34 & n134 ;
  assign n136 = n135 ^ x114 ^ x111 ;
  assign n137 = ( ~x75 & x81 ) | ( ~x75 & x110 ) | ( x81 & x110 ) ;
  assign n138 = x68 ^ x44 ^ 1'b0 ;
  assign n139 = x96 & n138 ;
  assign n140 = ( x122 & x123 ) | ( x122 & ~n139 ) | ( x123 & ~n139 ) ;
  assign n141 = x59 ^ x48 ^ x45 ;
  assign n142 = x61 & ~n141 ;
  assign n143 = n142 ^ x105 ^ 1'b0 ;
  assign n144 = n143 ^ x113 ^ x62 ;
  assign n145 = ( ~x7 & x20 ) | ( ~x7 & x95 ) | ( x20 & x95 ) ;
  assign n146 = ( x96 & x105 ) | ( x96 & n141 ) | ( x105 & n141 ) ;
  assign n147 = n129 ^ x115 ^ 1'b0 ;
  assign n148 = n146 & n147 ;
  assign n149 = ( x34 & ~x97 ) | ( x34 & x114 ) | ( ~x97 & x114 ) ;
  assign n150 = x58 & n149 ;
  assign n151 = ~x27 & n150 ;
  assign n152 = x94 & ~n151 ;
  assign n153 = ~x4 & n152 ;
  assign n154 = x110 ^ x73 ^ x29 ;
  assign n155 = x79 & ~n154 ;
  assign n156 = n155 ^ x127 ^ 1'b0 ;
  assign n157 = n156 ^ x119 ^ 1'b0 ;
  assign n158 = ~x118 & x122 ;
  assign n159 = ( x52 & n157 ) | ( x52 & n158 ) | ( n157 & n158 ) ;
  assign n160 = n129 ^ x126 ^ x90 ;
  assign n161 = x82 & ~n160 ;
  assign n162 = x6 & x47 ;
  assign n163 = n159 & n162 ;
  assign n164 = x33 ^ x26 ^ x13 ;
  assign n165 = ( ~x35 & x59 ) | ( ~x35 & x89 ) | ( x59 & x89 ) ;
  assign n166 = x13 & n165 ;
  assign n167 = n166 ^ x90 ^ 1'b0 ;
  assign n168 = ( x44 & x59 ) | ( x44 & ~x114 ) | ( x59 & ~x114 ) ;
  assign n169 = ( x5 & x69 ) | ( x5 & ~n168 ) | ( x69 & ~n168 ) ;
  assign n170 = n169 ^ x122 ^ x115 ;
  assign n171 = x95 ^ x8 ^ 1'b0 ;
  assign n172 = ~n170 & n171 ;
  assign n173 = x110 ^ x69 ^ 1'b0 ;
  assign n174 = n173 ^ x38 ^ 1'b0 ;
  assign n175 = x84 & n174 ;
  assign n176 = x58 & ~n175 ;
  assign n177 = n176 ^ x86 ^ x81 ;
  assign n178 = ( n131 & ~n151 ) | ( n131 & n177 ) | ( ~n151 & n177 ) ;
  assign n179 = ( x60 & ~x108 ) | ( x60 & n131 ) | ( ~x108 & n131 ) ;
  assign n180 = x120 ^ x88 ^ x65 ;
  assign n181 = x2 & ~n180 ;
  assign n182 = n181 ^ x84 ^ 1'b0 ;
  assign n183 = ( x2 & ~x4 ) | ( x2 & x47 ) | ( ~x4 & x47 ) ;
  assign n184 = n183 ^ x105 ^ x99 ;
  assign n185 = x31 & ~n184 ;
  assign n186 = n185 ^ x86 ^ 1'b0 ;
  assign n187 = ( x101 & n180 ) | ( x101 & n186 ) | ( n180 & n186 ) ;
  assign n188 = ( x75 & n173 ) | ( x75 & n187 ) | ( n173 & n187 ) ;
  assign n189 = n188 ^ x63 ^ 1'b0 ;
  assign n190 = ( ~n130 & n182 ) | ( ~n130 & n189 ) | ( n182 & n189 ) ;
  assign n191 = n133 ^ x68 ^ 1'b0 ;
  assign n192 = x64 & ~n191 ;
  assign n193 = x54 & ~n190 ;
  assign n194 = n193 ^ x92 ^ 1'b0 ;
  assign n195 = ( ~x6 & x53 ) | ( ~x6 & x119 ) | ( x53 & x119 ) ;
  assign n196 = n195 ^ x78 ^ x66 ;
  assign n197 = n196 ^ n154 ^ x75 ;
  assign n198 = x101 & n130 ;
  assign n199 = n198 ^ x57 ^ 1'b0 ;
  assign n200 = n199 ^ x102 ^ x69 ;
  assign n201 = x34 ^ x17 ^ x0 ;
  assign n202 = ( x52 & x54 ) | ( x52 & n201 ) | ( x54 & n201 ) ;
  assign n203 = n202 ^ x45 ^ x22 ;
  assign n207 = n140 ^ x93 ^ x53 ;
  assign n205 = ( x20 & x98 ) | ( x20 & n133 ) | ( x98 & n133 ) ;
  assign n204 = ( x76 & x87 ) | ( x76 & ~n183 ) | ( x87 & ~n183 ) ;
  assign n206 = n205 ^ n204 ^ n186 ;
  assign n208 = n207 ^ n206 ^ 1'b0 ;
  assign n209 = n203 | n208 ;
  assign n214 = ( x5 & x80 ) | ( x5 & n207 ) | ( x80 & n207 ) ;
  assign n215 = x78 & n183 ;
  assign n216 = ~x39 & n215 ;
  assign n217 = ( x112 & n214 ) | ( x112 & n216 ) | ( n214 & n216 ) ;
  assign n210 = x60 & x119 ;
  assign n211 = ~x113 & n210 ;
  assign n212 = x101 ^ x95 ^ x72 ;
  assign n213 = ( x86 & n211 ) | ( x86 & ~n212 ) | ( n211 & ~n212 ) ;
  assign n218 = n217 ^ n213 ^ 1'b0 ;
  assign n219 = x70 & n218 ;
  assign n220 = ~x120 & n219 ;
  assign n221 = x36 ^ x29 ^ 1'b0 ;
  assign n222 = x8 & n221 ;
  assign n223 = n222 ^ n145 ^ x126 ;
  assign n224 = n131 ^ x89 ^ 1'b0 ;
  assign n225 = ( x53 & x95 ) | ( x53 & n224 ) | ( x95 & n224 ) ;
  assign n226 = x83 ^ x37 ^ x33 ;
  assign n227 = n225 & ~n226 ;
  assign n228 = x16 ^ x4 ^ 1'b0 ;
  assign n229 = n227 & n228 ;
  assign n230 = ( n195 & n223 ) | ( n195 & ~n229 ) | ( n223 & ~n229 ) ;
  assign n231 = x64 ^ x53 ^ x15 ;
  assign n232 = n231 ^ n130 ^ x5 ;
  assign n233 = n232 ^ x123 ^ 1'b0 ;
  assign n235 = ( x43 & x110 ) | ( x43 & n176 ) | ( x110 & n176 ) ;
  assign n234 = n156 ^ x58 ^ x56 ;
  assign n236 = n235 ^ n234 ^ x28 ;
  assign n237 = n182 ^ x111 ^ x49 ;
  assign n238 = ( ~x89 & n227 ) | ( ~x89 & n237 ) | ( n227 & n237 ) ;
  assign n239 = x43 ^ x29 ^ x13 ;
  assign n240 = ( x39 & n226 ) | ( x39 & n239 ) | ( n226 & n239 ) ;
  assign n241 = ( ~x17 & x55 ) | ( ~x17 & n172 ) | ( x55 & n172 ) ;
  assign n242 = ( n184 & n240 ) | ( n184 & n241 ) | ( n240 & n241 ) ;
  assign n243 = x55 ^ x52 ^ x8 ;
  assign n244 = x78 & ~n243 ;
  assign n245 = n244 ^ n145 ^ 1'b0 ;
  assign n246 = x103 & ~n211 ;
  assign n247 = ~x3 & n246 ;
  assign n248 = n247 ^ n194 ^ x105 ;
  assign n249 = x63 & ~n248 ;
  assign n250 = ~x94 & n249 ;
  assign n251 = ( x53 & n245 ) | ( x53 & ~n250 ) | ( n245 & ~n250 ) ;
  assign n252 = ( x8 & x45 ) | ( x8 & ~x61 ) | ( x45 & ~x61 ) ;
  assign n253 = n252 ^ x41 ^ x9 ;
  assign n263 = x111 ^ x33 ^ 1'b0 ;
  assign n264 = x89 & n263 ;
  assign n262 = x34 & n237 ;
  assign n265 = n264 ^ n262 ^ 1'b0 ;
  assign n254 = x118 & n232 ;
  assign n255 = ~x13 & n254 ;
  assign n256 = ( x87 & n158 ) | ( x87 & n255 ) | ( n158 & n255 ) ;
  assign n257 = x51 ^ x9 ^ 1'b0 ;
  assign n258 = x96 & n257 ;
  assign n259 = ( n213 & n256 ) | ( n213 & n258 ) | ( n256 & n258 ) ;
  assign n260 = n259 ^ n182 ^ x70 ;
  assign n261 = n260 ^ n256 ^ n131 ;
  assign n266 = n265 ^ n261 ^ x43 ;
  assign n269 = ( ~n143 & n160 ) | ( ~n143 & n177 ) | ( n160 & n177 ) ;
  assign n267 = ( x31 & x76 ) | ( x31 & ~n237 ) | ( x76 & ~n237 ) ;
  assign n268 = n240 | n267 ;
  assign n270 = n269 ^ n268 ^ x48 ;
  assign n271 = ( x8 & x93 ) | ( x8 & ~n270 ) | ( x93 & ~n270 ) ;
  assign n272 = ( x76 & n205 ) | ( x76 & ~n270 ) | ( n205 & ~n270 ) ;
  assign n273 = ( x119 & x123 ) | ( x119 & n253 ) | ( x123 & n253 ) ;
  assign n274 = x87 & x96 ;
  assign n275 = n274 ^ x5 ^ 1'b0 ;
  assign n276 = x17 & x106 ;
  assign n277 = n276 ^ x70 ^ 1'b0 ;
  assign n278 = ( x54 & n201 ) | ( x54 & ~n277 ) | ( n201 & ~n277 ) ;
  assign n279 = x5 & n278 ;
  assign n280 = n275 & n279 ;
  assign n281 = n217 & ~n280 ;
  assign n282 = ~n204 & n281 ;
  assign n283 = x45 & ~n282 ;
  assign n284 = ~x57 & n283 ;
  assign n285 = n284 ^ n187 ^ x96 ;
  assign n288 = x118 ^ x94 ^ x72 ;
  assign n286 = ~n153 & n178 ;
  assign n287 = n190 & n286 ;
  assign n289 = n288 ^ n287 ^ 1'b0 ;
  assign n290 = ~x103 & n144 ;
  assign n291 = ( n132 & ~n140 ) | ( n132 & n290 ) | ( ~n140 & n290 ) ;
  assign n292 = n291 ^ x120 ^ 1'b0 ;
  assign n293 = x92 ^ x88 ^ x62 ;
  assign n294 = ( x58 & x89 ) | ( x58 & ~x97 ) | ( x89 & ~x97 ) ;
  assign n295 = n294 ^ n179 ^ x100 ;
  assign n296 = ( n140 & n293 ) | ( n140 & ~n295 ) | ( n293 & ~n295 ) ;
  assign n297 = x108 ^ x53 ^ 1'b0 ;
  assign n298 = x31 & n297 ;
  assign n299 = n298 ^ n227 ^ 1'b0 ;
  assign n300 = x102 & n299 ;
  assign n301 = x66 ^ x37 ^ x16 ;
  assign n302 = n238 & ~n301 ;
  assign n303 = ~x87 & n302 ;
  assign n304 = x19 | n265 ;
  assign n305 = ( x48 & n290 ) | ( x48 & ~n304 ) | ( n290 & ~n304 ) ;
  assign n306 = ( x49 & ~x98 ) | ( x49 & n148 ) | ( ~x98 & n148 ) ;
  assign n307 = x39 & x107 ;
  assign n308 = n307 ^ x74 ^ 1'b0 ;
  assign n309 = n292 & ~n308 ;
  assign n310 = ~x10 & n309 ;
  assign n311 = n306 & ~n310 ;
  assign n312 = ~x47 & n311 ;
  assign n313 = x55 & ~n132 ;
  assign n314 = n313 ^ n199 ^ x81 ;
  assign n315 = x124 ^ x116 ^ x55 ;
  assign n316 = x4 & ~n315 ;
  assign n317 = n211 & n316 ;
  assign n318 = x107 & ~n317 ;
  assign n319 = ~x29 & n318 ;
  assign n320 = x17 & n319 ;
  assign n321 = n136 ^ x99 ^ x46 ;
  assign n322 = ( n173 & n209 ) | ( n173 & n321 ) | ( n209 & n321 ) ;
  assign n323 = x85 & n322 ;
  assign n324 = n323 ^ x43 ^ 1'b0 ;
  assign n325 = ( x27 & n143 ) | ( x27 & ~n324 ) | ( n143 & ~n324 ) ;
  assign n326 = ( x32 & x105 ) | ( x32 & ~x108 ) | ( x105 & ~x108 ) ;
  assign n327 = n201 ^ n173 ^ 1'b0 ;
  assign n328 = n326 & ~n327 ;
  assign n329 = ( x95 & n156 ) | ( x95 & n328 ) | ( n156 & n328 ) ;
  assign n330 = ( x85 & n212 ) | ( x85 & ~n329 ) | ( n212 & ~n329 ) ;
  assign n334 = ( ~x6 & x95 ) | ( ~x6 & n237 ) | ( x95 & n237 ) ;
  assign n331 = ( ~x26 & x40 ) | ( ~x26 & x73 ) | ( x40 & x73 ) ;
  assign n332 = ( x9 & ~x103 ) | ( x9 & n331 ) | ( ~x103 & n331 ) ;
  assign n333 = ( ~x18 & x119 ) | ( ~x18 & n332 ) | ( x119 & n332 ) ;
  assign n335 = n334 ^ n333 ^ x120 ;
  assign n336 = n143 | n335 ;
  assign n337 = x106 & ~n336 ;
  assign n338 = ~n330 & n337 ;
  assign n339 = ~x92 & n338 ;
  assign n340 = n163 ^ n158 ^ x88 ;
  assign n341 = n151 ^ x98 ^ x57 ;
  assign n342 = n341 ^ n235 ^ x26 ;
  assign n343 = x45 & ~n342 ;
  assign n344 = ( n144 & n340 ) | ( n144 & n343 ) | ( n340 & n343 ) ;
  assign n345 = ( n183 & n234 ) | ( n183 & n293 ) | ( n234 & n293 ) ;
  assign n347 = n243 ^ n224 ^ n141 ;
  assign n348 = ( ~x65 & n190 ) | ( ~x65 & n347 ) | ( n190 & n347 ) ;
  assign n349 = ( n192 & ~n203 ) | ( n192 & n348 ) | ( ~n203 & n348 ) ;
  assign n346 = x67 & ~x124 ;
  assign n350 = n349 ^ n346 ^ x99 ;
  assign n354 = n226 ^ x88 ^ x58 ;
  assign n353 = n144 ^ x89 ^ x14 ;
  assign n355 = n354 ^ n353 ^ n294 ;
  assign n351 = x85 & ~n239 ;
  assign n352 = n176 & n351 ;
  assign n356 = n355 ^ n352 ^ n151 ;
  assign n357 = ( x123 & n131 ) | ( x123 & n356 ) | ( n131 & n356 ) ;
  assign n365 = n331 ^ n141 ^ x57 ;
  assign n363 = x14 & x85 ;
  assign n364 = ~x123 & n363 ;
  assign n358 = x44 & x69 ;
  assign n359 = ~n146 & n358 ;
  assign n360 = x70 ^ x50 ^ x35 ;
  assign n361 = n360 ^ x69 ^ 1'b0 ;
  assign n362 = n359 | n361 ;
  assign n366 = n365 ^ n364 ^ n362 ;
  assign n367 = n366 ^ n266 ^ n241 ;
  assign n368 = x26 & x28 ;
  assign n369 = n368 ^ x123 ^ 1'b0 ;
  assign n370 = n369 ^ n186 ^ x65 ;
  assign n371 = ( x91 & n148 ) | ( x91 & n370 ) | ( n148 & n370 ) ;
  assign n372 = x113 ^ x66 ^ x62 ;
  assign n373 = n372 ^ x89 ^ 1'b0 ;
  assign n374 = ( x31 & ~n371 ) | ( x31 & n373 ) | ( ~n371 & n373 ) ;
  assign n375 = x119 ^ x79 ^ x56 ;
  assign n376 = n234 & n326 ;
  assign n377 = n376 ^ n212 ^ 1'b0 ;
  assign n378 = ( n186 & ~n375 ) | ( n186 & n377 ) | ( ~n375 & n377 ) ;
  assign n379 = x99 ^ x50 ^ x34 ;
  assign n380 = x10 & ~n146 ;
  assign n381 = x104 & n326 ;
  assign n382 = ~x107 & n381 ;
  assign n383 = ( ~x48 & n189 ) | ( ~x48 & n382 ) | ( n189 & n382 ) ;
  assign n384 = n383 ^ n170 ^ x66 ;
  assign n385 = ( ~x7 & n252 ) | ( ~x7 & n384 ) | ( n252 & n384 ) ;
  assign n386 = ( n379 & ~n380 ) | ( n379 & n385 ) | ( ~n380 & n385 ) ;
  assign n388 = x106 & ~n167 ;
  assign n387 = n180 ^ x109 ^ x1 ;
  assign n389 = n388 ^ n387 ^ n369 ;
  assign n390 = ( x72 & x126 ) | ( x72 & n226 ) | ( x126 & n226 ) ;
  assign n391 = n347 & n390 ;
  assign n392 = n141 & n391 ;
  assign n393 = ( ~x24 & x110 ) | ( ~x24 & n154 ) | ( x110 & n154 ) ;
  assign n394 = n149 ^ x126 ^ x46 ;
  assign n395 = ( n177 & n393 ) | ( n177 & ~n394 ) | ( n393 & ~n394 ) ;
  assign n396 = n395 ^ x29 ^ 1'b0 ;
  assign n397 = ~n335 & n396 ;
  assign n398 = ( n233 & n369 ) | ( n233 & n397 ) | ( n369 & n397 ) ;
  assign n399 = ( x76 & x108 ) | ( x76 & ~x124 ) | ( x108 & ~x124 ) ;
  assign n400 = ( n392 & n398 ) | ( n392 & ~n399 ) | ( n398 & ~n399 ) ;
  assign n401 = n144 ^ n130 ^ 1'b0 ;
  assign n402 = x89 & n401 ;
  assign n403 = ( x45 & n237 ) | ( x45 & ~n402 ) | ( n237 & ~n402 ) ;
  assign n404 = x59 & n403 ;
  assign n405 = n400 & n404 ;
  assign n406 = ( ~n159 & n226 ) | ( ~n159 & n372 ) | ( n226 & n372 ) ;
  assign n407 = n406 ^ n202 ^ n153 ;
  assign n413 = n331 ^ n226 ^ x17 ;
  assign n408 = n157 ^ x19 ^ x0 ;
  assign n409 = x82 ^ x49 ^ x27 ;
  assign n410 = n408 & ~n409 ;
  assign n411 = ( ~x27 & x103 ) | ( ~x27 & n410 ) | ( x103 & n410 ) ;
  assign n412 = x67 & n411 ;
  assign n414 = n413 ^ n412 ^ 1'b0 ;
  assign n415 = ( x60 & n312 ) | ( x60 & n414 ) | ( n312 & n414 ) ;
  assign n416 = x116 ^ x34 ^ 1'b0 ;
  assign n417 = ( x56 & ~n143 ) | ( x56 & n416 ) | ( ~n143 & n416 ) ;
  assign n418 = n319 ^ n280 ^ x52 ;
  assign n419 = n418 ^ n242 ^ 1'b0 ;
  assign n420 = n417 & n419 ;
  assign n421 = x92 ^ x75 ^ x3 ;
  assign n422 = n379 | n421 ;
  assign n423 = x41 | n422 ;
  assign n424 = n293 & n423 ;
  assign n425 = n129 ^ x4 ^ 1'b0 ;
  assign n426 = ( n212 & n424 ) | ( n212 & n425 ) | ( n424 & n425 ) ;
  assign n427 = x117 & n417 ;
  assign n428 = n364 & n427 ;
  assign n429 = ( x65 & n392 ) | ( x65 & ~n428 ) | ( n392 & ~n428 ) ;
  assign n430 = ( n133 & ~n247 ) | ( n133 & n421 ) | ( ~n247 & n421 ) ;
  assign n431 = x48 & n195 ;
  assign n432 = n431 ^ n133 ^ 1'b0 ;
  assign n433 = n432 ^ x95 ^ 1'b0 ;
  assign n434 = ( n280 & n430 ) | ( n280 & n433 ) | ( n430 & n433 ) ;
  assign n435 = n260 ^ n141 ^ 1'b0 ;
  assign n436 = n435 ^ n408 ^ 1'b0 ;
  assign n440 = ( x100 & x112 ) | ( x100 & ~x115 ) | ( x112 & ~x115 ) ;
  assign n438 = n133 | n201 ;
  assign n439 = n438 ^ n214 ^ 1'b0 ;
  assign n441 = n440 ^ n439 ^ n348 ;
  assign n437 = x112 & n355 ;
  assign n442 = n441 ^ n437 ^ 1'b0 ;
  assign n443 = n175 ^ n137 ^ x45 ;
  assign n444 = ( x77 & n360 ) | ( x77 & n443 ) | ( n360 & n443 ) ;
  assign n445 = n444 ^ n424 ^ x54 ;
  assign n456 = ( x3 & ~n204 ) | ( x3 & n234 ) | ( ~n204 & n234 ) ;
  assign n457 = ~n372 & n456 ;
  assign n448 = n158 ^ x121 ^ 1'b0 ;
  assign n449 = n179 ^ x117 ^ x70 ;
  assign n450 = n449 ^ n225 ^ 1'b0 ;
  assign n451 = x70 & ~n450 ;
  assign n452 = n451 ^ n230 ^ 1'b0 ;
  assign n453 = n202 & ~n452 ;
  assign n454 = n453 ^ x78 ^ 1'b0 ;
  assign n455 = ~n448 & n454 ;
  assign n446 = x12 & x45 ;
  assign n447 = ~x85 & n446 ;
  assign n458 = n457 ^ n455 ^ n447 ;
  assign n459 = n232 ^ x125 ^ x123 ;
  assign n460 = ( x31 & ~n229 ) | ( x31 & n459 ) | ( ~n229 & n459 ) ;
  assign n461 = x62 | n369 ;
  assign n462 = n461 ^ n273 ^ 1'b0 ;
  assign n463 = ( x93 & n223 ) | ( x93 & n284 ) | ( n223 & n284 ) ;
  assign n464 = ( x44 & n385 ) | ( x44 & n463 ) | ( n385 & n463 ) ;
  assign n474 = x3 & ~n416 ;
  assign n475 = n277 & n474 ;
  assign n465 = ( x75 & n140 ) | ( x75 & ~n214 ) | ( n140 & ~n214 ) ;
  assign n466 = ( ~x36 & n216 ) | ( ~x36 & n365 ) | ( n216 & n365 ) ;
  assign n467 = n432 | n466 ;
  assign n469 = n239 ^ n157 ^ x42 ;
  assign n470 = n469 ^ x31 ^ 1'b0 ;
  assign n471 = x78 & ~n470 ;
  assign n468 = n421 ^ n220 ^ x119 ;
  assign n472 = n471 ^ n468 ^ x120 ;
  assign n473 = ( n465 & ~n467 ) | ( n465 & n472 ) | ( ~n467 & n472 ) ;
  assign n476 = n475 ^ n473 ^ x38 ;
  assign n477 = n334 & ~n456 ;
  assign n479 = ( x26 & n225 ) | ( x26 & n315 ) | ( n225 & n315 ) ;
  assign n478 = n132 & ~n377 ;
  assign n480 = n479 ^ n478 ^ n467 ;
  assign n481 = n140 ^ x121 ^ 1'b0 ;
  assign n482 = x79 & n481 ;
  assign n483 = x61 & ~n359 ;
  assign n484 = ~x51 & n483 ;
  assign n485 = ( x13 & ~x49 ) | ( x13 & x85 ) | ( ~x49 & x85 ) ;
  assign n486 = n485 ^ n342 ^ n217 ;
  assign n487 = n366 & n486 ;
  assign n488 = n487 ^ n399 ^ x13 ;
  assign n489 = ( n482 & n484 ) | ( n482 & n488 ) | ( n484 & n488 ) ;
  assign n490 = n365 ^ n234 ^ x30 ;
  assign n491 = ( n239 & n329 ) | ( n239 & ~n490 ) | ( n329 & ~n490 ) ;
  assign n492 = n334 ^ x82 ^ 1'b0 ;
  assign n493 = ~n153 & n492 ;
  assign n494 = n493 ^ n203 ^ 1'b0 ;
  assign n496 = n432 ^ n232 ^ x95 ;
  assign n495 = n451 ^ x69 ^ x53 ;
  assign n497 = n496 ^ n495 ^ 1'b0 ;
  assign n499 = x42 & ~n164 ;
  assign n498 = ( x10 & x113 ) | ( x10 & ~n183 ) | ( x113 & ~n183 ) ;
  assign n500 = n499 ^ n498 ^ n159 ;
  assign n501 = n192 & ~n461 ;
  assign n502 = n501 ^ n230 ^ 1'b0 ;
  assign n503 = x109 & n245 ;
  assign n504 = n502 & ~n503 ;
  assign n505 = ~n500 & n504 ;
  assign n506 = n304 ^ n240 ^ 1'b0 ;
  assign n507 = n505 | n506 ;
  assign n508 = ( ~n425 & n497 ) | ( ~n425 & n507 ) | ( n497 & n507 ) ;
  assign n509 = ( x38 & ~x39 ) | ( x38 & n369 ) | ( ~x39 & n369 ) ;
  assign n510 = ( n290 & ~n356 ) | ( n290 & n509 ) | ( ~n356 & n509 ) ;
  assign n511 = n510 ^ n271 ^ 1'b0 ;
  assign n512 = n268 ^ x59 ^ 1'b0 ;
  assign n513 = x47 & ~n512 ;
  assign n515 = x36 & x77 ;
  assign n516 = ~x116 & n515 ;
  assign n514 = n456 ^ x107 ^ x104 ;
  assign n517 = n516 ^ n514 ^ n240 ;
  assign n518 = ( n141 & n513 ) | ( n141 & n517 ) | ( n513 & n517 ) ;
  assign n526 = x101 ^ x41 ^ x19 ;
  assign n519 = n165 & n177 ;
  assign n520 = n519 ^ n326 ^ 1'b0 ;
  assign n521 = n520 ^ n432 ^ n359 ;
  assign n522 = x105 & ~n521 ;
  assign n523 = n522 ^ n255 ^ 1'b0 ;
  assign n524 = n523 ^ n471 ^ n207 ;
  assign n525 = ( n157 & ~n310 ) | ( n157 & n524 ) | ( ~n310 & n524 ) ;
  assign n527 = n526 ^ n525 ^ 1'b0 ;
  assign n528 = n518 & ~n527 ;
  assign n544 = n329 ^ x21 ^ 1'b0 ;
  assign n529 = x100 ^ x65 ^ 1'b0 ;
  assign n530 = ~n516 & n529 ;
  assign n531 = ~n453 & n530 ;
  assign n532 = n375 | n531 ;
  assign n533 = n220 & ~n532 ;
  assign n540 = n243 ^ n167 ^ x21 ;
  assign n541 = n163 & ~n540 ;
  assign n534 = n247 ^ x109 ^ 1'b0 ;
  assign n535 = x102 & ~n534 ;
  assign n536 = n146 & n535 ;
  assign n537 = n136 & n536 ;
  assign n538 = x91 | n537 ;
  assign n539 = x20 & ~n538 ;
  assign n542 = n541 ^ n539 ^ 1'b0 ;
  assign n543 = n533 & ~n542 ;
  assign n545 = n544 ^ n543 ^ x31 ;
  assign n546 = n545 ^ n378 ^ 1'b0 ;
  assign n547 = ~n141 & n546 ;
  assign n548 = ( x28 & ~n224 ) | ( x28 & n247 ) | ( ~n224 & n247 ) ;
  assign n549 = n548 ^ n187 ^ n156 ;
  assign n550 = n469 | n531 ;
  assign n551 = n550 ^ x52 ^ 1'b0 ;
  assign n552 = n551 ^ n386 ^ x52 ;
  assign n553 = ( x77 & n549 ) | ( x77 & ~n552 ) | ( n549 & ~n552 ) ;
  assign n554 = n203 ^ n140 ^ 1'b0 ;
  assign n555 = n146 & ~n554 ;
  assign n556 = n478 ^ n328 ^ x73 ;
  assign n557 = ~n131 & n556 ;
  assign n558 = ( ~x32 & n195 ) | ( ~x32 & n557 ) | ( n195 & n557 ) ;
  assign n559 = ( n139 & n319 ) | ( n139 & n558 ) | ( n319 & n558 ) ;
  assign n560 = n448 ^ x52 ^ 1'b0 ;
  assign n561 = n292 & ~n560 ;
  assign n562 = ( x53 & x89 ) | ( x53 & n275 ) | ( x89 & n275 ) ;
  assign n563 = ( ~n205 & n510 ) | ( ~n205 & n562 ) | ( n510 & n562 ) ;
  assign n570 = ~n243 & n272 ;
  assign n571 = n570 ^ n377 ^ 1'b0 ;
  assign n572 = n571 ^ x36 ^ x13 ;
  assign n569 = x39 & n192 ;
  assign n564 = ( x61 & ~x73 ) | ( x61 & x107 ) | ( ~x73 & x107 ) ;
  assign n565 = n564 ^ n417 ^ n410 ;
  assign n566 = n565 ^ n234 ^ n214 ;
  assign n567 = ( ~x97 & n255 ) | ( ~x97 & n566 ) | ( n255 & n566 ) ;
  assign n568 = n567 ^ n235 ^ x70 ;
  assign n573 = n572 ^ n569 ^ n568 ;
  assign n574 = n349 ^ n342 ^ 1'b0 ;
  assign n575 = n423 & ~n574 ;
  assign n576 = n575 ^ n354 ^ 1'b0 ;
  assign n577 = ( x94 & n573 ) | ( x94 & ~n576 ) | ( n573 & ~n576 ) ;
  assign n578 = ( ~x91 & n341 ) | ( ~x91 & n577 ) | ( n341 & n577 ) ;
  assign n587 = n493 ^ n202 ^ x44 ;
  assign n588 = ( n148 & n212 ) | ( n148 & ~n587 ) | ( n212 & ~n587 ) ;
  assign n589 = n588 ^ n368 ^ 1'b0 ;
  assign n590 = x40 & ~n549 ;
  assign n591 = n590 ^ n293 ^ 1'b0 ;
  assign n592 = n591 ^ n250 ^ x15 ;
  assign n593 = ( ~n487 & n589 ) | ( ~n487 & n592 ) | ( n589 & n592 ) ;
  assign n585 = ( x113 & n319 ) | ( x113 & n398 ) | ( n319 & n398 ) ;
  assign n580 = n199 ^ x44 ^ x20 ;
  assign n581 = n580 ^ n132 ^ x103 ;
  assign n582 = ( ~n180 & n192 ) | ( ~n180 & n421 ) | ( n192 & n421 ) ;
  assign n583 = ( n409 & n581 ) | ( n409 & n582 ) | ( n581 & n582 ) ;
  assign n579 = ~n346 & n439 ;
  assign n584 = n583 ^ n579 ^ 1'b0 ;
  assign n586 = n585 ^ n584 ^ 1'b0 ;
  assign n594 = n593 ^ n586 ^ 1'b0 ;
  assign n599 = x29 & n137 ;
  assign n600 = n379 & n599 ;
  assign n595 = x52 & n564 ;
  assign n596 = ~x30 & n595 ;
  assign n597 = n596 ^ n399 ^ 1'b0 ;
  assign n598 = ( ~x44 & n371 ) | ( ~x44 & n597 ) | ( n371 & n597 ) ;
  assign n601 = n600 ^ n598 ^ 1'b0 ;
  assign n602 = n223 | n601 ;
  assign n603 = n265 ^ n180 ^ x125 ;
  assign n604 = n603 ^ n294 ^ n202 ;
  assign n605 = n604 ^ n163 ^ x52 ;
  assign n607 = n580 ^ n288 ^ x119 ;
  assign n606 = x46 & x101 ;
  assign n608 = n607 ^ n606 ^ 1'b0 ;
  assign n609 = ~n133 & n608 ;
  assign n610 = ~n133 & n517 ;
  assign n611 = ~x32 & n610 ;
  assign n612 = n204 & ~n611 ;
  assign n613 = n612 ^ n305 ^ 1'b0 ;
  assign n614 = ( x112 & n609 ) | ( x112 & n613 ) | ( n609 & n613 ) ;
  assign n619 = n264 ^ n159 ^ 1'b0 ;
  assign n620 = n619 ^ n200 ^ n178 ;
  assign n621 = x18 & x78 ;
  assign n622 = n199 & n621 ;
  assign n623 = n238 ^ n172 ^ x122 ;
  assign n624 = n623 ^ n231 ^ n165 ;
  assign n625 = n622 | n624 ;
  assign n626 = n131 & ~n625 ;
  assign n627 = n411 ^ n341 ^ n243 ;
  assign n628 = ( n304 & n626 ) | ( n304 & n627 ) | ( n626 & n627 ) ;
  assign n629 = ( n478 & n620 ) | ( n478 & n628 ) | ( n620 & n628 ) ;
  assign n615 = x13 & ~n231 ;
  assign n616 = n615 ^ x41 ^ 1'b0 ;
  assign n617 = n616 ^ x84 ^ x6 ;
  assign n618 = ~n468 & n617 ;
  assign n630 = n629 ^ n618 ^ 1'b0 ;
  assign n632 = ( ~x12 & x54 ) | ( ~x12 & x80 ) | ( x54 & x80 ) ;
  assign n633 = n632 ^ x59 ^ 1'b0 ;
  assign n631 = n300 & n365 ;
  assign n634 = n633 ^ n631 ^ n319 ;
  assign n635 = ( ~n145 & n199 ) | ( ~n145 & n252 ) | ( n199 & n252 ) ;
  assign n636 = ( x0 & x50 ) | ( x0 & ~n402 ) | ( x50 & ~n402 ) ;
  assign n637 = ( n477 & n635 ) | ( n477 & n636 ) | ( n635 & n636 ) ;
  assign n643 = n130 ^ x93 ^ x75 ;
  assign n644 = n566 & n643 ;
  assign n638 = x78 ^ x75 ^ x31 ;
  assign n639 = ( n395 & ~n486 ) | ( n395 & n638 ) | ( ~n486 & n638 ) ;
  assign n640 = n322 | n639 ;
  assign n641 = ( n158 & n356 ) | ( n158 & n640 ) | ( n356 & n640 ) ;
  assign n642 = x21 & n641 ;
  assign n645 = n644 ^ n642 ^ n563 ;
  assign n647 = ( n151 & n175 ) | ( n151 & n493 ) | ( n175 & n493 ) ;
  assign n646 = ( n207 & n476 ) | ( n207 & ~n533 ) | ( n476 & ~n533 ) ;
  assign n648 = n647 ^ n646 ^ 1'b0 ;
  assign n649 = n417 ^ n184 ^ x43 ;
  assign n650 = n649 ^ n301 ^ n247 ;
  assign n651 = ( ~x78 & x113 ) | ( ~x78 & n129 ) | ( x113 & n129 ) ;
  assign n652 = x124 & ~n317 ;
  assign n653 = ~n222 & n652 ;
  assign n654 = n506 ^ x127 ^ 1'b0 ;
  assign n655 = n469 | n654 ;
  assign n656 = x47 & ~n616 ;
  assign n657 = n655 & n656 ;
  assign n663 = ( ~n132 & n184 ) | ( ~n132 & n321 ) | ( n184 & n321 ) ;
  assign n664 = n663 ^ n143 ^ x61 ;
  assign n658 = n432 ^ n291 ^ n231 ;
  assign n659 = n658 ^ n626 ^ n277 ;
  assign n660 = x15 & ~n659 ;
  assign n661 = ~n513 & n660 ;
  assign n662 = ( n347 & n624 ) | ( n347 & n661 ) | ( n624 & n661 ) ;
  assign n665 = n664 ^ n662 ^ n343 ;
  assign n666 = n270 | n665 ;
  assign n667 = ( n353 & n566 ) | ( n353 & ~n666 ) | ( n566 & ~n666 ) ;
  assign n668 = n667 ^ n455 ^ n199 ;
  assign n669 = n580 ^ n137 ^ x82 ;
  assign n670 = ( ~n214 & n439 ) | ( ~n214 & n503 ) | ( n439 & n503 ) ;
  assign n671 = n433 | n670 ;
  assign n672 = ~n669 & n671 ;
  assign n673 = ~x11 & n672 ;
  assign n674 = x108 & ~n163 ;
  assign n675 = n382 & n674 ;
  assign n676 = n273 | n466 ;
  assign n677 = ( n428 & n675 ) | ( n428 & n676 ) | ( n675 & n676 ) ;
  assign n678 = n377 ^ n328 ^ 1'b0 ;
  assign n679 = ~n677 & n678 ;
  assign n680 = n314 & ~n679 ;
  assign n681 = ( n242 & n359 ) | ( n242 & ~n418 ) | ( n359 & ~n418 ) ;
  assign n683 = n189 ^ x117 ^ 1'b0 ;
  assign n682 = n233 & ~n444 ;
  assign n684 = n683 ^ n682 ^ 1'b0 ;
  assign n685 = ( x14 & ~n133 ) | ( x14 & n684 ) | ( ~n133 & n684 ) ;
  assign n686 = ( n301 & n377 ) | ( n301 & ~n685 ) | ( n377 & ~n685 ) ;
  assign n687 = ( x90 & n267 ) | ( x90 & n538 ) | ( n267 & n538 ) ;
  assign n688 = ( n337 & n686 ) | ( n337 & n687 ) | ( n686 & n687 ) ;
  assign n689 = ( x62 & ~n681 ) | ( x62 & n688 ) | ( ~n681 & n688 ) ;
  assign n690 = n383 ^ x41 ^ 1'b0 ;
  assign n691 = ( n429 & n442 ) | ( n429 & ~n541 ) | ( n442 & ~n541 ) ;
  assign n692 = n467 & ~n508 ;
  assign n693 = n692 ^ x52 ^ 1'b0 ;
  assign n694 = n390 | n693 ;
  assign n695 = n691 | n694 ;
  assign n703 = x126 ^ x83 ^ x53 ;
  assign n702 = n435 ^ x15 ^ x11 ;
  assign n697 = ( x25 & ~x72 ) | ( x25 & n521 ) | ( ~x72 & n521 ) ;
  assign n698 = n580 ^ n290 ^ 1'b0 ;
  assign n699 = ( x84 & n290 ) | ( x84 & ~n698 ) | ( n290 & ~n698 ) ;
  assign n700 = ( n300 & n697 ) | ( n300 & n699 ) | ( n697 & n699 ) ;
  assign n696 = n319 ^ x46 ^ 1'b0 ;
  assign n701 = n700 ^ n696 ^ x47 ;
  assign n704 = n703 ^ n702 ^ n701 ;
  assign n708 = n375 ^ x68 ^ 1'b0 ;
  assign n705 = ( n408 & n542 ) | ( n408 & n580 ) | ( n542 & n580 ) ;
  assign n706 = n705 ^ n664 ^ 1'b0 ;
  assign n707 = n306 & ~n706 ;
  assign n709 = n708 ^ n707 ^ 1'b0 ;
  assign n710 = ( ~x5 & x113 ) | ( ~x5 & n206 ) | ( x113 & n206 ) ;
  assign n711 = ( n473 & ~n597 ) | ( n473 & n710 ) | ( ~n597 & n710 ) ;
  assign n713 = n343 ^ x88 ^ 1'b0 ;
  assign n714 = x59 & ~n211 ;
  assign n715 = ~n713 & n714 ;
  assign n712 = x109 & x127 ;
  assign n716 = n715 ^ n712 ^ 1'b0 ;
  assign n717 = n354 & n716 ;
  assign n718 = n717 ^ n559 ^ 1'b0 ;
  assign n721 = n328 & ~n496 ;
  assign n722 = ( x35 & n317 ) | ( x35 & ~n721 ) | ( n317 & ~n721 ) ;
  assign n719 = n600 ^ n397 ^ x39 ;
  assign n720 = n328 & n719 ;
  assign n723 = n722 ^ n720 ^ 1'b0 ;
  assign n724 = n723 ^ n348 ^ 1'b0 ;
  assign n725 = x48 & ~n503 ;
  assign n727 = n204 & n354 ;
  assign n728 = n727 ^ n499 ^ 1'b0 ;
  assign n726 = x49 & n636 ;
  assign n729 = n728 ^ n726 ^ 1'b0 ;
  assign n730 = n354 ^ n234 ^ 1'b0 ;
  assign n731 = ~n729 & n730 ;
  assign n732 = n418 | n603 ;
  assign n733 = n732 ^ n685 ^ 1'b0 ;
  assign n734 = n632 ^ n269 ^ x41 ;
  assign n735 = n734 ^ n650 ^ n390 ;
  assign n736 = n497 & n568 ;
  assign n737 = ~n408 & n736 ;
  assign n742 = ~x125 & n486 ;
  assign n743 = n742 ^ n409 ^ x30 ;
  assign n739 = n319 ^ x106 ^ x96 ;
  assign n740 = n739 ^ x11 ^ x2 ;
  assign n741 = n352 & ~n740 ;
  assign n738 = ( n180 & n399 ) | ( n180 & n665 ) | ( n399 & n665 ) ;
  assign n744 = n743 ^ n741 ^ n738 ;
  assign n745 = ( x16 & n277 ) | ( x16 & ~n298 ) | ( n277 & ~n298 ) ;
  assign n746 = ( x22 & n135 ) | ( x22 & n745 ) | ( n135 & n745 ) ;
  assign n747 = n746 ^ n265 ^ 1'b0 ;
  assign n748 = n441 & ~n747 ;
  assign n749 = ~n201 & n233 ;
  assign n750 = ~n627 & n749 ;
  assign n751 = n750 ^ n738 ^ x72 ;
  assign n752 = n751 ^ n448 ^ 1'b0 ;
  assign n753 = n748 & n752 ;
  assign n754 = ~n409 & n753 ;
  assign n757 = ( ~x14 & n190 ) | ( ~x14 & n341 ) | ( n190 & n341 ) ;
  assign n758 = n757 ^ x122 ^ x9 ;
  assign n755 = ( ~x57 & x125 ) | ( ~x57 & n183 ) | ( x125 & n183 ) ;
  assign n756 = ~n626 & n755 ;
  assign n759 = n758 ^ n756 ^ 1'b0 ;
  assign n765 = n225 & n294 ;
  assign n766 = ~n140 & n765 ;
  assign n761 = n132 ^ x14 ^ 1'b0 ;
  assign n760 = ( ~x14 & x81 ) | ( ~x14 & n278 ) | ( x81 & n278 ) ;
  assign n762 = n761 ^ n760 ^ n360 ;
  assign n763 = n461 ^ n133 ^ x36 ;
  assign n764 = n762 & ~n763 ;
  assign n767 = n766 ^ n764 ^ 1'b0 ;
  assign n768 = ( x21 & x116 ) | ( x21 & ~x122 ) | ( x116 & ~x122 ) ;
  assign n769 = n342 ^ n272 ^ 1'b0 ;
  assign n770 = n768 & ~n769 ;
  assign n771 = n770 ^ n426 ^ n407 ;
  assign n772 = n130 & ~n516 ;
  assign n773 = n211 & n772 ;
  assign n774 = n773 ^ n287 ^ x116 ;
  assign n776 = x81 & n214 ;
  assign n777 = n776 ^ x96 ^ 1'b0 ;
  assign n775 = n643 ^ n355 ^ x83 ;
  assign n778 = n777 ^ n775 ^ n206 ;
  assign n779 = ~n642 & n734 ;
  assign n780 = ( x54 & n265 ) | ( x54 & ~n572 ) | ( n265 & ~n572 ) ;
  assign n781 = ~n346 & n695 ;
  assign n782 = n780 & n781 ;
  assign n783 = n178 ^ x105 ^ x33 ;
  assign n784 = n207 | n783 ;
  assign n785 = n775 ^ n503 ^ n416 ;
  assign n786 = n768 ^ x54 ^ 1'b0 ;
  assign n787 = n241 & n786 ;
  assign n788 = n453 & n787 ;
  assign n789 = ~x52 & n788 ;
  assign n790 = x46 & x116 ;
  assign n791 = n790 ^ n387 ^ 1'b0 ;
  assign n792 = n465 & n588 ;
  assign n793 = n792 ^ x54 ^ 1'b0 ;
  assign n794 = ( n584 & ~n791 ) | ( n584 & n793 ) | ( ~n791 & n793 ) ;
  assign n795 = ( x23 & n304 ) | ( x23 & ~n713 ) | ( n304 & ~n713 ) ;
  assign n796 = n795 ^ x62 ^ 1'b0 ;
  assign n797 = n734 ^ n207 ^ 1'b0 ;
  assign n798 = x81 & n797 ;
  assign n805 = ( n206 & ~n278 ) | ( n206 & n379 ) | ( ~n278 & n379 ) ;
  assign n801 = n317 & ~n487 ;
  assign n799 = n616 ^ n398 ^ x50 ;
  assign n800 = n332 & n799 ;
  assign n802 = n801 ^ n800 ^ 1'b0 ;
  assign n803 = x34 & ~n449 ;
  assign n804 = ~n802 & n803 ;
  assign n806 = n805 ^ n804 ^ 1'b0 ;
  assign n807 = ~n301 & n806 ;
  assign n808 = ( n201 & n670 ) | ( n201 & n696 ) | ( n670 & n696 ) ;
  assign n809 = ~n807 & n808 ;
  assign n810 = x26 & ~n567 ;
  assign n811 = ~n514 & n585 ;
  assign n812 = ( x52 & n207 ) | ( x52 & n581 ) | ( n207 & n581 ) ;
  assign n813 = ( x15 & ~n540 ) | ( x15 & n812 ) | ( ~n540 & n812 ) ;
  assign n814 = ( ~n632 & n748 ) | ( ~n632 & n813 ) | ( n748 & n813 ) ;
  assign n815 = ~n449 & n814 ;
  assign n816 = n386 & n815 ;
  assign n817 = n160 | n816 ;
  assign n818 = n817 ^ n197 ^ 1'b0 ;
  assign n819 = n811 & ~n818 ;
  assign n820 = n819 ^ n697 ^ 1'b0 ;
  assign n821 = n820 ^ n562 ^ 1'b0 ;
  assign n822 = n500 & n821 ;
  assign n824 = n373 ^ n239 ^ 1'b0 ;
  assign n825 = n448 | n824 ;
  assign n823 = ( x51 & x73 ) | ( x51 & n780 ) | ( x73 & n780 ) ;
  assign n826 = n825 ^ n823 ^ x91 ;
  assign n827 = n558 ^ n386 ^ n183 ;
  assign n828 = ( x6 & x15 ) | ( x6 & n783 ) | ( x15 & n783 ) ;
  assign n829 = n828 ^ n771 ^ n169 ;
  assign n830 = n616 ^ x57 ^ 1'b0 ;
  assign n831 = n588 & ~n830 ;
  assign n832 = x14 & n831 ;
  assign n833 = n832 ^ n395 ^ 1'b0 ;
  assign n834 = n675 ^ n326 ^ 1'b0 ;
  assign n835 = n833 | n834 ;
  assign n836 = ~n250 & n591 ;
  assign n837 = n312 & n836 ;
  assign n838 = ( x81 & n285 ) | ( x81 & ~n497 ) | ( n285 & ~n497 ) ;
  assign n839 = ( ~n493 & n643 ) | ( ~n493 & n726 ) | ( n643 & n726 ) ;
  assign n840 = n290 ^ n183 ^ n154 ;
  assign n841 = n388 ^ x32 ^ x1 ;
  assign n842 = n841 ^ n414 ^ 1'b0 ;
  assign n843 = n486 & n842 ;
  assign n844 = ( n394 & ~n697 ) | ( n394 & n843 ) | ( ~n697 & n843 ) ;
  assign n845 = ( ~x114 & n840 ) | ( ~x114 & n844 ) | ( n840 & n844 ) ;
  assign n846 = n844 ^ n837 ^ n737 ;
  assign n847 = n557 & ~n584 ;
  assign n848 = ~n434 & n847 ;
  assign n850 = n746 ^ n644 ^ 1'b0 ;
  assign n851 = ( n688 & ~n760 ) | ( n688 & n850 ) | ( ~n760 & n850 ) ;
  assign n849 = ~n385 & n511 ;
  assign n852 = n851 ^ n849 ^ 1'b0 ;
  assign n853 = ~n301 & n809 ;
  assign n854 = ~x100 & n296 ;
  assign n855 = ~n201 & n854 ;
  assign n856 = n565 ^ n478 ^ n371 ;
  assign n857 = n856 ^ n441 ^ 1'b0 ;
  assign n858 = n857 ^ n517 ^ 1'b0 ;
  assign n859 = n465 ^ n390 ^ n319 ;
  assign n860 = ( ~n203 & n757 ) | ( ~n203 & n859 ) | ( n757 & n859 ) ;
  assign n861 = ( ~x102 & n646 ) | ( ~x102 & n659 ) | ( n646 & n659 ) ;
  assign n862 = ( ~x44 & x110 ) | ( ~x44 & n140 ) | ( x110 & n140 ) ;
  assign n863 = n862 ^ n556 ^ n183 ;
  assign n864 = n157 | n863 ;
  assign n865 = ( n533 & n799 ) | ( n533 & ~n864 ) | ( n799 & ~n864 ) ;
  assign n866 = ( n385 & ~n424 ) | ( n385 & n608 ) | ( ~n424 & n608 ) ;
  assign n867 = ( n253 & n578 ) | ( n253 & ~n866 ) | ( n578 & ~n866 ) ;
  assign n868 = n514 ^ n237 ^ 1'b0 ;
  assign n869 = n667 | n868 ;
  assign n870 = ( ~x90 & x92 ) | ( ~x90 & n267 ) | ( x92 & n267 ) ;
  assign n871 = ( ~x126 & n535 ) | ( ~x126 & n870 ) | ( n535 & n870 ) ;
  assign n872 = ~n236 & n871 ;
  assign n873 = n872 ^ x23 ^ 1'b0 ;
  assign n874 = n873 ^ n565 ^ 1'b0 ;
  assign n875 = ~n275 & n874 ;
  assign n876 = n494 & n875 ;
  assign n877 = n876 ^ n165 ^ 1'b0 ;
  assign n878 = n877 ^ x60 ^ 1'b0 ;
  assign n879 = x7 & ~n207 ;
  assign n880 = n879 ^ x14 ^ 1'b0 ;
  assign n881 = ( ~x70 & x76 ) | ( ~x70 & n303 ) | ( x76 & n303 ) ;
  assign n882 = n881 ^ x116 ^ 1'b0 ;
  assign n883 = n880 | n882 ;
  assign n884 = n190 | n670 ;
  assign n885 = n884 ^ x34 ^ 1'b0 ;
  assign n886 = ~n883 & n885 ;
  assign n887 = n886 ^ x89 ^ 1'b0 ;
  assign n888 = n195 & n332 ;
  assign n889 = n888 ^ n200 ^ 1'b0 ;
  assign n892 = ( ~x60 & n239 ) | ( ~x60 & n493 ) | ( n239 & n493 ) ;
  assign n890 = n250 ^ x115 ^ x72 ;
  assign n891 = ( x62 & n659 ) | ( x62 & ~n890 ) | ( n659 & ~n890 ) ;
  assign n893 = n892 ^ n891 ^ 1'b0 ;
  assign n894 = ~n889 & n893 ;
  assign n895 = ~n203 & n894 ;
  assign n896 = ~x41 & n895 ;
  assign n900 = n603 ^ n186 ^ x41 ;
  assign n898 = x17 & ~n341 ;
  assign n899 = n898 ^ n843 ^ 1'b0 ;
  assign n897 = n214 & n509 ;
  assign n901 = n900 ^ n899 ^ n897 ;
  assign n902 = x63 & n362 ;
  assign n903 = n197 | n902 ;
  assign n904 = n903 ^ n212 ^ 1'b0 ;
  assign n905 = ~x57 & n291 ;
  assign n906 = x52 & n905 ;
  assign n907 = ~x24 & n906 ;
  assign n908 = ( ~n153 & n867 ) | ( ~n153 & n907 ) | ( n867 & n907 ) ;
  assign n909 = n190 | n571 ;
  assign n910 = ~n300 & n322 ;
  assign n911 = n910 ^ n252 ^ 1'b0 ;
  assign n912 = n329 & ~n911 ;
  assign n913 = n909 & n912 ;
  assign n914 = ( x85 & n175 ) | ( x85 & n320 ) | ( n175 & n320 ) ;
  assign n915 = n347 & n636 ;
  assign n916 = ~n232 & n915 ;
  assign n917 = n226 ^ x25 ^ 1'b0 ;
  assign n918 = ( n151 & ~n372 ) | ( n151 & n687 ) | ( ~n372 & n687 ) ;
  assign n919 = ( n916 & n917 ) | ( n916 & n918 ) | ( n917 & n918 ) ;
  assign n920 = ( ~x48 & n914 ) | ( ~x48 & n919 ) | ( n914 & n919 ) ;
  assign n921 = ~n913 & n920 ;
  assign n922 = n567 ^ x123 ^ 1'b0 ;
  assign n923 = n379 | n922 ;
  assign n924 = n387 ^ x82 ^ x45 ;
  assign n925 = ( ~n479 & n604 ) | ( ~n479 & n639 ) | ( n604 & n639 ) ;
  assign n926 = ( n398 & n418 ) | ( n398 & ~n925 ) | ( n418 & ~n925 ) ;
  assign n927 = ( n696 & n924 ) | ( n696 & n926 ) | ( n924 & n926 ) ;
  assign n928 = ( x116 & ~n415 ) | ( x116 & n900 ) | ( ~n415 & n900 ) ;
  assign n930 = ( ~x87 & n496 ) | ( ~x87 & n859 ) | ( n496 & n859 ) ;
  assign n929 = n131 | n293 ;
  assign n931 = n930 ^ n929 ^ 1'b0 ;
  assign n932 = ~n211 & n482 ;
  assign n933 = n336 & n932 ;
  assign n941 = n187 | n366 ;
  assign n938 = n158 & n761 ;
  assign n934 = n175 & ~n746 ;
  assign n935 = n934 ^ n639 ^ n190 ;
  assign n936 = n349 & n935 ;
  assign n937 = ~n582 & n936 ;
  assign n939 = n938 ^ n937 ^ 1'b0 ;
  assign n940 = n823 & n939 ;
  assign n942 = n941 ^ n940 ^ n462 ;
  assign n943 = n942 ^ n653 ^ 1'b0 ;
  assign n944 = n476 & n943 ;
  assign n945 = n933 | n944 ;
  assign n949 = n443 ^ x2 ^ 1'b0 ;
  assign n950 = n944 & ~n949 ;
  assign n951 = ~n553 & n950 ;
  assign n952 = n951 ^ n514 ^ 1'b0 ;
  assign n946 = x66 & n467 ;
  assign n947 = n946 ^ n698 ^ 1'b0 ;
  assign n948 = n201 & ~n947 ;
  assign n953 = n952 ^ n948 ^ 1'b0 ;
  assign n961 = n332 ^ n319 ^ 1'b0 ;
  assign n962 = x114 & ~n961 ;
  assign n954 = ( ~x36 & x104 ) | ( ~x36 & n416 ) | ( x104 & n416 ) ;
  assign n955 = ( n272 & n588 ) | ( n272 & n954 ) | ( n588 & n954 ) ;
  assign n956 = ~n830 & n955 ;
  assign n957 = n956 ^ n202 ^ 1'b0 ;
  assign n958 = n252 | n818 ;
  assign n959 = n784 & ~n958 ;
  assign n960 = n957 | n959 ;
  assign n963 = n962 ^ n960 ^ 1'b0 ;
  assign n964 = n289 | n339 ;
  assign n965 = ( x113 & x123 ) | ( x113 & ~n365 ) | ( x123 & ~n365 ) ;
  assign n966 = n965 ^ n930 ^ n697 ;
  assign n967 = ( x109 & n141 ) | ( x109 & n432 ) | ( n141 & n432 ) ;
  assign n968 = x89 & n304 ;
  assign n969 = n209 & n968 ;
  assign n970 = ( n265 & n967 ) | ( n265 & ~n969 ) | ( n967 & ~n969 ) ;
  assign n971 = ( n436 & ~n966 ) | ( n436 & n970 ) | ( ~n966 & n970 ) ;
  assign n972 = n362 ^ x1 ^ 1'b0 ;
  assign n973 = n972 ^ n354 ^ x47 ;
  assign n974 = n394 ^ n331 ^ 1'b0 ;
  assign n975 = n461 | n974 ;
  assign n976 = ( x127 & n645 ) | ( x127 & ~n975 ) | ( n645 & ~n975 ) ;
  assign n977 = ( ~n200 & n328 ) | ( ~n200 & n855 ) | ( n328 & n855 ) ;
  assign n988 = ( x63 & ~n213 ) | ( x63 & n768 ) | ( ~n213 & n768 ) ;
  assign n985 = n217 & ~n638 ;
  assign n986 = n985 ^ n333 ^ 1'b0 ;
  assign n987 = n189 & ~n986 ;
  assign n989 = n988 ^ n987 ^ 1'b0 ;
  assign n980 = x65 ^ x23 ^ 1'b0 ;
  assign n981 = x89 & n980 ;
  assign n982 = x44 & n981 ;
  assign n983 = n982 ^ n334 ^ 1'b0 ;
  assign n978 = x25 & x126 ;
  assign n979 = n978 ^ n947 ^ 1'b0 ;
  assign n984 = n983 ^ n979 ^ x84 ;
  assign n990 = n989 ^ n984 ^ n937 ;
  assign n991 = n941 ^ n585 ^ n184 ;
  assign n992 = n991 ^ x85 ^ 1'b0 ;
  assign n993 = n992 ^ n973 ^ n291 ;
  assign n994 = ( n237 & ~n420 ) | ( n237 & n661 ) | ( ~n420 & n661 ) ;
  assign n995 = n994 ^ n941 ^ n564 ;
  assign n996 = n294 & ~n995 ;
  assign n997 = ( n177 & n247 ) | ( n177 & ~n742 ) | ( n247 & ~n742 ) ;
  assign n998 = ( ~n557 & n953 ) | ( ~n557 & n997 ) | ( n953 & n997 ) ;
  assign n1001 = x91 | n715 ;
  assign n1002 = n371 | n382 ;
  assign n1003 = n1002 ^ n383 ^ 1'b0 ;
  assign n1004 = ( n172 & n1001 ) | ( n172 & ~n1003 ) | ( n1001 & ~n1003 ) ;
  assign n999 = n306 & ~n669 ;
  assign n1000 = n999 ^ n665 ^ 1'b0 ;
  assign n1005 = n1004 ^ n1000 ^ 1'b0 ;
  assign n1006 = n702 ^ x122 ^ 1'b0 ;
  assign n1007 = ~n1005 & n1006 ;
  assign n1008 = ~n616 & n1007 ;
  assign n1009 = ~x51 & n1008 ;
  assign n1010 = n332 & ~n339 ;
  assign n1011 = n1010 ^ n418 ^ 1'b0 ;
  assign n1012 = ( ~n597 & n746 ) | ( ~n597 & n1011 ) | ( n746 & n1011 ) ;
  assign n1013 = n1012 ^ n957 ^ n650 ;
  assign n1014 = n335 | n624 ;
  assign n1015 = n1014 ^ n938 ^ 1'b0 ;
  assign n1016 = ( ~n383 & n740 ) | ( ~n383 & n760 ) | ( n740 & n760 ) ;
  assign n1017 = ( n290 & ~n548 ) | ( n290 & n1016 ) | ( ~n548 & n1016 ) ;
  assign n1018 = ( ~x94 & n389 ) | ( ~x94 & n1017 ) | ( n389 & n1017 ) ;
  assign n1019 = ( n420 & n1015 ) | ( n420 & n1018 ) | ( n1015 & n1018 ) ;
  assign n1020 = n887 ^ n873 ^ n725 ;
  assign n1021 = ( ~n273 & n555 ) | ( ~n273 & n694 ) | ( n555 & n694 ) ;
  assign n1022 = n733 & n1021 ;
  assign n1023 = ~n822 & n1022 ;
  assign n1026 = ~n187 & n607 ;
  assign n1027 = ~x53 & n1026 ;
  assign n1024 = ( n453 & ~n505 ) | ( n453 & n540 ) | ( ~n505 & n540 ) ;
  assign n1025 = n1024 ^ n565 ^ n149 ;
  assign n1028 = n1027 ^ n1025 ^ n909 ;
  assign n1035 = x104 & ~n315 ;
  assign n1034 = x59 & ~n475 ;
  assign n1032 = n482 ^ n334 ^ 1'b0 ;
  assign n1030 = x123 & ~n380 ;
  assign n1031 = n567 & n1030 ;
  assign n1029 = ( ~n241 & n284 ) | ( ~n241 & n562 ) | ( n284 & n562 ) ;
  assign n1033 = n1032 ^ n1031 ^ n1029 ;
  assign n1036 = n1035 ^ n1034 ^ n1033 ;
  assign n1037 = n643 ^ n498 ^ x86 ;
  assign n1038 = ( ~n710 & n880 ) | ( ~n710 & n1037 ) | ( n880 & n1037 ) ;
  assign n1039 = ( x86 & ~n802 ) | ( x86 & n1038 ) | ( ~n802 & n1038 ) ;
  assign n1044 = n197 ^ n179 ^ x4 ;
  assign n1041 = n593 ^ x9 ^ 1'b0 ;
  assign n1042 = x22 & n1041 ;
  assign n1040 = n663 ^ n636 ^ 1'b0 ;
  assign n1043 = n1042 ^ n1040 ^ n658 ;
  assign n1045 = n1044 ^ n1043 ^ n940 ;
  assign n1046 = x92 & ~n697 ;
  assign n1047 = n871 ^ n580 ^ n289 ;
  assign n1048 = ( ~x113 & n1046 ) | ( ~x113 & n1047 ) | ( n1046 & n1047 ) ;
  assign n1049 = n258 ^ n149 ^ 1'b0 ;
  assign n1050 = n135 & n1049 ;
  assign n1051 = ( ~n374 & n1048 ) | ( ~n374 & n1050 ) | ( n1048 & n1050 ) ;
  assign n1052 = n173 ^ x70 ^ x63 ;
  assign n1053 = n1052 ^ n272 ^ 1'b0 ;
  assign n1054 = n643 | n1053 ;
  assign n1055 = n1054 ^ n370 ^ n231 ;
  assign n1056 = n531 ^ n445 ^ x89 ;
  assign n1057 = ( ~n319 & n941 ) | ( ~n319 & n991 ) | ( n941 & n991 ) ;
  assign n1058 = ( n713 & ~n789 ) | ( n713 & n1057 ) | ( ~n789 & n1057 ) ;
  assign n1059 = n409 ^ x21 ^ 1'b0 ;
  assign n1060 = n1059 ^ n537 ^ 1'b0 ;
  assign n1061 = n1060 ^ n586 ^ 1'b0 ;
  assign n1062 = n243 & ~n653 ;
  assign n1063 = n304 & ~n380 ;
  assign n1064 = n1063 ^ n359 ^ 1'b0 ;
  assign n1065 = ~n496 & n760 ;
  assign n1066 = ~n252 & n1065 ;
  assign n1067 = ( x50 & ~n502 ) | ( x50 & n1066 ) | ( ~n502 & n1066 ) ;
  assign n1068 = n628 & ~n1067 ;
  assign n1084 = n523 ^ n304 ^ n151 ;
  assign n1083 = n232 & n679 ;
  assign n1085 = n1084 ^ n1083 ^ 1'b0 ;
  assign n1069 = ( ~x77 & n305 ) | ( ~x77 & n306 ) | ( n305 & n306 ) ;
  assign n1071 = n640 & ~n1032 ;
  assign n1070 = n199 | n243 ;
  assign n1072 = n1071 ^ n1070 ^ 1'b0 ;
  assign n1073 = n1069 & ~n1072 ;
  assign n1074 = ~x51 & n1073 ;
  assign n1075 = n1074 ^ x84 ^ 1'b0 ;
  assign n1077 = n204 ^ x51 ^ 1'b0 ;
  assign n1078 = n129 & n1077 ;
  assign n1076 = n833 ^ n722 ^ n294 ;
  assign n1079 = n1078 ^ n1076 ^ n409 ;
  assign n1080 = ~n663 & n778 ;
  assign n1081 = n1080 ^ n844 ^ 1'b0 ;
  assign n1082 = ( ~n1075 & n1079 ) | ( ~n1075 & n1081 ) | ( n1079 & n1081 ) ;
  assign n1086 = n1085 ^ n1082 ^ n370 ;
  assign n1091 = n272 & n905 ;
  assign n1092 = n1091 ^ n429 ^ 1'b0 ;
  assign n1089 = ( x16 & ~x27 ) | ( x16 & x94 ) | ( ~x27 & x94 ) ;
  assign n1087 = x124 & ~n750 ;
  assign n1088 = n1087 ^ n891 ^ 1'b0 ;
  assign n1090 = n1089 ^ n1088 ^ n256 ;
  assign n1093 = n1092 ^ n1090 ^ n933 ;
  assign n1094 = n908 | n1093 ;
  assign n1095 = x123 | n1094 ;
  assign n1099 = n195 | n426 ;
  assign n1097 = n1084 ^ n600 ^ n326 ;
  assign n1098 = ~n186 & n1097 ;
  assign n1096 = ( ~n614 & n624 ) | ( ~n614 & n636 ) | ( n624 & n636 ) ;
  assign n1100 = n1099 ^ n1098 ^ n1096 ;
  assign n1102 = ~x112 & n451 ;
  assign n1101 = ~n398 & n572 ;
  assign n1103 = n1102 ^ n1101 ^ 1'b0 ;
  assign n1104 = x52 & n1103 ;
  assign n1105 = n1104 ^ n475 ^ 1'b0 ;
  assign n1106 = n1100 | n1105 ;
  assign n1107 = ( ~x21 & x86 ) | ( ~x21 & n721 ) | ( x86 & n721 ) ;
  assign n1108 = ( n270 & ~n702 ) | ( n270 & n1107 ) | ( ~n702 & n1107 ) ;
  assign n1109 = n1108 ^ n1027 ^ 1'b0 ;
  assign n1110 = x63 | n571 ;
  assign n1111 = ~n131 & n1110 ;
  assign n1112 = ~n853 & n1111 ;
  assign n1113 = n177 ^ n131 ^ 1'b0 ;
  assign n1114 = ( n600 & n1112 ) | ( n600 & n1113 ) | ( n1112 & n1113 ) ;
  assign n1115 = x104 & n726 ;
  assign n1116 = n1114 & n1115 ;
  assign n1117 = ( n237 & ~n393 ) | ( n237 & n1116 ) | ( ~n393 & n1116 ) ;
  assign n1118 = n1117 ^ n935 ^ n825 ;
  assign n1119 = n636 ^ n271 ^ n157 ;
  assign n1120 = n1119 ^ n740 ^ x58 ;
  assign n1121 = ( n414 & ~n494 ) | ( n414 & n739 ) | ( ~n494 & n739 ) ;
  assign n1122 = ( ~n1110 & n1120 ) | ( ~n1110 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1123 = n1122 ^ n845 ^ 1'b0 ;
  assign n1125 = n479 ^ x83 ^ 1'b0 ;
  assign n1126 = n1125 ^ n507 ^ x34 ;
  assign n1124 = n349 ^ n326 ^ x17 ;
  assign n1127 = n1126 ^ n1124 ^ 1'b0 ;
  assign n1135 = ( n163 & n598 ) | ( n163 & ~n880 ) | ( n598 & ~n880 ) ;
  assign n1136 = n1135 ^ n719 ^ x69 ;
  assign n1137 = n409 | n1136 ;
  assign n1138 = n569 | n1137 ;
  assign n1132 = n156 ^ x114 ^ 1'b0 ;
  assign n1133 = x97 & ~n1132 ;
  assign n1131 = n1000 ^ n690 ^ n426 ;
  assign n1128 = n145 & n562 ;
  assign n1129 = n1128 ^ n414 ^ 1'b0 ;
  assign n1130 = n1129 ^ n787 ^ x109 ;
  assign n1134 = n1133 ^ n1131 ^ n1130 ;
  assign n1139 = n1138 ^ n1134 ^ x49 ;
  assign n1140 = n206 ^ n187 ^ 1'b0 ;
  assign n1141 = ( ~n435 & n1075 ) | ( ~n435 & n1140 ) | ( n1075 & n1140 ) ;
  assign n1144 = n856 ^ n189 ^ 1'b0 ;
  assign n1145 = n458 & ~n1144 ;
  assign n1146 = n1145 ^ n805 ^ n493 ;
  assign n1142 = ( x4 & x83 ) | ( x4 & ~n270 ) | ( x83 & ~n270 ) ;
  assign n1143 = ( n586 & ~n685 ) | ( n586 & n1142 ) | ( ~n685 & n1142 ) ;
  assign n1147 = n1146 ^ n1143 ^ 1'b0 ;
  assign n1148 = n828 & n1147 ;
  assign n1152 = ( n466 & ~n637 ) | ( n466 & n1047 ) | ( ~n637 & n1047 ) ;
  assign n1149 = n816 ^ n572 ^ n184 ;
  assign n1150 = n1149 ^ n457 ^ x1 ;
  assign n1151 = ( ~n264 & n514 ) | ( ~n264 & n1150 ) | ( n514 & n1150 ) ;
  assign n1153 = n1152 ^ n1151 ^ n494 ;
  assign n1154 = n988 & n1084 ;
  assign n1155 = ~x61 & n1154 ;
  assign n1156 = n402 & ~n933 ;
  assign n1157 = ~n296 & n1156 ;
  assign n1158 = ( n773 & n1155 ) | ( n773 & ~n1157 ) | ( n1155 & ~n1157 ) ;
  assign n1159 = ( ~x67 & n521 ) | ( ~x67 & n721 ) | ( n521 & n721 ) ;
  assign n1160 = n1159 ^ n1100 ^ 1'b0 ;
  assign n1161 = x110 & n1160 ;
  assign n1162 = ( x102 & n1158 ) | ( x102 & n1161 ) | ( n1158 & n1161 ) ;
  assign n1178 = x66 & ~n370 ;
  assign n1179 = n1178 ^ n225 ^ 1'b0 ;
  assign n1180 = n1179 ^ n728 ^ n277 ;
  assign n1181 = n1180 ^ n767 ^ n731 ;
  assign n1175 = n261 & ~n954 ;
  assign n1176 = ~n333 & n1175 ;
  assign n1171 = n1067 ^ n461 ^ n362 ;
  assign n1172 = ( ~x106 & n410 ) | ( ~x106 & n1171 ) | ( n410 & n1171 ) ;
  assign n1173 = n1172 ^ n1145 ^ x89 ;
  assign n1169 = n148 & ~n282 ;
  assign n1170 = ~x13 & n1169 ;
  assign n1174 = n1173 ^ n1170 ^ n807 ;
  assign n1164 = n230 ^ x13 ^ 1'b0 ;
  assign n1165 = n783 ^ n507 ^ 1'b0 ;
  assign n1166 = n1165 ^ n614 ^ n489 ;
  assign n1167 = ( ~n495 & n1164 ) | ( ~n495 & n1166 ) | ( n1164 & n1166 ) ;
  assign n1163 = ~n313 & n547 ;
  assign n1168 = n1167 ^ n1163 ^ x101 ;
  assign n1177 = n1176 ^ n1174 ^ n1168 ;
  assign n1182 = n1181 ^ n1177 ^ 1'b0 ;
  assign n1183 = n782 | n1182 ;
  assign n1184 = ( n282 & n328 ) | ( n282 & n1135 ) | ( n328 & n1135 ) ;
  assign n1185 = n1184 ^ n589 ^ x24 ;
  assign n1186 = ( n833 & ~n1101 ) | ( n833 & n1185 ) | ( ~n1101 & n1185 ) ;
  assign n1187 = ( n345 & n878 ) | ( n345 & n1186 ) | ( n878 & n1186 ) ;
  assign n1216 = n1059 ^ n457 ^ n230 ;
  assign n1215 = n505 ^ n479 ^ n167 ;
  assign n1217 = n1216 ^ n1215 ^ n494 ;
  assign n1218 = n1217 ^ n1042 ^ n835 ;
  assign n1188 = n1016 ^ n447 ^ x88 ;
  assign n1189 = ( x18 & ~n367 ) | ( x18 & n1188 ) | ( ~n367 & n1188 ) ;
  assign n1190 = ( x15 & n149 ) | ( x15 & ~n685 ) | ( n149 & ~n685 ) ;
  assign n1191 = ( x56 & ~x118 ) | ( x56 & n175 ) | ( ~x118 & n175 ) ;
  assign n1192 = n1191 ^ x56 ^ 1'b0 ;
  assign n1193 = n1192 ^ n1042 ^ n400 ;
  assign n1194 = n1193 ^ n721 ^ n472 ;
  assign n1195 = ( n687 & ~n1190 ) | ( n687 & n1194 ) | ( ~n1190 & n1194 ) ;
  assign n1196 = n270 & ~n1164 ;
  assign n1197 = n1196 ^ x50 ^ 1'b0 ;
  assign n1198 = x65 & ~n1197 ;
  assign n1199 = n1198 ^ n997 ^ 1'b0 ;
  assign n1200 = n1199 ^ n243 ^ 1'b0 ;
  assign n1201 = ~n974 & n1200 ;
  assign n1202 = n742 ^ n472 ^ x16 ;
  assign n1203 = n1202 ^ n336 ^ 1'b0 ;
  assign n1204 = ( n284 & n329 ) | ( n284 & n1203 ) | ( n329 & n1203 ) ;
  assign n1205 = n1204 ^ n509 ^ n303 ;
  assign n1206 = n1205 ^ n630 ^ n201 ;
  assign n1209 = n148 & ~n1170 ;
  assign n1210 = n369 & n1209 ;
  assign n1207 = n657 ^ n251 ^ 1'b0 ;
  assign n1208 = n1207 ^ n566 ^ n513 ;
  assign n1211 = n1210 ^ n1208 ^ x68 ;
  assign n1212 = ( n1201 & n1206 ) | ( n1201 & ~n1211 ) | ( n1206 & ~n1211 ) ;
  assign n1213 = ( n1189 & n1195 ) | ( n1189 & n1212 ) | ( n1195 & n1212 ) ;
  assign n1214 = ~n133 & n1213 ;
  assign n1219 = n1218 ^ n1214 ^ 1'b0 ;
  assign n1220 = ( x95 & n493 ) | ( x95 & n622 ) | ( n493 & n622 ) ;
  assign n1221 = ~n418 & n1220 ;
  assign n1222 = n972 ^ n328 ^ 1'b0 ;
  assign n1223 = ( n146 & ~n378 ) | ( n146 & n1222 ) | ( ~n378 & n1222 ) ;
  assign n1227 = ( x113 & n417 ) | ( x113 & n947 ) | ( n417 & n947 ) ;
  assign n1228 = n1227 ^ n540 ^ n284 ;
  assign n1229 = ( n160 & ~n1075 ) | ( n160 & n1228 ) | ( ~n1075 & n1228 ) ;
  assign n1224 = n213 & ~n643 ;
  assign n1225 = n1224 ^ n333 ^ 1'b0 ;
  assign n1226 = ( x48 & ~n541 ) | ( x48 & n1225 ) | ( ~n541 & n1225 ) ;
  assign n1230 = n1229 ^ n1226 ^ 1'b0 ;
  assign n1231 = ( n186 & ~n1206 ) | ( n186 & n1230 ) | ( ~n1206 & n1230 ) ;
  assign n1233 = ( x91 & ~n226 ) | ( x91 & n282 ) | ( ~n226 & n282 ) ;
  assign n1232 = n538 & ~n923 ;
  assign n1234 = n1233 ^ n1232 ^ n346 ;
  assign n1243 = n224 | n675 ;
  assign n1244 = x44 | n1243 ;
  assign n1245 = n743 ^ x98 ^ 1'b0 ;
  assign n1246 = n1244 & ~n1245 ;
  assign n1240 = n581 ^ n449 ^ n156 ;
  assign n1241 = n1240 ^ n252 ^ 1'b0 ;
  assign n1239 = ( x8 & n320 ) | ( x8 & n558 ) | ( n320 & n558 ) ;
  assign n1242 = n1241 ^ n1239 ^ n362 ;
  assign n1235 = n548 & n1199 ;
  assign n1236 = x47 | n1235 ;
  assign n1237 = x10 & n1236 ;
  assign n1238 = n1237 ^ n666 ^ 1'b0 ;
  assign n1247 = n1246 ^ n1242 ^ n1238 ;
  assign n1253 = n176 ^ x99 ^ x24 ;
  assign n1249 = n211 | n487 ;
  assign n1250 = n353 & ~n1249 ;
  assign n1251 = ( x9 & n1203 ) | ( x9 & n1250 ) | ( n1203 & n1250 ) ;
  assign n1252 = n1096 & n1251 ;
  assign n1254 = n1253 ^ n1252 ^ n321 ;
  assign n1248 = n763 ^ n709 ^ x11 ;
  assign n1255 = n1254 ^ n1248 ^ n718 ;
  assign n1256 = n201 & ~n659 ;
  assign n1257 = ( n791 & ~n839 ) | ( n791 & n1256 ) | ( ~n839 & n1256 ) ;
  assign n1258 = ( n216 & n264 ) | ( n216 & n1047 ) | ( n264 & n1047 ) ;
  assign n1259 = n1167 ^ n1033 ^ 1'b0 ;
  assign n1260 = n335 | n914 ;
  assign n1261 = n581 ^ n475 ^ x66 ;
  assign n1262 = n1261 ^ n924 ^ n371 ;
  assign n1263 = ( n1143 & n1260 ) | ( n1143 & n1262 ) | ( n1260 & n1262 ) ;
  assign n1264 = ( n252 & ~n490 ) | ( n252 & n684 ) | ( ~n490 & n684 ) ;
  assign n1265 = ( n393 & ~n622 ) | ( n393 & n850 ) | ( ~n622 & n850 ) ;
  assign n1266 = ( ~n1028 & n1254 ) | ( ~n1028 & n1265 ) | ( n1254 & n1265 ) ;
  assign n1272 = n356 ^ x24 ^ 1'b0 ;
  assign n1273 = n997 & ~n1272 ;
  assign n1267 = n154 | n770 ;
  assign n1268 = ( x122 & n144 ) | ( x122 & ~n290 ) | ( n144 & ~n290 ) ;
  assign n1269 = n1268 ^ n825 ^ n451 ;
  assign n1270 = n1269 ^ n742 ^ 1'b0 ;
  assign n1271 = n1267 & ~n1270 ;
  assign n1274 = n1273 ^ n1271 ^ n703 ;
  assign n1275 = n326 & ~n907 ;
  assign n1276 = ~n719 & n1275 ;
  assign n1277 = n1276 ^ n529 ^ 1'b0 ;
  assign n1278 = ( n173 & n627 ) | ( n173 & n835 ) | ( n627 & n835 ) ;
  assign n1279 = n400 ^ n277 ^ 1'b0 ;
  assign n1280 = x48 & n1279 ;
  assign n1281 = ~n738 & n1280 ;
  assign n1282 = ~n420 & n1281 ;
  assign n1283 = n509 ^ n506 ^ x36 ;
  assign n1284 = ( n466 & n802 ) | ( n466 & ~n890 ) | ( n802 & ~n890 ) ;
  assign n1285 = ( ~x46 & n354 ) | ( ~x46 & n761 ) | ( n354 & n761 ) ;
  assign n1286 = n1285 ^ n436 ^ x79 ;
  assign n1287 = n1286 ^ n344 ^ x18 ;
  assign n1288 = n1287 ^ n716 ^ n340 ;
  assign n1289 = n1234 ^ n957 ^ n723 ;
  assign n1300 = ~x126 & n1207 ;
  assign n1295 = n253 ^ n167 ^ 1'b0 ;
  assign n1296 = n1016 & ~n1179 ;
  assign n1297 = n1296 ^ n989 ^ 1'b0 ;
  assign n1298 = n1297 ^ n649 ^ n383 ;
  assign n1299 = ( ~x86 & n1295 ) | ( ~x86 & n1298 ) | ( n1295 & n1298 ) ;
  assign n1290 = n823 ^ n341 ^ 1'b0 ;
  assign n1291 = n1290 ^ n1028 ^ n847 ;
  assign n1292 = n333 & n1291 ;
  assign n1293 = ~n811 & n1292 ;
  assign n1294 = n1293 ^ n690 ^ n397 ;
  assign n1301 = n1300 ^ n1299 ^ n1294 ;
  assign n1302 = n490 ^ n260 ^ n240 ;
  assign n1303 = n1302 ^ n337 ^ n256 ;
  assign n1304 = ( x97 & n168 ) | ( x97 & ~n172 ) | ( n168 & ~n172 ) ;
  assign n1305 = n1304 ^ n667 ^ n291 ;
  assign n1306 = ( x48 & n1303 ) | ( x48 & n1305 ) | ( n1303 & n1305 ) ;
  assign n1307 = x33 | n665 ;
  assign n1308 = n1307 ^ n1099 ^ n598 ;
  assign n1309 = ( n189 & n510 ) | ( n189 & n538 ) | ( n510 & n538 ) ;
  assign n1310 = x36 & n399 ;
  assign n1311 = n1310 ^ n456 ^ 1'b0 ;
  assign n1312 = ( x78 & n1309 ) | ( x78 & n1311 ) | ( n1309 & n1311 ) ;
  assign n1313 = ( n1152 & n1269 ) | ( n1152 & n1312 ) | ( n1269 & n1312 ) ;
  assign n1314 = ( ~n357 & n364 ) | ( ~n357 & n898 ) | ( n364 & n898 ) ;
  assign n1315 = n243 & n1314 ;
  assign n1316 = x70 & n217 ;
  assign n1317 = ~x32 & n1316 ;
  assign n1318 = n988 ^ n243 ^ 1'b0 ;
  assign n1319 = x125 & ~n136 ;
  assign n1320 = n1318 & n1319 ;
  assign n1321 = ( n1059 & n1317 ) | ( n1059 & ~n1320 ) | ( n1317 & ~n1320 ) ;
  assign n1322 = n1321 ^ n1240 ^ n209 ;
  assign n1325 = n658 ^ n457 ^ n216 ;
  assign n1323 = n702 ^ n204 ^ 1'b0 ;
  assign n1324 = n1037 & ~n1323 ;
  assign n1326 = n1325 ^ n1324 ^ 1'b0 ;
  assign n1327 = n1326 ^ n622 ^ 1'b0 ;
  assign n1328 = n1107 & n1327 ;
  assign n1329 = n1328 ^ n1216 ^ 1'b0 ;
  assign n1330 = n268 ^ n218 ^ 1'b0 ;
  assign n1331 = n1199 ^ n863 ^ n558 ;
  assign n1332 = ( n762 & n1330 ) | ( n762 & ~n1331 ) | ( n1330 & ~n1331 ) ;
  assign n1333 = ( n659 & ~n1329 ) | ( n659 & n1332 ) | ( ~n1329 & n1332 ) ;
  assign n1334 = ( x67 & n506 ) | ( x67 & n941 ) | ( n506 & n941 ) ;
  assign n1340 = n542 ^ n293 ^ 1'b0 ;
  assign n1337 = n848 ^ n357 ^ n337 ;
  assign n1338 = n383 ^ n222 ^ 1'b0 ;
  assign n1339 = n1337 | n1338 ;
  assign n1335 = n510 ^ n242 ^ x38 ;
  assign n1336 = n1335 ^ n979 ^ n604 ;
  assign n1341 = n1340 ^ n1339 ^ n1336 ;
  assign n1342 = n619 ^ n204 ^ 1'b0 ;
  assign n1343 = ( x91 & ~n331 ) | ( x91 & n799 ) | ( ~n331 & n799 ) ;
  assign n1344 = ~n1342 & n1343 ;
  assign n1345 = n1344 ^ n1012 ^ 1'b0 ;
  assign n1346 = n1345 ^ n995 ^ n724 ;
  assign n1347 = n1346 ^ n633 ^ n200 ;
  assign n1348 = ( n395 & ~n826 ) | ( n395 & n1110 ) | ( ~n826 & n1110 ) ;
  assign n1349 = n1348 ^ n604 ^ n528 ;
  assign n1350 = ~n896 & n1349 ;
  assign n1351 = n1350 ^ x89 ^ 1'b0 ;
  assign n1352 = n1347 | n1351 ;
  assign n1353 = n805 ^ n588 ^ 1'b0 ;
  assign n1354 = n1232 ^ n1012 ^ n937 ;
  assign n1356 = n1108 ^ n582 ^ n352 ;
  assign n1355 = n1074 ^ n567 ^ x31 ;
  assign n1357 = n1356 ^ n1355 ^ 1'b0 ;
  assign n1358 = n255 ^ n227 ^ 1'b0 ;
  assign n1359 = n143 | n1358 ;
  assign n1360 = n135 ^ x36 ^ x9 ;
  assign n1361 = n1360 ^ n1210 ^ n1027 ;
  assign n1362 = n1361 ^ n600 ^ n352 ;
  assign n1363 = n1362 ^ n880 ^ n253 ;
  assign n1364 = n132 & ~n1363 ;
  assign n1365 = n1364 ^ x119 ^ 1'b0 ;
  assign n1366 = ( n229 & n498 ) | ( n229 & n1158 ) | ( n498 & n1158 ) ;
  assign n1367 = ( n1225 & ~n1365 ) | ( n1225 & n1366 ) | ( ~n1365 & n1366 ) ;
  assign n1368 = ~n1359 & n1367 ;
  assign n1369 = ~n1148 & n1368 ;
  assign n1370 = n1261 ^ n464 ^ n303 ;
  assign n1371 = n1370 ^ x99 ^ 1'b0 ;
  assign n1372 = ~n369 & n1069 ;
  assign n1373 = n1251 ^ n639 ^ n526 ;
  assign n1374 = ( ~n196 & n211 ) | ( ~n196 & n241 ) | ( n211 & n241 ) ;
  assign n1375 = n1374 ^ n671 ^ x105 ;
  assign n1376 = x79 ^ x36 ^ x33 ;
  assign n1377 = n1376 ^ n841 ^ x76 ;
  assign n1378 = ( n350 & ~n1375 ) | ( n350 & n1377 ) | ( ~n1375 & n1377 ) ;
  assign n1379 = n517 & n1378 ;
  assign n1380 = ( ~n1372 & n1373 ) | ( ~n1372 & n1379 ) | ( n1373 & n1379 ) ;
  assign n1381 = ( n270 & ~n552 ) | ( n270 & n557 ) | ( ~n552 & n557 ) ;
  assign n1382 = ( n535 & n751 ) | ( n535 & n1381 ) | ( n751 & n1381 ) ;
  assign n1383 = n328 & ~n608 ;
  assign n1384 = n1360 & n1383 ;
  assign n1385 = n1060 & ~n1384 ;
  assign n1386 = ~n1382 & n1385 ;
  assign n1395 = n722 ^ n562 ^ x85 ;
  assign n1392 = n647 ^ n218 ^ 1'b0 ;
  assign n1393 = ~n369 & n1392 ;
  assign n1394 = ( n336 & ~n385 ) | ( n336 & n1393 ) | ( ~n385 & n1393 ) ;
  assign n1389 = n1384 ^ n343 ^ n240 ;
  assign n1390 = n1389 ^ n1170 ^ n604 ;
  assign n1387 = n217 & ~n933 ;
  assign n1388 = n1387 ^ n204 ^ 1'b0 ;
  assign n1391 = n1390 ^ n1388 ^ n1376 ;
  assign n1396 = n1395 ^ n1394 ^ n1391 ;
  assign n1397 = n1396 ^ n811 ^ n213 ;
  assign n1398 = ~n445 & n1397 ;
  assign n1399 = n1398 ^ n889 ^ 1'b0 ;
  assign n1400 = n619 ^ n268 ^ x85 ;
  assign n1401 = n1400 ^ x18 ^ 1'b0 ;
  assign n1402 = n902 | n1401 ;
  assign n1403 = n1374 ^ n1131 ^ n317 ;
  assign n1404 = n1403 ^ n1114 ^ n934 ;
  assign n1405 = n581 ^ x83 ^ x64 ;
  assign n1406 = n1405 ^ n1232 ^ 1'b0 ;
  assign n1407 = n1404 & ~n1406 ;
  assign n1408 = ( ~n289 & n664 ) | ( ~n289 & n716 ) | ( n664 & n716 ) ;
  assign n1410 = n1059 ^ n912 ^ 1'b0 ;
  assign n1409 = ( x64 & n931 ) | ( x64 & n1301 ) | ( n931 & n1301 ) ;
  assign n1411 = n1410 ^ n1409 ^ n1000 ;
  assign n1412 = x126 & ~n136 ;
  assign n1413 = ~n1411 & n1412 ;
  assign n1414 = ( n342 & n642 ) | ( n342 & ~n990 ) | ( n642 & ~n990 ) ;
  assign n1415 = x13 & x62 ;
  assign n1416 = ~x79 & n1415 ;
  assign n1417 = n164 | n1416 ;
  assign n1418 = ( n542 & n822 ) | ( n542 & ~n1417 ) | ( n822 & ~n1417 ) ;
  assign n1419 = n300 & n914 ;
  assign n1420 = n461 & n1419 ;
  assign n1425 = n1136 ^ n305 ^ x55 ;
  assign n1421 = ( n478 & n503 ) | ( n478 & ~n600 ) | ( n503 & ~n600 ) ;
  assign n1422 = n1421 ^ n1179 ^ n312 ;
  assign n1423 = n394 | n643 ;
  assign n1424 = n1422 | n1423 ;
  assign n1426 = n1425 ^ n1424 ^ n857 ;
  assign n1427 = n629 & n1193 ;
  assign n1428 = n1427 ^ n479 ^ 1'b0 ;
  assign n1429 = n398 & ~n1428 ;
  assign n1430 = ~n1426 & n1429 ;
  assign n1431 = n1430 ^ n967 ^ x93 ;
  assign n1432 = n979 & ~n1360 ;
  assign n1433 = n537 & n1432 ;
  assign n1434 = ( x48 & ~x86 ) | ( x48 & n1069 ) | ( ~x86 & n1069 ) ;
  assign n1435 = n1042 & ~n1376 ;
  assign n1436 = ~n1190 & n1435 ;
  assign n1437 = n1436 ^ n538 ^ n217 ;
  assign n1438 = n1437 ^ n592 ^ 1'b0 ;
  assign n1439 = n1355 | n1438 ;
  assign n1440 = n1439 ^ n291 ^ 1'b0 ;
  assign n1441 = n1360 ^ n540 ^ n503 ;
  assign n1442 = n1441 ^ n340 ^ n204 ;
  assign n1443 = ( n557 & n862 ) | ( n557 & ~n1442 ) | ( n862 & ~n1442 ) ;
  assign n1444 = ( n466 & n547 ) | ( n466 & ~n967 ) | ( n547 & ~n967 ) ;
  assign n1445 = n1046 ^ n200 ^ n173 ;
  assign n1446 = n1445 ^ n1210 ^ 1'b0 ;
  assign n1447 = n1273 & n1446 ;
  assign n1448 = n1447 ^ n336 ^ 1'b0 ;
  assign n1449 = n1444 & ~n1448 ;
  assign n1450 = ( ~n1440 & n1443 ) | ( ~n1440 & n1449 ) | ( n1443 & n1449 ) ;
  assign n1451 = n631 & n1152 ;
  assign n1452 = n941 | n1451 ;
  assign n1453 = n271 | n1452 ;
  assign n1460 = n1417 ^ x27 ^ 1'b0 ;
  assign n1461 = n1460 ^ n950 ^ 1'b0 ;
  assign n1462 = n1461 ^ n979 ^ x110 ;
  assign n1456 = n214 & ~n1002 ;
  assign n1457 = ~n1025 & n1456 ;
  assign n1454 = n429 ^ x33 ^ 1'b0 ;
  assign n1455 = n1454 ^ n862 ^ n177 ;
  assign n1458 = n1457 ^ n1455 ^ 1'b0 ;
  assign n1459 = ~n1302 & n1458 ;
  assign n1463 = n1462 ^ n1459 ^ n1428 ;
  assign n1464 = n1121 ^ n551 ^ 1'b0 ;
  assign n1465 = n592 & ~n1464 ;
  assign n1466 = ( x8 & ~n326 ) | ( x8 & n1465 ) | ( ~n326 & n1465 ) ;
  assign n1467 = n1376 ^ n608 ^ x18 ;
  assign n1468 = n510 ^ n475 ^ x106 ;
  assign n1469 = ~n571 & n1468 ;
  assign n1470 = n669 & n1469 ;
  assign n1471 = n1470 ^ n168 ^ 1'b0 ;
  assign n1472 = n994 | n1471 ;
  assign n1473 = x71 & ~n1157 ;
  assign n1474 = n505 & n1473 ;
  assign n1475 = ( ~n847 & n1472 ) | ( ~n847 & n1474 ) | ( n1472 & n1474 ) ;
  assign n1476 = n689 ^ n664 ^ x48 ;
  assign n1477 = ~n352 & n1166 ;
  assign n1478 = n1477 ^ n679 ^ 1'b0 ;
  assign n1479 = n1478 ^ n858 ^ n525 ;
  assign n1480 = ( n133 & n1253 ) | ( n133 & n1273 ) | ( n1253 & n1273 ) ;
  assign n1481 = n1480 ^ n1299 ^ n1195 ;
  assign n1482 = ~n1291 & n1481 ;
  assign n1483 = ( n233 & n1479 ) | ( n233 & ~n1482 ) | ( n1479 & ~n1482 ) ;
  assign n1484 = n1483 ^ n211 ^ 1'b0 ;
  assign n1487 = n1416 ^ n609 ^ n253 ;
  assign n1486 = n1454 ^ n1253 ^ n508 ;
  assign n1488 = n1487 ^ n1486 ^ n871 ;
  assign n1485 = ( n209 & n367 ) | ( n209 & n865 ) | ( n367 & n865 ) ;
  assign n1489 = n1488 ^ n1485 ^ 1'b0 ;
  assign n1490 = x53 | n236 ;
  assign n1491 = n1490 ^ n1447 ^ 1'b0 ;
  assign n1492 = x125 & n1491 ;
  assign n1493 = n713 ^ n661 ^ x88 ;
  assign n1494 = ( x33 & x123 ) | ( x33 & ~n1493 ) | ( x123 & ~n1493 ) ;
  assign n1495 = ~n796 & n1494 ;
  assign n1496 = n383 ^ n137 ^ x102 ;
  assign n1497 = ~n324 & n1496 ;
  assign n1498 = n346 & n1497 ;
  assign n1499 = n1445 | n1498 ;
  assign n1500 = n156 & ~n1499 ;
  assign n1501 = n1381 ^ n728 ^ n553 ;
  assign n1502 = n418 | n1501 ;
  assign n1503 = n1500 & ~n1502 ;
  assign n1504 = n324 & ~n1503 ;
  assign n1506 = ( n168 & n330 ) | ( n168 & ~n436 ) | ( n330 & ~n436 ) ;
  assign n1505 = x13 & n921 ;
  assign n1507 = n1506 ^ n1505 ^ 1'b0 ;
  assign n1515 = n382 ^ n261 ^ n184 ;
  assign n1508 = n914 ^ n565 ^ n499 ;
  assign n1509 = n423 ^ x43 ^ 1'b0 ;
  assign n1510 = n1509 ^ n715 ^ x46 ;
  assign n1511 = ( n280 & n1203 ) | ( n280 & n1510 ) | ( n1203 & n1510 ) ;
  assign n1512 = n1511 ^ n510 ^ n348 ;
  assign n1513 = n1512 ^ n451 ^ n202 ;
  assign n1514 = ( n479 & ~n1508 ) | ( n479 & n1513 ) | ( ~n1508 & n1513 ) ;
  assign n1516 = n1515 ^ n1514 ^ x62 ;
  assign n1517 = n267 ^ n189 ^ x113 ;
  assign n1518 = n589 | n1517 ;
  assign n1519 = ( x1 & n220 ) | ( x1 & ~n1518 ) | ( n220 & ~n1518 ) ;
  assign n1520 = n1519 ^ x78 ^ 1'b0 ;
  assign n1521 = x60 & n1520 ;
  assign n1522 = n1256 ^ n561 ^ 1'b0 ;
  assign n1523 = ( ~x118 & n282 ) | ( ~x118 & n1522 ) | ( n282 & n1522 ) ;
  assign n1524 = ( ~n667 & n1248 ) | ( ~n667 & n1523 ) | ( n1248 & n1523 ) ;
  assign n1525 = n762 ^ n533 ^ 1'b0 ;
  assign n1526 = x123 & n592 ;
  assign n1527 = n230 & n1526 ;
  assign n1528 = n1527 ^ n937 ^ n793 ;
  assign n1529 = ( ~x100 & n135 ) | ( ~x100 & n1125 ) | ( n135 & n1125 ) ;
  assign n1530 = n1529 ^ n1525 ^ 1'b0 ;
  assign n1531 = n808 & ~n1530 ;
  assign n1532 = ( n1525 & n1528 ) | ( n1525 & n1531 ) | ( n1528 & n1531 ) ;
  assign n1533 = n1078 ^ n770 ^ n348 ;
  assign n1534 = n1533 ^ n1322 ^ n716 ;
  assign n1535 = ( ~n238 & n1341 ) | ( ~n238 & n1519 ) | ( n1341 & n1519 ) ;
  assign n1537 = n1031 ^ n705 ^ n442 ;
  assign n1536 = x97 & ~n675 ;
  assign n1538 = n1537 ^ n1536 ^ 1'b0 ;
  assign n1539 = n1129 & ~n1537 ;
  assign n1540 = n1539 ^ n1097 ^ 1'b0 ;
  assign n1542 = n511 ^ n337 ^ n133 ;
  assign n1543 = n1542 ^ n662 ^ x39 ;
  assign n1541 = ( x41 & ~n604 ) | ( x41 & n974 ) | ( ~n604 & n974 ) ;
  assign n1544 = n1543 ^ n1541 ^ n1298 ;
  assign n1545 = ( n355 & ~n1540 ) | ( n355 & n1544 ) | ( ~n1540 & n1544 ) ;
  assign n1547 = n440 ^ n428 ^ x17 ;
  assign n1548 = n322 & n1304 ;
  assign n1549 = n1548 ^ n883 ^ 1'b0 ;
  assign n1550 = ( n785 & ~n1547 ) | ( n785 & n1549 ) | ( ~n1547 & n1549 ) ;
  assign n1551 = n1550 ^ n808 ^ n578 ;
  assign n1546 = n863 ^ n131 ^ 1'b0 ;
  assign n1552 = n1551 ^ n1546 ^ n317 ;
  assign n1565 = ( n420 & n496 ) | ( n420 & n933 ) | ( n496 & n933 ) ;
  assign n1566 = ( n382 & n413 ) | ( n382 & n1565 ) | ( n413 & n1565 ) ;
  assign n1567 = ( n1280 & ~n1286 ) | ( n1280 & n1323 ) | ( ~n1286 & n1323 ) ;
  assign n1568 = n1567 ^ n655 ^ n375 ;
  assign n1569 = ( n294 & n1566 ) | ( n294 & ~n1568 ) | ( n1566 & ~n1568 ) ;
  assign n1553 = n685 | n791 ;
  assign n1554 = ~n706 & n1553 ;
  assign n1561 = n871 ^ n430 ^ 1'b0 ;
  assign n1556 = n919 ^ n204 ^ 1'b0 ;
  assign n1557 = n1556 ^ n1323 ^ n472 ;
  assign n1558 = n1557 ^ x31 ^ 1'b0 ;
  assign n1559 = n629 & ~n1558 ;
  assign n1560 = ( x125 & n755 ) | ( x125 & ~n1559 ) | ( n755 & ~n1559 ) ;
  assign n1555 = ( ~n490 & n663 ) | ( ~n490 & n839 ) | ( n663 & n839 ) ;
  assign n1562 = n1561 ^ n1560 ^ n1555 ;
  assign n1563 = n1562 ^ n945 ^ x113 ;
  assign n1564 = ~n1554 & n1563 ;
  assign n1570 = n1569 ^ n1564 ^ 1'b0 ;
  assign n1571 = ( ~n148 & n1552 ) | ( ~n148 & n1570 ) | ( n1552 & n1570 ) ;
  assign n1572 = ( ~n505 & n602 ) | ( ~n505 & n1513 ) | ( n602 & n1513 ) ;
  assign n1573 = ( x88 & n555 ) | ( x88 & ~n1269 ) | ( n555 & ~n1269 ) ;
  assign n1575 = x121 ^ x9 ^ x2 ;
  assign n1574 = n975 & ~n1550 ;
  assign n1576 = n1575 ^ n1574 ^ n1157 ;
  assign n1577 = ~n1573 & n1576 ;
  assign n1578 = ~n1572 & n1577 ;
  assign n1579 = n859 ^ n315 ^ 1'b0 ;
  assign n1580 = n1076 ^ n710 ^ n334 ;
  assign n1581 = ( n298 & n415 ) | ( n298 & n1580 ) | ( n415 & n1580 ) ;
  assign n1582 = ( ~n326 & n421 ) | ( ~n326 & n1581 ) | ( n421 & n1581 ) ;
  assign n1583 = ( ~n1386 & n1579 ) | ( ~n1386 & n1582 ) | ( n1579 & n1582 ) ;
  assign n1586 = ~n253 & n1494 ;
  assign n1587 = n1421 & n1586 ;
  assign n1588 = n1587 ^ n440 ^ x110 ;
  assign n1584 = ( n995 & ~n1046 ) | ( n995 & n1190 ) | ( ~n1046 & n1190 ) ;
  assign n1585 = n1325 & ~n1584 ;
  assign n1589 = n1588 ^ n1585 ^ 1'b0 ;
  assign n1594 = ( ~x0 & x110 ) | ( ~x0 & n217 ) | ( x110 & n217 ) ;
  assign n1590 = n271 & n329 ;
  assign n1591 = ~n1297 & n1590 ;
  assign n1592 = n1120 ^ n209 ^ x61 ;
  assign n1593 = ~n1591 & n1592 ;
  assign n1595 = n1594 ^ n1593 ^ 1'b0 ;
  assign n1596 = n1437 ^ n434 ^ 1'b0 ;
  assign n1597 = n453 & n1596 ;
  assign n1598 = n233 & n1597 ;
  assign n1599 = ~x62 & n1598 ;
  assign n1600 = n1599 ^ n1567 ^ x41 ;
  assign n1601 = n1325 ^ n1215 ^ n441 ;
  assign n1602 = ~n1331 & n1601 ;
  assign n1603 = n1602 ^ n1573 ^ 1'b0 ;
  assign n1604 = n582 & ~n1603 ;
  assign n1605 = n1600 & n1604 ;
  assign n1608 = n436 ^ n417 ^ 1'b0 ;
  assign n1606 = ( ~x64 & n178 ) | ( ~x64 & n493 ) | ( n178 & n493 ) ;
  assign n1607 = ( n199 & n229 ) | ( n199 & ~n1606 ) | ( n229 & ~n1606 ) ;
  assign n1609 = n1608 ^ n1607 ^ x3 ;
  assign n1610 = n1099 & n1609 ;
  assign n1617 = ( x22 & n199 ) | ( x22 & ~n367 ) | ( n199 & ~n367 ) ;
  assign n1611 = ( ~n691 & n701 ) | ( ~n691 & n1205 ) | ( n701 & n1205 ) ;
  assign n1612 = n456 ^ n196 ^ n144 ;
  assign n1613 = ( n230 & n1496 ) | ( n230 & ~n1612 ) | ( n1496 & ~n1612 ) ;
  assign n1614 = n1613 ^ n1047 ^ n746 ;
  assign n1615 = n1002 | n1614 ;
  assign n1616 = n1611 | n1615 ;
  assign n1618 = n1617 ^ n1616 ^ 1'b0 ;
  assign n1619 = ( ~n167 & n520 ) | ( ~n167 & n1618 ) | ( n520 & n1618 ) ;
  assign n1620 = ~n245 & n345 ;
  assign n1621 = n679 & n1620 ;
  assign n1622 = n969 ^ n529 ^ 1'b0 ;
  assign n1623 = x40 & ~n1622 ;
  assign n1624 = n1349 ^ n591 ^ n553 ;
  assign n1625 = ( ~n140 & n1623 ) | ( ~n140 & n1624 ) | ( n1623 & n1624 ) ;
  assign n1626 = ( x9 & n268 ) | ( x9 & ~n383 ) | ( n268 & ~n383 ) ;
  assign n1627 = ( ~n733 & n902 ) | ( ~n733 & n1626 ) | ( n902 & n1626 ) ;
  assign n1628 = n1625 & ~n1627 ;
  assign n1629 = ( n603 & n721 ) | ( n603 & ~n1285 ) | ( n721 & ~n1285 ) ;
  assign n1630 = ( ~x51 & n699 ) | ( ~x51 & n1629 ) | ( n699 & n1629 ) ;
  assign n1633 = n572 ^ n265 ^ x112 ;
  assign n1631 = x62 | n587 ;
  assign n1632 = n1631 ^ x126 ^ 1'b0 ;
  assign n1634 = n1633 ^ n1632 ^ n146 ;
  assign n1635 = ( n1007 & ~n1630 ) | ( n1007 & n1634 ) | ( ~n1630 & n1634 ) ;
  assign n1636 = n933 ^ n516 ^ 1'b0 ;
  assign n1637 = x50 & n1636 ;
  assign n1638 = n1635 & ~n1637 ;
  assign n1639 = n1470 ^ n604 ^ x46 ;
  assign n1643 = n1228 ^ n1024 ^ x14 ;
  assign n1640 = n870 ^ x72 ^ 1'b0 ;
  assign n1641 = x113 & n1640 ;
  assign n1642 = ~n802 & n1641 ;
  assign n1644 = n1643 ^ n1642 ^ n616 ;
  assign n1645 = ( ~x49 & n1639 ) | ( ~x49 & n1644 ) | ( n1639 & n1644 ) ;
  assign n1646 = n1204 ^ n784 ^ n611 ;
  assign n1647 = n1468 ^ n541 ^ x124 ;
  assign n1648 = ( n1345 & ~n1609 ) | ( n1345 & n1647 ) | ( ~n1609 & n1647 ) ;
  assign n1649 = n201 & n914 ;
  assign n1650 = n1649 ^ n352 ^ 1'b0 ;
  assign n1651 = ( x65 & ~n1494 ) | ( x65 & n1650 ) | ( ~n1494 & n1650 ) ;
  assign n1652 = ( ~x70 & n1362 ) | ( ~x70 & n1651 ) | ( n1362 & n1651 ) ;
  assign n1653 = n1652 ^ n1353 ^ n383 ;
  assign n1654 = x46 & ~n655 ;
  assign n1655 = n900 & n1654 ;
  assign n1656 = n977 | n1655 ;
  assign n1657 = n1656 ^ n544 ^ 1'b0 ;
  assign n1658 = n343 & ~n757 ;
  assign n1659 = ~n1657 & n1658 ;
  assign n1660 = ( n237 & n828 ) | ( n237 & ~n918 ) | ( n828 & ~n918 ) ;
  assign n1661 = ( n204 & ~n1606 ) | ( n204 & n1660 ) | ( ~n1606 & n1660 ) ;
  assign n1662 = ( n1213 & ~n1371 ) | ( n1213 & n1661 ) | ( ~n1371 & n1661 ) ;
  assign n1663 = n889 ^ x69 ^ x24 ;
  assign n1664 = n1663 ^ n787 ^ n693 ;
  assign n1665 = n1664 ^ n418 ^ n218 ;
  assign n1666 = n1665 ^ n997 ^ n755 ;
  assign n1667 = n1257 ^ n253 ^ 1'b0 ;
  assign n1668 = ( x3 & x54 ) | ( x3 & ~n1107 ) | ( x54 & ~n1107 ) ;
  assign n1669 = ( n135 & n1646 ) | ( n135 & ~n1668 ) | ( n1646 & ~n1668 ) ;
  assign n1670 = x14 & ~x56 ;
  assign n1671 = ( n334 & n918 ) | ( n334 & ~n1660 ) | ( n918 & ~n1660 ) ;
  assign n1672 = ~n1363 & n1671 ;
  assign n1673 = ( n622 & n633 ) | ( n622 & n1330 ) | ( n633 & n1330 ) ;
  assign n1674 = n214 & ~n1613 ;
  assign n1675 = n400 & n1674 ;
  assign n1676 = ( n935 & n1673 ) | ( n935 & ~n1675 ) | ( n1673 & ~n1675 ) ;
  assign n1677 = ~n780 & n1676 ;
  assign n1678 = n1677 ^ n365 ^ 1'b0 ;
  assign n1679 = ( ~x45 & n1373 ) | ( ~x45 & n1678 ) | ( n1373 & n1678 ) ;
  assign n1680 = ( x40 & n449 ) | ( x40 & n843 ) | ( n449 & n843 ) ;
  assign n1686 = n325 ^ x31 ^ 1'b0 ;
  assign n1684 = n1633 ^ n1079 ^ n1058 ;
  assign n1682 = n468 ^ n370 ^ n224 ;
  assign n1683 = ~n315 & n1682 ;
  assign n1685 = n1684 ^ n1683 ^ 1'b0 ;
  assign n1681 = n424 ^ n252 ^ x35 ;
  assign n1687 = n1686 ^ n1685 ^ n1681 ;
  assign n1688 = ( ~n771 & n1680 ) | ( ~n771 & n1687 ) | ( n1680 & n1687 ) ;
  assign n1693 = n706 ^ x98 ^ 1'b0 ;
  assign n1694 = n983 | n1693 ;
  assign n1689 = x101 & ~n153 ;
  assign n1690 = ~n580 & n1689 ;
  assign n1691 = n1005 | n1290 ;
  assign n1692 = n1690 & ~n1691 ;
  assign n1695 = n1694 ^ n1692 ^ n1459 ;
  assign n1698 = ( x28 & n439 ) | ( x28 & ~n811 ) | ( n439 & ~n811 ) ;
  assign n1701 = ( ~n165 & n689 ) | ( ~n165 & n1698 ) | ( n689 & n1698 ) ;
  assign n1699 = ( ~n183 & n686 ) | ( ~n183 & n1698 ) | ( n686 & n1698 ) ;
  assign n1702 = n1701 ^ n1699 ^ x123 ;
  assign n1703 = n1702 ^ n205 ^ n146 ;
  assign n1704 = n1703 ^ n1559 ^ x116 ;
  assign n1705 = x100 & n1071 ;
  assign n1706 = n508 | n1705 ;
  assign n1707 = n1706 ^ n494 ^ 1'b0 ;
  assign n1708 = ( n1498 & n1704 ) | ( n1498 & n1707 ) | ( n1704 & n1707 ) ;
  assign n1696 = n513 ^ n411 ^ x98 ;
  assign n1697 = n1696 ^ n1417 ^ n490 ;
  assign n1700 = n1699 ^ n1697 ^ n1123 ;
  assign n1709 = n1708 ^ n1700 ^ n1146 ;
  assign n1710 = n924 ^ n787 ^ n643 ;
  assign n1713 = n991 ^ x45 ^ x8 ;
  assign n1714 = ( n589 & ~n1248 ) | ( n589 & n1713 ) | ( ~n1248 & n1713 ) ;
  assign n1711 = n585 & n685 ;
  assign n1712 = n248 & n1711 ;
  assign n1715 = n1714 ^ n1712 ^ n200 ;
  assign n1716 = ( n1139 & ~n1710 ) | ( n1139 & n1715 ) | ( ~n1710 & n1715 ) ;
  assign n1717 = n342 | n1092 ;
  assign n1718 = n366 & ~n1717 ;
  assign n1719 = n1168 ^ n408 ^ 1'b0 ;
  assign n1720 = ~n485 & n1202 ;
  assign n1721 = ( x86 & n457 ) | ( x86 & n1720 ) | ( n457 & n1720 ) ;
  assign n1722 = ( n1072 & n1540 ) | ( n1072 & n1721 ) | ( n1540 & n1721 ) ;
  assign n1723 = n1365 ^ n1140 ^ n739 ;
  assign n1724 = n1723 ^ n950 ^ 1'b0 ;
  assign n1725 = n1655 | n1724 ;
  assign n1726 = n290 & ~n496 ;
  assign n1727 = n1726 ^ n397 ^ 1'b0 ;
  assign n1728 = n1727 ^ n1131 ^ n763 ;
  assign n1729 = ( n397 & n957 ) | ( n397 & n1194 ) | ( n957 & n1194 ) ;
  assign n1730 = n611 | n1729 ;
  assign n1731 = n1450 & ~n1730 ;
  assign n1733 = n285 | n854 ;
  assign n1734 = n1733 ^ n777 ^ 1'b0 ;
  assign n1732 = n1382 ^ n555 ^ n348 ;
  assign n1735 = n1734 ^ n1732 ^ 1'b0 ;
  assign n1736 = ( n186 & ~n278 ) | ( n186 & n429 ) | ( ~n278 & n429 ) ;
  assign n1737 = n168 & n347 ;
  assign n1738 = n1737 ^ n209 ^ 1'b0 ;
  assign n1739 = n1738 ^ n600 ^ n487 ;
  assign n1740 = n1736 | n1739 ;
  assign n1741 = n1012 ^ n668 ^ n194 ;
  assign n1742 = n875 & ~n1741 ;
  assign n1743 = n1742 ^ n1498 ^ 1'b0 ;
  assign n1744 = n540 & ~n1498 ;
  assign n1745 = n1744 ^ n253 ^ x115 ;
  assign n1746 = n586 & n1157 ;
  assign n1747 = ( n384 & n497 ) | ( n384 & n1075 ) | ( n497 & n1075 ) ;
  assign n1749 = ( n329 & ~n451 ) | ( n329 & n1129 ) | ( ~n451 & n1129 ) ;
  assign n1748 = ~n243 & n335 ;
  assign n1750 = n1749 ^ n1748 ^ n635 ;
  assign n1751 = ( x40 & n205 ) | ( x40 & n1342 ) | ( n205 & n1342 ) ;
  assign n1752 = n326 & n1751 ;
  assign n1753 = n1752 ^ n1095 ^ 1'b0 ;
  assign n1754 = n1753 ^ n1495 ^ n225 ;
  assign n1755 = n172 & n247 ;
  assign n1756 = n785 | n1755 ;
  assign n1757 = n1756 ^ n1549 ^ 1'b0 ;
  assign n1758 = ( n1750 & ~n1754 ) | ( n1750 & n1757 ) | ( ~n1754 & n1757 ) ;
  assign n1759 = ( n457 & n628 ) | ( n457 & n925 ) | ( n628 & n925 ) ;
  assign n1760 = n639 | n662 ;
  assign n1761 = n1759 | n1760 ;
  assign n1762 = n1761 ^ n952 ^ 1'b0 ;
  assign n1766 = x116 & n429 ;
  assign n1765 = n1067 ^ n780 ^ n321 ;
  assign n1767 = n1766 ^ n1765 ^ n551 ;
  assign n1764 = n696 ^ n688 ^ x122 ;
  assign n1763 = n1257 | n1318 ;
  assign n1768 = n1767 ^ n1764 ^ n1763 ;
  assign n1769 = ( n149 & ~n808 ) | ( n149 & n1768 ) | ( ~n808 & n1768 ) ;
  assign n1772 = n695 ^ n407 ^ n343 ;
  assign n1770 = n636 & n940 ;
  assign n1771 = ~n671 & n1770 ;
  assign n1773 = n1772 ^ n1771 ^ 1'b0 ;
  assign n1778 = n1226 ^ n1002 ^ n410 ;
  assign n1774 = n144 & n559 ;
  assign n1775 = ~x8 & n1774 ;
  assign n1776 = n1775 ^ n1158 ^ n640 ;
  assign n1777 = n1099 & ~n1776 ;
  assign n1779 = n1778 ^ n1777 ^ 1'b0 ;
  assign n1780 = n1197 ^ n1042 ^ n549 ;
  assign n1781 = n1780 ^ n617 ^ x16 ;
  assign n1785 = ( n129 & n526 ) | ( n129 & ~n1527 ) | ( n526 & ~n1527 ) ;
  assign n1786 = n1785 ^ x37 ^ 1'b0 ;
  assign n1787 = x10 & n1786 ;
  assign n1782 = n379 | n1326 ;
  assign n1783 = n569 | n1782 ;
  assign n1784 = n1783 ^ n471 ^ 1'b0 ;
  assign n1788 = n1787 ^ n1784 ^ 1'b0 ;
  assign n1789 = n1613 ^ n1521 ^ n1388 ;
  assign n1790 = n1707 ^ n535 ^ 1'b0 ;
  assign n1791 = n371 & ~n1790 ;
  assign n1792 = ~n1021 & n1791 ;
  assign n1793 = ( ~n661 & n1789 ) | ( ~n661 & n1792 ) | ( n1789 & n1792 ) ;
  assign n1795 = n645 ^ n186 ^ x17 ;
  assign n1796 = n1795 ^ n667 ^ n211 ;
  assign n1794 = x112 & n1370 ;
  assign n1797 = n1796 ^ n1794 ^ n883 ;
  assign n1799 = ( n871 & n902 ) | ( n871 & ~n965 ) | ( n902 & ~n965 ) ;
  assign n1798 = n1078 ^ n988 ^ x95 ;
  assign n1800 = n1799 ^ n1798 ^ n1223 ;
  assign n1801 = ( n201 & n380 ) | ( n201 & ~n930 ) | ( n380 & ~n930 ) ;
  assign n1804 = n1686 ^ n897 ^ 1'b0 ;
  assign n1802 = n243 | n1199 ;
  assign n1803 = x7 & ~n1802 ;
  assign n1805 = n1804 ^ n1803 ^ 1'b0 ;
  assign n1806 = ( n1184 & ~n1213 ) | ( n1184 & n1805 ) | ( ~n1213 & n1805 ) ;
  assign n1814 = n270 & ~n571 ;
  assign n1815 = ~x125 & n1814 ;
  assign n1816 = n862 & ~n1815 ;
  assign n1817 = n1816 ^ n704 ^ 1'b0 ;
  assign n1809 = ( n189 & n301 ) | ( n189 & n326 ) | ( n301 & n326 ) ;
  assign n1810 = ( ~n331 & n909 ) | ( ~n331 & n1809 ) | ( n909 & n1809 ) ;
  assign n1808 = n697 ^ x111 ^ x38 ;
  assign n1811 = n1810 ^ n1808 ^ 1'b0 ;
  assign n1812 = n975 | n1811 ;
  assign n1807 = n1069 & ~n1495 ;
  assign n1813 = n1812 ^ n1807 ^ 1'b0 ;
  assign n1818 = n1817 ^ n1813 ^ n680 ;
  assign n1819 = ( n1307 & ~n1716 ) | ( n1307 & n1818 ) | ( ~n1716 & n1818 ) ;
  assign n1820 = n585 ^ n406 ^ x92 ;
  assign n1821 = ~n194 & n390 ;
  assign n1822 = n1821 ^ x80 ^ 1'b0 ;
  assign n1823 = n178 & ~n1822 ;
  assign n1824 = ~n914 & n1823 ;
  assign n1825 = n632 & ~n684 ;
  assign n1826 = n1825 ^ n346 ^ 1'b0 ;
  assign n1827 = n1655 ^ n287 ^ 1'b0 ;
  assign n1828 = n1826 & n1827 ;
  assign n1829 = n1828 ^ n1588 ^ n537 ;
  assign n1830 = ~n1824 & n1829 ;
  assign n1831 = n1830 ^ n1120 ^ 1'b0 ;
  assign n1832 = n1820 & n1831 ;
  assign n1833 = n1572 ^ n1193 ^ n375 ;
  assign n1834 = ( n469 & n1269 ) | ( n469 & ~n1495 ) | ( n1269 & ~n1495 ) ;
  assign n1835 = n139 & ~n356 ;
  assign n1836 = ~x72 & n1835 ;
  assign n1837 = x110 & ~n190 ;
  assign n1838 = n1836 & n1837 ;
  assign n1839 = ( ~n192 & n336 ) | ( ~n192 & n1233 ) | ( n336 & n1233 ) ;
  assign n1840 = n1496 ^ n924 ^ x110 ;
  assign n1841 = n698 & n1840 ;
  assign n1842 = n1839 & n1841 ;
  assign n1843 = ( n1402 & n1838 ) | ( n1402 & ~n1842 ) | ( n1838 & ~n1842 ) ;
  assign n1844 = n529 & n905 ;
  assign n1845 = ~n130 & n1844 ;
  assign n1846 = n1845 ^ n1206 ^ 1'b0 ;
  assign n1847 = ~n1703 & n1846 ;
  assign n1855 = n1454 ^ n235 ^ 1'b0 ;
  assign n1856 = ~n1261 & n1855 ;
  assign n1857 = ( n487 & ~n1685 ) | ( n487 & n1856 ) | ( ~n1685 & n1856 ) ;
  assign n1852 = n1253 ^ x127 ^ 1'b0 ;
  assign n1853 = ( x92 & ~n907 ) | ( x92 & n1852 ) | ( ~n907 & n1852 ) ;
  assign n1849 = ( n484 & n559 ) | ( n484 & ~n757 ) | ( n559 & ~n757 ) ;
  assign n1850 = n1849 ^ n1317 ^ n571 ;
  assign n1851 = n1850 ^ n1382 ^ n762 ;
  assign n1848 = ( n416 & ~n1681 ) | ( n416 & n1713 ) | ( ~n1681 & n1713 ) ;
  assign n1854 = n1853 ^ n1851 ^ n1848 ;
  assign n1858 = n1857 ^ n1854 ^ n1428 ;
  assign n1859 = ( n434 & n1069 ) | ( n434 & n1420 ) | ( n1069 & n1420 ) ;
  assign n1860 = n633 & n1698 ;
  assign n1861 = ( n223 & ~n296 ) | ( n223 & n698 ) | ( ~n296 & n698 ) ;
  assign n1862 = ~n242 & n1861 ;
  assign n1863 = n1862 ^ n1475 ^ x75 ;
  assign n1864 = n972 ^ n275 ^ n139 ;
  assign n1865 = ( n357 & ~n841 ) | ( n357 & n1864 ) | ( ~n841 & n1864 ) ;
  assign n1866 = x112 ^ x30 ^ 1'b0 ;
  assign n1867 = n557 & n1866 ;
  assign n1868 = ( n441 & ~n945 ) | ( n441 & n1867 ) | ( ~n945 & n1867 ) ;
  assign n1869 = ( n952 & n1865 ) | ( n952 & ~n1868 ) | ( n1865 & ~n1868 ) ;
  assign n1870 = ( x0 & ~n1809 ) | ( x0 & n1869 ) | ( ~n1809 & n1869 ) ;
  assign n1871 = n1575 ^ n204 ^ 1'b0 ;
  assign n1872 = n1871 ^ n1761 ^ 1'b0 ;
  assign n1873 = x113 & ~n1872 ;
  assign n1874 = ( ~x119 & n168 ) | ( ~x119 & n870 ) | ( n168 & n870 ) ;
  assign n1875 = n1754 & n1874 ;
  assign n1876 = n1875 ^ n528 ^ 1'b0 ;
  assign n1879 = n411 & ~n426 ;
  assign n1880 = n1879 ^ n837 ^ 1'b0 ;
  assign n1877 = ( ~n655 & n740 ) | ( ~n655 & n780 ) | ( n740 & n780 ) ;
  assign n1878 = ( n555 & n1441 ) | ( n555 & n1877 ) | ( n1441 & n1877 ) ;
  assign n1881 = n1880 ^ n1878 ^ 1'b0 ;
  assign n1882 = ~n1876 & n1881 ;
  assign n1886 = n575 ^ n544 ^ n239 ;
  assign n1887 = n1886 ^ n925 ^ n826 ;
  assign n1883 = n1790 ^ n1470 ^ 1'b0 ;
  assign n1884 = ( x11 & n1804 ) | ( x11 & ~n1883 ) | ( n1804 & ~n1883 ) ;
  assign n1885 = ( x76 & x105 ) | ( x76 & n1884 ) | ( x105 & n1884 ) ;
  assign n1888 = n1887 ^ n1885 ^ 1'b0 ;
  assign n1889 = ( x43 & n1159 ) | ( x43 & ~n1218 ) | ( n1159 & ~n1218 ) ;
  assign n1890 = n1889 ^ n1092 ^ n1002 ;
  assign n1897 = n840 ^ n416 ^ 1'b0 ;
  assign n1898 = n924 | n1897 ;
  assign n1894 = n1125 ^ n998 ^ 1'b0 ;
  assign n1895 = n196 | n1894 ;
  assign n1896 = ( n744 & n1009 ) | ( n744 & n1895 ) | ( n1009 & n1895 ) ;
  assign n1891 = n278 & ~n1027 ;
  assign n1892 = ~n253 & n1891 ;
  assign n1893 = ~n486 & n1892 ;
  assign n1899 = n1898 ^ n1896 ^ n1893 ;
  assign n1904 = n1624 ^ n222 ^ 1'b0 ;
  assign n1900 = n1378 & ~n1790 ;
  assign n1901 = n846 ^ n838 ^ n303 ;
  assign n1902 = n1021 & ~n1901 ;
  assign n1903 = n1900 & ~n1902 ;
  assign n1905 = n1904 ^ n1903 ^ 1'b0 ;
  assign n1906 = n1260 ^ n469 ^ 1'b0 ;
  assign n1907 = ( ~n139 & n194 ) | ( ~n139 & n912 ) | ( n194 & n912 ) ;
  assign n1908 = n1907 ^ n1176 ^ n577 ;
  assign n1910 = n663 ^ n426 ^ n355 ;
  assign n1909 = n914 & n1549 ;
  assign n1911 = n1910 ^ n1909 ^ 1'b0 ;
  assign n1912 = ( n1287 & n1576 ) | ( n1287 & n1700 ) | ( n1576 & n1700 ) ;
  assign n1913 = n1606 ^ n768 ^ n596 ;
  assign n1914 = n1734 ^ n1410 ^ n213 ;
  assign n1915 = ( n1508 & n1913 ) | ( n1508 & ~n1914 ) | ( n1913 & ~n1914 ) ;
  assign n1916 = n1256 ^ n619 ^ n187 ;
  assign n1918 = ~n247 & n1254 ;
  assign n1919 = ~n411 & n1918 ;
  assign n1917 = n1331 ^ n1059 ^ x108 ;
  assign n1920 = n1919 ^ n1917 ^ n1676 ;
  assign n1921 = ( n326 & n1000 ) | ( n326 & n1518 ) | ( n1000 & n1518 ) ;
  assign n1922 = n1921 ^ n934 ^ 1'b0 ;
  assign n1923 = n373 & ~n857 ;
  assign n1924 = ~n1922 & n1923 ;
  assign n1925 = ( n1776 & ~n1920 ) | ( n1776 & n1924 ) | ( ~n1920 & n1924 ) ;
  assign n1926 = n1916 | n1925 ;
  assign n1927 = n1699 & ~n1926 ;
  assign n1928 = n1524 | n1927 ;
  assign n1929 = n1928 ^ n591 ^ 1'b0 ;
  assign n1930 = n1759 ^ n306 ^ n226 ;
  assign n1931 = ( ~n710 & n867 ) | ( ~n710 & n1930 ) | ( n867 & n1930 ) ;
  assign n1932 = n751 ^ n459 ^ 1'b0 ;
  assign n1933 = x95 & n1932 ;
  assign n1934 = n1933 ^ n1703 ^ 1'b0 ;
  assign n1935 = ( ~n1159 & n1931 ) | ( ~n1159 & n1934 ) | ( n1931 & n1934 ) ;
  assign n1936 = n1632 ^ x96 ^ x76 ;
  assign n1937 = n738 | n1936 ;
  assign n1938 = n1935 | n1937 ;
  assign n1939 = n1938 ^ n1110 ^ x124 ;
  assign n1940 = n940 & ~n1682 ;
  assign n1941 = ( n1016 & n1488 ) | ( n1016 & ~n1940 ) | ( n1488 & ~n1940 ) ;
  assign n1942 = ( n137 & n1325 ) | ( n137 & n1815 ) | ( n1325 & n1815 ) ;
  assign n1943 = n525 & n1942 ;
  assign n1944 = n1943 ^ n189 ^ 1'b0 ;
  assign n1945 = n643 ^ n202 ^ x50 ;
  assign n1946 = n1945 ^ n417 ^ 1'b0 ;
  assign n1947 = n1946 ^ n866 ^ n559 ;
  assign n1948 = n1947 ^ n1097 ^ n223 ;
  assign n1949 = n1493 ^ n392 ^ 1'b0 ;
  assign n1950 = ( n520 & ~n1215 ) | ( n520 & n1949 ) | ( ~n1215 & n1949 ) ;
  assign n1951 = ( n204 & n430 ) | ( n204 & ~n1231 ) | ( n430 & ~n1231 ) ;
  assign n1952 = n1951 ^ n630 ^ 1'b0 ;
  assign n1958 = ( x109 & n357 ) | ( x109 & n545 ) | ( n357 & n545 ) ;
  assign n1959 = n1958 ^ n1317 ^ x40 ;
  assign n1960 = n332 & ~n384 ;
  assign n1961 = ~n1959 & n1960 ;
  assign n1957 = n1254 ^ n941 ^ n811 ;
  assign n1954 = ( ~n176 & n346 ) | ( ~n176 & n748 ) | ( n346 & n748 ) ;
  assign n1953 = n979 ^ n704 ^ n460 ;
  assign n1955 = n1954 ^ n1953 ^ n137 ;
  assign n1956 = n1955 ^ n1016 ^ n782 ;
  assign n1962 = n1961 ^ n1957 ^ n1956 ;
  assign n1963 = ( n581 & ~n738 ) | ( n581 & n755 ) | ( ~n738 & n755 ) ;
  assign n1964 = n1963 ^ n1551 ^ n1352 ;
  assign n1966 = n1032 ^ n255 ^ n165 ;
  assign n1965 = ( n557 & n1764 ) | ( n557 & ~n1891 ) | ( n1764 & ~n1891 ) ;
  assign n1967 = n1966 ^ n1965 ^ n967 ;
  assign n1968 = n270 & n1291 ;
  assign n1969 = ~n935 & n1968 ;
  assign n1970 = x39 & ~n287 ;
  assign n1971 = n1970 ^ n640 ^ 1'b0 ;
  assign n1972 = n755 ^ n600 ^ n362 ;
  assign n1973 = ( n508 & n1971 ) | ( n508 & n1972 ) | ( n1971 & n1972 ) ;
  assign n1974 = n1973 ^ n506 ^ 1'b0 ;
  assign n1975 = x83 & n1974 ;
  assign n1976 = n1579 | n1975 ;
  assign n1977 = ( n1134 & n1546 ) | ( n1134 & ~n1976 ) | ( n1546 & ~n1976 ) ;
  assign n1978 = n398 ^ x55 ^ 1'b0 ;
  assign n1979 = ~n613 & n1978 ;
  assign n1980 = ~n1145 & n1979 ;
  assign n1983 = n1374 ^ n685 ^ n684 ;
  assign n1982 = ( n317 & n517 ) | ( n317 & ~n854 ) | ( n517 & ~n854 ) ;
  assign n1981 = ( x18 & ~n343 ) | ( x18 & n386 ) | ( ~n343 & n386 ) ;
  assign n1984 = n1983 ^ n1982 ^ n1981 ;
  assign n1985 = n1984 ^ n1360 ^ 1'b0 ;
  assign n1986 = n1980 | n1985 ;
  assign n1987 = n794 ^ n758 ^ x4 ;
  assign n1988 = x33 & x111 ;
  assign n1989 = n1988 ^ n167 ^ 1'b0 ;
  assign n1990 = n1989 ^ n855 ^ n745 ;
  assign n1991 = n1990 ^ n1023 ^ n467 ;
  assign n1992 = ( ~x66 & n269 ) | ( ~x66 & n1991 ) | ( n269 & n1991 ) ;
  assign n1999 = n1062 & n1327 ;
  assign n2000 = n510 | n1999 ;
  assign n1993 = ~n163 & n439 ;
  assign n1994 = ( n284 & n1422 ) | ( n284 & ~n1993 ) | ( n1422 & ~n1993 ) ;
  assign n1995 = n1815 ^ n1496 ^ 1'b0 ;
  assign n1996 = n780 | n1995 ;
  assign n1997 = n1001 | n1996 ;
  assign n1998 = ( n1246 & n1994 ) | ( n1246 & ~n1997 ) | ( n1994 & ~n1997 ) ;
  assign n2001 = n2000 ^ n1998 ^ 1'b0 ;
  assign n2002 = n1898 | n2001 ;
  assign n2003 = ( n553 & ~n846 ) | ( n553 & n1513 ) | ( ~n846 & n1513 ) ;
  assign n2004 = n2003 ^ n1179 ^ 1'b0 ;
  assign n2005 = n2002 | n2004 ;
  assign n2006 = ~n255 & n1661 ;
  assign n2007 = n2006 ^ n898 ^ 1'b0 ;
  assign n2008 = n1883 ^ n487 ^ n375 ;
  assign n2009 = n440 ^ n169 ^ x102 ;
  assign n2010 = x117 & ~n638 ;
  assign n2011 = n2009 & n2010 ;
  assign n2012 = ~n312 & n456 ;
  assign n2013 = n2011 & n2012 ;
  assign n2014 = n1840 ^ n1813 ^ n646 ;
  assign n2015 = ~n2013 & n2014 ;
  assign n2016 = n1591 ^ n1411 ^ n1081 ;
  assign n2017 = n2016 ^ n1799 ^ n1533 ;
  assign n2018 = n293 | n529 ;
  assign n2019 = ( n292 & n354 ) | ( n292 & ~n814 ) | ( n354 & ~n814 ) ;
  assign n2020 = n2019 ^ n1101 ^ n1099 ;
  assign n2021 = x64 & n2020 ;
  assign n2022 = n268 & n2021 ;
  assign n2023 = ~x62 & n398 ;
  assign n2024 = ( n634 & ~n2022 ) | ( n634 & n2023 ) | ( ~n2022 & n2023 ) ;
  assign n2025 = ( n1046 & ~n2018 ) | ( n1046 & n2024 ) | ( ~n2018 & n2024 ) ;
  assign n2027 = n332 & n489 ;
  assign n2028 = n816 & n2027 ;
  assign n2029 = n2028 ^ x57 ^ 1'b0 ;
  assign n2026 = n188 & n852 ;
  assign n2030 = n2029 ^ n2026 ^ n1627 ;
  assign n2031 = ( n357 & n877 ) | ( n357 & n979 ) | ( n877 & n979 ) ;
  assign n2032 = n2031 ^ n1347 ^ n1020 ;
  assign n2038 = ( x110 & n321 ) | ( x110 & ~n541 ) | ( n321 & ~n541 ) ;
  assign n2039 = n1241 ^ n837 ^ n477 ;
  assign n2040 = ( n1074 & n2038 ) | ( n1074 & ~n2039 ) | ( n2038 & ~n2039 ) ;
  assign n2041 = n1133 ^ n508 ^ 1'b0 ;
  assign n2042 = n445 | n2041 ;
  assign n2043 = n2040 | n2042 ;
  assign n2044 = n2043 ^ n373 ^ 1'b0 ;
  assign n2045 = n526 ^ n506 ^ n432 ;
  assign n2046 = n543 | n2045 ;
  assign n2047 = n942 & ~n2046 ;
  assign n2048 = x112 & ~n2047 ;
  assign n2049 = ~n2044 & n2048 ;
  assign n2050 = n195 & n256 ;
  assign n2051 = n1482 | n2050 ;
  assign n2052 = n2049 & ~n2051 ;
  assign n2033 = ~n880 & n1303 ;
  assign n2034 = n2033 ^ n657 ^ n272 ;
  assign n2035 = n2034 ^ n1498 ^ 1'b0 ;
  assign n2036 = n2034 ^ n1697 ^ n928 ;
  assign n2037 = ~n2035 & n2036 ;
  assign n2053 = n2052 ^ n2037 ^ 1'b0 ;
  assign n2054 = n356 ^ n291 ^ x26 ;
  assign n2055 = n2054 ^ n1054 ^ n993 ;
  assign n2056 = n639 ^ x52 ^ 1'b0 ;
  assign n2057 = n425 & ~n2056 ;
  assign n2058 = n2057 ^ n1613 ^ x40 ;
  assign n2059 = ( x45 & n2055 ) | ( x45 & n2058 ) | ( n2055 & n2058 ) ;
  assign n2060 = n1584 | n1630 ;
  assign n2064 = n218 & ~n670 ;
  assign n2065 = n2064 ^ n1349 ^ 1'b0 ;
  assign n2066 = n2065 ^ n853 ^ x35 ;
  assign n2061 = n643 ^ x14 ^ x0 ;
  assign n2062 = n1702 ^ n1207 ^ 1'b0 ;
  assign n2063 = n2061 & n2062 ;
  assign n2067 = n2066 ^ n2063 ^ 1'b0 ;
  assign n2068 = n2060 | n2067 ;
  assign n2069 = ( n300 & ~n664 ) | ( n300 & n681 ) | ( ~n664 & n681 ) ;
  assign n2070 = n1887 ^ n1265 ^ n1021 ;
  assign n2071 = ( n913 & n2069 ) | ( n913 & ~n2070 ) | ( n2069 & ~n2070 ) ;
  assign n2072 = n588 ^ n420 ^ 1'b0 ;
  assign n2073 = ( n259 & n459 ) | ( n259 & n646 ) | ( n459 & n646 ) ;
  assign n2074 = ( n430 & n451 ) | ( n430 & n1749 ) | ( n451 & n1749 ) ;
  assign n2075 = ( n898 & ~n1904 ) | ( n898 & n2074 ) | ( ~n1904 & n2074 ) ;
  assign n2076 = n242 | n763 ;
  assign n2077 = n573 & ~n2076 ;
  assign n2078 = ( ~n176 & n2075 ) | ( ~n176 & n2077 ) | ( n2075 & n2077 ) ;
  assign n2079 = ( ~n2072 & n2073 ) | ( ~n2072 & n2078 ) | ( n2073 & n2078 ) ;
  assign n2084 = n377 & n594 ;
  assign n2085 = n2084 ^ n429 ^ 1'b0 ;
  assign n2080 = n505 ^ n341 ^ x98 ;
  assign n2081 = ( n1247 & n1706 ) | ( n1247 & ~n1776 ) | ( n1706 & ~n1776 ) ;
  assign n2082 = n2081 ^ n1451 ^ 1'b0 ;
  assign n2083 = n2080 & ~n2082 ;
  assign n2086 = n2085 ^ n2083 ^ n1413 ;
  assign n2087 = ( n926 & n1417 ) | ( n926 & ~n1599 ) | ( n1417 & ~n1599 ) ;
  assign n2088 = n1751 & n2087 ;
  assign n2089 = n2088 ^ n525 ^ 1'b0 ;
  assign n2090 = ( x110 & n216 ) | ( x110 & n1042 ) | ( n216 & n1042 ) ;
  assign n2091 = ( x109 & ~n1865 ) | ( x109 & n2090 ) | ( ~n1865 & n2090 ) ;
  assign n2096 = n354 & ~n369 ;
  assign n2097 = n382 & n2096 ;
  assign n2092 = n1490 ^ n716 ^ n553 ;
  assign n2093 = n2092 ^ n1629 ^ 1'b0 ;
  assign n2094 = n1437 | n2093 ;
  assign n2095 = x74 & ~n2094 ;
  assign n2098 = n2097 ^ n2095 ^ 1'b0 ;
  assign n2099 = ( x62 & n2091 ) | ( x62 & ~n2098 ) | ( n2091 & ~n2098 ) ;
  assign n2101 = n320 ^ x103 ^ x72 ;
  assign n2100 = n367 & ~n1541 ;
  assign n2102 = n2101 ^ n2100 ^ 1'b0 ;
  assign n2103 = ( x14 & n659 ) | ( x14 & ~n1289 ) | ( n659 & ~n1289 ) ;
  assign n2110 = ( x73 & n149 ) | ( x73 & n466 ) | ( n149 & n466 ) ;
  assign n2109 = ( x8 & ~n694 ) | ( x8 & n902 ) | ( ~n694 & n902 ) ;
  assign n2111 = n2110 ^ n2109 ^ x105 ;
  assign n2112 = n2111 ^ n1038 ^ 1'b0 ;
  assign n2113 = n902 | n2112 ;
  assign n2108 = ( n551 & n759 ) | ( n551 & ~n1129 ) | ( n759 & ~n1129 ) ;
  assign n2104 = ~n757 & n1378 ;
  assign n2105 = ~x95 & n2104 ;
  assign n2106 = n2105 ^ n498 ^ 1'b0 ;
  assign n2107 = n170 | n2106 ;
  assign n2114 = n2113 ^ n2108 ^ n2107 ;
  assign n2115 = ( n1326 & n1660 ) | ( n1326 & n1715 ) | ( n1660 & n1715 ) ;
  assign n2117 = n1768 ^ n561 ^ n473 ;
  assign n2116 = ( n132 & ~n1085 ) | ( n132 & n1321 ) | ( ~n1085 & n1321 ) ;
  assign n2118 = n2117 ^ n2116 ^ n1349 ;
  assign n2119 = n823 & ~n2118 ;
  assign n2120 = n2119 ^ n1978 ^ 1'b0 ;
  assign n2121 = n1422 ^ n1195 ^ n662 ;
  assign n2122 = n2121 ^ n1692 ^ n642 ;
  assign n2123 = n912 ^ n348 ^ 1'b0 ;
  assign n2124 = n378 & ~n2123 ;
  assign n2125 = ~n284 & n2124 ;
  assign n2126 = n1335 ^ n1108 ^ n200 ;
  assign n2127 = n2126 ^ n847 ^ 1'b0 ;
  assign n2128 = x64 & n2127 ;
  assign n2129 = ( ~n1140 & n1206 ) | ( ~n1140 & n2128 ) | ( n1206 & n2128 ) ;
  assign n2130 = n2129 ^ n2061 ^ n798 ;
  assign n2131 = n2125 & ~n2130 ;
  assign n2132 = ~n2122 & n2131 ;
  assign n2133 = x59 & ~n1567 ;
  assign n2134 = n2133 ^ n389 ^ 1'b0 ;
  assign n2138 = x37 & x57 ;
  assign n2137 = n778 ^ n455 ^ 1'b0 ;
  assign n2139 = n2138 ^ n2137 ^ n1220 ;
  assign n2140 = ( n799 & ~n1228 ) | ( n799 & n2139 ) | ( ~n1228 & n2139 ) ;
  assign n2136 = n426 | n1191 ;
  assign n2141 = n2140 ^ n2136 ^ n1054 ;
  assign n2135 = n380 | n1668 ;
  assign n2142 = n2141 ^ n2135 ^ n280 ;
  assign n2143 = ( ~n2052 & n2134 ) | ( ~n2052 & n2142 ) | ( n2134 & n2142 ) ;
  assign n2152 = n1349 ^ n970 ^ 1'b0 ;
  assign n2148 = n942 ^ n195 ^ 1'b0 ;
  assign n2149 = n695 & ~n2148 ;
  assign n2150 = n1138 & n2149 ;
  assign n2151 = ~x12 & n2150 ;
  assign n2145 = n698 | n974 ;
  assign n2146 = ( n675 & ~n1480 ) | ( n675 & n2145 ) | ( ~n1480 & n2145 ) ;
  assign n2147 = n643 | n2146 ;
  assign n2153 = n2152 ^ n2151 ^ n2147 ;
  assign n2154 = ( x29 & n2054 ) | ( x29 & n2153 ) | ( n2054 & n2153 ) ;
  assign n2144 = n1820 ^ n441 ^ n226 ;
  assign n2155 = n2154 ^ n2144 ^ n1710 ;
  assign n2156 = n2070 ^ n1958 ^ n1365 ;
  assign n2157 = ( n1285 & n1767 ) | ( n1285 & n2156 ) | ( n1767 & n2156 ) ;
  assign n2158 = n2157 ^ n1587 ^ n133 ;
  assign n2159 = n2158 ^ n1311 ^ 1'b0 ;
  assign n2160 = n838 | n1223 ;
  assign n2161 = n981 & n1904 ;
  assign n2162 = n2160 & n2161 ;
  assign n2168 = n2070 ^ n1828 ^ x55 ;
  assign n2169 = n2168 ^ n1739 ^ n217 ;
  assign n2164 = ( n223 & ~n256 ) | ( n223 & n365 ) | ( ~n256 & n365 ) ;
  assign n2165 = n2164 ^ n418 ^ n130 ;
  assign n2166 = n2165 ^ n1042 ^ n202 ;
  assign n2163 = n2087 ^ n1451 ^ n252 ;
  assign n2167 = n2166 ^ n2163 ^ 1'b0 ;
  assign n2170 = n2169 ^ n2167 ^ n603 ;
  assign n2171 = ~n611 & n1633 ;
  assign n2172 = n2171 ^ n494 ^ 1'b0 ;
  assign n2173 = n2172 ^ n374 ^ 1'b0 ;
  assign n2174 = n2173 ^ n398 ^ n225 ;
  assign n2175 = ( ~n352 & n563 ) | ( ~n352 & n600 ) | ( n563 & n600 ) ;
  assign n2176 = n2175 ^ n853 ^ n545 ;
  assign n2177 = n1110 & ~n1203 ;
  assign n2178 = n2176 & n2177 ;
  assign n2179 = ( n250 & n1889 ) | ( n250 & n2178 ) | ( n1889 & n2178 ) ;
  assign n2180 = x61 & n558 ;
  assign n2181 = ~x104 & n2180 ;
  assign n2182 = n264 & n973 ;
  assign n2183 = ~n597 & n2182 ;
  assign n2184 = ( n289 & n594 ) | ( n289 & ~n1982 ) | ( n594 & ~n1982 ) ;
  assign n2185 = n2184 ^ n1627 ^ 1'b0 ;
  assign n2187 = n809 ^ n252 ^ n188 ;
  assign n2186 = x63 & ~n553 ;
  assign n2188 = n2187 ^ n2186 ^ 1'b0 ;
  assign n2189 = n1009 ^ x97 ^ 1'b0 ;
  assign n2190 = n2188 | n2189 ;
  assign n2191 = ( n2183 & ~n2185 ) | ( n2183 & n2190 ) | ( ~n2185 & n2190 ) ;
  assign n2192 = ( n725 & ~n2181 ) | ( n725 & n2191 ) | ( ~n2181 & n2191 ) ;
  assign n2193 = n1619 ^ n580 ^ 1'b0 ;
  assign n2194 = ~n1457 & n2193 ;
  assign n2195 = n357 ^ n203 ^ 1'b0 ;
  assign n2196 = n2194 & n2195 ;
  assign n2197 = ( x8 & x111 ) | ( x8 & n224 ) | ( x111 & n224 ) ;
  assign n2198 = ( x18 & n1173 ) | ( x18 & n2197 ) | ( n1173 & n2197 ) ;
  assign n2199 = n578 | n2139 ;
  assign n2200 = n2198 | n2199 ;
  assign n2201 = n2200 ^ n992 ^ n909 ;
  assign n2202 = n1592 ^ n651 ^ 1'b0 ;
  assign n2203 = n775 & ~n1428 ;
  assign n2204 = n2203 ^ n463 ^ 1'b0 ;
  assign n2205 = ~n267 & n935 ;
  assign n2206 = n921 ^ n538 ^ x83 ;
  assign n2207 = n844 & n2206 ;
  assign n2208 = n2207 ^ n1680 ^ 1'b0 ;
  assign n2209 = ~n873 & n2208 ;
  assign n2210 = n1765 ^ n310 ^ 1'b0 ;
  assign n2211 = n2210 ^ n1444 ^ 1'b0 ;
  assign n2212 = ( n1489 & n1723 ) | ( n1489 & ~n2211 ) | ( n1723 & ~n2211 ) ;
  assign n2213 = ( n1054 & n2162 ) | ( n1054 & ~n2212 ) | ( n2162 & ~n2212 ) ;
  assign n2216 = n1376 ^ x79 ^ 1'b0 ;
  assign n2217 = n2216 ^ x16 ^ 1'b0 ;
  assign n2218 = n232 & ~n2217 ;
  assign n2219 = ( n1023 & n1227 ) | ( n1023 & ~n2218 ) | ( n1227 & ~n2218 ) ;
  assign n2214 = n1064 ^ n436 ^ 1'b0 ;
  assign n2215 = n1337 & n2214 ;
  assign n2220 = n2219 ^ n2215 ^ 1'b0 ;
  assign n2222 = n1362 ^ n1226 ^ x91 ;
  assign n2223 = n2031 ^ n380 ^ 1'b0 ;
  assign n2224 = n2222 & n2223 ;
  assign n2225 = n991 & n2224 ;
  assign n2221 = ( ~n845 & n1700 ) | ( ~n845 & n2198 ) | ( n1700 & n2198 ) ;
  assign n2226 = n2225 ^ n2221 ^ n1635 ;
  assign n2228 = ( n156 & n241 ) | ( n156 & ~n1723 ) | ( n241 & ~n1723 ) ;
  assign n2229 = n2228 ^ n646 ^ 1'b0 ;
  assign n2230 = ~n154 & n2229 ;
  assign n2227 = ( x22 & x121 ) | ( x22 & ~n482 ) | ( x121 & ~n482 ) ;
  assign n2231 = n2230 ^ n2227 ^ n1778 ;
  assign n2232 = x20 & n2231 ;
  assign n2233 = x11 & n1097 ;
  assign n2234 = n2233 ^ n1331 ^ 1'b0 ;
  assign n2235 = n2234 ^ n1668 ^ 1'b0 ;
  assign n2236 = n1079 ^ n1043 ^ x112 ;
  assign n2237 = n2228 ^ n894 ^ 1'b0 ;
  assign n2238 = ( ~x80 & n2236 ) | ( ~x80 & n2237 ) | ( n2236 & n2237 ) ;
  assign n2239 = ( ~n466 & n797 ) | ( ~n466 & n1302 ) | ( n797 & n1302 ) ;
  assign n2240 = ( n429 & ~n440 ) | ( n429 & n663 ) | ( ~n440 & n663 ) ;
  assign n2241 = n2239 & ~n2240 ;
  assign n2242 = n2241 ^ n913 ^ 1'b0 ;
  assign n2243 = ( n285 & n1048 ) | ( n285 & ~n1428 ) | ( n1048 & ~n1428 ) ;
  assign n2244 = ( n1242 & ~n2242 ) | ( n1242 & n2243 ) | ( ~n2242 & n2243 ) ;
  assign n2245 = n988 ^ n375 ^ 1'b0 ;
  assign n2246 = n460 | n2245 ;
  assign n2247 = ( x120 & n1023 ) | ( x120 & n2246 ) | ( n1023 & n2246 ) ;
  assign n2248 = ( n315 & ~n928 ) | ( n315 & n1560 ) | ( ~n928 & n1560 ) ;
  assign n2249 = ( n1366 & n2247 ) | ( n1366 & ~n2248 ) | ( n2247 & ~n2248 ) ;
  assign n2250 = n1947 ^ n1579 ^ n737 ;
  assign n2251 = n1627 ^ n1519 ^ n497 ;
  assign n2252 = n1027 ^ n622 ^ x110 ;
  assign n2253 = ( n696 & n1818 ) | ( n696 & n2252 ) | ( n1818 & n2252 ) ;
  assign n2257 = ( ~n132 & n366 ) | ( ~n132 & n1297 ) | ( n366 & n1297 ) ;
  assign n2258 = n2257 ^ n333 ^ x45 ;
  assign n2255 = n458 ^ n357 ^ n214 ;
  assign n2254 = n583 | n1204 ;
  assign n2256 = n2255 ^ n2254 ^ 1'b0 ;
  assign n2259 = n2258 ^ n2256 ^ 1'b0 ;
  assign n2260 = n2232 & n2259 ;
  assign n2261 = n2178 ^ n1952 ^ n1475 ;
  assign n2264 = n2252 ^ n1411 ^ n478 ;
  assign n2262 = ( ~x39 & n799 ) | ( ~x39 & n1606 ) | ( n799 & n1606 ) ;
  assign n2263 = ~n1566 & n2262 ;
  assign n2265 = n2264 ^ n2263 ^ 1'b0 ;
  assign n2266 = n1078 ^ n758 ^ 1'b0 ;
  assign n2267 = n341 & n2266 ;
  assign n2268 = n2230 & n2267 ;
  assign n2269 = ~n459 & n2268 ;
  assign n2270 = ( n1644 & n2265 ) | ( n1644 & ~n2269 ) | ( n2265 & ~n2269 ) ;
  assign n2271 = n1436 ^ n1173 ^ n393 ;
  assign n2272 = n310 ^ n247 ^ 1'b0 ;
  assign n2273 = n241 & n2272 ;
  assign n2274 = ( n222 & n1309 ) | ( n222 & ~n2273 ) | ( n1309 & ~n2273 ) ;
  assign n2275 = n2274 ^ n2239 ^ n1668 ;
  assign n2276 = ( n485 & n1942 ) | ( n485 & n2275 ) | ( n1942 & n2275 ) ;
  assign n2277 = n2138 & n2276 ;
  assign n2278 = n2277 ^ n1277 ^ 1'b0 ;
  assign n2279 = n855 ^ n738 ^ n187 ;
  assign n2280 = ( n436 & ~n1698 ) | ( n436 & n2279 ) | ( ~n1698 & n2279 ) ;
  assign n2281 = n1542 ^ n894 ^ n460 ;
  assign n2282 = ( n497 & n635 ) | ( n497 & ~n2281 ) | ( n635 & ~n2281 ) ;
  assign n2283 = ( ~n282 & n458 ) | ( ~n282 & n2282 ) | ( n458 & n2282 ) ;
  assign n2291 = n2273 ^ n151 ^ 1'b0 ;
  assign n2292 = x3 & ~n2291 ;
  assign n2293 = ( n1069 & n1421 ) | ( n1069 & n2292 ) | ( n1421 & n2292 ) ;
  assign n2294 = ( x96 & ~n1201 ) | ( x96 & n2293 ) | ( ~n1201 & n2293 ) ;
  assign n2288 = n902 | n1537 ;
  assign n2289 = n2288 ^ n1454 ^ 1'b0 ;
  assign n2290 = n591 & n2289 ;
  assign n2295 = n2294 ^ n2290 ^ 1'b0 ;
  assign n2284 = n1614 ^ x84 ^ 1'b0 ;
  assign n2285 = n271 & ~n2284 ;
  assign n2286 = n2285 ^ n1013 ^ 1'b0 ;
  assign n2287 = n2286 ^ n1122 ^ 1'b0 ;
  assign n2296 = n2295 ^ n2287 ^ n2073 ;
  assign n2300 = x117 & n1510 ;
  assign n2301 = ~n476 & n2300 ;
  assign n2297 = x98 & ~n159 ;
  assign n2298 = n900 & n2297 ;
  assign n2299 = n2298 ^ n1591 ^ n945 ;
  assign n2302 = n2301 ^ n2299 ^ n1917 ;
  assign n2303 = ( n2283 & n2296 ) | ( n2283 & ~n2302 ) | ( n2296 & ~n2302 ) ;
  assign n2305 = n1428 ^ n580 ^ 1'b0 ;
  assign n2306 = n2305 ^ n468 ^ 1'b0 ;
  assign n2307 = ( n643 & n2286 ) | ( n643 & n2306 ) | ( n2286 & n2306 ) ;
  assign n2304 = n953 | n2070 ;
  assign n2308 = n2307 ^ n2304 ^ 1'b0 ;
  assign n2309 = ( n163 & n1490 ) | ( n163 & n1980 ) | ( n1490 & n1980 ) ;
  assign n2311 = n1836 ^ n779 ^ n748 ;
  assign n2310 = n410 & n1004 ;
  assign n2312 = n2311 ^ n2310 ^ 1'b0 ;
  assign n2313 = n2312 ^ n2049 ^ n639 ;
  assign n2315 = n580 & ~n780 ;
  assign n2314 = ( x98 & ~n767 ) | ( x98 & n941 ) | ( ~n767 & n941 ) ;
  assign n2316 = n2315 ^ n2314 ^ n1034 ;
  assign n2317 = ( ~x28 & n2313 ) | ( ~x28 & n2316 ) | ( n2313 & n2316 ) ;
  assign n2318 = n468 | n2317 ;
  assign n2319 = n2309 & ~n2318 ;
  assign n2325 = ( n802 & ~n1267 ) | ( n802 & n2039 ) | ( ~n1267 & n2039 ) ;
  assign n2320 = n2112 ^ x122 ^ 1'b0 ;
  assign n2321 = ( n365 & ~n535 ) | ( n365 & n1329 ) | ( ~n535 & n1329 ) ;
  assign n2322 = n2321 ^ n986 ^ n900 ;
  assign n2323 = ( n140 & ~n716 ) | ( n140 & n2322 ) | ( ~n716 & n2322 ) ;
  assign n2324 = ( n924 & n2320 ) | ( n924 & ~n2323 ) | ( n2320 & ~n2323 ) ;
  assign n2326 = n2325 ^ n2324 ^ n213 ;
  assign n2327 = n1762 ^ n1012 ^ x85 ;
  assign n2329 = n1634 ^ n360 ^ x122 ;
  assign n2328 = n352 ^ n314 ^ x31 ;
  assign n2330 = n2329 ^ n2328 ^ x71 ;
  assign n2334 = ( n324 & ~n816 ) | ( n324 & n2172 ) | ( ~n816 & n2172 ) ;
  assign n2331 = ( ~n814 & n1120 ) | ( ~n814 & n1126 ) | ( n1120 & n1126 ) ;
  assign n2332 = n2331 ^ n668 ^ n524 ;
  assign n2333 = ( n226 & n2023 ) | ( n226 & n2332 ) | ( n2023 & n2332 ) ;
  assign n2335 = n2334 ^ n2333 ^ n1374 ;
  assign n2336 = n1437 ^ n1202 ^ 1'b0 ;
  assign n2337 = n2336 ^ n694 ^ n344 ;
  assign n2338 = n407 | n2337 ;
  assign n2339 = ( n2330 & n2335 ) | ( n2330 & n2338 ) | ( n2335 & n2338 ) ;
  assign n2340 = n1966 ^ n919 ^ n728 ;
  assign n2341 = n2340 ^ x112 ^ x23 ;
  assign n2342 = n768 & n1510 ;
  assign n2343 = n2342 ^ n774 ^ 1'b0 ;
  assign n2344 = ~n1858 & n2214 ;
  assign n2345 = n2344 ^ n1273 ^ 1'b0 ;
  assign n2346 = ( n609 & n2343 ) | ( n609 & ~n2345 ) | ( n2343 & ~n2345 ) ;
  assign n2347 = n854 | n1599 ;
  assign n2348 = n2347 ^ n1544 ^ 1'b0 ;
  assign n2349 = ( x79 & ~n1673 ) | ( x79 & n1707 ) | ( ~n1673 & n1707 ) ;
  assign n2350 = ( n2169 & n2348 ) | ( n2169 & n2349 ) | ( n2348 & n2349 ) ;
  assign n2351 = ( n393 & ~n489 ) | ( n393 & n762 ) | ( ~n489 & n762 ) ;
  assign n2352 = x43 & ~n2351 ;
  assign n2353 = n2352 ^ n577 ^ 1'b0 ;
  assign n2360 = n1100 | n1490 ;
  assign n2357 = ( n387 & n698 ) | ( n387 & n889 ) | ( n698 & n889 ) ;
  assign n2358 = n2357 ^ n628 ^ n473 ;
  assign n2354 = n1356 & ~n1461 ;
  assign n2355 = n2354 ^ n835 ^ 1'b0 ;
  assign n2356 = ~n462 & n2355 ;
  assign n2359 = n2358 ^ n2356 ^ n1356 ;
  assign n2361 = n2360 ^ n2359 ^ 1'b0 ;
  assign n2362 = n2353 & n2361 ;
  assign n2363 = n2362 ^ n1367 ^ n413 ;
  assign n2364 = ( ~n383 & n2350 ) | ( ~n383 & n2363 ) | ( n2350 & n2363 ) ;
  assign n2365 = ~n301 & n386 ;
  assign n2366 = n1183 & n2365 ;
  assign n2367 = n1258 & ~n2366 ;
  assign n2368 = ( ~n1567 & n2101 ) | ( ~n1567 & n2367 ) | ( n2101 & n2367 ) ;
  assign n2370 = n1236 ^ n553 ^ n270 ;
  assign n2369 = n507 | n1989 ;
  assign n2371 = n2370 ^ n2369 ^ n935 ;
  assign n2372 = n1317 ^ n1256 ^ 1'b0 ;
  assign n2373 = n2372 ^ n1001 ^ n545 ;
  assign n2374 = ~n2085 & n2373 ;
  assign n2375 = n2374 ^ x11 ^ 1'b0 ;
  assign n2376 = n710 & ~n2375 ;
  assign n2377 = n277 & ~n855 ;
  assign n2378 = n2377 ^ n1635 ^ 1'b0 ;
  assign n2379 = n1055 & ~n2378 ;
  assign n2385 = n1250 ^ x48 ^ x32 ;
  assign n2386 = n271 & ~n2385 ;
  assign n2380 = n631 ^ n608 ^ n160 ;
  assign n2381 = n773 | n1799 ;
  assign n2382 = x29 & ~n2381 ;
  assign n2383 = n2380 & n2382 ;
  assign n2384 = x50 & ~n2383 ;
  assign n2387 = n2386 ^ n2384 ^ n1584 ;
  assign n2388 = n1919 ^ n1895 ^ n1817 ;
  assign n2389 = ( ~n411 & n2273 ) | ( ~n411 & n2388 ) | ( n2273 & n2388 ) ;
  assign n2390 = n2343 ^ n2163 ^ 1'b0 ;
  assign n2392 = ( n596 & n684 ) | ( n596 & ~n1377 ) | ( n684 & ~n1377 ) ;
  assign n2393 = n2392 ^ n801 ^ 1'b0 ;
  assign n2391 = ~n405 & n1647 ;
  assign n2394 = n2393 ^ n2391 ^ x66 ;
  assign n2395 = n2394 ^ n1576 ^ 1'b0 ;
  assign n2396 = n1376 | n2395 ;
  assign n2397 = n1257 ^ n402 ^ 1'b0 ;
  assign n2398 = n1762 & n2397 ;
  assign n2399 = n1327 ^ n807 ^ 1'b0 ;
  assign n2400 = n1110 & n2399 ;
  assign n2401 = n924 ^ n478 ^ 1'b0 ;
  assign n2402 = ( n259 & ~n2400 ) | ( n259 & n2401 ) | ( ~n2400 & n2401 ) ;
  assign n2403 = ( ~n750 & n2193 ) | ( ~n750 & n2402 ) | ( n2193 & n2402 ) ;
  assign n2410 = n1129 ^ n767 ^ n462 ;
  assign n2404 = n2255 ^ n489 ^ n373 ;
  assign n2405 = ( ~n232 & n238 ) | ( ~n232 & n854 ) | ( n238 & n854 ) ;
  assign n2406 = n2405 ^ n1703 ^ x117 ;
  assign n2407 = n2406 ^ n587 ^ 1'b0 ;
  assign n2408 = ~n2404 & n2407 ;
  assign n2409 = ( n1108 & n1784 ) | ( n1108 & n2408 ) | ( n1784 & n2408 ) ;
  assign n2411 = n2410 ^ n2409 ^ n2153 ;
  assign n2412 = n2403 & ~n2411 ;
  assign n2416 = ~n153 & n408 ;
  assign n2417 = n2416 ^ n312 ^ 1'b0 ;
  assign n2418 = n2417 ^ n1696 ^ n641 ;
  assign n2413 = ~n1360 & n1519 ;
  assign n2414 = n2413 ^ n2097 ^ 1'b0 ;
  assign n2415 = n2149 & n2414 ;
  assign n2419 = n2418 ^ n2415 ^ 1'b0 ;
  assign n2420 = n544 & ~n2419 ;
  assign n2424 = n1796 ^ n1611 ^ x43 ;
  assign n2421 = ( x75 & ~n808 ) | ( x75 & n1011 ) | ( ~n808 & n1011 ) ;
  assign n2422 = x123 ^ x0 ^ 1'b0 ;
  assign n2423 = n2421 & n2422 ;
  assign n2425 = n2424 ^ n2423 ^ n362 ;
  assign n2426 = n421 ^ n184 ^ 1'b0 ;
  assign n2427 = n2426 ^ n1603 ^ 1'b0 ;
  assign n2428 = ( ~n434 & n479 ) | ( ~n434 & n2139 ) | ( n479 & n2139 ) ;
  assign n2429 = ( x35 & ~n716 ) | ( x35 & n1227 ) | ( ~n716 & n1227 ) ;
  assign n2430 = n710 ^ n689 ^ n433 ;
  assign n2431 = n2430 ^ n686 ^ 1'b0 ;
  assign n2432 = n2429 & n2431 ;
  assign n2433 = ~n2428 & n2432 ;
  assign n2435 = n448 | n1517 ;
  assign n2436 = n400 & ~n2435 ;
  assign n2434 = n593 ^ n476 ^ 1'b0 ;
  assign n2437 = n2436 ^ n2434 ^ x33 ;
  assign n2438 = n1436 ^ n1417 ^ 1'b0 ;
  assign n2439 = ~n708 & n2438 ;
  assign n2440 = n2439 ^ n1704 ^ x63 ;
  assign n2441 = n523 | n1871 ;
  assign n2442 = x43 & n592 ;
  assign n2443 = ~n1304 & n2442 ;
  assign n2444 = n2443 ^ n667 ^ 1'b0 ;
  assign n2445 = n2441 & n2444 ;
  assign n2446 = n2445 ^ n1692 ^ 1'b0 ;
  assign n2447 = ( n2437 & n2440 ) | ( n2437 & n2446 ) | ( n2440 & n2446 ) ;
  assign n2448 = n1393 ^ n186 ^ 1'b0 ;
  assign n2449 = ( x36 & n306 ) | ( x36 & n2448 ) | ( n306 & n2448 ) ;
  assign n2450 = ( x115 & n686 ) | ( x115 & n2449 ) | ( n686 & n2449 ) ;
  assign n2451 = n2450 ^ n344 ^ 1'b0 ;
  assign n2452 = ~n1416 & n2451 ;
  assign n2453 = n453 & n2452 ;
  assign n2454 = n2453 ^ n340 ^ 1'b0 ;
  assign n2455 = ~n686 & n2454 ;
  assign n2457 = n1703 ^ n1451 ^ n226 ;
  assign n2456 = n1278 & ~n1449 ;
  assign n2458 = n2457 ^ n2456 ^ 1'b0 ;
  assign n2459 = n1757 ^ n753 ^ 1'b0 ;
  assign n2460 = ( n317 & n1813 ) | ( n317 & n2459 ) | ( n1813 & n2459 ) ;
  assign n2468 = n1976 ^ n762 ^ 1'b0 ;
  assign n2469 = ~n277 & n2468 ;
  assign n2465 = ( n457 & n1486 ) | ( n457 & n2013 ) | ( n1486 & n2013 ) ;
  assign n2466 = n2465 ^ n622 ^ 1'b0 ;
  assign n2467 = n537 | n2466 ;
  assign n2464 = n839 ^ n571 ^ 1'b0 ;
  assign n2470 = n2469 ^ n2467 ^ n2464 ;
  assign n2461 = n2176 ^ n634 ^ 1'b0 ;
  assign n2462 = n693 | n2461 ;
  assign n2463 = n2439 | n2462 ;
  assign n2471 = n2470 ^ n2463 ^ n1337 ;
  assign n2472 = x96 ^ x18 ^ 1'b0 ;
  assign n2473 = ~n2246 & n2472 ;
  assign n2475 = ( n459 & ~n1106 ) | ( n459 & n1442 ) | ( ~n1106 & n1442 ) ;
  assign n2474 = n494 & n809 ;
  assign n2476 = n2475 ^ n2474 ^ n608 ;
  assign n2477 = x10 & x43 ;
  assign n2478 = ~n304 & n2477 ;
  assign n2479 = ( n300 & ~n355 ) | ( n300 & n2478 ) | ( ~n355 & n2478 ) ;
  assign n2480 = n1410 & ~n2479 ;
  assign n2481 = ~n1054 & n2480 ;
  assign n2482 = n2481 ^ n1345 ^ 1'b0 ;
  assign n2483 = n2482 ^ n1763 ^ 1'b0 ;
  assign n2484 = n2483 ^ n1597 ^ 1'b0 ;
  assign n2485 = n2035 ^ n1327 ^ n1322 ;
  assign n2486 = n2485 ^ n1570 ^ n346 ;
  assign n2487 = n214 & ~n1877 ;
  assign n2488 = n1047 & n2487 ;
  assign n2489 = ( n1184 & n1761 ) | ( n1184 & n2488 ) | ( n1761 & n2488 ) ;
  assign n2490 = ( n285 & ~n1024 ) | ( n285 & n1840 ) | ( ~n1024 & n1840 ) ;
  assign n2491 = n2490 ^ n2201 ^ n397 ;
  assign n2492 = n140 & n561 ;
  assign n2493 = n1417 & n2492 ;
  assign n2495 = ( x84 & n1069 ) | ( x84 & n1376 ) | ( n1069 & n1376 ) ;
  assign n2496 = ~n774 & n2495 ;
  assign n2497 = ~n885 & n2496 ;
  assign n2498 = n2497 ^ x95 ^ 1'b0 ;
  assign n2499 = n928 & ~n2498 ;
  assign n2500 = n2499 ^ n1699 ^ 1'b0 ;
  assign n2494 = ~n1238 & n2285 ;
  assign n2501 = n2500 ^ n2494 ^ 1'b0 ;
  assign n2502 = ( n1493 & n2493 ) | ( n1493 & n2501 ) | ( n2493 & n2501 ) ;
  assign n2508 = ( n1342 & ~n1836 ) | ( n1342 & n2033 ) | ( ~n1836 & n2033 ) ;
  assign n2503 = n1018 & n1225 ;
  assign n2504 = n1680 ^ n566 ^ 1'b0 ;
  assign n2505 = n2504 ^ n432 ^ 1'b0 ;
  assign n2506 = ~n2503 & n2505 ;
  assign n2507 = ~n1285 & n2506 ;
  assign n2509 = n2508 ^ n2507 ^ x5 ;
  assign n2510 = ( n205 & n641 ) | ( n205 & ~n2509 ) | ( n641 & ~n2509 ) ;
  assign n2513 = ( n385 & ~n448 ) | ( n385 & n718 ) | ( ~n448 & n718 ) ;
  assign n2514 = n2513 ^ n924 ^ n555 ;
  assign n2515 = n2514 ^ n1738 ^ n1170 ;
  assign n2511 = n315 ^ n239 ^ x68 ;
  assign n2512 = n2511 ^ n1678 ^ n1020 ;
  assign n2516 = n2515 ^ n2512 ^ n144 ;
  assign n2517 = ( n600 & n856 ) | ( n600 & n1046 ) | ( n856 & n1046 ) ;
  assign n2518 = n2517 ^ n1650 ^ 1'b0 ;
  assign n2519 = n2003 ^ n1551 ^ n1525 ;
  assign n2520 = x78 & ~n2519 ;
  assign n2522 = n1556 ^ n1143 ^ 1'b0 ;
  assign n2523 = n571 | n2522 ;
  assign n2521 = n1664 ^ n1001 ^ n331 ;
  assign n2524 = n2523 ^ n2521 ^ 1'b0 ;
  assign n2525 = n2520 & n2524 ;
  assign n2526 = n2194 & n2525 ;
  assign n2533 = n272 & ~n1259 ;
  assign n2534 = ~n1623 & n2533 ;
  assign n2527 = n2434 ^ n1131 ^ n734 ;
  assign n2528 = n2527 ^ n1917 ^ n1162 ;
  assign n2529 = n1159 & ~n2028 ;
  assign n2530 = n2529 ^ x107 ^ 1'b0 ;
  assign n2531 = n2530 ^ n1047 ^ 1'b0 ;
  assign n2532 = n2528 | n2531 ;
  assign n2535 = n2534 ^ n2532 ^ 1'b0 ;
  assign n2536 = n2449 ^ n1238 ^ n1146 ;
  assign n2537 = ( ~x41 & n1052 ) | ( ~x41 & n2536 ) | ( n1052 & n2536 ) ;
  assign n2538 = ( ~n1311 & n1503 ) | ( ~n1311 & n2537 ) | ( n1503 & n2537 ) ;
  assign n2539 = ( n729 & n798 ) | ( n729 & n865 ) | ( n798 & n865 ) ;
  assign n2540 = n580 & n1543 ;
  assign n2541 = n864 & n2540 ;
  assign n2542 = ( ~n708 & n2539 ) | ( ~n708 & n2541 ) | ( n2539 & n2541 ) ;
  assign n2543 = n2542 ^ n143 ^ 1'b0 ;
  assign n2544 = n826 ^ n212 ^ 1'b0 ;
  assign n2545 = n1953 | n2544 ;
  assign n2546 = n203 ^ x97 ^ 1'b0 ;
  assign n2547 = ( ~n2543 & n2545 ) | ( ~n2543 & n2546 ) | ( n2545 & n2546 ) ;
  assign n2548 = n1299 & n2547 ;
  assign n2549 = n2509 ^ n2246 ^ n1461 ;
  assign n2550 = n2287 ^ n2280 ^ 1'b0 ;
  assign n2551 = ( ~x114 & n143 ) | ( ~x114 & n875 ) | ( n143 & n875 ) ;
  assign n2552 = n2551 ^ n1549 ^ n186 ;
  assign n2553 = n557 & ~n2552 ;
  assign n2554 = n2553 ^ n1293 ^ 1'b0 ;
  assign n2555 = n2436 ^ n1522 ^ x12 ;
  assign n2556 = n510 ^ x36 ^ 1'b0 ;
  assign n2557 = n1231 & n2556 ;
  assign n2558 = ~n2098 & n2557 ;
  assign n2559 = ( n420 & ~n760 ) | ( n420 & n2558 ) | ( ~n760 & n2558 ) ;
  assign n2560 = n1713 ^ n1323 ^ 1'b0 ;
  assign n2561 = n2560 ^ n1084 ^ 1'b0 ;
  assign n2562 = ( n1042 & ~n2437 ) | ( n1042 & n2561 ) | ( ~n2437 & n2561 ) ;
  assign n2563 = ( ~n203 & n416 ) | ( ~n203 & n853 ) | ( n416 & n853 ) ;
  assign n2564 = n321 & n2563 ;
  assign n2565 = n2564 ^ n386 ^ 1'b0 ;
  assign n2566 = n2565 ^ n1288 ^ 1'b0 ;
  assign n2567 = x70 & ~n1725 ;
  assign n2568 = n2567 ^ n253 ^ 1'b0 ;
  assign n2569 = n1793 & n2568 ;
  assign n2572 = ( n186 & n1390 ) | ( n186 & ~n2041 ) | ( n1390 & ~n2041 ) ;
  assign n2570 = n1120 ^ n918 ^ n295 ;
  assign n2571 = n1958 & n2570 ;
  assign n2573 = n2572 ^ n2571 ^ 1'b0 ;
  assign n2574 = ( n1680 & n2569 ) | ( n1680 & n2573 ) | ( n2569 & n2573 ) ;
  assign n2575 = n2574 ^ n2465 ^ n204 ;
  assign n2576 = n2014 ^ n1800 ^ 1'b0 ;
  assign n2577 = n1769 & ~n2576 ;
  assign n2578 = n2577 ^ n2524 ^ 1'b0 ;
  assign n2579 = ( n1251 & n2475 ) | ( n1251 & ~n2578 ) | ( n2475 & ~n2578 ) ;
  assign n2580 = ( n976 & n2575 ) | ( n976 & n2579 ) | ( n2575 & n2579 ) ;
  assign n2581 = n1773 ^ n1560 ^ n571 ;
  assign n2582 = ( ~n1170 & n2450 ) | ( ~n1170 & n2581 ) | ( n2450 & n2581 ) ;
  assign n2583 = n594 & n1840 ;
  assign n2584 = n1796 ^ n650 ^ 1'b0 ;
  assign n2585 = n1019 & ~n2584 ;
  assign n2586 = n1544 ^ n1362 ^ n1038 ;
  assign n2587 = ( n844 & ~n2585 ) | ( n844 & n2586 ) | ( ~n2585 & n2586 ) ;
  assign n2588 = n1630 ^ n1624 ^ 1'b0 ;
  assign n2589 = n2588 ^ x87 ^ 1'b0 ;
  assign n2590 = ~n1005 & n2589 ;
  assign n2591 = n1365 | n1472 ;
  assign n2592 = n641 & ~n2591 ;
  assign n2593 = n1149 | n2089 ;
  assign n2594 = ( n465 & ~n1407 ) | ( n465 & n2593 ) | ( ~n1407 & n2593 ) ;
  assign n2600 = ( n667 & ~n1509 ) | ( n667 & n2197 ) | ( ~n1509 & n2197 ) ;
  assign n2595 = n1304 & n2373 ;
  assign n2596 = n2595 ^ n1176 ^ 1'b0 ;
  assign n2597 = n2596 ^ n1501 ^ n957 ;
  assign n2598 = n1990 | n2597 ;
  assign n2599 = n2390 & ~n2598 ;
  assign n2601 = n2600 ^ n2599 ^ 1'b0 ;
  assign n2602 = n2090 ^ n238 ^ 1'b0 ;
  assign n2603 = n2602 ^ n1708 ^ n547 ;
  assign n2604 = n1763 ^ n1127 ^ 1'b0 ;
  assign n2605 = n2603 | n2604 ;
  assign n2606 = n2188 & ~n2605 ;
  assign n2607 = ( n1242 & ~n1652 ) | ( n1242 & n1738 ) | ( ~n1652 & n1738 ) ;
  assign n2608 = ( ~n1194 & n2497 ) | ( ~n1194 & n2607 ) | ( n2497 & n2607 ) ;
  assign n2609 = ( n917 & n1673 ) | ( n917 & ~n2608 ) | ( n1673 & ~n2608 ) ;
  assign n2610 = n337 ^ n329 ^ 1'b0 ;
  assign n2611 = ( n140 & n596 ) | ( n140 & ~n2610 ) | ( n596 & ~n2610 ) ;
  assign n2612 = n1600 ^ n1430 ^ n1056 ;
  assign n2613 = n2612 ^ n2018 ^ n1529 ;
  assign n2614 = ( x96 & n616 ) | ( x96 & ~n1285 ) | ( n616 & ~n1285 ) ;
  assign n2615 = ( n2611 & n2613 ) | ( n2611 & ~n2614 ) | ( n2613 & ~n2614 ) ;
  assign n2616 = n2542 ^ n762 ^ n239 ;
  assign n2617 = n2616 ^ n386 ^ 1'b0 ;
  assign n2618 = ( n187 & ~n1354 ) | ( n187 & n1716 ) | ( ~n1354 & n1716 ) ;
  assign n2619 = n1194 & n1513 ;
  assign n2620 = ( n1192 & n1732 ) | ( n1192 & n2619 ) | ( n1732 & n2619 ) ;
  assign n2621 = ( n440 & ~n1055 ) | ( n440 & n2169 ) | ( ~n1055 & n2169 ) ;
  assign n2622 = ( ~n235 & n2620 ) | ( ~n235 & n2621 ) | ( n2620 & n2621 ) ;
  assign n2623 = n2195 ^ n510 ^ 1'b0 ;
  assign n2624 = ~n426 & n2623 ;
  assign n2625 = n1818 & ~n2624 ;
  assign n2626 = n1713 & ~n2625 ;
  assign n2627 = n2626 ^ n663 ^ 1'b0 ;
  assign n2628 = n567 ^ n397 ^ 1'b0 ;
  assign n2629 = n2627 & ~n2628 ;
  assign n2630 = n1537 ^ n245 ^ 1'b0 ;
  assign n2631 = ( ~n168 & n414 ) | ( ~n168 & n2630 ) | ( n414 & n2630 ) ;
  assign n2632 = n1116 | n2631 ;
  assign n2633 = ~n243 & n2227 ;
  assign n2634 = n1998 & n2633 ;
  assign n2635 = ( n418 & n1236 ) | ( n418 & ~n2634 ) | ( n1236 & ~n2634 ) ;
  assign n2636 = x98 & ~n1659 ;
  assign n2641 = n805 | n2600 ;
  assign n2642 = n2641 ^ n295 ^ 1'b0 ;
  assign n2643 = n632 & n1262 ;
  assign n2644 = n2642 | n2643 ;
  assign n2645 = n1673 ^ n1027 ^ 1'b0 ;
  assign n2646 = n2645 ^ n1695 ^ n799 ;
  assign n2647 = n149 & n2646 ;
  assign n2648 = n2644 & n2647 ;
  assign n2639 = ( n329 & n352 ) | ( n329 & n1295 ) | ( n352 & n1295 ) ;
  assign n2637 = n2169 ^ n1963 ^ 1'b0 ;
  assign n2638 = n2637 ^ n1867 ^ n475 ;
  assign n2640 = n2639 ^ n2638 ^ n1594 ;
  assign n2649 = n2648 ^ n2640 ^ 1'b0 ;
  assign n2650 = n2636 & n2649 ;
  assign n2651 = n1853 & n2072 ;
  assign n2652 = ~n1668 & n2651 ;
  assign n2653 = n1472 ^ n1126 ^ 1'b0 ;
  assign n2654 = n2653 ^ n1044 ^ 1'b0 ;
  assign n2655 = n1850 | n2654 ;
  assign n2656 = n2103 | n2655 ;
  assign n2657 = n2445 ^ n366 ^ 1'b0 ;
  assign n2658 = n525 & ~n2657 ;
  assign n2659 = n2228 ^ n1953 ^ 1'b0 ;
  assign n2660 = x67 & ~n2659 ;
  assign n2661 = n840 & n1829 ;
  assign n2662 = n2661 ^ n2130 ^ 1'b0 ;
  assign n2663 = n2662 ^ n2192 ^ n136 ;
  assign n2664 = ( ~n1522 & n2660 ) | ( ~n1522 & n2663 ) | ( n2660 & n2663 ) ;
  assign n2666 = n496 ^ n468 ^ 1'b0 ;
  assign n2667 = n1177 & n2666 ;
  assign n2665 = n1118 ^ n580 ^ 1'b0 ;
  assign n2668 = n2667 ^ n2665 ^ n2355 ;
  assign n2674 = ( n135 & ~n605 ) | ( n135 & n1191 ) | ( ~n605 & n1191 ) ;
  assign n2670 = n640 ^ n429 ^ x121 ;
  assign n2671 = n2670 ^ n1664 ^ 1'b0 ;
  assign n2669 = ~n933 & n1051 ;
  assign n2672 = n2671 ^ n2669 ^ 1'b0 ;
  assign n2673 = ( n280 & ~n2144 ) | ( n280 & n2672 ) | ( ~n2144 & n2672 ) ;
  assign n2675 = n2674 ^ n2673 ^ n252 ;
  assign n2676 = ( n400 & ~n514 ) | ( n400 & n2675 ) | ( ~n514 & n2675 ) ;
  assign n2678 = ~n861 & n1871 ;
  assign n2677 = n1164 ^ n1032 ^ n937 ;
  assign n2679 = n2678 ^ n2677 ^ n1546 ;
  assign n2680 = n2448 ^ n2047 ^ x90 ;
  assign n2681 = n2680 ^ n2179 ^ 1'b0 ;
  assign n2688 = n1652 ^ n1356 ^ n977 ;
  assign n2682 = ~n240 & n1799 ;
  assign n2683 = n1220 & ~n2523 ;
  assign n2684 = ~n1804 & n2683 ;
  assign n2685 = ~n2682 & n2684 ;
  assign n2686 = ( n2234 & n2669 ) | ( n2234 & n2685 ) | ( n2669 & n2685 ) ;
  assign n2687 = n1225 | n2686 ;
  assign n2689 = n2688 ^ n2687 ^ 1'b0 ;
  assign n2690 = n2551 ^ n2437 ^ n1574 ;
  assign n2695 = ( n1244 & ~n1633 ) | ( n1244 & n1682 ) | ( ~n1633 & n1682 ) ;
  assign n2691 = n1582 ^ n1318 ^ 1'b0 ;
  assign n2692 = ~n780 & n2691 ;
  assign n2693 = n2692 ^ n598 ^ n348 ;
  assign n2694 = n2693 ^ n2513 ^ n2184 ;
  assign n2696 = n2695 ^ n2694 ^ n894 ;
  assign n2704 = n367 & n1126 ;
  assign n2705 = n2704 ^ n2038 ^ 1'b0 ;
  assign n2706 = n2705 ^ n2414 ^ n1101 ;
  assign n2700 = n1754 ^ n1668 ^ n659 ;
  assign n2701 = n2613 ^ n1557 ^ 1'b0 ;
  assign n2702 = ( ~n1216 & n2700 ) | ( ~n1216 & n2701 ) | ( n2700 & n2701 ) ;
  assign n2697 = n577 ^ n289 ^ x1 ;
  assign n2698 = ( x72 & n1205 ) | ( x72 & ~n2697 ) | ( n1205 & ~n2697 ) ;
  assign n2699 = ~n268 & n2698 ;
  assign n2703 = n2702 ^ n2699 ^ 1'b0 ;
  assign n2707 = n2706 ^ n2703 ^ n2079 ;
  assign n2708 = ( n175 & n346 ) | ( n175 & n1597 ) | ( n346 & n1597 ) ;
  assign n2709 = n587 & n2708 ;
  assign n2710 = n2709 ^ n2024 ^ 1'b0 ;
  assign n2711 = ~n265 & n390 ;
  assign n2712 = n2711 ^ n270 ^ 1'b0 ;
  assign n2713 = ( n844 & ~n1171 ) | ( n844 & n2712 ) | ( ~n1171 & n2712 ) ;
  assign n2714 = ( n2218 & n2394 ) | ( n2218 & n2713 ) | ( n2394 & n2713 ) ;
  assign n2715 = n2072 & ~n2181 ;
  assign n2716 = n2715 ^ n2163 ^ 1'b0 ;
  assign n2717 = n1707 ^ n1559 ^ n977 ;
  assign n2718 = n172 & ~n1040 ;
  assign n2719 = n2718 ^ x5 ^ 1'b0 ;
  assign n2720 = n1180 ^ n927 ^ n916 ;
  assign n2721 = ~n1967 & n2720 ;
  assign n2722 = ( n741 & n2719 ) | ( n741 & ~n2721 ) | ( n2719 & ~n2721 ) ;
  assign n2723 = n2483 ^ n2459 ^ 1'b0 ;
  assign n2724 = n2722 & n2723 ;
  assign n2725 = ( n2092 & n2717 ) | ( n2092 & n2724 ) | ( n2717 & n2724 ) ;
  assign n2727 = ( n397 & n661 ) | ( n397 & ~n1295 ) | ( n661 & ~n1295 ) ;
  assign n2726 = n480 & n950 ;
  assign n2728 = n2727 ^ n2726 ^ 1'b0 ;
  assign n2729 = ( x41 & n1360 ) | ( x41 & n2539 ) | ( n1360 & n2539 ) ;
  assign n2730 = n2728 & n2729 ;
  assign n2731 = n2730 ^ n2253 ^ 1'b0 ;
  assign n2732 = ~n2609 & n2731 ;
  assign n2739 = n2228 ^ n942 ^ n691 ;
  assign n2734 = n2080 ^ n1204 ^ 1'b0 ;
  assign n2735 = n394 | n2734 ;
  assign n2736 = n1922 | n2735 ;
  assign n2737 = n2736 ^ n2139 ^ 1'b0 ;
  assign n2738 = n2563 & ~n2737 ;
  assign n2733 = ( ~n1597 & n1868 ) | ( ~n1597 & n2339 ) | ( n1868 & n2339 ) ;
  assign n2740 = n2739 ^ n2738 ^ n2733 ;
  assign n2741 = ( ~n133 & n339 ) | ( ~n133 & n2740 ) | ( n339 & n2740 ) ;
  assign n2742 = ( n724 & ~n1219 ) | ( n724 & n1552 ) | ( ~n1219 & n1552 ) ;
  assign n2743 = n2742 ^ n1492 ^ 1'b0 ;
  assign n2744 = ( n1101 & n2643 ) | ( n1101 & ~n2743 ) | ( n2643 & ~n2743 ) ;
  assign n2745 = ( n544 & n581 ) | ( n544 & n1699 ) | ( n581 & n1699 ) ;
  assign n2746 = n184 | n1428 ;
  assign n2747 = n2746 ^ n167 ^ 1'b0 ;
  assign n2748 = x43 & ~n1052 ;
  assign n2749 = n708 & n2748 ;
  assign n2750 = n414 | n2749 ;
  assign n2751 = ( n2138 & n2747 ) | ( n2138 & n2750 ) | ( n2747 & n2750 ) ;
  assign n2752 = n270 & ~n2751 ;
  assign n2753 = n1789 ^ x53 ^ 1'b0 ;
  assign n2754 = n1611 ^ n1482 ^ n891 ;
  assign n2755 = n2754 ^ n1369 ^ 1'b0 ;
  assign n2756 = ~n1457 & n2755 ;
  assign n2757 = ~n2753 & n2756 ;
  assign n2766 = n1978 ^ n992 ^ 1'b0 ;
  assign n2767 = n670 | n2766 ;
  assign n2759 = n551 & ~n822 ;
  assign n2760 = n1575 ^ x91 ^ 1'b0 ;
  assign n2761 = n1550 ^ n813 ^ x62 ;
  assign n2762 = n2761 ^ n1004 ^ n979 ;
  assign n2763 = ( n924 & ~n1772 ) | ( n924 & n2762 ) | ( ~n1772 & n2762 ) ;
  assign n2764 = n2760 | n2763 ;
  assign n2765 = n2759 & ~n2764 ;
  assign n2758 = n1616 ^ x103 ^ 1'b0 ;
  assign n2768 = n2767 ^ n2765 ^ n2758 ;
  assign n2769 = ( ~x26 & n335 ) | ( ~x26 & n433 ) | ( n335 & n433 ) ;
  assign n2770 = ( n223 & ~n1527 ) | ( n223 & n2769 ) | ( ~n1527 & n2769 ) ;
  assign n2771 = ( ~n334 & n799 ) | ( ~n334 & n2770 ) | ( n799 & n2770 ) ;
  assign n2772 = n2771 ^ n1480 ^ n1369 ;
  assign n2773 = n1164 ^ n1002 ^ 1'b0 ;
  assign n2780 = n1360 ^ n577 ^ n541 ;
  assign n2779 = ( ~x40 & x86 ) | ( ~x40 & n1058 ) | ( x86 & n1058 ) ;
  assign n2778 = n1665 ^ n1493 ^ n520 ;
  assign n2781 = n2780 ^ n2779 ^ n2778 ;
  assign n2783 = n2642 ^ n2047 ^ n317 ;
  assign n2782 = ~n211 & n724 ;
  assign n2784 = n2783 ^ n2782 ^ 1'b0 ;
  assign n2785 = n2784 ^ n1240 ^ n878 ;
  assign n2786 = n2785 ^ n1318 ^ 1'b0 ;
  assign n2787 = n2781 & n2786 ;
  assign n2774 = n1124 ^ n1099 ^ n132 ;
  assign n2775 = ( n366 & ~n2218 ) | ( n366 & n2774 ) | ( ~n2218 & n2774 ) ;
  assign n2776 = ~n1317 & n1720 ;
  assign n2777 = ( ~n2005 & n2775 ) | ( ~n2005 & n2776 ) | ( n2775 & n2776 ) ;
  assign n2788 = n2787 ^ n2777 ^ x120 ;
  assign n2789 = ( ~n2359 & n2773 ) | ( ~n2359 & n2788 ) | ( n2773 & n2788 ) ;
  assign n2790 = n2357 ^ n1913 ^ n1021 ;
  assign n2791 = n2790 ^ n1312 ^ n350 ;
  assign n2792 = n2508 ^ n2157 ^ n2069 ;
  assign n2793 = n649 & ~n2792 ;
  assign n2794 = ~n544 & n2793 ;
  assign n2795 = n870 & n1921 ;
  assign n2796 = n2795 ^ n328 ^ 1'b0 ;
  assign n2797 = n2794 | n2796 ;
  assign n2798 = n2791 | n2797 ;
  assign n2799 = n1643 ^ n1037 ^ n773 ;
  assign n2800 = n2799 ^ n697 ^ 1'b0 ;
  assign n2801 = ( x109 & ~n1624 ) | ( x109 & n2800 ) | ( ~n1624 & n2800 ) ;
  assign n2802 = n2801 ^ n1011 ^ 1'b0 ;
  assign n2803 = n633 ^ n291 ^ n255 ;
  assign n2804 = n2784 ^ n1838 ^ n1168 ;
  assign n2810 = n1110 ^ n647 ^ x18 ;
  assign n2811 = x24 & ~n2810 ;
  assign n2805 = n2498 ^ n1257 ^ 1'b0 ;
  assign n2806 = ~n334 & n2805 ;
  assign n2807 = ~n1145 & n2806 ;
  assign n2808 = n2807 ^ n2178 ^ 1'b0 ;
  assign n2809 = x91 & n2808 ;
  assign n2812 = n2811 ^ n2809 ^ n2400 ;
  assign n2813 = ( n568 & ~n844 ) | ( n568 & n853 ) | ( ~n844 & n853 ) ;
  assign n2814 = ( ~n542 & n665 ) | ( ~n542 & n1498 ) | ( n665 & n1498 ) ;
  assign n2815 = n2495 ^ n954 ^ 1'b0 ;
  assign n2816 = n2814 | n2815 ;
  assign n2817 = n1140 ^ x5 ^ 1'b0 ;
  assign n2818 = n871 | n2817 ;
  assign n2819 = n2816 & n2818 ;
  assign n2820 = ~n742 & n2819 ;
  assign n2821 = n2120 ^ n377 ^ n275 ;
  assign n2822 = ( x41 & n908 ) | ( x41 & n2391 ) | ( n908 & n2391 ) ;
  assign n2823 = n2165 ^ n639 ^ n594 ;
  assign n2824 = ~n2436 & n2823 ;
  assign n2825 = n2824 ^ n1222 ^ 1'b0 ;
  assign n2826 = n2825 ^ n2298 ^ n1047 ;
  assign n2828 = n2022 ^ n1547 ^ n1342 ;
  assign n2827 = n455 & n2129 ;
  assign n2829 = n2828 ^ n2827 ^ 1'b0 ;
  assign n2830 = n2826 | n2829 ;
  assign n2832 = n1480 ^ n1379 ^ 1'b0 ;
  assign n2833 = n2832 ^ n1114 ^ 1'b0 ;
  assign n2834 = n1107 & ~n2833 ;
  assign n2831 = x98 & ~n942 ;
  assign n2835 = n2834 ^ n2831 ^ 1'b0 ;
  assign n2836 = n1680 & n1809 ;
  assign n2837 = n825 & n2836 ;
  assign n2838 = ( n372 & n1568 ) | ( n372 & ~n1908 ) | ( n1568 & ~n1908 ) ;
  assign n2839 = ~n2837 & n2838 ;
  assign n2840 = ( n380 & n760 ) | ( n380 & n2069 ) | ( n760 & n2069 ) ;
  assign n2841 = n636 & n2840 ;
  assign n2842 = n2841 ^ n1705 ^ 1'b0 ;
  assign n2843 = n1798 ^ n1019 ^ 1'b0 ;
  assign n2844 = n273 & ~n2843 ;
  assign n2845 = n2844 ^ n1889 ^ 1'b0 ;
  assign n2846 = n2842 & n2845 ;
  assign n2847 = n2210 ^ n270 ^ 1'b0 ;
  assign n2848 = n1562 | n2847 ;
  assign n2851 = ( n335 & n975 ) | ( n335 & n2449 ) | ( n975 & n2449 ) ;
  assign n2852 = n2851 ^ n1189 ^ n1104 ;
  assign n2849 = ( ~n742 & n1443 ) | ( ~n742 & n2216 ) | ( n1443 & n2216 ) ;
  assign n2850 = n2849 ^ n833 ^ n464 ;
  assign n2853 = n2852 ^ n2850 ^ n634 ;
  assign n2854 = ( n684 & ~n2529 ) | ( n684 & n2627 ) | ( ~n2529 & n2627 ) ;
  assign n2859 = n2045 ^ n840 ^ n165 ;
  assign n2860 = n2859 ^ n342 ^ n256 ;
  assign n2858 = ( n464 & ~n1058 ) | ( n464 & n1983 ) | ( ~n1058 & n1983 ) ;
  assign n2855 = n2124 ^ n418 ^ 1'b0 ;
  assign n2856 = n2844 & n2855 ;
  assign n2857 = ( n367 & ~n2565 ) | ( n367 & n2856 ) | ( ~n2565 & n2856 ) ;
  assign n2861 = n2860 ^ n2858 ^ n2857 ;
  assign n2863 = n2859 ^ n1330 ^ n637 ;
  assign n2864 = ~n1523 & n2262 ;
  assign n2865 = n2863 & n2864 ;
  assign n2862 = ~n411 & n545 ;
  assign n2866 = n2865 ^ n2862 ^ n428 ;
  assign n2867 = ~n1384 & n2164 ;
  assign n2868 = ~n1466 & n2867 ;
  assign n2869 = n2219 ^ n1906 ^ n1721 ;
  assign n2870 = n1702 ^ n513 ^ 1'b0 ;
  assign n2871 = n591 & n679 ;
  assign n2872 = n2870 & n2871 ;
  assign n2873 = n1887 & ~n2872 ;
  assign n2874 = x4 & n277 ;
  assign n2875 = n2874 ^ n282 ^ 1'b0 ;
  assign n2876 = n2873 | n2875 ;
  assign n2877 = n1670 ^ n1645 ^ n1443 ;
  assign n2882 = ( x49 & n989 ) | ( x49 & ~n1031 ) | ( n989 & ~n1031 ) ;
  assign n2883 = n2882 ^ x93 ^ 1'b0 ;
  assign n2884 = ~n409 & n2883 ;
  assign n2885 = n2884 ^ n1981 ^ n897 ;
  assign n2878 = n571 & n1298 ;
  assign n2879 = ~n567 & n1186 ;
  assign n2880 = n2879 ^ n1524 ^ 1'b0 ;
  assign n2881 = ~n2878 & n2880 ;
  assign n2886 = n2885 ^ n2881 ^ 1'b0 ;
  assign n2894 = ( x70 & n507 ) | ( x70 & n989 ) | ( n507 & n989 ) ;
  assign n2895 = ( x83 & n1384 ) | ( x83 & ~n2894 ) | ( n1384 & ~n2894 ) ;
  assign n2896 = n2895 ^ n1677 ^ 1'b0 ;
  assign n2897 = ( n1390 & n2509 ) | ( n1390 & n2896 ) | ( n2509 & n2896 ) ;
  assign n2890 = ~n353 & n525 ;
  assign n2891 = n2890 ^ n240 ^ 1'b0 ;
  assign n2892 = n2891 ^ n2256 ^ n1450 ;
  assign n2893 = n2892 ^ n2372 ^ n2247 ;
  assign n2887 = n1543 ^ n1011 ^ 1'b0 ;
  assign n2888 = ~n514 & n2887 ;
  assign n2889 = n2888 ^ n2872 ^ n1624 ;
  assign n2898 = n2897 ^ n2893 ^ n2889 ;
  assign n2899 = n1425 & n1694 ;
  assign n2900 = n2899 ^ n2421 ^ n1430 ;
  assign n2901 = ( n671 & ~n2488 ) | ( n671 & n2900 ) | ( ~n2488 & n2900 ) ;
  assign n2907 = n1551 ^ n810 ^ n608 ;
  assign n2908 = x52 & n1914 ;
  assign n2909 = ( n2767 & ~n2907 ) | ( n2767 & n2908 ) | ( ~n2907 & n2908 ) ;
  assign n2902 = ( x46 & ~n1509 ) | ( x46 & n1676 ) | ( ~n1509 & n1676 ) ;
  assign n2903 = ( n1780 & ~n2630 ) | ( n1780 & n2902 ) | ( ~n2630 & n2902 ) ;
  assign n2904 = ( ~x75 & n464 ) | ( ~x75 & n500 ) | ( n464 & n500 ) ;
  assign n2905 = n2904 ^ n2620 ^ 1'b0 ;
  assign n2906 = n2903 | n2905 ;
  assign n2910 = n2909 ^ n2906 ^ n1989 ;
  assign n2911 = n810 & ~n1990 ;
  assign n2912 = n2911 ^ n2771 ^ 1'b0 ;
  assign n2913 = n159 ^ x110 ^ 1'b0 ;
  assign n2914 = n1510 & ~n2913 ;
  assign n2915 = n2914 ^ n853 ^ n775 ;
  assign n2916 = n2915 ^ n2000 ^ 1'b0 ;
  assign n2917 = ( n840 & n2912 ) | ( n840 & ~n2916 ) | ( n2912 & ~n2916 ) ;
  assign n2918 = n2216 ^ n1032 ^ n158 ;
  assign n2919 = ( ~n1176 & n1413 ) | ( ~n1176 & n2918 ) | ( n1413 & n2918 ) ;
  assign n2920 = n2919 ^ n974 ^ 1'b0 ;
  assign n2921 = n900 & n2920 ;
  assign n2922 = n2921 ^ n1058 ^ n758 ;
  assign n2923 = ( n2357 & n2491 ) | ( n2357 & n2922 ) | ( n2491 & n2922 ) ;
  assign n2924 = x37 & n918 ;
  assign n2925 = n2924 ^ x89 ^ 1'b0 ;
  assign n2926 = n2925 ^ n1159 ^ x65 ;
  assign n2927 = ( n2779 & ~n2852 ) | ( n2779 & n2926 ) | ( ~n2852 & n2926 ) ;
  assign n2935 = n1020 ^ n782 ^ 1'b0 ;
  assign n2933 = n1640 ^ n1556 ^ n976 ;
  assign n2928 = ( n211 & n1208 ) | ( n211 & n1325 ) | ( n1208 & n1325 ) ;
  assign n2929 = n145 ^ x123 ^ 1'b0 ;
  assign n2930 = ~n2928 & n2929 ;
  assign n2931 = n2930 ^ n1765 ^ n524 ;
  assign n2932 = ( n771 & n1266 ) | ( n771 & n2931 ) | ( n1266 & n2931 ) ;
  assign n2934 = n2933 ^ n2932 ^ n1753 ;
  assign n2936 = n2935 ^ n2934 ^ n1773 ;
  assign n2937 = ( n337 & n2733 ) | ( n337 & n2936 ) | ( n2733 & n2936 ) ;
  assign n2938 = n136 | n2031 ;
  assign n2939 = n1288 & ~n2938 ;
  assign n2940 = n1519 | n2939 ;
  assign n2941 = x104 & ~n1290 ;
  assign n2942 = n1331 ^ n616 ^ 1'b0 ;
  assign n2943 = n305 & ~n2942 ;
  assign n2944 = n1013 ^ n638 ^ n352 ;
  assign n2945 = n1295 & ~n2112 ;
  assign n2946 = ~n733 & n2945 ;
  assign n2947 = n1616 & ~n2946 ;
  assign n2948 = ~n2944 & n2947 ;
  assign n2949 = n509 | n2948 ;
  assign n2950 = n2312 ^ n634 ^ n131 ;
  assign n2951 = ( ~n305 & n2949 ) | ( ~n305 & n2950 ) | ( n2949 & n2950 ) ;
  assign n2952 = n2951 ^ n1972 ^ 1'b0 ;
  assign n2953 = ( ~n2941 & n2943 ) | ( ~n2941 & n2952 ) | ( n2943 & n2952 ) ;
  assign n2954 = ~n812 & n1617 ;
  assign n2955 = n2128 ^ n1785 ^ n989 ;
  assign n2956 = n2955 ^ n1561 ^ 1'b0 ;
  assign n2957 = n2139 | n2956 ;
  assign n2961 = n2329 ^ n1836 ^ n129 ;
  assign n2958 = n2907 ^ n644 ^ n471 ;
  assign n2959 = n2958 ^ n1533 ^ n963 ;
  assign n2960 = n2959 ^ n697 ^ n645 ;
  assign n2962 = n2961 ^ n2960 ^ 1'b0 ;
  assign n2963 = n420 ^ x85 ^ 1'b0 ;
  assign n2964 = n2963 ^ n2835 ^ n1314 ;
  assign n2965 = ( x57 & ~x106 ) | ( x57 & n187 ) | ( ~x106 & n187 ) ;
  assign n2966 = ( ~n1148 & n1762 ) | ( ~n1148 & n2039 ) | ( n1762 & n2039 ) ;
  assign n2967 = n1565 ^ n459 ^ 1'b0 ;
  assign n2968 = n725 & ~n2967 ;
  assign n2969 = n2968 ^ n2108 ^ n347 ;
  assign n2970 = n2969 ^ n2519 ^ n1617 ;
  assign n2971 = ( ~n897 & n2966 ) | ( ~n897 & n2970 ) | ( n2966 & n2970 ) ;
  assign n2972 = n1566 ^ n1493 ^ n814 ;
  assign n2973 = n196 ^ x84 ^ x6 ;
  assign n2974 = n2973 ^ n2780 ^ n2024 ;
  assign n2975 = x27 & n1920 ;
  assign n2976 = ( ~n2972 & n2974 ) | ( ~n2972 & n2975 ) | ( n2974 & n2975 ) ;
  assign n2977 = n1643 ^ n1228 ^ x110 ;
  assign n2978 = ( n609 & ~n2258 ) | ( n609 & n2977 ) | ( ~n2258 & n2977 ) ;
  assign n2979 = n2898 | n2978 ;
  assign n2980 = n2979 ^ x118 ^ 1'b0 ;
  assign n2981 = ( ~x98 & n407 ) | ( ~x98 & n1808 ) | ( n407 & n1808 ) ;
  assign n2982 = n1688 ^ x62 ^ 1'b0 ;
  assign n2983 = n2982 ^ n1241 ^ n1126 ;
  assign n2984 = ( ~n643 & n1226 ) | ( ~n643 & n2406 ) | ( n1226 & n2406 ) ;
  assign n2985 = n533 | n2984 ;
  assign n2986 = n593 | n2985 ;
  assign n2987 = n2983 & n2986 ;
  assign n2988 = ~n1459 & n2987 ;
  assign n2989 = ( x0 & ~n405 ) | ( x0 & n1333 ) | ( ~n405 & n1333 ) ;
  assign n2990 = ( n2981 & ~n2988 ) | ( n2981 & n2989 ) | ( ~n2988 & n2989 ) ;
  assign n2991 = ~n2280 & n2725 ;
  assign n2992 = n2991 ^ n662 ^ 1'b0 ;
  assign n2993 = x11 & ~n2448 ;
  assign n2994 = n2993 ^ n1504 ^ 1'b0 ;
  assign n2995 = n2111 ^ n1705 ^ 1'b0 ;
  assign n2996 = n2995 ^ n1480 ^ 1'b0 ;
  assign n2997 = n928 ^ n429 ^ n370 ;
  assign n2998 = n1159 ^ n1029 ^ n235 ;
  assign n2999 = ( n2168 & ~n2380 ) | ( n2168 & n2998 ) | ( ~n2380 & n2998 ) ;
  assign n3000 = n2999 ^ n280 ^ 1'b0 ;
  assign n3001 = ( ~n306 & n2103 ) | ( ~n306 & n3000 ) | ( n2103 & n3000 ) ;
  assign n3002 = ( n2996 & n2997 ) | ( n2996 & n3001 ) | ( n2997 & n3001 ) ;
  assign n3003 = n2994 & ~n3002 ;
  assign n3004 = ~n1276 & n2285 ;
  assign n3005 = n3004 ^ n2305 ^ 1'b0 ;
  assign n3007 = ~n409 & n2324 ;
  assign n3006 = n2774 ^ n1703 ^ n178 ;
  assign n3008 = n3007 ^ n3006 ^ n1096 ;
  assign n3009 = n2712 ^ n655 ^ 1'b0 ;
  assign n3010 = n1055 & n1989 ;
  assign n3011 = n3010 ^ n1524 ^ 1'b0 ;
  assign n3012 = ( n269 & n3009 ) | ( n269 & ~n3011 ) | ( n3009 & ~n3011 ) ;
  assign n3013 = n278 & ~n2086 ;
  assign n3014 = n443 & n3013 ;
  assign n3015 = n1531 & ~n2205 ;
  assign n3016 = n3014 & n3015 ;
  assign n3017 = ~n233 & n814 ;
  assign n3018 = n278 & n1910 ;
  assign n3019 = n3018 ^ n2643 ^ 1'b0 ;
  assign n3020 = n3019 ^ n1671 ^ 1'b0 ;
  assign n3021 = n2768 | n3020 ;
  assign n3022 = n600 ^ n445 ^ n159 ;
  assign n3023 = n3022 ^ n881 ^ n287 ;
  assign n3024 = n2075 ^ n1595 ^ x72 ;
  assign n3026 = n379 ^ x119 ^ x28 ;
  assign n3025 = x63 ^ x21 ^ 1'b0 ;
  assign n3027 = n3026 ^ n3025 ^ n1416 ;
  assign n3028 = n3027 ^ n1176 ^ 1'b0 ;
  assign n3029 = x28 & n3028 ;
  assign n3030 = n3024 & n3029 ;
  assign n3031 = n3030 ^ n723 ^ 1'b0 ;
  assign n3032 = ( n523 & ~n3023 ) | ( n523 & n3031 ) | ( ~n3023 & n3031 ) ;
  assign n3033 = n482 & ~n3003 ;
  assign n3034 = ~n889 & n1594 ;
  assign n3035 = n3034 ^ x117 ^ 1'b0 ;
  assign n3036 = n1913 ^ n1454 ^ 1'b0 ;
  assign n3037 = ( n971 & n1699 ) | ( n971 & n3036 ) | ( n1699 & n3036 ) ;
  assign n3038 = n2762 ^ n691 ^ x121 ;
  assign n3039 = n3038 ^ n2998 ^ n2771 ;
  assign n3040 = n3039 ^ n1942 ^ n476 ;
  assign n3041 = n3040 ^ n2251 ^ 1'b0 ;
  assign n3042 = n235 & n787 ;
  assign n3043 = n3042 ^ n870 ^ 1'b0 ;
  assign n3044 = n920 ^ n694 ^ 1'b0 ;
  assign n3045 = n2620 & ~n3044 ;
  assign n3046 = ( n146 & n738 ) | ( n146 & ~n808 ) | ( n738 & ~n808 ) ;
  assign n3047 = n3046 ^ n697 ^ x37 ;
  assign n3048 = n2169 ^ n334 ^ 1'b0 ;
  assign n3049 = n3047 | n3048 ;
  assign n3050 = ( n3043 & n3045 ) | ( n3043 & ~n3049 ) | ( n3045 & ~n3049 ) ;
  assign n3053 = n2469 ^ n1221 ^ 1'b0 ;
  assign n3051 = n796 ^ n164 ^ 1'b0 ;
  assign n3052 = x36 & ~n3051 ;
  assign n3054 = n3053 ^ n3052 ^ 1'b0 ;
  assign n3056 = n355 & ~n2247 ;
  assign n3055 = n2607 ^ n1766 ^ n1003 ;
  assign n3057 = n3056 ^ n3055 ^ n1003 ;
  assign n3058 = n3038 ^ n2420 ^ n1659 ;
  assign n3059 = n934 ^ n211 ^ n205 ;
  assign n3060 = ( ~n533 & n1314 ) | ( ~n533 & n3059 ) | ( n1314 & n3059 ) ;
  assign n3061 = n1289 & n1829 ;
  assign n3062 = n3061 ^ n2840 ^ 1'b0 ;
  assign n3063 = ( n1029 & ~n3060 ) | ( n1029 & n3062 ) | ( ~n3060 & n3062 ) ;
  assign n3065 = ( n204 & n326 ) | ( n204 & n448 ) | ( n326 & n448 ) ;
  assign n3064 = n2479 ^ n300 ^ 1'b0 ;
  assign n3066 = n3065 ^ n3064 ^ 1'b0 ;
  assign n3067 = n3066 ^ n2552 ^ x70 ;
  assign n3068 = x87 ^ x12 ^ 1'b0 ;
  assign n3069 = n1510 ^ n600 ^ x76 ;
  assign n3070 = n3069 ^ n1157 ^ n487 ;
  assign n3071 = ~n284 & n2646 ;
  assign n3072 = ~n1271 & n3071 ;
  assign n3073 = ( n334 & n1864 ) | ( n334 & ~n2859 ) | ( n1864 & ~n2859 ) ;
  assign n3074 = n3073 ^ n2739 ^ n1317 ;
  assign n3075 = ( n2899 & ~n3072 ) | ( n2899 & n3074 ) | ( ~n3072 & n3074 ) ;
  assign n3076 = ( n3068 & n3070 ) | ( n3068 & ~n3075 ) | ( n3070 & ~n3075 ) ;
  assign n3081 = n1153 ^ n288 ^ x107 ;
  assign n3082 = n3081 ^ n1624 ^ 1'b0 ;
  assign n3077 = n979 ^ n238 ^ 1'b0 ;
  assign n3078 = ( x19 & n1745 ) | ( x19 & n3077 ) | ( n1745 & n3077 ) ;
  assign n3079 = ~n2618 & n3078 ;
  assign n3080 = n3079 ^ n2621 ^ n2582 ;
  assign n3083 = n3082 ^ n3080 ^ n1016 ;
  assign n3084 = n2249 ^ n2065 ^ n1309 ;
  assign n3085 = n375 & n1267 ;
  assign n3086 = n3084 | n3085 ;
  assign n3087 = n3086 ^ n1579 ^ 1'b0 ;
  assign n3088 = n897 | n1858 ;
  assign n3089 = n3088 ^ n1470 ^ 1'b0 ;
  assign n3090 = n169 & n2097 ;
  assign n3091 = n1864 ^ n526 ^ 1'b0 ;
  assign n3092 = n2222 & n3091 ;
  assign n3093 = n2257 ^ n489 ^ 1'b0 ;
  assign n3094 = n2273 & n3093 ;
  assign n3095 = ( n2919 & n3092 ) | ( n2919 & ~n3094 ) | ( n3092 & ~n3094 ) ;
  assign n3096 = x83 & ~n616 ;
  assign n3097 = n1422 ^ n508 ^ x8 ;
  assign n3098 = ( n365 & n825 ) | ( n365 & ~n3097 ) | ( n825 & ~n3097 ) ;
  assign n3099 = n3098 ^ n2014 ^ n1997 ;
  assign n3100 = ( n1431 & ~n3096 ) | ( n1431 & n3099 ) | ( ~n3096 & n3099 ) ;
  assign n3101 = n3008 ^ n1019 ^ 1'b0 ;
  assign n3102 = ( n236 & n350 ) | ( n236 & ~n1076 ) | ( n350 & ~n1076 ) ;
  assign n3103 = ( n399 & n1239 ) | ( n399 & ~n3102 ) | ( n1239 & ~n3102 ) ;
  assign n3104 = x46 | n2172 ;
  assign n3105 = n3103 & n3104 ;
  assign n3106 = n3105 ^ n3017 ^ 1'b0 ;
  assign n3108 = n974 ^ n211 ^ x63 ;
  assign n3109 = n967 & ~n3108 ;
  assign n3110 = n3109 ^ n443 ^ 1'b0 ;
  assign n3107 = ~n2105 & n3074 ;
  assign n3111 = n3110 ^ n3107 ^ 1'b0 ;
  assign n3112 = n966 ^ n924 ^ 1'b0 ;
  assign n3113 = n544 & n3112 ;
  assign n3114 = x39 & ~n160 ;
  assign n3115 = ~n3113 & n3114 ;
  assign n3116 = n2111 & ~n3115 ;
  assign n3117 = ~n2214 & n3116 ;
  assign n3118 = ( n2024 & ~n2392 ) | ( n2024 & n3117 ) | ( ~n2392 & n3117 ) ;
  assign n3120 = n1898 ^ n1287 ^ x58 ;
  assign n3119 = n444 | n774 ;
  assign n3121 = n3120 ^ n3119 ^ n158 ;
  assign n3122 = ( n212 & n593 ) | ( n212 & ~n851 ) | ( n593 & ~n851 ) ;
  assign n3123 = n1748 ^ n1676 ^ n1284 ;
  assign n3124 = n334 ^ n314 ^ 1'b0 ;
  assign n3125 = x100 & ~n3124 ;
  assign n3126 = ( n201 & ~n293 ) | ( n201 & n3125 ) | ( ~n293 & n3125 ) ;
  assign n3127 = ( n1121 & ~n3123 ) | ( n1121 & n3126 ) | ( ~n3123 & n3126 ) ;
  assign n3128 = n2667 ^ n373 ^ 1'b0 ;
  assign n3129 = n3127 & n3128 ;
  assign n3131 = ( n443 & n459 ) | ( n443 & n2563 ) | ( n459 & n2563 ) ;
  assign n3132 = n3131 ^ n2671 ^ 1'b0 ;
  assign n3130 = n2951 ^ n1833 ^ n952 ;
  assign n3133 = n3132 ^ n3130 ^ n2321 ;
  assign n3134 = ( n3122 & n3129 ) | ( n3122 & ~n3133 ) | ( n3129 & ~n3133 ) ;
  assign n3135 = n3023 ^ n2313 ^ n1840 ;
  assign n3136 = n1052 | n1612 ;
  assign n3137 = x20 & ~n1994 ;
  assign n3138 = n3137 ^ n366 ^ 1'b0 ;
  assign n3139 = ( n529 & ~n1769 ) | ( n529 & n3138 ) | ( ~n1769 & n3138 ) ;
  assign n3140 = n3136 & n3139 ;
  assign n3141 = ( n477 & n967 ) | ( n477 & ~n975 ) | ( n967 & ~n975 ) ;
  assign n3142 = n199 & n3141 ;
  assign n3143 = n1546 & ~n3142 ;
  assign n3144 = n3143 ^ n565 ^ 1'b0 ;
  assign n3145 = ( n944 & n1680 ) | ( n944 & ~n1698 ) | ( n1680 & ~n1698 ) ;
  assign n3146 = ( ~n908 & n1479 ) | ( ~n908 & n3145 ) | ( n1479 & n3145 ) ;
  assign n3147 = ( ~n344 & n1998 ) | ( ~n344 & n3146 ) | ( n1998 & n3146 ) ;
  assign n3148 = n3147 ^ n1106 ^ n774 ;
  assign n3149 = x27 & ~n2013 ;
  assign n3150 = n3149 ^ n1216 ^ 1'b0 ;
  assign n3151 = ( n2121 & n2350 ) | ( n2121 & ~n3150 ) | ( n2350 & ~n3150 ) ;
  assign n3152 = n2670 ^ n2216 ^ 1'b0 ;
  assign n3153 = ~n1232 & n3152 ;
  assign n3154 = ~n445 & n3153 ;
  assign n3155 = ~n1849 & n3154 ;
  assign n3156 = n3155 ^ n1424 ^ 1'b0 ;
  assign n3157 = ( ~n387 & n1488 ) | ( ~n387 & n2072 ) | ( n1488 & n2072 ) ;
  assign n3158 = ( n1185 & ~n2367 ) | ( n1185 & n3157 ) | ( ~n2367 & n3157 ) ;
  assign n3159 = n3158 ^ n2518 ^ n1037 ;
  assign n3160 = n1302 | n1509 ;
  assign n3161 = ( ~n846 & n1409 ) | ( ~n846 & n3160 ) | ( n1409 & n3160 ) ;
  assign n3162 = n459 & n1248 ;
  assign n3163 = n2712 ^ n1036 ^ 1'b0 ;
  assign n3164 = n734 | n3163 ;
  assign n3165 = n3164 ^ n2939 ^ n901 ;
  assign n3166 = n3165 ^ n826 ^ n580 ;
  assign n3167 = n2049 ^ n783 ^ 1'b0 ;
  assign n3168 = ( ~n665 & n3043 ) | ( ~n665 & n3167 ) | ( n3043 & n3167 ) ;
  assign n3169 = ( n992 & ~n1382 ) | ( n992 & n3168 ) | ( ~n1382 & n3168 ) ;
  assign n3170 = ( ~n3034 & n3166 ) | ( ~n3034 & n3169 ) | ( n3166 & n3169 ) ;
  assign n3171 = n265 | n2358 ;
  assign n3172 = n497 | n3171 ;
  assign n3175 = n1035 ^ n934 ^ 1'b0 ;
  assign n3173 = n288 | n349 ;
  assign n3174 = ( n371 & n2256 ) | ( n371 & ~n3173 ) | ( n2256 & ~n3173 ) ;
  assign n3176 = n3175 ^ n3174 ^ 1'b0 ;
  assign n3177 = n3172 & ~n3176 ;
  assign n3178 = ~n1785 & n3177 ;
  assign n3179 = n3178 ^ n272 ^ n161 ;
  assign n3180 = n1817 ^ n699 ^ 1'b0 ;
  assign n3181 = n813 & n3180 ;
  assign n3182 = ~n1723 & n3181 ;
  assign n3183 = n3182 ^ n575 ^ 1'b0 ;
  assign n3184 = n3183 ^ n2767 ^ n1563 ;
  assign n3185 = n3184 ^ n2733 ^ n643 ;
  assign n3186 = ( n269 & n1808 ) | ( n269 & ~n2428 ) | ( n1808 & ~n2428 ) ;
  assign n3187 = ( n738 & n2950 ) | ( n738 & ~n3186 ) | ( n2950 & ~n3186 ) ;
  assign n3193 = n2503 ^ n2137 ^ n1547 ;
  assign n3188 = ( ~x10 & n1000 ) | ( ~x10 & n2139 ) | ( n1000 & n2139 ) ;
  assign n3189 = n1088 & n2682 ;
  assign n3190 = n3188 & n3189 ;
  assign n3191 = ( n635 & ~n3131 ) | ( n635 & n3190 ) | ( ~n3131 & n3190 ) ;
  assign n3192 = n3191 ^ n2932 ^ n1297 ;
  assign n3194 = n3193 ^ n3192 ^ n2940 ;
  assign n3195 = ( ~n544 & n1376 ) | ( ~n544 & n1989 ) | ( n1376 & n1989 ) ;
  assign n3196 = n1953 ^ n1117 ^ 1'b0 ;
  assign n3197 = n3196 ^ n2669 ^ n1108 ;
  assign n3198 = x15 & n805 ;
  assign n3199 = n1472 & ~n1582 ;
  assign n3200 = ( n414 & n1626 ) | ( n414 & ~n3199 ) | ( n1626 & ~n3199 ) ;
  assign n3201 = ( n3197 & n3198 ) | ( n3197 & ~n3200 ) | ( n3198 & ~n3200 ) ;
  assign n3202 = ( n551 & ~n3195 ) | ( n551 & n3201 ) | ( ~n3195 & n3201 ) ;
  assign n3203 = n722 ^ n165 ^ 1'b0 ;
  assign n3204 = n728 | n3203 ;
  assign n3205 = n1353 & ~n3204 ;
  assign n3206 = ( ~n1826 & n3202 ) | ( ~n1826 & n3205 ) | ( n3202 & n3205 ) ;
  assign n3210 = n913 ^ n486 ^ x106 ;
  assign n3207 = ( n564 & n857 ) | ( n564 & ~n860 ) | ( n857 & ~n860 ) ;
  assign n3208 = n2968 ^ n1470 ^ 1'b0 ;
  assign n3209 = ( n429 & ~n3207 ) | ( n429 & n3208 ) | ( ~n3207 & n3208 ) ;
  assign n3211 = n3210 ^ n3209 ^ n1201 ;
  assign n3212 = n2495 & n3211 ;
  assign n3213 = ~n280 & n535 ;
  assign n3214 = ~n337 & n3213 ;
  assign n3215 = ~n1136 & n1258 ;
  assign n3216 = n545 & ~n2928 ;
  assign n3217 = n3216 ^ n883 ^ 1'b0 ;
  assign n3218 = n451 ^ n313 ^ 1'b0 ;
  assign n3219 = ~n743 & n3218 ;
  assign n3220 = ~n1407 & n3219 ;
  assign n3221 = ( n3198 & ~n3217 ) | ( n3198 & n3220 ) | ( ~n3217 & n3220 ) ;
  assign n3226 = ( n1540 & n1550 ) | ( n1540 & n1601 ) | ( n1550 & n1601 ) ;
  assign n3227 = n3226 ^ n1578 ^ n741 ;
  assign n3222 = n1707 ^ n1374 ^ 1'b0 ;
  assign n3223 = n801 ^ n285 ^ n264 ;
  assign n3224 = n2410 & ~n3223 ;
  assign n3225 = ( n278 & ~n3222 ) | ( n278 & n3224 ) | ( ~n3222 & n3224 ) ;
  assign n3228 = n3227 ^ n3225 ^ n785 ;
  assign n3229 = ( ~n3215 & n3221 ) | ( ~n3215 & n3228 ) | ( n3221 & n3228 ) ;
  assign n3230 = n2139 ^ n731 ^ 1'b0 ;
  assign n3231 = n589 ^ n330 ^ 1'b0 ;
  assign n3232 = ~n370 & n3231 ;
  assign n3233 = n3232 ^ n1355 ^ n1285 ;
  assign n3234 = n3233 ^ n844 ^ n386 ;
  assign n3235 = n372 | n986 ;
  assign n3236 = n3235 ^ n146 ^ 1'b0 ;
  assign n3237 = ( n728 & ~n1356 ) | ( n728 & n3236 ) | ( ~n1356 & n3236 ) ;
  assign n3241 = n129 & n1647 ;
  assign n3242 = n1663 & ~n3241 ;
  assign n3238 = n1710 ^ n969 ^ n582 ;
  assign n3239 = n3238 ^ n345 ^ 1'b0 ;
  assign n3240 = n3239 ^ n2146 ^ n723 ;
  assign n3243 = n3242 ^ n3240 ^ n831 ;
  assign n3244 = n3237 | n3243 ;
  assign n3245 = n253 | n1687 ;
  assign n3246 = n278 | n3245 ;
  assign n3247 = n3246 ^ n3093 ^ n2385 ;
  assign n3248 = n3247 ^ n2882 ^ n1476 ;
  assign n3259 = x12 & ~n1362 ;
  assign n3260 = ~n930 & n3259 ;
  assign n3261 = n3260 ^ n1620 ^ 1'b0 ;
  assign n3262 = n433 & ~n3261 ;
  assign n3263 = ~n1347 & n3262 ;
  assign n3249 = n725 ^ x102 ^ 1'b0 ;
  assign n3253 = n1858 ^ n1332 ^ 1'b0 ;
  assign n3254 = n3138 & ~n3253 ;
  assign n3255 = n3254 ^ n1062 ^ 1'b0 ;
  assign n3256 = n2860 | n3255 ;
  assign n3250 = ( n477 & ~n688 ) | ( n477 & n965 ) | ( ~n688 & n965 ) ;
  assign n3251 = n2999 | n3250 ;
  assign n3252 = ( n1309 & ~n1984 ) | ( n1309 & n3251 ) | ( ~n1984 & n3251 ) ;
  assign n3257 = n3256 ^ n3252 ^ n1362 ;
  assign n3258 = n3249 & n3257 ;
  assign n3264 = n3263 ^ n3258 ^ 1'b0 ;
  assign n3265 = n1508 ^ n794 ^ n222 ;
  assign n3266 = ~n2513 & n3265 ;
  assign n3267 = n1919 ^ n1534 ^ x93 ;
  assign n3268 = n3267 ^ n609 ^ n165 ;
  assign n3274 = n641 ^ n367 ^ 1'b0 ;
  assign n3275 = n2840 & ~n3274 ;
  assign n3269 = n1199 ^ n671 ^ n326 ;
  assign n3270 = n777 | n3269 ;
  assign n3271 = n3270 ^ n1347 ^ n379 ;
  assign n3272 = n635 | n3000 ;
  assign n3273 = n3271 & ~n3272 ;
  assign n3276 = n3275 ^ n3273 ^ 1'b0 ;
  assign n3277 = ( ~n222 & n557 ) | ( ~n222 & n2164 ) | ( n557 & n2164 ) ;
  assign n3278 = ( ~n711 & n1745 ) | ( ~n711 & n2695 ) | ( n1745 & n2695 ) ;
  assign n3279 = ( ~n820 & n3277 ) | ( ~n820 & n3278 ) | ( n3277 & n3278 ) ;
  assign n3280 = n3279 ^ n2933 ^ 1'b0 ;
  assign n3281 = n3276 | n3280 ;
  assign n3282 = n2069 ^ n333 ^ 1'b0 ;
  assign n3283 = ~n2448 & n2570 ;
  assign n3284 = ~n2738 & n3283 ;
  assign n3285 = n3282 & n3284 ;
  assign n3286 = n3285 ^ n3266 ^ n2972 ;
  assign n3287 = ~n840 & n2349 ;
  assign n3288 = n3287 ^ n1421 ^ 1'b0 ;
  assign n3289 = n676 & n2968 ;
  assign n3290 = ~n3288 & n3289 ;
  assign n3295 = n2328 ^ n1303 ^ 1'b0 ;
  assign n3296 = n3295 ^ n2645 ^ n132 ;
  assign n3292 = ( x5 & n330 ) | ( x5 & ~n490 ) | ( n330 & ~n490 ) ;
  assign n3293 = n3292 ^ n461 ^ n339 ;
  assign n3294 = ( ~x110 & n2943 ) | ( ~x110 & n3293 ) | ( n2943 & n3293 ) ;
  assign n3291 = n2091 ^ n1990 ^ 1'b0 ;
  assign n3297 = n3296 ^ n3294 ^ n3291 ;
  assign n3298 = n823 ^ n611 ^ n496 ;
  assign n3299 = n233 & ~n3298 ;
  assign n3300 = n1773 & n3299 ;
  assign n3301 = n3222 ^ n390 ^ 1'b0 ;
  assign n3302 = n1574 | n2314 ;
  assign n3303 = n203 | n2264 ;
  assign n3304 = n1106 & ~n3303 ;
  assign n3305 = ( n552 & n1173 ) | ( n552 & ~n1353 ) | ( n1173 & ~n1353 ) ;
  assign n3306 = n2019 ^ n1015 ^ x85 ;
  assign n3307 = ( n809 & n3305 ) | ( n809 & ~n3306 ) | ( n3305 & ~n3306 ) ;
  assign n3308 = ( ~n3302 & n3304 ) | ( ~n3302 & n3307 ) | ( n3304 & n3307 ) ;
  assign n3311 = n3295 ^ n2517 ^ 1'b0 ;
  assign n3309 = n658 | n681 ;
  assign n3310 = n3309 ^ n1204 ^ n543 ;
  assign n3312 = n3311 ^ n3310 ^ n145 ;
  assign n3313 = n3312 ^ n3078 ^ 1'b0 ;
  assign n3314 = n2287 | n3313 ;
  assign n3315 = ( ~n333 & n551 ) | ( ~n333 & n1210 ) | ( n551 & n1210 ) ;
  assign n3316 = x26 | n3315 ;
  assign n3317 = ( n1187 & n2221 ) | ( n1187 & ~n3316 ) | ( n2221 & ~n3316 ) ;
  assign n3318 = n1101 ^ n386 ^ x111 ;
  assign n3319 = ( x87 & ~n494 ) | ( x87 & n3318 ) | ( ~n494 & n3318 ) ;
  assign n3320 = ~n810 & n2495 ;
  assign n3321 = ~n3319 & n3320 ;
  assign n3322 = ( x126 & n2156 ) | ( x126 & ~n3321 ) | ( n2156 & ~n3321 ) ;
  assign n3323 = n1267 ^ n423 ^ x102 ;
  assign n3324 = n591 & n1560 ;
  assign n3325 = ~n3323 & n3324 ;
  assign n3326 = n3325 ^ n1957 ^ 1'b0 ;
  assign n3327 = ( n1421 & n3113 ) | ( n1421 & ~n3326 ) | ( n3113 & ~n3326 ) ;
  assign n3328 = n3327 ^ n486 ^ 1'b0 ;
  assign n3330 = ( x62 & ~x106 ) | ( x62 & n680 ) | ( ~x106 & n680 ) ;
  assign n3329 = n2383 ^ n2083 ^ 1'b0 ;
  assign n3331 = n3330 ^ n3329 ^ n1616 ;
  assign n3332 = n1528 ^ n867 ^ 1'b0 ;
  assign n3333 = n2246 | n3332 ;
  assign n3334 = ~n3331 & n3333 ;
  assign n3335 = ( n859 & n1229 ) | ( n859 & ~n1518 ) | ( n1229 & ~n1518 ) ;
  assign n3336 = ( n1845 & n2358 ) | ( n1845 & n3335 ) | ( n2358 & n3335 ) ;
  assign n3337 = n3336 ^ n2524 ^ n1032 ;
  assign n3338 = x83 & ~n3337 ;
  assign n3339 = n3338 ^ n3307 ^ x115 ;
  assign n3340 = ( n154 & n2020 ) | ( n154 & ~n2402 ) | ( n2020 & ~n2402 ) ;
  assign n3341 = n3129 & n3248 ;
  assign n3342 = n3340 & n3341 ;
  assign n3343 = n291 & ~n1017 ;
  assign n3344 = n3343 ^ n3024 ^ n1876 ;
  assign n3346 = n914 & n2639 ;
  assign n3347 = n1603 & n3346 ;
  assign n3348 = n394 | n1047 ;
  assign n3349 = n3348 ^ n1061 ^ 1'b0 ;
  assign n3350 = n3347 | n3349 ;
  assign n3345 = n2185 ^ n1413 ^ n503 ;
  assign n3351 = n3350 ^ n3345 ^ 1'b0 ;
  assign n3352 = n1889 ^ n881 ^ x108 ;
  assign n3353 = ( ~n362 & n1066 ) | ( ~n362 & n3352 ) | ( n1066 & n3352 ) ;
  assign n3354 = ~n423 & n3353 ;
  assign n3355 = n1632 ^ n669 ^ 1'b0 ;
  assign n3356 = n3355 ^ n2467 ^ n2312 ;
  assign n3357 = ( x55 & ~n1190 ) | ( x55 & n3356 ) | ( ~n1190 & n3356 ) ;
  assign n3358 = ( n2144 & n3354 ) | ( n2144 & n3357 ) | ( n3354 & n3357 ) ;
  assign n3359 = n2414 & ~n3358 ;
  assign n3360 = ~n2783 & n3359 ;
  assign n3372 = n535 & n1248 ;
  assign n3373 = ~n225 & n3372 ;
  assign n3374 = n1051 ^ n658 ^ 1'b0 ;
  assign n3375 = n3373 | n3374 ;
  assign n3369 = n608 | n1517 ;
  assign n3370 = n132 | n3369 ;
  assign n3371 = ~n3315 & n3370 ;
  assign n3376 = n3375 ^ n3371 ^ 1'b0 ;
  assign n3361 = ( n823 & n2097 ) | ( n823 & ~n2727 ) | ( n2097 & ~n2727 ) ;
  assign n3362 = ( n577 & ~n1646 ) | ( n577 & n3361 ) | ( ~n1646 & n3361 ) ;
  assign n3363 = n187 | n1384 ;
  assign n3364 = n378 | n3363 ;
  assign n3365 = ( n1097 & n1591 ) | ( n1097 & n3364 ) | ( n1591 & n3364 ) ;
  assign n3366 = n3365 ^ n3053 ^ 1'b0 ;
  assign n3367 = n3362 | n3366 ;
  assign n3368 = n3367 ^ n663 ^ 1'b0 ;
  assign n3377 = n3376 ^ n3368 ^ 1'b0 ;
  assign n3386 = ~n667 & n1166 ;
  assign n3387 = n3386 ^ n1971 ^ 1'b0 ;
  assign n3388 = n553 & n3387 ;
  assign n3378 = n2950 ^ n1763 ^ 1'b0 ;
  assign n3379 = n1560 & n3378 ;
  assign n3380 = n3379 ^ n3306 ^ x5 ;
  assign n3381 = n2760 ^ n1840 ^ n997 ;
  assign n3382 = n494 & n617 ;
  assign n3383 = n3381 & n3382 ;
  assign n3384 = n3383 ^ n1991 ^ 1'b0 ;
  assign n3385 = ( n2846 & ~n3380 ) | ( n2846 & n3384 ) | ( ~n3380 & n3384 ) ;
  assign n3389 = n3388 ^ n3385 ^ x74 ;
  assign n3390 = n2826 ^ n2804 ^ n1540 ;
  assign n3391 = ~n1302 & n2423 ;
  assign n3399 = ( n820 & n1191 ) | ( n820 & n2918 ) | ( n1191 & n2918 ) ;
  assign n3400 = n3399 ^ n3094 ^ 1'b0 ;
  assign n3401 = n2110 & n3400 ;
  assign n3392 = n1808 ^ n1314 ^ 1'b0 ;
  assign n3393 = ( n1518 & n2479 ) | ( n1518 & n3392 ) | ( n2479 & n3392 ) ;
  assign n3394 = n3393 ^ n742 ^ 1'b0 ;
  assign n3395 = ~n583 & n3394 ;
  assign n3396 = ( ~n770 & n1114 ) | ( ~n770 & n3395 ) | ( n1114 & n3395 ) ;
  assign n3397 = n1468 & ~n3396 ;
  assign n3398 = ~n2193 & n3397 ;
  assign n3402 = n3401 ^ n3398 ^ 1'b0 ;
  assign n3404 = n2497 ^ n750 ^ 1'b0 ;
  assign n3403 = n460 | n3354 ;
  assign n3405 = n3404 ^ n3403 ^ 1'b0 ;
  assign n3406 = x112 & n2353 ;
  assign n3407 = n3405 & n3406 ;
  assign n3408 = n2185 | n2548 ;
  assign n3410 = ( n516 & n997 ) | ( n516 & n3232 ) | ( n997 & n3232 ) ;
  assign n3409 = x3 & ~n2616 ;
  assign n3411 = n3410 ^ n3409 ^ n2385 ;
  assign n3415 = ( ~n892 & n2168 ) | ( ~n892 & n3208 ) | ( n2168 & n3208 ) ;
  assign n3416 = n3415 ^ n236 ^ n157 ;
  assign n3412 = ~n611 & n1626 ;
  assign n3413 = n1810 & n3412 ;
  assign n3414 = n2784 | n3413 ;
  assign n3417 = n3416 ^ n3414 ^ 1'b0 ;
  assign n3418 = ~n2701 & n3417 ;
  assign n3419 = n2175 ^ x97 ^ 1'b0 ;
  assign n3420 = x62 & n3419 ;
  assign n3421 = n3420 ^ n1626 ^ n292 ;
  assign n3422 = n2840 ^ n1616 ^ n320 ;
  assign n3423 = ( ~x15 & n3421 ) | ( ~x15 & n3422 ) | ( n3421 & n3422 ) ;
  assign n3424 = n3423 ^ n1211 ^ 1'b0 ;
  assign n3425 = n3424 ^ n2135 ^ 1'b0 ;
  assign n3433 = n1632 ^ n1459 ^ n831 ;
  assign n3434 = ( n487 & ~n2009 ) | ( n487 & n3433 ) | ( ~n2009 & n3433 ) ;
  assign n3436 = ~n406 & n1269 ;
  assign n3437 = n3436 ^ n238 ^ 1'b0 ;
  assign n3438 = ( n533 & n739 ) | ( n533 & n1246 ) | ( n739 & n1246 ) ;
  assign n3439 = ( n673 & n3437 ) | ( n673 & n3438 ) | ( n3437 & n3438 ) ;
  assign n3435 = n970 & ~n1741 ;
  assign n3440 = n3439 ^ n3435 ^ 1'b0 ;
  assign n3441 = ( n2149 & n3434 ) | ( n2149 & n3440 ) | ( n3434 & n3440 ) ;
  assign n3430 = n1366 ^ n690 ^ 1'b0 ;
  assign n3429 = n2920 & ~n3393 ;
  assign n3431 = n3430 ^ n3429 ^ 1'b0 ;
  assign n3426 = x104 & n2081 ;
  assign n3427 = ~n2944 & n3426 ;
  assign n3428 = n291 & n3427 ;
  assign n3432 = n3431 ^ n3428 ^ n1190 ;
  assign n3442 = n3441 ^ n3432 ^ 1'b0 ;
  assign n3443 = n298 & ~n1061 ;
  assign n3445 = x46 & n2138 ;
  assign n3446 = ~n165 & n3445 ;
  assign n3444 = n3420 ^ n2517 ^ n870 ;
  assign n3447 = n3446 ^ n3444 ^ 1'b0 ;
  assign n3448 = n3443 | n3447 ;
  assign n3449 = ( n447 & n1069 ) | ( n447 & n3448 ) | ( n1069 & n3448 ) ;
  assign n3459 = n1525 ^ n667 ^ 1'b0 ;
  assign n3460 = n2070 | n3459 ;
  assign n3455 = n2730 ^ n334 ^ 1'b0 ;
  assign n3456 = ~n1780 & n3455 ;
  assign n3457 = n2826 ^ n2305 ^ 1'b0 ;
  assign n3458 = n3456 & n3457 ;
  assign n3450 = n583 ^ n333 ^ x32 ;
  assign n3451 = n3450 ^ n132 ^ 1'b0 ;
  assign n3452 = n139 & n3451 ;
  assign n3453 = ~n2712 & n3452 ;
  assign n3454 = n3453 ^ n3132 ^ 1'b0 ;
  assign n3461 = n3460 ^ n3458 ^ n3454 ;
  assign n3462 = ( ~n204 & n523 ) | ( ~n204 & n559 ) | ( n523 & n559 ) ;
  assign n3463 = n499 & n3462 ;
  assign n3464 = ( n478 & ~n670 ) | ( n478 & n1705 ) | ( ~n670 & n1705 ) ;
  assign n3465 = ( n1396 & n3463 ) | ( n1396 & n3464 ) | ( n3463 & n3464 ) ;
  assign n3466 = n2079 & n3084 ;
  assign n3467 = ( n1686 & n1900 ) | ( n1686 & ~n3466 ) | ( n1900 & ~n3466 ) ;
  assign n3468 = ~n881 & n3093 ;
  assign n3469 = n1176 & n3468 ;
  assign n3470 = n3469 ^ n2747 ^ n2515 ;
  assign n3471 = n3470 ^ n2059 ^ x1 ;
  assign n3472 = n1131 ^ n320 ^ n293 ;
  assign n3473 = n2925 | n3472 ;
  assign n3474 = n3473 ^ n1806 ^ n1326 ;
  assign n3475 = ( n870 & n2412 ) | ( n870 & ~n3474 ) | ( n2412 & ~n3474 ) ;
  assign n3476 = n3475 ^ n462 ^ 1'b0 ;
  assign n3477 = n3471 | n3476 ;
  assign n3478 = n1402 ^ n684 ^ n310 ;
  assign n3479 = ~n783 & n3478 ;
  assign n3480 = ~n3236 & n3479 ;
  assign n3481 = n3480 ^ n2503 ^ n1573 ;
  assign n3482 = ( ~n1780 & n2308 ) | ( ~n1780 & n3481 ) | ( n2308 & n3481 ) ;
  assign n3483 = n1690 ^ n822 ^ n392 ;
  assign n3484 = ( n2089 & n2388 ) | ( n2089 & ~n3483 ) | ( n2388 & ~n3483 ) ;
  assign n3485 = ( n190 & n1972 ) | ( n190 & n2443 ) | ( n1972 & n2443 ) ;
  assign n3486 = ( n287 & ~n293 ) | ( n287 & n742 ) | ( ~n293 & n742 ) ;
  assign n3487 = ~n506 & n1425 ;
  assign n3488 = n3486 & n3487 ;
  assign n3489 = ( x7 & n1079 ) | ( x7 & n3488 ) | ( n1079 & n3488 ) ;
  assign n3490 = n3489 ^ n2996 ^ n887 ;
  assign n3491 = ( n1046 & n3485 ) | ( n1046 & n3490 ) | ( n3485 & n3490 ) ;
  assign n3493 = n2019 & n3141 ;
  assign n3494 = ~n1166 & n3493 ;
  assign n3495 = n3494 ^ n3421 ^ n2031 ;
  assign n3492 = n1131 | n2978 ;
  assign n3496 = n3495 ^ n3492 ^ 1'b0 ;
  assign n3497 = n433 & ~n848 ;
  assign n3498 = n3497 ^ n897 ^ 1'b0 ;
  assign n3499 = n3498 ^ n3424 ^ n2893 ;
  assign n3500 = ( n3491 & ~n3496 ) | ( n3491 & n3499 ) | ( ~n3496 & n3499 ) ;
  assign n3501 = ( n897 & n1688 ) | ( n897 & ~n3225 ) | ( n1688 & ~n3225 ) ;
  assign n3502 = n261 ^ n226 ^ 1'b0 ;
  assign n3503 = n255 | n3502 ;
  assign n3504 = n3034 ^ n2539 ^ 1'b0 ;
  assign n3505 = ~n3503 & n3504 ;
  assign n3506 = n3505 ^ n2935 ^ n1632 ;
  assign n3507 = n2622 ^ n1686 ^ n826 ;
  assign n3508 = n3219 ^ n1961 ^ n385 ;
  assign n3509 = n2708 ^ n2504 ^ n1075 ;
  assign n3510 = x55 | n673 ;
  assign n3511 = n572 & ~n1925 ;
  assign n3512 = n3511 ^ n1127 ^ 1'b0 ;
  assign n3513 = n3510 | n3512 ;
  assign n3514 = n3509 & n3513 ;
  assign n3515 = n533 ^ n379 ^ n231 ;
  assign n3516 = n704 & ~n1164 ;
  assign n3518 = n2436 ^ n2292 ^ n1216 ;
  assign n3517 = ( ~n403 & n799 ) | ( ~n403 & n1917 ) | ( n799 & n1917 ) ;
  assign n3519 = n3518 ^ n3517 ^ 1'b0 ;
  assign n3520 = n3516 & n3519 ;
  assign n3521 = n3515 & n3520 ;
  assign n3522 = n3228 | n3521 ;
  assign n3523 = ( n1493 & n1685 ) | ( n1493 & ~n2436 ) | ( n1685 & ~n2436 ) ;
  assign n3524 = n3523 ^ n2386 ^ 1'b0 ;
  assign n3525 = n3524 ^ n1836 ^ n490 ;
  assign n3526 = ( ~n1981 & n2147 ) | ( ~n1981 & n3525 ) | ( n2147 & n3525 ) ;
  assign n3527 = ( ~n607 & n1345 ) | ( ~n607 & n3526 ) | ( n1345 & n3526 ) ;
  assign n3528 = ( n613 & n1697 ) | ( n613 & n2933 ) | ( n1697 & n2933 ) ;
  assign n3529 = n3528 ^ n1929 ^ n186 ;
  assign n3530 = n496 ^ n222 ^ 1'b0 ;
  assign n3531 = ( ~n233 & n2450 ) | ( ~n233 & n2958 ) | ( n2450 & n2958 ) ;
  assign n3532 = ( n1294 & n3530 ) | ( n1294 & ~n3531 ) | ( n3530 & ~n3531 ) ;
  assign n3533 = n1935 & ~n3532 ;
  assign n3534 = n3529 & n3533 ;
  assign n3535 = ( ~n729 & n1792 ) | ( ~n729 & n2928 ) | ( n1792 & n2928 ) ;
  assign n3536 = ( n784 & ~n1054 ) | ( n784 & n2063 ) | ( ~n1054 & n2063 ) ;
  assign n3537 = n3536 ^ n2234 ^ n2124 ;
  assign n3538 = n3537 ^ n2512 ^ 1'b0 ;
  assign n3539 = n2400 ^ x3 ^ 1'b0 ;
  assign n3540 = x73 & n3539 ;
  assign n3542 = ~n1566 & n2218 ;
  assign n3543 = n1512 & n3542 ;
  assign n3544 = n1139 & ~n1294 ;
  assign n3545 = ~n3543 & n3544 ;
  assign n3546 = n196 & n3545 ;
  assign n3541 = n3081 ^ n600 ^ n243 ;
  assign n3547 = n3546 ^ n3541 ^ 1'b0 ;
  assign n3548 = n503 | n3547 ;
  assign n3549 = n3548 ^ n1553 ^ 1'b0 ;
  assign n3550 = n3540 & n3549 ;
  assign n3551 = n2412 ^ n1054 ^ x48 ;
  assign n3552 = n2581 ^ n1538 ^ n1320 ;
  assign n3553 = ~n160 & n484 ;
  assign n3554 = n3553 ^ n3305 ^ n1052 ;
  assign n3555 = x80 & ~n738 ;
  assign n3556 = n3555 ^ n591 ^ 1'b0 ;
  assign n3557 = ~n3259 & n3556 ;
  assign n3558 = n3557 ^ n1207 ^ n370 ;
  assign n3559 = ( ~n2296 & n3554 ) | ( ~n2296 & n3558 ) | ( n3554 & n3558 ) ;
  assign n3560 = n2025 & n3559 ;
  assign n3561 = n3560 ^ n496 ^ 1'b0 ;
  assign n3562 = ~n342 & n2736 ;
  assign n3563 = n3562 ^ n589 ^ 1'b0 ;
  assign n3564 = ( ~n500 & n1991 ) | ( ~n500 & n2561 ) | ( n1991 & n2561 ) ;
  assign n3565 = n3564 ^ n3097 ^ 1'b0 ;
  assign n3566 = n3565 ^ n1955 ^ n950 ;
  assign n3575 = ( x49 & n250 ) | ( x49 & n870 ) | ( n250 & n870 ) ;
  assign n3576 = n1515 | n3575 ;
  assign n3570 = n1749 ^ n1117 ^ 1'b0 ;
  assign n3567 = n1078 & ~n1484 ;
  assign n3568 = ~n753 & n3567 ;
  assign n3569 = ~n1170 & n3568 ;
  assign n3571 = n3570 ^ n3569 ^ n2185 ;
  assign n3572 = ( n1000 & n1515 ) | ( n1000 & n3571 ) | ( n1515 & n3571 ) ;
  assign n3573 = n3572 ^ n3395 ^ x108 ;
  assign n3574 = n3573 ^ n1715 ^ n472 ;
  assign n3577 = n3576 ^ n3574 ^ n1583 ;
  assign n3580 = ( n581 & n1210 ) | ( n581 & ~n1910 ) | ( n1210 & ~n1910 ) ;
  assign n3578 = n1099 & ~n3319 ;
  assign n3579 = n3578 ^ n1953 ^ 1'b0 ;
  assign n3581 = n3580 ^ n3579 ^ n3145 ;
  assign n3582 = n2870 ^ n2335 ^ n913 ;
  assign n3583 = n3582 ^ n3336 ^ n3333 ;
  assign n3584 = ( n1646 & n3296 ) | ( n1646 & n3583 ) | ( n3296 & n3583 ) ;
  assign n3585 = ~n1293 & n3584 ;
  assign n3586 = ~n3581 & n3585 ;
  assign n3587 = n760 ^ n565 ^ x78 ;
  assign n3588 = n1522 ^ n1130 ^ n914 ;
  assign n3589 = ( n686 & n780 ) | ( n686 & n3364 ) | ( n780 & n3364 ) ;
  assign n3590 = n3589 ^ n322 ^ 1'b0 ;
  assign n3591 = n3588 & ~n3590 ;
  assign n3592 = n3591 ^ n2434 ^ n778 ;
  assign n3593 = ( ~n1131 & n3587 ) | ( ~n1131 & n3592 ) | ( n3587 & n3592 ) ;
  assign n3594 = n3593 ^ n2483 ^ n356 ;
  assign n3598 = n2211 ^ n2039 ^ n1474 ;
  assign n3595 = n642 ^ n383 ^ n366 ;
  assign n3596 = ( n462 & ~n2513 ) | ( n462 & n2750 ) | ( ~n2513 & n2750 ) ;
  assign n3597 = ( n1442 & ~n3595 ) | ( n1442 & n3596 ) | ( ~n3595 & n3596 ) ;
  assign n3599 = n3598 ^ n3597 ^ n883 ;
  assign n3600 = n3599 ^ n2907 ^ 1'b0 ;
  assign n3601 = ( n517 & n1597 ) | ( n517 & ~n3370 ) | ( n1597 & ~n3370 ) ;
  assign n3602 = ( n1699 & ~n1944 ) | ( n1699 & n3601 ) | ( ~n1944 & n3601 ) ;
  assign n3603 = n2452 ^ n933 ^ n705 ;
  assign n3604 = n3603 ^ n2248 ^ 1'b0 ;
  assign n3605 = n329 & ~n3604 ;
  assign n3606 = n3605 ^ n2019 ^ 1'b0 ;
  assign n3607 = n3606 ^ n2848 ^ n2493 ;
  assign n3608 = n3607 ^ n139 ^ 1'b0 ;
  assign n3609 = n1967 & ~n3608 ;
  assign n3611 = ( x122 & n859 ) | ( x122 & ~n1191 ) | ( n859 & ~n1191 ) ;
  assign n3610 = n2461 ^ n2282 ^ n1436 ;
  assign n3612 = n3611 ^ n3610 ^ n835 ;
  assign n3618 = ~n487 & n1104 ;
  assign n3619 = n3618 ^ n312 ^ 1'b0 ;
  assign n3613 = n1480 ^ x59 ^ x18 ;
  assign n3614 = n267 & ~n3613 ;
  assign n3615 = n3614 ^ n2405 ^ 1'b0 ;
  assign n3616 = n2011 ^ n2003 ^ n480 ;
  assign n3617 = ( n3361 & n3615 ) | ( n3361 & ~n3616 ) | ( n3615 & ~n3616 ) ;
  assign n3620 = n3619 ^ n3617 ^ n1042 ;
  assign n3623 = ~n744 & n2057 ;
  assign n3621 = ( n290 & ~n1556 ) | ( n290 & n3265 ) | ( ~n1556 & n3265 ) ;
  assign n3622 = ( n1402 & n3006 ) | ( n1402 & ~n3621 ) | ( n3006 & ~n3621 ) ;
  assign n3624 = n3623 ^ n3622 ^ n2984 ;
  assign n3629 = ~n341 & n828 ;
  assign n3625 = n889 | n1059 ;
  assign n3626 = n421 & ~n3625 ;
  assign n3627 = n3626 ^ n830 ^ x45 ;
  assign n3628 = n1695 | n3627 ;
  assign n3630 = n3629 ^ n3628 ^ 1'b0 ;
  assign n3631 = ( ~n355 & n569 ) | ( ~n355 & n3065 ) | ( n569 & n3065 ) ;
  assign n3632 = n540 & n871 ;
  assign n3633 = n1869 ^ n1686 ^ n1599 ;
  assign n3634 = ~n2105 & n3379 ;
  assign n3635 = n3634 ^ n1189 ^ 1'b0 ;
  assign n3636 = n3635 ^ n2554 ^ n1044 ;
  assign n3637 = ( n214 & n575 ) | ( n214 & n1967 ) | ( n575 & n1967 ) ;
  assign n3638 = ( n2594 & n3636 ) | ( n2594 & ~n3637 ) | ( n3636 & ~n3637 ) ;
  assign n3639 = ~n549 & n2403 ;
  assign n3640 = n3380 & n3639 ;
  assign n3641 = n3115 ^ n247 ^ x96 ;
  assign n3642 = ( n1032 & ~n2740 ) | ( n1032 & n3027 ) | ( ~n2740 & n3027 ) ;
  assign n3643 = ( ~n1905 & n1932 ) | ( ~n1905 & n3642 ) | ( n1932 & n3642 ) ;
  assign n3644 = ~n3641 & n3643 ;
  assign n3651 = x29 & n917 ;
  assign n3652 = n1082 & n3651 ;
  assign n3650 = n252 & n1187 ;
  assign n3653 = n3652 ^ n3650 ^ 1'b0 ;
  assign n3645 = n238 & n1573 ;
  assign n3646 = ~n870 & n3645 ;
  assign n3647 = n1100 ^ n253 ^ 1'b0 ;
  assign n3648 = n3647 ^ n1470 ^ n1339 ;
  assign n3649 = n3646 | n3648 ;
  assign n3654 = n3653 ^ n3649 ^ 1'b0 ;
  assign n3655 = ( n627 & n1374 ) | ( n627 & n2372 ) | ( n1374 & n2372 ) ;
  assign n3656 = ( n308 & ~n3654 ) | ( n308 & n3655 ) | ( ~n3654 & n3655 ) ;
  assign n3657 = n1475 | n3482 ;
  assign n3661 = n3595 ^ n1488 ^ x125 ;
  assign n3658 = ( n441 & n828 ) | ( n441 & n1199 ) | ( n828 & n1199 ) ;
  assign n3659 = n2380 ^ n1321 ^ n600 ;
  assign n3660 = ( n477 & ~n3658 ) | ( n477 & n3659 ) | ( ~n3658 & n3659 ) ;
  assign n3662 = n3661 ^ n3660 ^ n2212 ;
  assign n3664 = ( n1120 & n1199 ) | ( n1120 & n2089 ) | ( n1199 & n2089 ) ;
  assign n3663 = ~n284 & n914 ;
  assign n3665 = n3664 ^ n3663 ^ 1'b0 ;
  assign n3666 = n2252 ^ n981 ^ n750 ;
  assign n3667 = n3666 ^ n3431 ^ n2264 ;
  assign n3668 = n3667 ^ n3323 ^ n2339 ;
  assign n3669 = x28 & ~n779 ;
  assign n3670 = n3669 ^ n1011 ^ 1'b0 ;
  assign n3671 = n3670 ^ n1718 ^ x54 ;
  assign n3672 = ( n1787 & n1925 ) | ( n1787 & n3671 ) | ( n1925 & n3671 ) ;
  assign n3673 = n3672 ^ n329 ^ 1'b0 ;
  assign n3674 = n3673 ^ n2386 ^ n1009 ;
  assign n3676 = x6 & x57 ;
  assign n3675 = ( n334 & n1476 ) | ( n334 & n3188 ) | ( n1476 & n3188 ) ;
  assign n3677 = n3676 ^ n3675 ^ x108 ;
  assign n3678 = ~n3185 & n3677 ;
  assign n3679 = n3678 ^ n2242 ^ 1'b0 ;
  assign n3680 = n2724 ^ n780 ^ n169 ;
  assign n3681 = ~x126 & n3680 ;
  assign n3682 = ( n359 & n1393 ) | ( n359 & n1673 ) | ( n1393 & n1673 ) ;
  assign n3683 = n2778 | n3682 ;
  assign n3684 = n2061 ^ x34 ^ 1'b0 ;
  assign n3685 = n3684 ^ n2434 ^ 1'b0 ;
  assign n3686 = ( ~x61 & n626 ) | ( ~x61 & n709 ) | ( n626 & n709 ) ;
  assign n3687 = n1191 & ~n3686 ;
  assign n3688 = ( n783 & n2998 ) | ( n783 & n3687 ) | ( n2998 & n3687 ) ;
  assign n3689 = ( ~n3683 & n3685 ) | ( ~n3683 & n3688 ) | ( n3685 & n3688 ) ;
  assign n3690 = n1016 & n1695 ;
  assign n3691 = n3690 ^ n2968 ^ n1832 ;
  assign n3692 = n2942 ^ n1570 ^ n1283 ;
  assign n3693 = ( n850 & ~n1805 ) | ( n850 & n3692 ) | ( ~n1805 & n3692 ) ;
  assign n3694 = n1714 | n3693 ;
  assign n3695 = n3691 | n3694 ;
  assign n3696 = ( ~n409 & n484 ) | ( ~n409 & n902 ) | ( n484 & n902 ) ;
  assign n3697 = n1557 | n3696 ;
  assign n3698 = n1040 ^ n491 ^ 1'b0 ;
  assign n3699 = ( n1056 & n1150 ) | ( n1056 & n2479 ) | ( n1150 & n2479 ) ;
  assign n3700 = n3676 ^ n3516 ^ 1'b0 ;
  assign n3701 = ( n2750 & n3409 ) | ( n2750 & n3700 ) | ( n3409 & n3700 ) ;
  assign n3702 = n3699 | n3701 ;
  assign n3703 = ( n330 & n482 ) | ( n330 & ~n3702 ) | ( n482 & ~n3702 ) ;
  assign n3704 = ( ~n2706 & n3698 ) | ( ~n2706 & n3703 ) | ( n3698 & n3703 ) ;
  assign n3705 = ( n562 & n1953 ) | ( n562 & n3704 ) | ( n1953 & n3704 ) ;
  assign n3706 = ( n2231 & ~n2379 ) | ( n2231 & n3248 ) | ( ~n2379 & n3248 ) ;
  assign n3707 = ( n1567 & n2620 ) | ( n1567 & ~n3172 ) | ( n2620 & ~n3172 ) ;
  assign n3711 = n1382 & ~n1895 ;
  assign n3712 = n3711 ^ n2904 ^ n569 ;
  assign n3713 = ( n319 & ~n750 ) | ( n319 & n3712 ) | ( ~n750 & n3712 ) ;
  assign n3710 = n686 ^ n509 ^ n192 ;
  assign n3714 = n3713 ^ n3710 ^ 1'b0 ;
  assign n3715 = n1348 & n2053 ;
  assign n3716 = n3714 & n3715 ;
  assign n3708 = n2569 ^ n1643 ^ n1389 ;
  assign n3709 = n1509 & ~n3708 ;
  assign n3717 = n3716 ^ n3709 ^ 1'b0 ;
  assign n3718 = ( n447 & n3707 ) | ( n447 & n3717 ) | ( n3707 & n3717 ) ;
  assign n3719 = n988 & ~n2040 ;
  assign n3720 = n1190 & ~n3719 ;
  assign n3721 = n3720 ^ n186 ^ 1'b0 ;
  assign n3722 = n665 | n2275 ;
  assign n3723 = n3721 | n3722 ;
  assign n3724 = n3723 ^ n3421 ^ 1'b0 ;
  assign n3725 = n667 | n3724 ;
  assign n3729 = ( ~n197 & n1384 ) | ( ~n197 & n2645 ) | ( n1384 & n2645 ) ;
  assign n3727 = x79 & ~n2247 ;
  assign n3728 = ~n2281 & n3727 ;
  assign n3726 = n3485 ^ n3018 ^ n731 ;
  assign n3730 = n3729 ^ n3728 ^ n3726 ;
  assign n3731 = n3730 ^ n508 ^ x45 ;
  assign n3732 = ~n3725 & n3731 ;
  assign n3733 = n3732 ^ n1388 ^ 1'b0 ;
  assign n3734 = ~n3718 & n3733 ;
  assign n3735 = ( n609 & ~n1599 ) | ( n609 & n2108 ) | ( ~n1599 & n2108 ) ;
  assign n3736 = n3735 ^ n2124 ^ n434 ;
  assign n3737 = ( n1303 & n2219 ) | ( n1303 & n3422 ) | ( n2219 & n3422 ) ;
  assign n3738 = n3737 ^ n2994 ^ 1'b0 ;
  assign n3739 = n3736 & ~n3738 ;
  assign n3740 = n2513 ^ n1669 ^ n994 ;
  assign n3741 = n3740 ^ n3668 ^ n445 ;
  assign n3742 = ~n359 & n1088 ;
  assign n3743 = n3742 ^ n941 ^ 1'b0 ;
  assign n3744 = n1606 & n3743 ;
  assign n3745 = n746 & n1044 ;
  assign n3746 = n3745 ^ n3222 ^ 1'b0 ;
  assign n3747 = n984 & ~n1219 ;
  assign n3748 = n3747 ^ n2034 ^ n379 ;
  assign n3749 = n3746 | n3748 ;
  assign n3750 = n3749 ^ n2521 ^ 1'b0 ;
  assign n3751 = n3750 ^ n3203 ^ n2817 ;
  assign n3756 = n1721 & n2054 ;
  assign n3757 = ~n2058 & n3756 ;
  assign n3758 = ( n555 & ~n698 ) | ( n555 & n3757 ) | ( ~n698 & n3757 ) ;
  assign n3759 = ( n567 & n2154 ) | ( n567 & ~n3758 ) | ( n2154 & ~n3758 ) ;
  assign n3752 = n1667 ^ n1648 ^ 1'b0 ;
  assign n3753 = n1230 ^ n525 ^ 1'b0 ;
  assign n3754 = ( n2151 & n3752 ) | ( n2151 & ~n3753 ) | ( n3752 & ~n3753 ) ;
  assign n3755 = n2880 & ~n3754 ;
  assign n3760 = n3759 ^ n3755 ^ 1'b0 ;
  assign n3766 = ( n526 & n1201 ) | ( n526 & n2792 ) | ( n1201 & n2792 ) ;
  assign n3767 = n485 & ~n3766 ;
  assign n3764 = n1467 | n2424 ;
  assign n3765 = n3764 ^ n1201 ^ 1'b0 ;
  assign n3768 = n3767 ^ n3765 ^ n1802 ;
  assign n3761 = ~n218 & n2779 ;
  assign n3762 = n3761 ^ n2581 ^ n1203 ;
  assign n3763 = n1167 & n3762 ;
  assign n3769 = n3768 ^ n3763 ^ 1'b0 ;
  assign n3777 = n1589 ^ n212 ^ 1'b0 ;
  assign n3778 = n355 & n3777 ;
  assign n3779 = ( n330 & ~n1642 ) | ( n330 & n3778 ) | ( ~n1642 & n3778 ) ;
  assign n3770 = n1186 ^ x49 ^ 1'b0 ;
  assign n3771 = n813 ^ x110 ^ 1'b0 ;
  assign n3772 = n2020 & n3771 ;
  assign n3773 = ( n1274 & n2009 ) | ( n1274 & n3772 ) | ( n2009 & n3772 ) ;
  assign n3774 = n3773 ^ n3651 ^ 1'b0 ;
  assign n3775 = n566 & n3774 ;
  assign n3776 = ( ~x76 & n3770 ) | ( ~x76 & n3775 ) | ( n3770 & n3775 ) ;
  assign n3780 = n3779 ^ n3776 ^ n1599 ;
  assign n3781 = n3090 ^ n2044 ^ n301 ;
  assign n3782 = n140 & ~n2480 ;
  assign n3783 = n3259 ^ n2218 ^ n977 ;
  assign n3784 = n3387 & ~n3783 ;
  assign n3785 = ~n998 & n3784 ;
  assign n3786 = n2914 ^ n2401 ^ n1029 ;
  assign n3787 = ( n2511 & ~n3785 ) | ( n2511 & n3786 ) | ( ~n3785 & n3786 ) ;
  assign n3788 = ( n928 & n1694 ) | ( n928 & ~n2816 ) | ( n1694 & ~n2816 ) ;
  assign n3789 = n3788 ^ n1092 ^ n743 ;
  assign n3790 = ( n403 & ~n965 ) | ( n403 & n1220 ) | ( ~n965 & n1220 ) ;
  assign n3791 = n681 | n3790 ;
  assign n3792 = n3789 | n3791 ;
  assign n3793 = n3162 & n3792 ;
  assign n3794 = ~n2103 & n3793 ;
  assign n3795 = ( n2151 & n3582 ) | ( n2151 & ~n3794 ) | ( n3582 & ~n3794 ) ;
  assign n3796 = n2645 ^ n1258 ^ 1'b0 ;
  assign n3797 = n425 & ~n1015 ;
  assign n3798 = n3797 ^ x93 ^ 1'b0 ;
  assign n3799 = n3798 ^ n1129 ^ n1076 ;
  assign n3800 = n3799 ^ n1850 ^ n645 ;
  assign n3801 = ( ~n2232 & n2642 ) | ( ~n2232 & n3800 ) | ( n2642 & n3800 ) ;
  assign n3802 = n1068 & ~n3801 ;
  assign n3803 = n3802 ^ n1915 ^ 1'b0 ;
  assign n3804 = n1644 ^ n974 ^ 1'b0 ;
  assign n3805 = n1212 & ~n3804 ;
  assign n3806 = n2849 & ~n3805 ;
  assign n3807 = n2028 & n3806 ;
  assign n3808 = n317 | n1294 ;
  assign n3809 = n994 & ~n3808 ;
  assign n3810 = n3809 ^ n2606 ^ 1'b0 ;
  assign n3811 = n1254 ^ n523 ^ n403 ;
  assign n3812 = n2358 ^ n1437 ^ n894 ;
  assign n3813 = n395 & ~n3812 ;
  assign n3814 = n3813 ^ n2234 ^ 1'b0 ;
  assign n3815 = ( n1066 & ~n1916 ) | ( n1066 & n3814 ) | ( ~n1916 & n3814 ) ;
  assign n3816 = ( n343 & ~n2648 ) | ( n343 & n3815 ) | ( ~n2648 & n3815 ) ;
  assign n3817 = ( n2301 & n3495 ) | ( n2301 & n3816 ) | ( n3495 & n3816 ) ;
  assign n3818 = ~n3811 & n3817 ;
  assign n3819 = ~n3810 & n3818 ;
  assign n3820 = n3792 ^ n3432 ^ n2847 ;
  assign n3821 = n2373 ^ n1438 ^ n1007 ;
  assign n3822 = n3821 ^ n3115 ^ 1'b0 ;
  assign n3823 = n3215 ^ n2153 ^ n1282 ;
  assign n3824 = n2950 ^ n2807 ^ n1901 ;
  assign n3825 = n2779 ^ n1428 ^ n1345 ;
  assign n3826 = n2925 ^ n400 ^ 1'b0 ;
  assign n3827 = ~n3825 & n3826 ;
  assign n3828 = ~n3322 & n3827 ;
  assign n3829 = n3824 & n3828 ;
  assign n3830 = n3047 & n3829 ;
  assign n3831 = ( n1352 & n1367 ) | ( n1352 & ~n1684 ) | ( n1367 & ~n1684 ) ;
  assign n3832 = n2392 ^ n2163 ^ 1'b0 ;
  assign n3833 = ~n2860 & n3832 ;
  assign n3834 = n3833 ^ n3291 ^ n521 ;
  assign n3835 = n3834 ^ n2405 ^ 1'b0 ;
  assign n3836 = ( x63 & n296 ) | ( x63 & n3531 ) | ( n296 & n3531 ) ;
  assign n3837 = ( n2433 & ~n2511 ) | ( n2433 & n3836 ) | ( ~n2511 & n3836 ) ;
  assign n3838 = ( n3831 & n3835 ) | ( n3831 & n3837 ) | ( n3835 & n3837 ) ;
  assign n3839 = n2754 | n3785 ;
  assign n3840 = n1112 ^ n801 ^ n149 ;
  assign n3841 = n1107 & ~n3840 ;
  assign n3842 = n3841 ^ n440 ^ 1'b0 ;
  assign n3843 = n3842 ^ n3161 ^ n1124 ;
  assign n3844 = x10 & ~n641 ;
  assign n3845 = n589 & n3844 ;
  assign n3846 = n545 | n2107 ;
  assign n3847 = n3845 & ~n3846 ;
  assign n3848 = n3847 ^ n2479 ^ 1'b0 ;
  assign n3851 = n1972 ^ n697 ^ n303 ;
  assign n3852 = n3851 ^ n2734 ^ n2669 ;
  assign n3849 = n811 & ~n957 ;
  assign n3850 = n3849 ^ n2747 ^ n1219 ;
  assign n3853 = n3852 ^ n3850 ^ n1994 ;
  assign n3854 = n1919 ^ n1318 ^ x36 ;
  assign n3855 = n2302 & n3854 ;
  assign n3856 = ( n175 & ~n1138 ) | ( n175 & n1334 ) | ( ~n1138 & n1334 ) ;
  assign n3857 = n3856 ^ n1060 ^ n418 ;
  assign n3858 = n2497 & ~n3857 ;
  assign n3859 = n420 & n2239 ;
  assign n3860 = n3859 ^ n799 ^ 1'b0 ;
  assign n3861 = ( n1238 & n3002 ) | ( n1238 & ~n3860 ) | ( n3002 & ~n3860 ) ;
  assign n3869 = n3845 ^ n1900 ^ n1229 ;
  assign n3868 = n2768 ^ n898 ^ n763 ;
  assign n3862 = ( x56 & n226 ) | ( x56 & ~n1659 ) | ( n226 & ~n1659 ) ;
  assign n3863 = n3241 ^ x119 ^ 1'b0 ;
  assign n3864 = n1669 & ~n3863 ;
  assign n3865 = n3862 & n3864 ;
  assign n3866 = ~n1253 & n3865 ;
  assign n3867 = ( ~n213 & n2901 ) | ( ~n213 & n3866 ) | ( n2901 & n3866 ) ;
  assign n3870 = n3869 ^ n3868 ^ n3867 ;
  assign n3871 = ( n455 & ~n944 ) | ( n455 & n2121 ) | ( ~n944 & n2121 ) ;
  assign n3872 = n651 & n3871 ;
  assign n3873 = n3783 ^ n1886 ^ 1'b0 ;
  assign n3874 = ~n3872 & n3873 ;
  assign n3875 = n3874 ^ n1941 ^ n1457 ;
  assign n3876 = ( n1563 & n2314 ) | ( n1563 & ~n3062 ) | ( n2314 & ~n3062 ) ;
  assign n3877 = ( n1465 & ~n3026 ) | ( n1465 & n3876 ) | ( ~n3026 & n3876 ) ;
  assign n3878 = n2919 & ~n3877 ;
  assign n3879 = ( n763 & ~n1264 ) | ( n763 & n2298 ) | ( ~n1264 & n2298 ) ;
  assign n3880 = n3879 ^ n2206 ^ n1633 ;
  assign n3881 = n3880 ^ n3611 ^ n205 ;
  assign n3882 = ~n3340 & n3881 ;
  assign n3885 = n2424 ^ n1635 ^ n823 ;
  assign n3883 = ( ~n1294 & n1394 ) | ( ~n1294 & n1744 ) | ( n1394 & n1744 ) ;
  assign n3884 = n2709 & n3883 ;
  assign n3886 = n3885 ^ n3884 ^ n1650 ;
  assign n3887 = n1325 ^ n796 ^ n525 ;
  assign n3888 = n3887 ^ n1399 ^ 1'b0 ;
  assign n3889 = ( ~n2665 & n3424 ) | ( ~n2665 & n3888 ) | ( n3424 & n3888 ) ;
  assign n3890 = ( ~n1486 & n1712 ) | ( ~n1486 & n2969 ) | ( n1712 & n2969 ) ;
  assign n3891 = ( n1167 & n2050 ) | ( n1167 & n2125 ) | ( n2050 & n2125 ) ;
  assign n3892 = ( n2674 & n3890 ) | ( n2674 & ~n3891 ) | ( n3890 & ~n3891 ) ;
  assign n3893 = n3840 ^ n1003 ^ n445 ;
  assign n3894 = n440 & ~n1485 ;
  assign n3895 = ( n840 & n3893 ) | ( n840 & ~n3894 ) | ( n3893 & ~n3894 ) ;
  assign n3896 = n2065 ^ n603 ^ 1'b0 ;
  assign n3897 = n957 | n3896 ;
  assign n3898 = n1210 | n3897 ;
  assign n3899 = n3898 ^ n1519 ^ n259 ;
  assign n3900 = ( n1790 & n2942 ) | ( n1790 & ~n3899 ) | ( n2942 & ~n3899 ) ;
  assign n3901 = n698 & ~n1059 ;
  assign n3902 = ( x62 & n1019 ) | ( x62 & n3901 ) | ( n1019 & n3901 ) ;
  assign n3903 = ~n1159 & n1560 ;
  assign n3904 = ~n3902 & n3903 ;
  assign n3905 = ( n1102 & n3900 ) | ( n1102 & n3904 ) | ( n3900 & n3904 ) ;
  assign n3906 = ( ~n1448 & n1579 ) | ( ~n1448 & n2754 ) | ( n1579 & n2754 ) ;
  assign n3907 = ( n683 & ~n750 ) | ( n683 & n1416 ) | ( ~n750 & n1416 ) ;
  assign n3908 = ( n787 & n1254 ) | ( n787 & ~n3907 ) | ( n1254 & ~n3907 ) ;
  assign n3909 = n1193 ^ n881 ^ 1'b0 ;
  assign n3910 = n294 & ~n3909 ;
  assign n3911 = n3910 ^ n3897 ^ n1592 ;
  assign n3912 = n1838 ^ n399 ^ 1'b0 ;
  assign n3913 = ( n1574 & ~n2281 ) | ( n1574 & n2891 ) | ( ~n2281 & n2891 ) ;
  assign n3914 = n3913 ^ n1954 ^ n236 ;
  assign n3915 = ( n176 & ~n3912 ) | ( n176 & n3914 ) | ( ~n3912 & n3914 ) ;
  assign n3916 = ( ~n3207 & n3911 ) | ( ~n3207 & n3915 ) | ( n3911 & n3915 ) ;
  assign n3917 = ( n485 & n3908 ) | ( n485 & ~n3916 ) | ( n3908 & ~n3916 ) ;
  assign n3918 = n3917 ^ n3765 ^ n1796 ;
  assign n3919 = ( n3073 & n3906 ) | ( n3073 & ~n3918 ) | ( n3906 & ~n3918 ) ;
  assign n3920 = n3430 ^ n1709 ^ 1'b0 ;
  assign n3921 = n3444 & n3920 ;
  assign n3922 = n3866 & n3921 ;
  assign n3923 = n3395 & ~n3922 ;
  assign n3924 = n3919 & n3923 ;
  assign n3927 = n1099 ^ n619 ^ n304 ;
  assign n3928 = ( n1874 & n2383 ) | ( n1874 & n3927 ) | ( n2383 & n3927 ) ;
  assign n3929 = ( n312 & ~n1449 ) | ( n312 & n3670 ) | ( ~n1449 & n3670 ) ;
  assign n3930 = n3388 & ~n3929 ;
  assign n3931 = ~n3928 & n3930 ;
  assign n3925 = n3438 ^ n3219 ^ n2772 ;
  assign n3926 = ( n2948 & n3053 ) | ( n2948 & ~n3925 ) | ( n3053 & ~n3925 ) ;
  assign n3932 = n3931 ^ n3926 ^ n1625 ;
  assign n3933 = n3265 ^ n1337 ^ 1'b0 ;
  assign n3934 = n2152 & n3933 ;
  assign n3935 = n3199 ^ n923 ^ n743 ;
  assign n3936 = n3934 & n3935 ;
  assign n3937 = n3936 ^ n1075 ^ 1'b0 ;
  assign n3938 = x119 & n3101 ;
  assign n3943 = n2454 & ~n2467 ;
  assign n3944 = n3943 ^ n1624 ^ 1'b0 ;
  assign n3941 = n748 & n2810 ;
  assign n3939 = n1339 & ~n1850 ;
  assign n3940 = n3939 ^ n2502 ^ 1'b0 ;
  assign n3942 = n3941 ^ n3940 ^ 1'b0 ;
  assign n3945 = n3944 ^ n3942 ^ n914 ;
  assign n3947 = ~n964 & n3857 ;
  assign n3946 = n2360 ^ n1991 ^ 1'b0 ;
  assign n3948 = n3947 ^ n3946 ^ n3210 ;
  assign n3949 = ( n831 & n1354 ) | ( n831 & n2674 ) | ( n1354 & n2674 ) ;
  assign n3950 = ( ~n432 & n1124 ) | ( ~n432 & n3949 ) | ( n1124 & n3949 ) ;
  assign n3951 = ( ~x83 & n1826 ) | ( ~x83 & n2934 ) | ( n1826 & n2934 ) ;
  assign n3952 = n382 & ~n3951 ;
  assign n3953 = n2398 & n3952 ;
  assign n3954 = n3953 ^ n827 ^ x115 ;
  assign n3955 = n2729 ^ n1798 ^ n486 ;
  assign n3956 = n609 | n1059 ;
  assign n3957 = n826 & ~n3956 ;
  assign n3958 = n2934 | n3957 ;
  assign n3959 = n3955 | n3958 ;
  assign n3960 = n1983 & n2790 ;
  assign n3961 = n3138 & n3960 ;
  assign n3962 = n2158 & n3961 ;
  assign n3963 = n3962 ^ n2169 ^ n1040 ;
  assign n3964 = ( n3954 & ~n3959 ) | ( n3954 & n3963 ) | ( ~n3959 & n3963 ) ;
  assign n3965 = n3130 ^ n2868 ^ n2236 ;
  assign n3966 = ( n540 & n1236 ) | ( n540 & n2814 ) | ( n1236 & n2814 ) ;
  assign n3967 = n1703 ^ n671 ^ n214 ;
  assign n3968 = n1669 & n3967 ;
  assign n3969 = n3968 ^ n410 ^ 1'b0 ;
  assign n3970 = ( n1661 & n3966 ) | ( n1661 & ~n3969 ) | ( n3966 & ~n3969 ) ;
  assign n3971 = n3198 ^ n1164 ^ n211 ;
  assign n3972 = n3971 ^ n2264 ^ 1'b0 ;
  assign n3973 = ~n1252 & n3972 ;
  assign n3974 = ~n1741 & n2585 ;
  assign n3975 = n3974 ^ n1157 ^ 1'b0 ;
  assign n3976 = n860 & ~n1024 ;
  assign n3977 = n3976 ^ n2157 ^ n1158 ;
  assign n3978 = x76 & ~n3977 ;
  assign n3979 = n3978 ^ n2728 ^ 1'b0 ;
  assign n3980 = n1975 & ~n3531 ;
  assign n3981 = n1778 & n3980 ;
  assign n3982 = ( n2669 & ~n3979 ) | ( n2669 & n3981 ) | ( ~n3979 & n3981 ) ;
  assign n3983 = n3975 & n3982 ;
  assign n3984 = ( ~x78 & n317 ) | ( ~x78 & n1494 ) | ( n317 & n1494 ) ;
  assign n3985 = n3984 ^ n928 ^ 1'b0 ;
  assign n3986 = n828 ^ n337 ^ 1'b0 ;
  assign n3987 = n3986 ^ n2285 ^ 1'b0 ;
  assign n3988 = n1989 & n3987 ;
  assign n3989 = ( n456 & n3985 ) | ( n456 & n3988 ) | ( n3985 & n3988 ) ;
  assign n3995 = x29 & n1100 ;
  assign n3996 = ( n1568 & ~n2541 ) | ( n1568 & n3995 ) | ( ~n2541 & n3995 ) ;
  assign n3990 = n2551 ^ n2080 ^ n184 ;
  assign n3991 = n3990 ^ n436 ^ n377 ;
  assign n3992 = n3991 ^ x16 ^ 1'b0 ;
  assign n3993 = n1947 & ~n3992 ;
  assign n3994 = n2396 & n3993 ;
  assign n3997 = n3996 ^ n3994 ^ 1'b0 ;
  assign n3998 = ( n966 & n1409 ) | ( n966 & n3790 ) | ( n1409 & n3790 ) ;
  assign n3999 = n3998 ^ n1356 ^ 1'b0 ;
  assign n4000 = n986 | n1778 ;
  assign n4001 = ~n1537 & n4000 ;
  assign n4002 = n2224 ^ n1255 ^ n321 ;
  assign n4003 = ( n2108 & n2712 ) | ( n2108 & n4002 ) | ( n2712 & n4002 ) ;
  assign n4004 = ( n345 & n3238 ) | ( n345 & ~n4003 ) | ( n3238 & ~n4003 ) ;
  assign n4005 = n4004 ^ n667 ^ 1'b0 ;
  assign n4006 = ~n1444 & n4005 ;
  assign n4008 = n146 | n600 ;
  assign n4007 = n1056 ^ n644 ^ 1'b0 ;
  assign n4009 = n4008 ^ n4007 ^ 1'b0 ;
  assign n4010 = n4006 & n4009 ;
  assign n4011 = ( ~n2251 & n2278 ) | ( ~n2251 & n4010 ) | ( n2278 & n4010 ) ;
  assign n4012 = n4011 ^ n2410 ^ n1826 ;
  assign n4013 = ( ~n1917 & n2176 ) | ( ~n1917 & n4012 ) | ( n2176 & n4012 ) ;
  assign n4014 = n1840 ^ n904 ^ n835 ;
  assign n4015 = n4014 ^ n2862 ^ n1978 ;
  assign n4016 = n3310 ^ n1510 ^ 1'b0 ;
  assign n4017 = n1162 & n4016 ;
  assign n4018 = n1663 & ~n3871 ;
  assign n4019 = n4018 ^ n2982 ^ 1'b0 ;
  assign n4020 = n4019 ^ n2848 ^ 1'b0 ;
  assign n4021 = ( n830 & n2441 ) | ( n830 & ~n2653 ) | ( n2441 & ~n2653 ) ;
  assign n4022 = n810 ^ x8 ^ 1'b0 ;
  assign n4023 = n828 & ~n4022 ;
  assign n4030 = n3591 ^ n1623 ^ n735 ;
  assign n4031 = n2255 & n4030 ;
  assign n4032 = n3338 & n4031 ;
  assign n4026 = n1171 & n2997 ;
  assign n4027 = n4026 ^ n305 ^ 1'b0 ;
  assign n4028 = n4027 ^ n3833 ^ n1425 ;
  assign n4029 = n3992 | n4028 ;
  assign n4024 = n1360 ^ n1309 ^ 1'b0 ;
  assign n4025 = ( x77 & n2052 ) | ( x77 & n4024 ) | ( n2052 & n4024 ) ;
  assign n4033 = n4032 ^ n4029 ^ n4025 ;
  assign n4034 = ~n1303 & n1875 ;
  assign n4035 = n4034 ^ n2155 ^ 1'b0 ;
  assign n4036 = ~n2952 & n3138 ;
  assign n4037 = n1377 & n4036 ;
  assign n4038 = n4037 ^ n3773 ^ 1'b0 ;
  assign n4039 = n2611 ^ n1122 ^ n667 ;
  assign n4040 = n2118 ^ n1931 ^ x2 ;
  assign n4041 = ( x12 & ~n285 ) | ( x12 & n1470 ) | ( ~n285 & n1470 ) ;
  assign n4042 = ~n1461 & n2771 ;
  assign n4043 = ~n1930 & n4042 ;
  assign n4044 = ( n1492 & ~n2912 ) | ( n1492 & n4043 ) | ( ~n2912 & n4043 ) ;
  assign n4045 = ( n496 & ~n2353 ) | ( n496 & n4044 ) | ( ~n2353 & n4044 ) ;
  assign n4046 = n4041 & n4045 ;
  assign n4047 = n4022 & n4046 ;
  assign n4048 = n4040 & n4047 ;
  assign n4049 = n902 | n1836 ;
  assign n4050 = n3667 & ~n4049 ;
  assign n4071 = n3770 ^ x69 ^ 1'b0 ;
  assign n4072 = n3173 & n4071 ;
  assign n4073 = n852 & n2301 ;
  assign n4074 = ( n1116 & n4072 ) | ( n1116 & ~n4073 ) | ( n4072 & ~n4073 ) ;
  assign n4051 = n2224 ^ n1684 ^ n1478 ;
  assign n4052 = n4051 ^ n1792 ^ n1707 ;
  assign n4053 = n1453 & n4052 ;
  assign n4054 = n2463 & ~n2915 ;
  assign n4055 = n697 & n4054 ;
  assign n4056 = n3215 ^ n2145 ^ n852 ;
  assign n4057 = n1305 ^ n1206 ^ 1'b0 ;
  assign n4058 = n4056 & ~n4057 ;
  assign n4059 = n3849 ^ n694 ^ 1'b0 ;
  assign n4060 = n3789 & n4059 ;
  assign n4061 = n475 & n4060 ;
  assign n4062 = ( n433 & ~n1034 ) | ( n433 & n1627 ) | ( ~n1034 & n1627 ) ;
  assign n4063 = n1365 | n4062 ;
  assign n4064 = n4061 & ~n4063 ;
  assign n4065 = n4064 ^ n2574 ^ 1'b0 ;
  assign n4066 = x126 & ~n4065 ;
  assign n4067 = ( n4055 & n4058 ) | ( n4055 & ~n4066 ) | ( n4058 & ~n4066 ) ;
  assign n4068 = n4053 | n4067 ;
  assign n4069 = n2504 | n4068 ;
  assign n4070 = n4069 ^ n3831 ^ n3501 ;
  assign n4075 = n4074 ^ n4070 ^ 1'b0 ;
  assign n4076 = ~n4050 & n4075 ;
  assign n4077 = ( ~n793 & n1709 ) | ( ~n793 & n2333 ) | ( n1709 & n2333 ) ;
  assign n4078 = n4077 ^ n2258 ^ n1369 ;
  assign n4079 = n4078 ^ n2147 ^ x102 ;
  assign n4080 = ( ~n342 & n1138 ) | ( ~n342 & n4079 ) | ( n1138 & n4079 ) ;
  assign n4081 = n4080 ^ x87 ^ 1'b0 ;
  assign n4082 = n4081 ^ n3942 ^ n591 ;
  assign n4084 = n799 & ~n900 ;
  assign n4085 = ~n389 & n4084 ;
  assign n4086 = ( n1205 & n1594 ) | ( n1205 & n4085 ) | ( n1594 & n4085 ) ;
  assign n4083 = ( n188 & n1524 ) | ( n188 & n3074 ) | ( n1524 & n3074 ) ;
  assign n4087 = n4086 ^ n4083 ^ n3019 ;
  assign n4107 = n3985 ^ n3174 ^ n2230 ;
  assign n4088 = n3450 ^ n779 ^ 1'b0 ;
  assign n4089 = n2817 ^ n203 ^ 1'b0 ;
  assign n4090 = ~n462 & n4089 ;
  assign n4091 = n4090 ^ x45 ^ 1'b0 ;
  assign n4092 = n397 & n4091 ;
  assign n4093 = ( n4002 & n4088 ) | ( n4002 & n4092 ) | ( n4088 & n4092 ) ;
  assign n4101 = n2181 ^ n374 ^ 1'b0 ;
  assign n4099 = x124 & n617 ;
  assign n4100 = n4099 ^ n1318 ^ 1'b0 ;
  assign n4102 = n4101 ^ n4100 ^ n2436 ;
  assign n4103 = n4102 ^ n2358 ^ n975 ;
  assign n4094 = n2882 & n3277 ;
  assign n4095 = n1562 & n4094 ;
  assign n4096 = ~n1488 & n3009 ;
  assign n4097 = n4095 & n4096 ;
  assign n4098 = ( n1728 & n2865 ) | ( n1728 & ~n4097 ) | ( n2865 & ~n4097 ) ;
  assign n4104 = n4103 ^ n4098 ^ n2832 ;
  assign n4105 = ( n3439 & n4093 ) | ( n3439 & ~n4104 ) | ( n4093 & ~n4104 ) ;
  assign n4106 = n1453 & n4105 ;
  assign n4108 = n4107 ^ n4106 ^ 1'b0 ;
  assign n4109 = ( ~n374 & n1523 ) | ( ~n374 & n1743 ) | ( n1523 & n1743 ) ;
  assign n4110 = n3931 ^ n1748 ^ n1371 ;
  assign n4111 = n2258 ^ n1274 ^ 1'b0 ;
  assign n4112 = n3814 | n4111 ;
  assign n4113 = x107 | n303 ;
  assign n4114 = ~n4112 & n4113 ;
  assign n4120 = n2514 ^ n1875 ^ n217 ;
  assign n4117 = n3293 ^ n1638 ^ n711 ;
  assign n4118 = n1468 & n3202 ;
  assign n4119 = n4117 & n4118 ;
  assign n4115 = n3099 ^ n1878 ^ 1'b0 ;
  assign n4116 = n1016 & ~n4115 ;
  assign n4121 = n4120 ^ n4119 ^ n4116 ;
  assign n4122 = n3256 ^ n1967 ^ n576 ;
  assign n4123 = ~n203 & n2141 ;
  assign n4124 = n4123 ^ n3659 ^ 1'b0 ;
  assign n4125 = n4124 ^ n3478 ^ x45 ;
  assign n4126 = n3924 ^ n2667 ^ 1'b0 ;
  assign n4127 = n913 | n2068 ;
  assign n4128 = n1854 & ~n4127 ;
  assign n4129 = n3684 ^ n3279 ^ n941 ;
  assign n4133 = n1317 ^ n131 ^ 1'b0 ;
  assign n4130 = ( n1125 & n3097 ) | ( n1125 & n3845 ) | ( n3097 & n3845 ) ;
  assign n4131 = ~n236 & n4130 ;
  assign n4132 = n4131 ^ n1595 ^ 1'b0 ;
  assign n4134 = n4133 ^ n4132 ^ n2311 ;
  assign n4135 = n1922 ^ n1490 ^ n587 ;
  assign n4136 = n4135 ^ n2662 ^ n385 ;
  assign n4137 = n3692 ^ n1902 ^ n979 ;
  assign n4138 = ( ~n443 & n3483 ) | ( ~n443 & n3591 ) | ( n3483 & n3591 ) ;
  assign n4139 = n2686 ^ n1042 ^ n526 ;
  assign n4140 = n3103 & n4139 ;
  assign n4141 = n1228 & n4140 ;
  assign n4143 = n2928 ^ n780 ^ n628 ;
  assign n4142 = ( n838 & ~n854 ) | ( n838 & n2551 ) | ( ~n854 & n2551 ) ;
  assign n4144 = n4143 ^ n4142 ^ n805 ;
  assign n4145 = n4144 ^ n3928 ^ n2868 ;
  assign n4146 = ~n428 & n1304 ;
  assign n4147 = n4146 ^ n1750 ^ 1'b0 ;
  assign n4148 = n4147 ^ n1601 ^ n459 ;
  assign n4149 = ( ~n2805 & n4145 ) | ( ~n2805 & n4148 ) | ( n4145 & n4148 ) ;
  assign n4155 = x52 & ~n216 ;
  assign n4156 = n4155 ^ n1362 ^ n1223 ;
  assign n4157 = ( n319 & n455 ) | ( n319 & ~n4156 ) | ( n455 & ~n4156 ) ;
  assign n4158 = n4157 ^ n2155 ^ 1'b0 ;
  assign n4159 = n2515 | n4158 ;
  assign n4160 = n3872 | n4159 ;
  assign n4161 = n3635 & ~n4160 ;
  assign n4151 = ( n972 & n1441 ) | ( n972 & n3068 ) | ( n1441 & n3068 ) ;
  assign n4150 = n1701 ^ n1048 ^ n581 ;
  assign n4152 = n4151 ^ n4150 ^ n2287 ;
  assign n4153 = n4078 ^ n3157 ^ n1017 ;
  assign n4154 = ( x105 & n4152 ) | ( x105 & ~n4153 ) | ( n4152 & ~n4153 ) ;
  assign n4162 = n4161 ^ n4154 ^ n2058 ;
  assign n4164 = n671 & n2036 ;
  assign n4165 = n4164 ^ n151 ^ 1'b0 ;
  assign n4166 = n1790 | n4165 ;
  assign n4167 = n2948 & ~n4166 ;
  assign n4163 = ~n1208 & n3126 ;
  assign n4168 = n4167 ^ n4163 ^ 1'b0 ;
  assign n4169 = n4168 ^ n2594 ^ 1'b0 ;
  assign n4170 = n2916 ^ n1727 ^ n336 ;
  assign n4171 = n3388 & n4170 ;
  assign n4172 = n4171 ^ n928 ^ 1'b0 ;
  assign n4177 = ( n850 & ~n1917 ) | ( n850 & n2919 ) | ( ~n1917 & n2919 ) ;
  assign n4178 = ( n476 & n1776 ) | ( n476 & n4177 ) | ( n1776 & n4177 ) ;
  assign n4175 = ( n214 & n487 ) | ( n214 & ~n2295 ) | ( n487 & ~n2295 ) ;
  assign n4173 = n1054 | n2669 ;
  assign n4174 = n2385 | n4173 ;
  assign n4176 = n4175 ^ n4174 ^ n1779 ;
  assign n4179 = n4178 ^ n4176 ^ n2975 ;
  assign n4180 = n1828 & n4179 ;
  assign n4181 = ~n687 & n4180 ;
  assign n4182 = n926 & n1543 ;
  assign n4183 = ~x1 & n4182 ;
  assign n4184 = n4183 ^ n406 ^ 1'b0 ;
  assign n4185 = n467 & n4184 ;
  assign n4186 = ~n374 & n4185 ;
  assign n4187 = n460 & ~n4186 ;
  assign n4188 = n2009 ^ n1367 ^ n380 ;
  assign n4189 = ~n867 & n2294 ;
  assign n4190 = ( n1101 & ~n4188 ) | ( n1101 & n4189 ) | ( ~n4188 & n4189 ) ;
  assign n4191 = ( ~n4041 & n4168 ) | ( ~n4041 & n4190 ) | ( n4168 & n4190 ) ;
  assign n4192 = ( ~n385 & n3571 ) | ( ~n385 & n4191 ) | ( n3571 & n4191 ) ;
  assign n4193 = ( n3072 & n3557 ) | ( n3072 & ~n4109 ) | ( n3557 & ~n4109 ) ;
  assign n4199 = n2955 ^ n2927 ^ n2111 ;
  assign n4195 = ( n2454 & n3034 ) | ( n2454 & ~n3113 ) | ( n3034 & ~n3113 ) ;
  assign n4196 = ( n2620 & n3032 ) | ( n2620 & ~n3798 ) | ( n3032 & ~n3798 ) ;
  assign n4197 = ~n1381 & n4196 ;
  assign n4198 = n4195 & ~n4197 ;
  assign n4200 = n4199 ^ n4198 ^ 1'b0 ;
  assign n4194 = x62 & n3490 ;
  assign n4201 = n4200 ^ n4194 ^ 1'b0 ;
  assign n4205 = ( n293 & n2050 ) | ( n293 & n2216 ) | ( n2050 & n2216 ) ;
  assign n4206 = n1366 & ~n2486 ;
  assign n4207 = n4205 & n4206 ;
  assign n4208 = n2818 ^ n883 ^ 1'b0 ;
  assign n4209 = n4207 | n4208 ;
  assign n4202 = ( n1326 & n2384 ) | ( n1326 & ~n2697 ) | ( n2384 & ~n2697 ) ;
  assign n4203 = n3145 ^ n3017 ^ 1'b0 ;
  assign n4204 = n4202 | n4203 ;
  assign n4210 = n4209 ^ n4204 ^ n1713 ;
  assign n4216 = n2949 ^ n1455 ^ n1258 ;
  assign n4214 = n3026 ^ n2972 ^ n563 ;
  assign n4215 = n1804 | n4214 ;
  assign n4217 = n4216 ^ n4215 ^ 1'b0 ;
  assign n4212 = ( n2009 & ~n2246 ) | ( n2009 & n2312 ) | ( ~n2246 & n2312 ) ;
  assign n4211 = ~n538 & n1382 ;
  assign n4213 = n4212 ^ n4211 ^ 1'b0 ;
  assign n4218 = n4217 ^ n4213 ^ n2694 ;
  assign n4219 = ( ~n667 & n4195 ) | ( ~n667 & n4218 ) | ( n4195 & n4218 ) ;
  assign n4220 = n3396 ^ n2394 ^ n525 ;
  assign n4221 = ( n233 & n4024 ) | ( n233 & n4220 ) | ( n4024 & n4220 ) ;
  assign n4222 = ( ~n164 & n3068 ) | ( ~n164 & n4221 ) | ( n3068 & n4221 ) ;
  assign n4223 = n1342 ^ x46 ^ 1'b0 ;
  assign n4224 = n1935 & ~n4223 ;
  assign n4225 = n4224 ^ n1829 ^ 1'b0 ;
  assign n4226 = n3321 & ~n3798 ;
  assign n4227 = ~n2450 & n4226 ;
  assign n4228 = ~n2425 & n4227 ;
  assign n4229 = ( n377 & n2792 ) | ( n377 & ~n4228 ) | ( n2792 & ~n4228 ) ;
  assign n4230 = ( x12 & x47 ) | ( x12 & n743 ) | ( x47 & n743 ) ;
  assign n4231 = n3387 ^ n3271 ^ n1282 ;
  assign n4232 = ( ~n2508 & n4230 ) | ( ~n2508 & n4231 ) | ( n4230 & n4231 ) ;
  assign n4233 = ( ~n853 & n1019 ) | ( ~n853 & n4232 ) | ( n1019 & n4232 ) ;
  assign n4238 = n178 & ~n989 ;
  assign n4239 = n4238 ^ n1052 ^ 1'b0 ;
  assign n4240 = n4239 ^ n3423 ^ 1'b0 ;
  assign n4241 = n3591 ^ n2870 ^ n131 ;
  assign n4242 = ( n1517 & n3845 ) | ( n1517 & n4241 ) | ( n3845 & n4241 ) ;
  assign n4243 = n4242 ^ n241 ^ 1'b0 ;
  assign n4244 = n4240 | n4243 ;
  assign n4234 = ~n1511 & n3814 ;
  assign n4235 = n1188 & ~n1801 ;
  assign n4236 = n841 & n4235 ;
  assign n4237 = n4234 | n4236 ;
  assign n4245 = n4244 ^ n4237 ^ 1'b0 ;
  assign n4251 = n1388 | n2320 ;
  assign n4252 = n4251 ^ n1481 ^ 1'b0 ;
  assign n4246 = n1317 & ~n3350 ;
  assign n4247 = n4246 ^ n3582 ^ n1159 ;
  assign n4248 = n1677 & ~n4247 ;
  assign n4249 = n4248 ^ n2423 ^ 1'b0 ;
  assign n4250 = n4249 ^ x27 ^ 1'b0 ;
  assign n4253 = n4252 ^ n4250 ^ n3155 ;
  assign n4254 = n4245 | n4253 ;
  assign n4255 = n937 & ~n4254 ;
  assign n4256 = ( n265 & n457 ) | ( n265 & ~n2885 ) | ( n457 & ~n2885 ) ;
  assign n4257 = n4256 ^ n1781 ^ n344 ;
  assign n4258 = n317 | n1403 ;
  assign n4259 = n4258 ^ n3350 ^ 1'b0 ;
  assign n4260 = n2898 | n4259 ;
  assign n4261 = n4260 ^ n1140 ^ 1'b0 ;
  assign n4262 = n3090 | n3835 ;
  assign n4263 = n3957 & ~n4262 ;
  assign n4264 = n1781 ^ n364 ^ 1'b0 ;
  assign n4265 = ( ~n804 & n3068 ) | ( ~n804 & n4264 ) | ( n3068 & n4264 ) ;
  assign n4266 = ~n3887 & n4265 ;
  assign n4267 = ~n1280 & n4266 ;
  assign n4268 = n3754 ^ n3607 ^ n2367 ;
  assign n4269 = ( n983 & n2370 ) | ( n983 & n2749 ) | ( n2370 & n2749 ) ;
  assign n4270 = n1533 | n4269 ;
  assign n4274 = ~n1246 & n1891 ;
  assign n4272 = n3955 ^ n3621 ^ n2040 ;
  assign n4271 = n3236 ^ n2063 ^ n1924 ;
  assign n4273 = n4272 ^ n4271 ^ n1876 ;
  assign n4275 = n4274 ^ n4273 ^ n346 ;
  assign n4276 = ( n1661 & n2676 ) | ( n1661 & n4275 ) | ( n2676 & n4275 ) ;
  assign n4277 = x120 & ~n880 ;
  assign n4278 = n608 & n4277 ;
  assign n4279 = n4278 ^ n1867 ^ 1'b0 ;
  assign n4280 = n4279 ^ n2279 ^ n1329 ;
  assign n4282 = n688 ^ n633 ^ n248 ;
  assign n4281 = n3158 ^ n1518 ^ x27 ;
  assign n4283 = n4282 ^ n4281 ^ n791 ;
  assign n4284 = n2355 ^ n1024 ^ 1'b0 ;
  assign n4290 = n1767 ^ n424 ^ 1'b0 ;
  assign n4291 = n2138 ^ n1708 ^ n861 ;
  assign n4292 = n4290 & ~n4291 ;
  assign n4293 = n4102 ^ n223 ^ 1'b0 ;
  assign n4294 = n4292 & n4293 ;
  assign n4285 = ( n317 & n1836 ) | ( n317 & ~n2166 ) | ( n1836 & ~n2166 ) ;
  assign n4286 = n4285 ^ n1301 ^ 1'b0 ;
  assign n4287 = ~n3430 & n4286 ;
  assign n4288 = n4287 ^ n3450 ^ n372 ;
  assign n4289 = ( ~n971 & n2110 ) | ( ~n971 & n4288 ) | ( n2110 & n4288 ) ;
  assign n4295 = n4294 ^ n4289 ^ 1'b0 ;
  assign n4296 = n4284 & n4295 ;
  assign n4297 = n256 | n659 ;
  assign n4298 = n3254 | n4297 ;
  assign n4303 = n3986 ^ n1481 ^ n1184 ;
  assign n4304 = n1568 ^ n1301 ^ n813 ;
  assign n4305 = ( ~n1470 & n4303 ) | ( ~n1470 & n4304 ) | ( n4303 & n4304 ) ;
  assign n4301 = n629 & ~n2179 ;
  assign n4302 = n4301 ^ n3792 ^ 1'b0 ;
  assign n4299 = n628 & ~n925 ;
  assign n4300 = n4299 ^ n511 ^ 1'b0 ;
  assign n4306 = n4305 ^ n4302 ^ n4300 ;
  assign n4307 = ( n1500 & n1785 ) | ( n1500 & ~n1887 ) | ( n1785 & ~n1887 ) ;
  assign n4308 = n4307 ^ n2103 ^ 1'b0 ;
  assign n4309 = n2819 ^ n2713 ^ 1'b0 ;
  assign n4310 = ~n2790 & n4309 ;
  assign n4311 = ~x21 & n1016 ;
  assign n4312 = n2552 | n4311 ;
  assign n4313 = n4310 | n4312 ;
  assign n4318 = n976 ^ n887 ^ n573 ;
  assign n4316 = ( n459 & n2622 ) | ( n459 & ~n2805 ) | ( n2622 & ~n2805 ) ;
  assign n4314 = n3387 ^ n3239 ^ n2781 ;
  assign n4315 = n2994 & n4314 ;
  assign n4317 = n4316 ^ n4315 ^ 1'b0 ;
  assign n4319 = n4318 ^ n4317 ^ n3707 ;
  assign n4320 = ( n434 & n2959 ) | ( n434 & n4165 ) | ( n2959 & n4165 ) ;
  assign n4321 = n2882 & n3817 ;
  assign n4322 = n4320 & n4321 ;
  assign n4324 = ~n661 & n3658 ;
  assign n4325 = n4324 ^ n602 ^ 1'b0 ;
  assign n4323 = ~n1112 & n3244 ;
  assign n4326 = n4325 ^ n4323 ^ 1'b0 ;
  assign n4327 = ( n1753 & n2761 ) | ( n1753 & ~n4326 ) | ( n2761 & ~n4326 ) ;
  assign n4328 = n434 | n3746 ;
  assign n4329 = n4328 ^ n2643 ^ 1'b0 ;
  assign n4330 = ( n197 & n1796 ) | ( n197 & n4329 ) | ( n1796 & n4329 ) ;
  assign n4331 = n4330 ^ n944 ^ n921 ;
  assign n4332 = n4331 ^ n2299 ^ n2140 ;
  assign n4333 = n2087 ^ n2034 ^ n1375 ;
  assign n4334 = n4191 & n4333 ;
  assign n4335 = ~n1989 & n4334 ;
  assign n4336 = ( ~n1269 & n1568 ) | ( ~n1269 & n3093 ) | ( n1568 & n3093 ) ;
  assign n4337 = n3361 & n4336 ;
  assign n4338 = n4337 ^ n1768 ^ 1'b0 ;
  assign n4339 = n473 & ~n4338 ;
  assign n4340 = ( ~n1274 & n1434 ) | ( ~n1274 & n2646 ) | ( n1434 & n2646 ) ;
  assign n4341 = n1389 ^ n1290 ^ n313 ;
  assign n4342 = n339 & ~n4341 ;
  assign n4343 = ( n251 & ~n1718 ) | ( n251 & n4342 ) | ( ~n1718 & n4342 ) ;
  assign n4344 = n4223 ^ n2908 ^ n1064 ;
  assign n4345 = ( n846 & n4343 ) | ( n846 & ~n4344 ) | ( n4343 & ~n4344 ) ;
  assign n4353 = ( n357 & ~n1185 ) | ( n357 & n1253 ) | ( ~n1185 & n1253 ) ;
  assign n4346 = ( ~n234 & n878 ) | ( ~n234 & n1305 ) | ( n878 & n1305 ) ;
  assign n4347 = n4346 ^ n2794 ^ 1'b0 ;
  assign n4348 = ~n1712 & n4347 ;
  assign n4349 = n785 ^ n723 ^ 1'b0 ;
  assign n4350 = ( n791 & n1568 ) | ( n791 & ~n4349 ) | ( n1568 & ~n4349 ) ;
  assign n4351 = n4348 & n4350 ;
  assign n4352 = n4351 ^ n2652 ^ 1'b0 ;
  assign n4354 = n4353 ^ n4352 ^ n626 ;
  assign n4355 = n1719 | n2817 ;
  assign n4356 = n4354 & ~n4355 ;
  assign n4357 = ( x64 & n2982 ) | ( x64 & ~n3682 ) | ( n2982 & ~n3682 ) ;
  assign n4358 = ( ~n541 & n1938 ) | ( ~n541 & n2287 ) | ( n1938 & n2287 ) ;
  assign n4359 = ( n1749 & n4357 ) | ( n1749 & n4358 ) | ( n4357 & n4358 ) ;
  assign n4360 = ( ~x65 & n984 ) | ( ~x65 & n4129 ) | ( n984 & n4129 ) ;
  assign n4361 = ( n1916 & ~n2543 ) | ( n1916 & n3293 ) | ( ~n2543 & n3293 ) ;
  assign n4362 = n4361 ^ n3326 ^ n2028 ;
  assign n4363 = ( ~n1723 & n2928 ) | ( ~n1723 & n4362 ) | ( n2928 & n4362 ) ;
  assign n4364 = ~n1322 & n2401 ;
  assign n4365 = ~x8 & n4364 ;
  assign n4366 = n4365 ^ n2357 ^ n925 ;
  assign n4367 = n4366 ^ n4088 ^ n2606 ;
  assign n4368 = n4367 ^ n2863 ^ 1'b0 ;
  assign n4369 = n2823 & ~n4368 ;
  assign n4375 = n2258 ^ n1709 ^ 1'b0 ;
  assign n4370 = n658 & n1025 ;
  assign n4371 = n4370 ^ n900 ^ 1'b0 ;
  assign n4372 = n913 ^ n521 ^ 1'b0 ;
  assign n4373 = ~n2545 & n4372 ;
  assign n4374 = ( n1378 & n4371 ) | ( n1378 & ~n4373 ) | ( n4371 & ~n4373 ) ;
  assign n4376 = n4375 ^ n4374 ^ x111 ;
  assign n4377 = n1158 ^ n791 ^ n306 ;
  assign n4378 = ( n2197 & n4143 ) | ( n2197 & ~n4377 ) | ( n4143 & ~n4377 ) ;
  assign n4379 = n2321 & n4378 ;
  assign n4380 = n783 & n4379 ;
  assign n4381 = ( n3430 & n4376 ) | ( n3430 & n4380 ) | ( n4376 & n4380 ) ;
  assign n4382 = ~n160 & n1286 ;
  assign n4383 = n4382 ^ n2727 ^ 1'b0 ;
  assign n4384 = n4383 ^ n2636 ^ n1833 ;
  assign n4385 = n4384 ^ n857 ^ n582 ;
  assign n4386 = n2510 ^ n1818 ^ 1'b0 ;
  assign n4387 = ( x89 & ~n2928 ) | ( x89 & n4386 ) | ( ~n2928 & n4386 ) ;
  assign n4388 = n4362 ^ x7 ^ 1'b0 ;
  assign n4389 = n4388 ^ n2763 ^ n1374 ;
  assign n4390 = n4389 ^ n275 ^ x4 ;
  assign n4391 = ~n1195 & n2703 ;
  assign n4392 = n4391 ^ n2512 ^ 1'b0 ;
  assign n4393 = n3151 | n3265 ;
  assign n4394 = n4392 | n4393 ;
  assign n4395 = ~n812 & n2463 ;
  assign n4396 = n4395 ^ n1129 ^ 1'b0 ;
  assign n4397 = n3571 | n4396 ;
  assign n4398 = n4397 ^ n2930 ^ 1'b0 ;
  assign n4399 = n1133 & n2079 ;
  assign n4400 = ( n963 & ~n1004 ) | ( n963 & n4399 ) | ( ~n1004 & n4399 ) ;
  assign n4401 = ( ~n135 & n2122 ) | ( ~n135 & n2159 ) | ( n2122 & n2159 ) ;
  assign n4402 = n4400 & ~n4401 ;
  assign n4403 = n4402 ^ x125 ^ x21 ;
  assign n4404 = n4403 ^ n3005 ^ n2351 ;
  assign n4405 = ~n146 & n1405 ;
  assign n4406 = n2739 ^ n2500 ^ n1366 ;
  assign n4407 = n4406 ^ n1518 ^ 1'b0 ;
  assign n4408 = n4405 | n4407 ;
  assign n4409 = n754 & ~n4049 ;
  assign n4410 = n1072 & n4409 ;
  assign n4411 = n1610 | n4410 ;
  assign n4412 = n4411 ^ n3788 ^ 1'b0 ;
  assign n4413 = ( n677 & n2044 ) | ( n677 & n4336 ) | ( n2044 & n4336 ) ;
  assign n4414 = n3175 ^ n1749 ^ n623 ;
  assign n4415 = n3347 & ~n4414 ;
  assign n4416 = n4415 ^ n2970 ^ n1990 ;
  assign n4417 = ( ~n723 & n4413 ) | ( ~n723 & n4416 ) | ( n4413 & n4416 ) ;
  assign n4418 = ( n1465 & n4412 ) | ( n1465 & ~n4417 ) | ( n4412 & ~n4417 ) ;
  assign n4419 = n1183 | n3203 ;
  assign n4420 = n1761 | n4419 ;
  assign n4421 = n2073 & ~n3905 ;
  assign n4422 = ( n697 & n4420 ) | ( n697 & ~n4421 ) | ( n4420 & ~n4421 ) ;
  assign n4423 = x39 & ~n2817 ;
  assign n4424 = n4423 ^ n436 ^ 1'b0 ;
  assign n4425 = n4424 ^ n2457 ^ n399 ;
  assign n4426 = n2236 & ~n4425 ;
  assign n4427 = ~n2364 & n4426 ;
  assign n4429 = n4133 ^ n2693 ^ x35 ;
  assign n4428 = n1519 & ~n4201 ;
  assign n4430 = n4429 ^ n4428 ^ 1'b0 ;
  assign n4431 = n716 & ~n2144 ;
  assign n4433 = ( n538 & ~n1870 ) | ( n538 & n2015 ) | ( ~n1870 & n2015 ) ;
  assign n4432 = ~n1599 & n2876 ;
  assign n4434 = n4433 ^ n4432 ^ 1'b0 ;
  assign n4435 = ~n706 & n4434 ;
  assign n4436 = ( n440 & n1570 ) | ( n440 & ~n3122 ) | ( n1570 & ~n3122 ) ;
  assign n4437 = n881 ^ n558 ^ x72 ;
  assign n4438 = n4437 ^ n3957 ^ n1516 ;
  assign n4439 = n1934 ^ n592 ^ 1'b0 ;
  assign n4440 = ~n4438 & n4439 ;
  assign n4441 = n1400 & n3849 ;
  assign n4444 = n472 ^ x51 ^ 1'b0 ;
  assign n4445 = n4444 ^ n2328 ^ 1'b0 ;
  assign n4442 = ~n2146 & n3498 ;
  assign n4443 = n2908 & n4442 ;
  assign n4446 = n4445 ^ n4443 ^ 1'b0 ;
  assign n4447 = ( n1750 & ~n4441 ) | ( n1750 & n4446 ) | ( ~n4441 & n4446 ) ;
  assign n4448 = n4447 ^ n1535 ^ 1'b0 ;
  assign n4449 = n4448 ^ n2652 ^ n639 ;
  assign n4453 = ~n207 & n1340 ;
  assign n4450 = n2282 ^ n420 ^ 1'b0 ;
  assign n4451 = n463 | n4450 ;
  assign n4452 = ( n588 & ~n2506 ) | ( n588 & n4451 ) | ( ~n2506 & n4451 ) ;
  assign n4454 = n4453 ^ n4452 ^ 1'b0 ;
  assign n4455 = ( n2170 & n4234 ) | ( n2170 & n4454 ) | ( n4234 & n4454 ) ;
  assign n4456 = n3165 ^ n1503 ^ 1'b0 ;
  assign n4457 = ( n1490 & ~n1630 ) | ( n1490 & n4456 ) | ( ~n1630 & n4456 ) ;
  assign n4458 = n4455 | n4457 ;
  assign n4463 = n1021 & ~n3682 ;
  assign n4464 = n2970 & n4463 ;
  assign n4465 = ( ~x41 & n188 ) | ( ~x41 & n4464 ) | ( n188 & n4464 ) ;
  assign n4459 = n165 | n2406 ;
  assign n4460 = n4459 ^ n1339 ^ 1'b0 ;
  assign n4461 = n1792 | n4460 ;
  assign n4462 = n3712 & ~n4461 ;
  assign n4466 = n4465 ^ n4462 ^ 1'b0 ;
  assign n4467 = n3906 ^ n1386 ^ 1'b0 ;
  assign n4468 = n4467 ^ n1734 ^ 1'b0 ;
  assign n4473 = ~n343 & n1166 ;
  assign n4474 = n1165 | n4473 ;
  assign n4475 = ( n1614 & ~n2450 ) | ( n1614 & n4474 ) | ( ~n2450 & n4474 ) ;
  assign n4472 = n349 & ~n2739 ;
  assign n4476 = n4475 ^ n4472 ^ 1'b0 ;
  assign n4469 = n2969 | n3446 ;
  assign n4470 = n4469 ^ n2972 ^ n2695 ;
  assign n4471 = n695 & ~n4470 ;
  assign n4477 = n4476 ^ n4471 ^ 1'b0 ;
  assign n4478 = n3025 ^ n2230 ^ n1372 ;
  assign n4479 = n4478 ^ n2011 ^ 1'b0 ;
  assign n4480 = n775 & ~n4479 ;
  assign n4481 = ( n242 & ~n247 ) | ( n242 & n4480 ) | ( ~n247 & n4480 ) ;
  assign n4482 = n4481 ^ n2210 ^ n1350 ;
  assign n4485 = n1046 ^ n207 ^ x49 ;
  assign n4483 = n831 | n1555 ;
  assign n4484 = ~x90 & n4483 ;
  assign n4486 = n4485 ^ n4484 ^ n1186 ;
  assign n4487 = n3598 | n4486 ;
  assign n4492 = ( n472 & n986 ) | ( n472 & n1360 ) | ( n986 & n1360 ) ;
  assign n4488 = ( n163 & n909 ) | ( n163 & n1034 ) | ( n909 & n1034 ) ;
  assign n4489 = n1714 ^ n1542 ^ n1018 ;
  assign n4490 = ( ~n1057 & n4488 ) | ( ~n1057 & n4489 ) | ( n4488 & n4489 ) ;
  assign n4491 = ( n581 & n2599 ) | ( n581 & n4490 ) | ( n2599 & n4490 ) ;
  assign n4493 = n4492 ^ n4491 ^ 1'b0 ;
  assign n4496 = ( n791 & n1203 ) | ( n791 & n1684 ) | ( n1203 & n1684 ) ;
  assign n4494 = n572 & n3446 ;
  assign n4495 = n4494 ^ n2545 ^ x122 ;
  assign n4497 = n4496 ^ n4495 ^ 1'b0 ;
  assign n4498 = n375 | n1176 ;
  assign n4499 = n4498 ^ n3902 ^ 1'b0 ;
  assign n4500 = ( n2410 & n4497 ) | ( n2410 & n4499 ) | ( n4497 & n4499 ) ;
  assign n4509 = ~n900 & n2267 ;
  assign n4510 = n4509 ^ n1274 ^ 1'b0 ;
  assign n4501 = n4062 | n4285 ;
  assign n4502 = n3023 | n4501 ;
  assign n4503 = ( n1474 & n2195 ) | ( n1474 & n4502 ) | ( n2195 & n4502 ) ;
  assign n4504 = x80 & ~n2410 ;
  assign n4505 = n4504 ^ n1633 ^ n1410 ;
  assign n4506 = n4505 ^ n2228 ^ 1'b0 ;
  assign n4507 = n4503 & ~n4506 ;
  assign n4508 = n2400 & n4507 ;
  assign n4511 = n4510 ^ n4508 ^ n1219 ;
  assign n4512 = x85 & n4511 ;
  assign n4513 = n4512 ^ n807 ^ 1'b0 ;
  assign n4514 = n2644 ^ n782 ^ n266 ;
  assign n4515 = n4514 ^ n328 ^ 1'b0 ;
  assign n4516 = n1135 ^ n451 ^ 1'b0 ;
  assign n4517 = ~n2744 & n4516 ;
  assign n4518 = n3905 ^ n2971 ^ 1'b0 ;
  assign n4519 = ( n955 & ~n1120 ) | ( n955 & n1436 ) | ( ~n1120 & n1436 ) ;
  assign n4520 = n1651 ^ n926 ^ n614 ;
  assign n4521 = ( n604 & ~n700 ) | ( n604 & n4520 ) | ( ~n700 & n4520 ) ;
  assign n4522 = n3439 ^ n2362 ^ 1'b0 ;
  assign n4523 = n2753 & ~n4522 ;
  assign n4524 = ( ~n2059 & n4521 ) | ( ~n2059 & n4523 ) | ( n4521 & n4523 ) ;
  assign n4525 = ( ~n411 & n4519 ) | ( ~n411 & n4524 ) | ( n4519 & n4524 ) ;
  assign n4534 = n2302 & ~n2849 ;
  assign n4535 = n441 & ~n4534 ;
  assign n4536 = n4535 ^ n2708 ^ 1'b0 ;
  assign n4528 = n1785 ^ n1701 ^ n180 ;
  assign n4526 = n3040 & n3759 ;
  assign n4527 = n2759 & n4526 ;
  assign n4529 = n4528 ^ n4527 ^ n1190 ;
  assign n4530 = ( ~n2431 & n3876 ) | ( ~n2431 & n4529 ) | ( n3876 & n4529 ) ;
  assign n4531 = ( x62 & ~n424 ) | ( x62 & n3333 ) | ( ~n424 & n3333 ) ;
  assign n4532 = n4531 ^ n696 ^ 1'b0 ;
  assign n4533 = n4530 | n4532 ;
  assign n4537 = n4536 ^ n4533 ^ 1'b0 ;
  assign n4538 = n3219 ^ n3181 ^ n2524 ;
  assign n4539 = ( n696 & n2504 ) | ( n696 & n4538 ) | ( n2504 & n4538 ) ;
  assign n4547 = ( n207 & n1449 ) | ( n207 & ~n3084 ) | ( n1449 & ~n3084 ) ;
  assign n4540 = ( n495 & n877 ) | ( n495 & ~n3354 ) | ( n877 & ~n3354 ) ;
  assign n4541 = ( n3544 & ~n4406 ) | ( n3544 & n4540 ) | ( ~n4406 & n4540 ) ;
  assign n4542 = n453 & n4383 ;
  assign n4543 = n4542 ^ n2920 ^ 1'b0 ;
  assign n4544 = n4543 ^ n4373 ^ n1320 ;
  assign n4545 = ( n820 & ~n4541 ) | ( n820 & n4544 ) | ( ~n4541 & n4544 ) ;
  assign n4546 = n2849 & n4545 ;
  assign n4548 = n4547 ^ n4546 ^ 1'b0 ;
  assign n4564 = n1380 ^ n1035 ^ n697 ;
  assign n4563 = n1694 ^ n1361 ^ n1262 ;
  assign n4565 = n4564 ^ n4563 ^ n3711 ;
  assign n4566 = ( n325 & n1072 ) | ( n325 & ~n3061 ) | ( n1072 & ~n3061 ) ;
  assign n4567 = n4566 ^ n1321 ^ 1'b0 ;
  assign n4568 = ~n4565 & n4567 ;
  assign n4562 = n2471 ^ n604 ^ 1'b0 ;
  assign n4556 = n2771 ^ n2025 ^ n164 ;
  assign n4557 = ( ~x0 & n201 ) | ( ~x0 & n1971 ) | ( n201 & n1971 ) ;
  assign n4558 = n4557 ^ n2644 ^ 1'b0 ;
  assign n4559 = n4556 & n4558 ;
  assign n4550 = n593 ^ n145 ^ 1'b0 ;
  assign n4551 = n967 & n4550 ;
  assign n4552 = n688 ^ x3 ^ 1'b0 ;
  assign n4553 = ~n1895 & n4552 ;
  assign n4554 = n4551 & n4553 ;
  assign n4555 = n4554 ^ n3788 ^ 1'b0 ;
  assign n4549 = ( n1349 & ~n2677 ) | ( n1349 & n2763 ) | ( ~n2677 & n2763 ) ;
  assign n4560 = n4559 ^ n4555 ^ n4549 ;
  assign n4561 = ( ~n805 & n3982 ) | ( ~n805 & n4560 ) | ( n3982 & n4560 ) ;
  assign n4569 = n4568 ^ n4562 ^ n4561 ;
  assign n4570 = n2762 ^ n1112 ^ 1'b0 ;
  assign n4571 = n4570 ^ n1798 ^ 1'b0 ;
  assign n4572 = n4360 | n4475 ;
  assign n4573 = n4572 ^ n778 ^ 1'b0 ;
  assign n4574 = n3279 ^ n2306 ^ x67 ;
  assign n4575 = n4574 ^ n620 ^ n205 ;
  assign n4576 = n4575 ^ n4067 ^ n3638 ;
  assign n4577 = n1817 & n3907 ;
  assign n4578 = ~n2126 & n3125 ;
  assign n4579 = ~n4577 & n4578 ;
  assign n4580 = n1206 ^ n417 ^ 1'b0 ;
  assign n4581 = ( n891 & n2369 ) | ( n891 & ~n2426 ) | ( n2369 & ~n2426 ) ;
  assign n4582 = n2246 | n4581 ;
  assign n4583 = n4582 ^ n1741 ^ 1'b0 ;
  assign n4584 = n4583 ^ n4551 ^ n1569 ;
  assign n4585 = ( n4579 & n4580 ) | ( n4579 & ~n4584 ) | ( n4580 & ~n4584 ) ;
  assign n4586 = n4585 ^ n581 ^ 1'b0 ;
  assign n4587 = n2900 ^ n496 ^ x60 ;
  assign n4588 = n1228 | n3269 ;
  assign n4590 = ( n139 & ~n187 ) | ( n139 & n1168 ) | ( ~n187 & n1168 ) ;
  assign n4591 = ( n1424 & n1732 ) | ( n1424 & n2816 ) | ( n1732 & n2816 ) ;
  assign n4592 = ( n285 & ~n4590 ) | ( n285 & n4591 ) | ( ~n4590 & n4591 ) ;
  assign n4589 = n1859 ^ n1342 ^ n1015 ;
  assign n4593 = n4592 ^ n4589 ^ n2548 ;
  assign n4594 = n877 | n4593 ;
  assign n4595 = n4588 | n4594 ;
  assign n4596 = n444 | n784 ;
  assign n4597 = n4596 ^ n1290 ^ 1'b0 ;
  assign n4598 = n4597 ^ n2662 ^ n2200 ;
  assign n4599 = n4598 ^ n805 ^ 1'b0 ;
  assign n4600 = n4595 & ~n4599 ;
  assign n4601 = ( ~n2912 & n4587 ) | ( ~n2912 & n4600 ) | ( n4587 & n4600 ) ;
  assign n4606 = ( n611 & n676 ) | ( n611 & n1628 ) | ( n676 & n1628 ) ;
  assign n4607 = n4606 ^ n4271 ^ n1671 ;
  assign n4608 = ( x116 & n1433 ) | ( x116 & ~n4607 ) | ( n1433 & ~n4607 ) ;
  assign n4602 = ( n1238 & ~n1366 ) | ( n1238 & n2779 ) | ( ~n1366 & n2779 ) ;
  assign n4603 = n1107 & ~n4602 ;
  assign n4604 = n4603 ^ n409 ^ 1'b0 ;
  assign n4605 = n4604 ^ n3254 ^ n256 ;
  assign n4609 = n4608 ^ n4605 ^ n305 ;
  assign n4610 = n2614 ^ n2459 ^ n1621 ;
  assign n4611 = n3138 ^ n926 ^ x80 ;
  assign n4612 = n1645 & ~n4611 ;
  assign n4613 = n4610 & ~n4612 ;
  assign n4614 = n2209 & n4613 ;
  assign n4615 = n4523 ^ n2115 ^ 1'b0 ;
  assign n4622 = n1799 ^ n1290 ^ n643 ;
  assign n4623 = ( n545 & ~n3736 ) | ( n545 & n4622 ) | ( ~n3736 & n4622 ) ;
  assign n4621 = x113 & ~n3929 ;
  assign n4624 = n4623 ^ n4621 ^ 1'b0 ;
  assign n4616 = n2262 ^ n1174 ^ 1'b0 ;
  assign n4617 = n336 | n4616 ;
  assign n4618 = n410 & ~n2066 ;
  assign n4619 = ~n3145 & n4618 ;
  assign n4620 = n4617 | n4619 ;
  assign n4625 = n4624 ^ n4620 ^ 1'b0 ;
  assign n4640 = ( x94 & ~n1650 ) | ( x94 & n3646 ) | ( ~n1650 & n3646 ) ;
  assign n4631 = n3330 ^ n2449 ^ 1'b0 ;
  assign n4632 = n1543 & ~n4631 ;
  assign n4634 = n1360 ^ n255 ^ n169 ;
  assign n4635 = n188 ^ x42 ^ 1'b0 ;
  assign n4636 = ~n4634 & n4635 ;
  assign n4633 = n4290 ^ n902 ^ x113 ;
  assign n4637 = n4636 ^ n4633 ^ n2008 ;
  assign n4638 = n4632 & n4637 ;
  assign n4639 = ~n1819 & n4638 ;
  assign n4626 = ( ~n571 & n1982 ) | ( ~n571 & n2770 ) | ( n1982 & n2770 ) ;
  assign n4627 = n3456 ^ n2121 ^ n289 ;
  assign n4628 = n4371 ^ n992 ^ n562 ;
  assign n4629 = n709 & n4628 ;
  assign n4630 = ( n4626 & n4627 ) | ( n4626 & ~n4629 ) | ( n4627 & ~n4629 ) ;
  assign n4641 = n4640 ^ n4639 ^ n4630 ;
  assign n4642 = n4302 ^ n2216 ^ n372 ;
  assign n4643 = n3770 ^ n846 ^ 1'b0 ;
  assign n4644 = n3123 | n4643 ;
  assign n4645 = ( n663 & n1199 ) | ( n663 & n1440 ) | ( n1199 & n1440 ) ;
  assign n4646 = n4007 ^ n3438 ^ 1'b0 ;
  assign n4647 = ( x42 & n4645 ) | ( x42 & ~n4646 ) | ( n4645 & ~n4646 ) ;
  assign n4648 = n305 & n2779 ;
  assign n4649 = ~n1084 & n4648 ;
  assign n4652 = ( n523 & n1715 ) | ( n523 & ~n2689 ) | ( n1715 & ~n2689 ) ;
  assign n4653 = n4652 ^ n2097 ^ n1990 ;
  assign n4650 = n3319 ^ n1567 ^ x87 ;
  assign n4651 = n4650 ^ n2886 ^ n388 ;
  assign n4654 = n4653 ^ n4651 ^ n3740 ;
  assign n4655 = ( n2146 & ~n4649 ) | ( n2146 & n4654 ) | ( ~n4649 & n4654 ) ;
  assign n4656 = ~n1240 & n1611 ;
  assign n4657 = n4656 ^ n3651 ^ n1698 ;
  assign n4658 = n3573 & ~n3904 ;
  assign n4659 = n4658 ^ n1451 ^ 1'b0 ;
  assign n4660 = n4659 ^ n2801 ^ x122 ;
  assign n4661 = n2047 ^ n305 ^ 1'b0 ;
  assign n4662 = n332 & ~n4661 ;
  assign n4663 = ( ~x68 & n2122 ) | ( ~x68 & n4662 ) | ( n2122 & n4662 ) ;
  assign n4664 = n4663 ^ n4291 ^ n1361 ;
  assign n4665 = n2031 ^ n139 ^ 1'b0 ;
  assign n4666 = n3136 & ~n4665 ;
  assign n4670 = n1286 ^ n967 ^ n885 ;
  assign n4669 = n4055 ^ n2514 ^ n2498 ;
  assign n4667 = ( n1911 & n2018 ) | ( n1911 & n2625 ) | ( n2018 & n2625 ) ;
  assign n4668 = ( n1323 & n2476 ) | ( n1323 & n4667 ) | ( n2476 & n4667 ) ;
  assign n4671 = n4670 ^ n4669 ^ n4668 ;
  assign n4675 = n2256 ^ n2147 ^ 1'b0 ;
  assign n4676 = n4675 ^ n1283 ^ n851 ;
  assign n4677 = ( x59 & ~n4044 ) | ( x59 & n4676 ) | ( ~n4044 & n4676 ) ;
  assign n4672 = n814 & n1468 ;
  assign n4673 = n4672 ^ n216 ^ 1'b0 ;
  assign n4674 = ( ~n1465 & n4113 ) | ( ~n1465 & n4673 ) | ( n4113 & n4673 ) ;
  assign n4678 = n4677 ^ n4674 ^ n1617 ;
  assign n4679 = ( n616 & ~n4671 ) | ( n616 & n4678 ) | ( ~n4671 & n4678 ) ;
  assign n4680 = ( n694 & n3247 ) | ( n694 & ~n3772 ) | ( n3247 & ~n3772 ) ;
  assign n4681 = ( n156 & ~n2202 ) | ( n156 & n2813 ) | ( ~n2202 & n2813 ) ;
  assign n4682 = ~n226 & n3582 ;
  assign n4683 = ~n4681 & n4682 ;
  assign n4684 = n434 ^ n399 ^ 1'b0 ;
  assign n4685 = n2895 & n4684 ;
  assign n4686 = ~n447 & n585 ;
  assign n4687 = ~n1410 & n4686 ;
  assign n4688 = ~n1748 & n2457 ;
  assign n4689 = n475 & n4688 ;
  assign n4690 = n4689 ^ n3849 ^ n880 ;
  assign n4691 = n1795 | n4690 ;
  assign n4692 = n4687 & ~n4691 ;
  assign n4693 = n4692 ^ n3462 ^ n843 ;
  assign n4694 = n4685 & n4693 ;
  assign n4695 = n3800 ^ n513 ^ 1'b0 ;
  assign n4696 = n4376 & n4695 ;
  assign n4697 = n4696 ^ n3622 ^ n1954 ;
  assign n4698 = n1951 ^ n331 ^ 1'b0 ;
  assign n4699 = n4150 | n4698 ;
  assign n4700 = x50 & n1298 ;
  assign n4701 = n609 & n4700 ;
  assign n4702 = ( n339 & ~n2464 ) | ( n339 & n4701 ) | ( ~n2464 & n4701 ) ;
  assign n4703 = n1102 | n4702 ;
  assign n4704 = n4703 ^ n2452 ^ 1'b0 ;
  assign n4705 = n984 & n2811 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4707 = ( ~n4134 & n4699 ) | ( ~n4134 & n4706 ) | ( n4699 & n4706 ) ;
  assign n4708 = n2785 ^ n156 ^ 1'b0 ;
  assign n4709 = ~n3408 & n4708 ;
  assign n4710 = n2102 & n4709 ;
  assign n4711 = ( ~n1157 & n3078 ) | ( ~n1157 & n3485 ) | ( n3078 & n3485 ) ;
  assign n4712 = n4711 ^ n4338 ^ n2155 ;
  assign n4713 = n782 & ~n1207 ;
  assign n4714 = ~n3319 & n4317 ;
  assign n4715 = ~n4713 & n4714 ;
  assign n4716 = n3322 ^ n129 ^ 1'b0 ;
  assign n4717 = n4453 & ~n4716 ;
  assign n4718 = n2151 | n4671 ;
  assign n4719 = n4717 | n4718 ;
  assign n4720 = ( x56 & n718 ) | ( x56 & n3437 ) | ( n718 & n3437 ) ;
  assign n4721 = ( x116 & n1470 ) | ( x116 & n3306 ) | ( n1470 & n3306 ) ;
  assign n4722 = ( n1428 & n2034 ) | ( n1428 & ~n2054 ) | ( n2034 & ~n2054 ) ;
  assign n4723 = ( n1700 & n4721 ) | ( n1700 & n4722 ) | ( n4721 & n4722 ) ;
  assign n4725 = x47 & n230 ;
  assign n4724 = n4566 ^ n434 ^ 1'b0 ;
  assign n4726 = n4725 ^ n4724 ^ n899 ;
  assign n4727 = ~n2193 & n2717 ;
  assign n4728 = n3437 ^ n1775 ^ n1331 ;
  assign n4729 = n2394 & n4728 ;
  assign n4730 = ( n347 & n858 ) | ( n347 & n1761 ) | ( n858 & n1761 ) ;
  assign n4731 = n3901 & ~n4730 ;
  assign n4732 = ( n1867 & ~n2448 ) | ( n1867 & n4318 ) | ( ~n2448 & n4318 ) ;
  assign n4739 = ( ~n1262 & n1318 ) | ( ~n1262 & n1629 ) | ( n1318 & n1629 ) ;
  assign n4736 = ~n991 & n3728 ;
  assign n4737 = n4736 ^ n1551 ^ 1'b0 ;
  assign n4738 = ~n2470 & n4737 ;
  assign n4733 = n2227 ^ n2201 ^ 1'b0 ;
  assign n4734 = n890 & ~n4733 ;
  assign n4735 = n4734 ^ n3671 ^ x115 ;
  assign n4740 = n4739 ^ n4738 ^ n4735 ;
  assign n4741 = n2495 ^ n402 ^ 1'b0 ;
  assign n4742 = n4740 & n4741 ;
  assign n4743 = ( n3574 & ~n4732 ) | ( n3574 & n4742 ) | ( ~n4732 & n4742 ) ;
  assign n4744 = ( ~n4081 & n4731 ) | ( ~n4081 & n4743 ) | ( n4731 & n4743 ) ;
  assign n4745 = n1556 | n2323 ;
  assign n4746 = n3619 | n4745 ;
  assign n4747 = x107 & n3370 ;
  assign n4748 = n974 & n4747 ;
  assign n4750 = ( ~n509 & n913 ) | ( ~n509 & n1421 ) | ( n913 & n1421 ) ;
  assign n4749 = n613 | n4461 ;
  assign n4751 = n4750 ^ n4749 ^ n3833 ;
  assign n4752 = n4751 ^ n4034 ^ 1'b0 ;
  assign n4753 = ~n4748 & n4752 ;
  assign n4754 = ~n4746 & n4753 ;
  assign n4755 = n2708 ^ n1629 ^ n700 ;
  assign n4756 = ( ~n1370 & n3952 ) | ( ~n1370 & n4755 ) | ( n3952 & n4755 ) ;
  assign n4757 = n4754 & ~n4756 ;
  assign n4758 = ( n489 & n1090 ) | ( n489 & ~n2294 ) | ( n1090 & ~n2294 ) ;
  assign n4759 = n1233 & n1948 ;
  assign n4760 = n4759 ^ n4430 ^ 1'b0 ;
  assign n4761 = ( ~n1687 & n2385 ) | ( ~n1687 & n3553 ) | ( n2385 & n3553 ) ;
  assign n4762 = n2931 ^ n558 ^ n319 ;
  assign n4763 = ~n916 & n4762 ;
  assign n4764 = ~n4761 & n4763 ;
  assign n4765 = ( x119 & ~n4197 ) | ( x119 & n4764 ) | ( ~n4197 & n4764 ) ;
  assign n4782 = n3912 ^ n2520 ^ 1'b0 ;
  assign n4780 = ( n657 & ~n909 ) | ( n657 & n2728 ) | ( ~n909 & n2728 ) ;
  assign n4781 = n1651 & ~n4780 ;
  assign n4766 = n189 & ~n3226 ;
  assign n4767 = ~n2033 & n4766 ;
  assign n4768 = ( n1046 & ~n1184 ) | ( n1046 & n3305 ) | ( ~n1184 & n3305 ) ;
  assign n4771 = ( ~n332 & n458 ) | ( ~n332 & n516 ) | ( n458 & n516 ) ;
  assign n4772 = n562 & ~n4771 ;
  assign n4773 = ~x120 & n4772 ;
  assign n4769 = n675 | n1114 ;
  assign n4770 = n2282 & ~n4769 ;
  assign n4774 = n4773 ^ n4770 ^ n3247 ;
  assign n4775 = ( n1618 & n2738 ) | ( n1618 & n3041 ) | ( n2738 & n3041 ) ;
  assign n4776 = n4775 ^ n3568 ^ 1'b0 ;
  assign n4777 = ( n4527 & ~n4774 ) | ( n4527 & n4776 ) | ( ~n4774 & n4776 ) ;
  assign n4778 = n4777 ^ n4240 ^ n161 ;
  assign n4779 = ( ~n4767 & n4768 ) | ( ~n4767 & n4778 ) | ( n4768 & n4778 ) ;
  assign n4783 = n4782 ^ n4781 ^ n4779 ;
  assign n4787 = ( ~n245 & n1545 ) | ( ~n245 & n1653 ) | ( n1545 & n1653 ) ;
  assign n4785 = ( n141 & n594 ) | ( n141 & ~n2218 ) | ( n594 & ~n2218 ) ;
  assign n4786 = ( n1239 & ~n2433 ) | ( n1239 & n4785 ) | ( ~n2433 & n4785 ) ;
  assign n4784 = n3811 ^ n2488 ^ n1862 ;
  assign n4788 = n4787 ^ n4786 ^ n4784 ;
  assign n4796 = n816 ^ n676 ^ n556 ;
  assign n4797 = n4796 ^ n861 ^ x17 ;
  assign n4798 = n4797 ^ n2820 ^ n2538 ;
  assign n4793 = n591 ^ x58 ^ 1'b0 ;
  assign n4794 = n235 & n4793 ;
  assign n4795 = ( n1447 & n1723 ) | ( n1447 & ~n4794 ) | ( n1723 & ~n4794 ) ;
  assign n4789 = n4234 ^ n1833 ^ x90 ;
  assign n4790 = n4789 ^ n3845 ^ n1843 ;
  assign n4791 = n3781 & n4093 ;
  assign n4792 = ( ~n1905 & n4790 ) | ( ~n1905 & n4791 ) | ( n4790 & n4791 ) ;
  assign n4799 = n4798 ^ n4795 ^ n4792 ;
  assign n4801 = ( x98 & n529 ) | ( x98 & ~n1000 ) | ( n529 & ~n1000 ) ;
  assign n4800 = ( n457 & ~n1362 ) | ( n457 & n3090 ) | ( ~n1362 & n3090 ) ;
  assign n4802 = n4801 ^ n4800 ^ n1704 ;
  assign n4803 = n1031 ^ x106 ^ 1'b0 ;
  assign n4804 = n154 | n4803 ;
  assign n4805 = ( n2097 & n3986 ) | ( n2097 & n4804 ) | ( n3986 & n4804 ) ;
  assign n4806 = n4805 ^ n3413 ^ 1'b0 ;
  assign n4807 = ~n520 & n760 ;
  assign n4808 = n4807 ^ n4386 ^ 1'b0 ;
  assign n4809 = ~n1595 & n1883 ;
  assign n4810 = ~n4808 & n4809 ;
  assign n4811 = n4806 | n4810 ;
  assign n4813 = ( ~n582 & n2779 ) | ( ~n582 & n3075 ) | ( n2779 & n3075 ) ;
  assign n4812 = n4354 ^ n1989 ^ n230 ;
  assign n4814 = n4813 ^ n4812 ^ n1375 ;
  assign n4815 = n1403 ^ n1367 ^ 1'b0 ;
  assign n4816 = ( ~n2193 & n2747 ) | ( ~n2193 & n3072 ) | ( n2747 & n3072 ) ;
  assign n4817 = ( n3032 & n4815 ) | ( n3032 & n4816 ) | ( n4815 & n4816 ) ;
  assign n4818 = n4817 ^ n2887 ^ n1634 ;
  assign n4819 = n2508 ^ n2097 ^ n1071 ;
  assign n4820 = n3234 ^ n2645 ^ n1930 ;
  assign n4821 = n4820 ^ n4483 ^ n1035 ;
  assign n4822 = n919 & n4821 ;
  assign n4823 = ~n4819 & n4822 ;
  assign n4824 = n237 & n4310 ;
  assign n4825 = n4824 ^ n3975 ^ 1'b0 ;
  assign n4826 = n1768 & n4629 ;
  assign n4827 = n4826 ^ n825 ^ 1'b0 ;
  assign n4828 = n4827 ^ n4623 ^ n1663 ;
  assign n4829 = ( n232 & ~n4825 ) | ( n232 & n4828 ) | ( ~n4825 & n4828 ) ;
  assign n4832 = n737 ^ n561 ^ 1'b0 ;
  assign n4833 = n4832 ^ n3275 ^ n603 ;
  assign n4834 = ( n339 & n3811 ) | ( n339 & ~n4833 ) | ( n3811 & ~n4833 ) ;
  assign n4830 = n2697 & ~n3595 ;
  assign n4831 = ( ~n573 & n1912 ) | ( ~n573 & n4830 ) | ( n1912 & n4830 ) ;
  assign n4835 = n4834 ^ n4831 ^ 1'b0 ;
  assign n4836 = ( n3711 & n4008 ) | ( n3711 & ~n4216 ) | ( n4008 & ~n4216 ) ;
  assign n4837 = ( n2172 & n3197 ) | ( n2172 & n4836 ) | ( n3197 & n4836 ) ;
  assign n4838 = n4837 ^ n4352 ^ 1'b0 ;
  assign n4839 = n2899 | n4838 ;
  assign n4840 = n1273 & ~n1511 ;
  assign n4841 = n4840 ^ n2244 ^ 1'b0 ;
  assign n4847 = n1017 & ~n1753 ;
  assign n4848 = n4847 ^ n778 ^ 1'b0 ;
  assign n4842 = ~n1288 & n3874 ;
  assign n4843 = n4842 ^ n3217 ^ 1'b0 ;
  assign n4844 = ( ~n1528 & n3525 ) | ( ~n1528 & n4843 ) | ( n3525 & n4843 ) ;
  assign n4845 = n1166 & ~n4844 ;
  assign n4846 = ( ~n909 & n4831 ) | ( ~n909 & n4845 ) | ( n4831 & n4845 ) ;
  assign n4849 = n4848 ^ n4846 ^ 1'b0 ;
  assign n4850 = n4841 & ~n4849 ;
  assign n4851 = n3541 & ~n4850 ;
  assign n4855 = ( n295 & ~n1300 ) | ( n295 & n3158 ) | ( ~n1300 & n3158 ) ;
  assign n4856 = ( ~n1833 & n4392 ) | ( ~n1833 & n4855 ) | ( n4392 & n4855 ) ;
  assign n4852 = n4085 ^ n835 ^ 1'b0 ;
  assign n4853 = n778 & n4852 ;
  assign n4854 = n4853 ^ n2379 ^ n1146 ;
  assign n4857 = n4856 ^ n4854 ^ n2110 ;
  assign n4866 = n549 | n2234 ;
  assign n4867 = n4866 ^ n3637 ^ n661 ;
  assign n4858 = n3324 ^ n1504 ^ n1191 ;
  assign n4859 = n3486 ^ n1100 ^ n462 ;
  assign n4860 = ( x29 & n1557 ) | ( x29 & ~n4859 ) | ( n1557 & ~n4859 ) ;
  assign n4861 = ( n2279 & ~n4858 ) | ( n2279 & n4860 ) | ( ~n4858 & n4860 ) ;
  assign n4862 = n4861 ^ n4556 ^ n2634 ;
  assign n4863 = n2668 | n4862 ;
  assign n4864 = n4863 ^ n472 ^ 1'b0 ;
  assign n4865 = n593 & n4864 ;
  assign n4868 = n4867 ^ n4865 ^ 1'b0 ;
  assign n4869 = n3721 ^ n1218 ^ x58 ;
  assign n4870 = n4869 ^ n2215 ^ 1'b0 ;
  assign n4871 = n4870 ^ n2225 ^ n1824 ;
  assign n4872 = n4871 ^ n3106 ^ n382 ;
  assign n4873 = n1251 | n3292 ;
  assign n4874 = ( n343 & n377 ) | ( n343 & ~n865 ) | ( n377 & ~n865 ) ;
  assign n4875 = n1767 & n4874 ;
  assign n4876 = n1500 & n4875 ;
  assign n4877 = n4873 & ~n4876 ;
  assign n4878 = n1393 ^ n741 ^ n426 ;
  assign n4879 = n4878 ^ n2733 ^ x102 ;
  assign n4880 = n4120 ^ n1644 ^ n1067 ;
  assign n4881 = ( n500 & ~n2356 ) | ( n500 & n4497 ) | ( ~n2356 & n4497 ) ;
  assign n4882 = n4444 ^ n2787 ^ n1138 ;
  assign n4883 = n4882 ^ n2208 ^ n1681 ;
  assign n4884 = n3355 ^ n1731 ^ n335 ;
  assign n4885 = n2115 ^ n1466 ^ 1'b0 ;
  assign n4886 = n3552 | n4885 ;
  assign n4887 = n4884 & ~n4886 ;
  assign n4888 = ~x33 & n4887 ;
  assign n4894 = n1253 ^ n608 ^ 1'b0 ;
  assign n4893 = ( ~n319 & n2066 ) | ( ~n319 & n2755 ) | ( n2066 & n2755 ) ;
  assign n4895 = n4894 ^ n4893 ^ 1'b0 ;
  assign n4890 = n4626 ^ n1940 ^ 1'b0 ;
  assign n4889 = ( n1162 & n1801 ) | ( n1162 & n3413 ) | ( n1801 & n3413 ) ;
  assign n4891 = n4890 ^ n4889 ^ 1'b0 ;
  assign n4892 = ~n4205 & n4891 ;
  assign n4896 = n4895 ^ n4892 ^ 1'b0 ;
  assign n4897 = ( ~n2000 & n2408 ) | ( ~n2000 & n3708 ) | ( n2408 & n3708 ) ;
  assign n4907 = ( ~n1901 & n1924 ) | ( ~n1901 & n3316 ) | ( n1924 & n3316 ) ;
  assign n4905 = ( n1393 & n3164 ) | ( n1393 & ~n3259 ) | ( n3164 & ~n3259 ) ;
  assign n4903 = n2769 & ~n4684 ;
  assign n4904 = n1919 | n4903 ;
  assign n4906 = n4905 ^ n4904 ^ 1'b0 ;
  assign n4898 = n3928 ^ n1085 ^ 1'b0 ;
  assign n4899 = n2683 & ~n4898 ;
  assign n4900 = n2809 ^ n2474 ^ 1'b0 ;
  assign n4901 = ( n686 & n4899 ) | ( n686 & ~n4900 ) | ( n4899 & ~n4900 ) ;
  assign n4902 = n4901 ^ n2341 ^ n898 ;
  assign n4908 = n4907 ^ n4906 ^ n4902 ;
  assign n4909 = n277 & ~n1732 ;
  assign n4910 = n2611 ^ n639 ^ 1'b0 ;
  assign n4911 = ( x127 & n600 ) | ( x127 & n4910 ) | ( n600 & n4910 ) ;
  assign n4912 = ( ~n1601 & n3153 ) | ( ~n1601 & n4911 ) | ( n3153 & n4911 ) ;
  assign n4921 = ( n553 & n1478 ) | ( n553 & n4467 ) | ( n1478 & n4467 ) ;
  assign n4922 = n4921 ^ n1685 ^ 1'b0 ;
  assign n4916 = n995 | n2085 ;
  assign n4917 = n4916 ^ n543 ^ 1'b0 ;
  assign n4918 = n1594 & n4917 ;
  assign n4914 = ( ~n280 & n878 ) | ( ~n280 & n1834 ) | ( n878 & n1834 ) ;
  assign n4915 = n4914 ^ n1768 ^ n1521 ;
  assign n4919 = n4918 ^ n4915 ^ n558 ;
  assign n4913 = n1630 & n2429 ;
  assign n4920 = n4919 ^ n4913 ^ n4184 ;
  assign n4923 = n4922 ^ n4920 ^ n680 ;
  assign n4924 = ( n397 & n1235 ) | ( n397 & ~n1961 ) | ( n1235 & ~n1961 ) ;
  assign n4929 = n728 | n1342 ;
  assign n4930 = n2035 & ~n4929 ;
  assign n4931 = n4930 ^ n4910 ^ x125 ;
  assign n4925 = n1309 ^ n1242 ^ n312 ;
  assign n4926 = n4925 ^ n3977 ^ 1'b0 ;
  assign n4927 = ( ~n275 & n3350 ) | ( ~n275 & n4926 ) | ( n3350 & n4926 ) ;
  assign n4928 = n2420 | n4927 ;
  assign n4932 = n4931 ^ n4928 ^ 1'b0 ;
  assign n4933 = ( ~n3040 & n4924 ) | ( ~n3040 & n4932 ) | ( n4924 & n4932 ) ;
  assign n4934 = ( ~n447 & n488 ) | ( ~n447 & n1323 ) | ( n488 & n1323 ) ;
  assign n4935 = n4934 ^ n1712 ^ n1573 ;
  assign n4936 = n3976 ^ n3576 ^ n3155 ;
  assign n4937 = ( n1833 & n4935 ) | ( n1833 & ~n4936 ) | ( n4935 & ~n4936 ) ;
  assign n4940 = ( ~x34 & n272 ) | ( ~x34 & n3773 ) | ( n272 & n3773 ) ;
  assign n4941 = n4940 ^ n2749 ^ n251 ;
  assign n4938 = n4911 ^ n393 ^ 1'b0 ;
  assign n4939 = n2930 & n4938 ;
  assign n4942 = n4941 ^ n4939 ^ 1'b0 ;
  assign n4943 = n3603 & n4942 ;
  assign n4944 = n3489 ^ n2678 ^ n1725 ;
  assign n4945 = ( ~x26 & n4943 ) | ( ~x26 & n4944 ) | ( n4943 & n4944 ) ;
  assign n4946 = ~n1136 & n1648 ;
  assign n4947 = n4946 ^ n1167 ^ 1'b0 ;
  assign n4948 = ( n505 & ~n1605 ) | ( n505 & n4947 ) | ( ~n1605 & n4947 ) ;
  assign n4949 = n2863 ^ n399 ^ 1'b0 ;
  assign n4950 = n287 | n4949 ;
  assign n4952 = n205 & ~n2240 ;
  assign n4953 = n4952 ^ n2409 ^ n1366 ;
  assign n4951 = n3439 ^ n2424 ^ n143 ;
  assign n4954 = n4953 ^ n4951 ^ n2038 ;
  assign n4955 = ~n4950 & n4954 ;
  assign n4956 = ~n1442 & n4955 ;
  assign n4957 = n4948 | n4956 ;
  assign n4958 = n4153 & ~n4957 ;
  assign n4959 = ( ~n2188 & n2774 ) | ( ~n2188 & n4815 ) | ( n2774 & n4815 ) ;
  assign n4960 = ( n505 & n1174 ) | ( n505 & n4959 ) | ( n1174 & n4959 ) ;
  assign n4961 = n3604 ^ n1190 ^ n667 ;
  assign n4962 = ( ~x10 & n378 ) | ( ~x10 & n4190 ) | ( n378 & n4190 ) ;
  assign n4963 = n4961 & n4962 ;
  assign n4964 = ~n691 & n1072 ;
  assign n4965 = ( n130 & ~n226 ) | ( n130 & n2367 ) | ( ~n226 & n2367 ) ;
  assign n4966 = n4965 ^ n1875 ^ n289 ;
  assign n4967 = ( ~n260 & n4964 ) | ( ~n260 & n4966 ) | ( n4964 & n4966 ) ;
  assign n4968 = ( n611 & n4230 ) | ( n611 & ~n4967 ) | ( n4230 & ~n4967 ) ;
  assign n4969 = n3991 ^ n542 ^ 1'b0 ;
  assign n4970 = n4968 & n4969 ;
  assign n4971 = ( n1299 & n2181 ) | ( n1299 & ~n2239 ) | ( n2181 & ~n2239 ) ;
  assign n4972 = n4971 ^ n2402 ^ 1'b0 ;
  assign n4973 = n710 ^ n379 ^ 1'b0 ;
  assign n4974 = ( ~n1233 & n3288 ) | ( ~n1233 & n4973 ) | ( n3288 & n4973 ) ;
  assign n4975 = n4974 ^ n2000 ^ 1'b0 ;
  assign n4976 = n4972 | n4975 ;
  assign n4977 = n4976 ^ n2853 ^ n1833 ;
  assign n4978 = x123 & n2692 ;
  assign n4979 = ~n146 & n4978 ;
  assign n4980 = ( ~n3209 & n4241 ) | ( ~n3209 & n4979 ) | ( n4241 & n4979 ) ;
  assign n4981 = n4980 ^ n3575 ^ 1'b0 ;
  assign n4982 = n4977 & ~n4981 ;
  assign n4987 = ( n944 & n2022 ) | ( n944 & n3431 ) | ( n2022 & n3431 ) ;
  assign n4983 = ( n436 & ~n1074 ) | ( n436 & n3139 ) | ( ~n1074 & n3139 ) ;
  assign n4984 = n4983 ^ n1396 ^ n1020 ;
  assign n4985 = n4984 ^ n3700 ^ 1'b0 ;
  assign n4986 = n4862 | n4985 ;
  assign n4988 = n4987 ^ n4986 ^ 1'b0 ;
  assign n4989 = n4988 ^ n4247 ^ n3027 ;
  assign n4990 = ~n1092 & n1236 ;
  assign n4991 = n4990 ^ n2728 ^ n201 ;
  assign n4992 = ( n3726 & n4729 ) | ( n3726 & ~n4991 ) | ( n4729 & ~n4991 ) ;
  assign n4996 = ( n768 & ~n1009 ) | ( n768 & n2009 ) | ( ~n1009 & n2009 ) ;
  assign n4993 = ( ~n2356 & n3254 ) | ( ~n2356 & n3423 ) | ( n3254 & n3423 ) ;
  assign n4994 = ( x68 & n3510 ) | ( x68 & ~n4384 ) | ( n3510 & ~n4384 ) ;
  assign n4995 = ~n4993 & n4994 ;
  assign n4997 = n4996 ^ n4995 ^ 1'b0 ;
  assign n4998 = n3872 ^ n2599 ^ 1'b0 ;
  assign n4999 = n3168 & n4998 ;
  assign n5000 = n4999 ^ n3680 ^ 1'b0 ;
  assign n5001 = ( n1887 & ~n3178 ) | ( n1887 & n4615 ) | ( ~n3178 & n4615 ) ;
  assign n5002 = ( ~n2827 & n3922 ) | ( ~n2827 & n4941 ) | ( n3922 & n4941 ) ;
  assign n5003 = n3319 ^ n1542 ^ n1527 ;
  assign n5004 = ( ~n2081 & n2933 ) | ( ~n2081 & n5003 ) | ( n2933 & n5003 ) ;
  assign n5005 = n553 | n4819 ;
  assign n5006 = n5005 ^ n693 ^ 1'b0 ;
  assign n5007 = n5004 | n5006 ;
  assign n5008 = n1859 ^ n1490 ^ 1'b0 ;
  assign n5009 = ( n265 & n1886 ) | ( n265 & n5008 ) | ( n1886 & n5008 ) ;
  assign n5010 = n4076 ^ n3817 ^ 1'b0 ;
  assign n5011 = ~n2761 & n5010 ;
  assign n5020 = n3223 ^ n1573 ^ 1'b0 ;
  assign n5019 = ( n202 & n2662 ) | ( n202 & ~n3713 ) | ( n2662 & ~n3713 ) ;
  assign n5021 = n5020 ^ n5019 ^ n1917 ;
  assign n5012 = n4474 ^ n2398 ^ n1163 ;
  assign n5013 = n5012 ^ n3337 ^ n758 ;
  assign n5014 = n2294 & n5013 ;
  assign n5015 = n1097 & ~n5014 ;
  assign n5016 = n4336 ^ n2036 ^ n896 ;
  assign n5017 = ~n3278 & n5016 ;
  assign n5018 = n5015 & n5017 ;
  assign n5022 = n5021 ^ n5018 ^ 1'b0 ;
  assign n5027 = n2140 ^ n1887 ^ x4 ;
  assign n5023 = n2041 ^ n1348 ^ x47 ;
  assign n5024 = n5023 ^ n1335 ^ n816 ;
  assign n5025 = n5024 ^ n3224 ^ n1510 ;
  assign n5026 = x19 & ~n5025 ;
  assign n5028 = n5027 ^ n5026 ^ 1'b0 ;
  assign n5029 = n5028 ^ n1250 ^ 1'b0 ;
  assign n5030 = ~n4823 & n5029 ;
  assign n5031 = n670 & n3498 ;
  assign n5032 = x121 | n1840 ;
  assign n5033 = n5032 ^ n1771 ^ 1'b0 ;
  assign n5034 = n5033 ^ n4373 ^ n2094 ;
  assign n5035 = ( n4600 & n5031 ) | ( n4600 & n5034 ) | ( n5031 & n5034 ) ;
  assign n5036 = ( n480 & ~n981 ) | ( n480 & n1303 ) | ( ~n981 & n1303 ) ;
  assign n5037 = ( n928 & n3644 ) | ( n928 & n5036 ) | ( n3644 & n5036 ) ;
  assign n5038 = n3354 ^ n1599 ^ n659 ;
  assign n5039 = n5038 ^ n3464 ^ n3434 ;
  assign n5040 = n4947 ^ n2319 ^ n2306 ;
  assign n5041 = ( n313 & n543 ) | ( n313 & ~n3714 ) | ( n543 & ~n3714 ) ;
  assign n5042 = ~n1540 & n5041 ;
  assign n5043 = ~n962 & n5042 ;
  assign n5050 = x97 | n3176 ;
  assign n5046 = n2234 ^ n1748 ^ n578 ;
  assign n5047 = n4288 ^ n3947 ^ 1'b0 ;
  assign n5048 = n1887 | n5047 ;
  assign n5049 = ~n5046 & n5048 ;
  assign n5051 = n5050 ^ n5049 ^ n4907 ;
  assign n5052 = n5051 ^ n4853 ^ n2184 ;
  assign n5044 = n1046 ^ n962 ^ n837 ;
  assign n5045 = n5044 ^ n1263 ^ n1207 ;
  assign n5053 = n5052 ^ n5045 ^ n2683 ;
  assign n5055 = n620 & ~n3423 ;
  assign n5056 = n5055 ^ n1627 ^ 1'b0 ;
  assign n5054 = ( x9 & ~n222 ) | ( x9 & n2977 ) | ( ~n222 & n2977 ) ;
  assign n5057 = n5056 ^ n5054 ^ n3192 ;
  assign n5058 = n3203 ^ n1767 ^ n426 ;
  assign n5059 = n5058 ^ n676 ^ 1'b0 ;
  assign n5060 = ( x60 & n1692 ) | ( x60 & ~n3238 ) | ( n1692 & ~n3238 ) ;
  assign n5061 = n169 & ~n5060 ;
  assign n5062 = ( n1262 & ~n2301 ) | ( n1262 & n2607 ) | ( ~n2301 & n2607 ) ;
  assign n5063 = n5062 ^ n4634 ^ n4062 ;
  assign n5064 = n2568 & n4015 ;
  assign n5065 = n2541 & n5064 ;
  assign n5066 = ( ~x25 & n1402 ) | ( ~x25 & n2000 ) | ( n1402 & n2000 ) ;
  assign n5067 = n5066 ^ n2179 ^ n865 ;
  assign n5068 = n2103 ^ n1232 ^ 1'b0 ;
  assign n5069 = n5068 ^ n2060 ^ 1'b0 ;
  assign n5070 = n2270 ^ n1893 ^ n1518 ;
  assign n5071 = n1320 | n5070 ;
  assign n5072 = n5069 | n5071 ;
  assign n5073 = n5072 ^ n386 ^ 1'b0 ;
  assign n5074 = n405 ^ x89 ^ 1'b0 ;
  assign n5075 = ( ~x25 & x83 ) | ( ~x25 & n384 ) | ( x83 & n384 ) ;
  assign n5076 = n502 & n820 ;
  assign n5077 = ~n1190 & n5076 ;
  assign n5078 = ( ~n608 & n1112 ) | ( ~n608 & n5077 ) | ( n1112 & n5077 ) ;
  assign n5079 = n1929 ^ n927 ^ n624 ;
  assign n5080 = ( n1239 & n5078 ) | ( n1239 & n5079 ) | ( n5078 & n5079 ) ;
  assign n5081 = ( n5074 & n5075 ) | ( n5074 & n5080 ) | ( n5075 & n5080 ) ;
  assign n5082 = n5081 ^ n4451 ^ n2078 ;
  assign n5083 = ( n681 & n2058 ) | ( n681 & ~n4405 ) | ( n2058 & ~n4405 ) ;
  assign n5084 = n5083 ^ n1350 ^ n1247 ;
  assign n5088 = ~n1067 & n1594 ;
  assign n5089 = ~n2087 & n5088 ;
  assign n5090 = ( n2622 & ~n3483 ) | ( n2622 & n5089 ) | ( ~n3483 & n5089 ) ;
  assign n5091 = n967 & ~n5090 ;
  assign n5085 = n1326 ^ n548 ^ 1'b0 ;
  assign n5086 = n724 & ~n5085 ;
  assign n5087 = n5086 ^ n4699 ^ 1'b0 ;
  assign n5092 = n5091 ^ n5087 ^ 1'b0 ;
  assign n5093 = ~n5084 & n5092 ;
  assign n5094 = n3045 | n3464 ;
  assign n5095 = n5094 ^ n1021 ^ 1'b0 ;
  assign n5096 = n2274 & n5095 ;
  assign n5097 = n5096 ^ x44 ^ 1'b0 ;
  assign n5098 = ( ~n2992 & n4626 ) | ( ~n2992 & n4882 ) | ( n4626 & n4882 ) ;
  assign n5111 = ~n1403 & n4704 ;
  assign n5112 = n164 & n5111 ;
  assign n5108 = n2513 ^ n2449 ^ n1382 ;
  assign n5100 = n1409 ^ n1183 ^ n614 ;
  assign n5101 = n5100 ^ n3196 ^ 1'b0 ;
  assign n5102 = n2299 | n5101 ;
  assign n5103 = n287 & ~n5102 ;
  assign n5104 = ( n1797 & n2309 ) | ( n1797 & ~n5103 ) | ( n2309 & ~n5103 ) ;
  assign n5105 = n591 & n2165 ;
  assign n5106 = ~n5104 & n5105 ;
  assign n5107 = n5106 ^ n4767 ^ n2886 ;
  assign n5109 = n5108 ^ n5107 ^ 1'b0 ;
  assign n5110 = n3501 | n5109 ;
  assign n5099 = ( n710 & n1295 ) | ( n710 & n1607 ) | ( n1295 & n1607 ) ;
  assign n5113 = n5112 ^ n5110 ^ n5099 ;
  assign n5114 = n3165 ^ n1566 ^ x121 ;
  assign n5115 = n5114 ^ n4503 ^ n2250 ;
  assign n5116 = n5115 ^ n4815 ^ 1'b0 ;
  assign n5117 = ( n1917 & ~n4270 ) | ( n1917 & n5116 ) | ( ~n4270 & n5116 ) ;
  assign n5118 = n505 | n2224 ;
  assign n5119 = ~n1822 & n5118 ;
  assign n5120 = ( n631 & n2686 ) | ( n631 & ~n5119 ) | ( n2686 & ~n5119 ) ;
  assign n5121 = n2449 ^ n1519 ^ n1417 ;
  assign n5122 = n5121 ^ n3641 ^ 1'b0 ;
  assign n5123 = ~n4502 & n4939 ;
  assign n5124 = n1973 ^ n1242 ^ x23 ;
  assign n5125 = n4796 ^ n739 ^ n468 ;
  assign n5126 = ( n2491 & n5124 ) | ( n2491 & ~n5125 ) | ( n5124 & ~n5125 ) ;
  assign n5127 = ~n5123 & n5126 ;
  assign n5128 = x106 & ~n1840 ;
  assign n5129 = ( n1738 & n3534 ) | ( n1738 & n5128 ) | ( n3534 & n5128 ) ;
  assign n5130 = n273 & ~n1741 ;
  assign n5131 = n5130 ^ n4593 ^ 1'b0 ;
  assign n5132 = n4117 ^ n1356 ^ n291 ;
  assign n5133 = n5132 ^ n3079 ^ x104 ;
  assign n5134 = n3094 & n5133 ;
  assign n5135 = ~n5131 & n5134 ;
  assign n5136 = n3410 ^ n2791 ^ n324 ;
  assign n5137 = n2414 & n5136 ;
  assign n5138 = n5135 & n5137 ;
  assign n5139 = ( n1732 & n3098 ) | ( n1732 & ~n3805 ) | ( n3098 & ~n3805 ) ;
  assign n5140 = n4377 ^ n3284 ^ 1'b0 ;
  assign n5141 = ~n190 & n5140 ;
  assign n5146 = n1078 & ~n1297 ;
  assign n5145 = n729 | n924 ;
  assign n5147 = n5146 ^ n5145 ^ 1'b0 ;
  assign n5142 = n2137 ^ n1776 ^ n635 ;
  assign n5143 = n1873 & ~n5142 ;
  assign n5144 = ~n3382 & n5143 ;
  assign n5148 = n5147 ^ n5144 ^ n2364 ;
  assign n5149 = n3798 ^ n722 ^ n643 ;
  assign n5150 = n5149 ^ n2066 ^ 1'b0 ;
  assign n5151 = n548 & ~n5150 ;
  assign n5152 = ( n3408 & n3952 ) | ( n3408 & ~n4860 ) | ( n3952 & ~n4860 ) ;
  assign n5153 = ( ~n561 & n3653 ) | ( ~n561 & n3735 ) | ( n3653 & n3735 ) ;
  assign n5154 = n5038 & ~n5153 ;
  assign n5155 = n5152 & n5154 ;
  assign n5156 = n5155 ^ n4595 ^ n176 ;
  assign n5157 = n5156 ^ n4202 ^ n3428 ;
  assign n5158 = n5157 ^ n260 ^ 1'b0 ;
  assign n5159 = n811 & n5158 ;
  assign n5160 = ( n1228 & n4056 ) | ( n1228 & n5025 ) | ( n4056 & n5025 ) ;
  assign n5161 = x28 & n2943 ;
  assign n5162 = ~n1125 & n5161 ;
  assign n5163 = n3269 ^ n1400 ^ n830 ;
  assign n5164 = n5163 ^ n2569 ^ 1'b0 ;
  assign n5165 = n5162 | n5164 ;
  assign n5166 = n5165 ^ n4148 ^ 1'b0 ;
  assign n5167 = ~n2000 & n5166 ;
  assign n5168 = ( n529 & n1315 ) | ( n529 & ~n2138 ) | ( n1315 & ~n2138 ) ;
  assign n5169 = ( ~x99 & n1529 ) | ( ~x99 & n5168 ) | ( n1529 & n5168 ) ;
  assign n5170 = ( n1075 & n1307 ) | ( n1075 & n5169 ) | ( n1307 & n5169 ) ;
  assign n5171 = n1779 & ~n1822 ;
  assign n5172 = ~n2033 & n5171 ;
  assign n5173 = n5172 ^ n3334 ^ 1'b0 ;
  assign n5174 = n5170 | n5173 ;
  assign n5175 = n1796 & ~n5174 ;
  assign n5176 = n5175 ^ n1361 ^ 1'b0 ;
  assign n5177 = n2385 & ~n4561 ;
  assign n5179 = n1253 & ~n2110 ;
  assign n5178 = ( n634 & n1644 ) | ( n634 & n1871 ) | ( n1644 & n1871 ) ;
  assign n5180 = n5179 ^ n5178 ^ n3413 ;
  assign n5181 = ( ~n1393 & n2029 ) | ( ~n1393 & n5180 ) | ( n2029 & n5180 ) ;
  assign n5182 = n4704 & ~n5181 ;
  assign n5183 = n1553 & n5182 ;
  assign n5184 = n878 | n4719 ;
  assign n5193 = ( n405 & n2621 ) | ( n405 & n4406 ) | ( n2621 & n4406 ) ;
  assign n5185 = x71 & ~n1203 ;
  assign n5186 = ~n337 & n5185 ;
  assign n5187 = n5186 ^ n2092 ^ 1'b0 ;
  assign n5188 = n3145 ^ n2778 ^ 1'b0 ;
  assign n5189 = ~n5187 & n5188 ;
  assign n5190 = n3198 & n5189 ;
  assign n5191 = n5190 ^ n902 ^ 1'b0 ;
  assign n5192 = n5191 ^ n3609 ^ n3219 ;
  assign n5194 = n5193 ^ n5192 ^ n4085 ;
  assign n5195 = n1963 ^ n1396 ^ n1366 ;
  assign n5196 = n5195 ^ n4331 ^ 1'b0 ;
  assign n5197 = n5196 ^ n1532 ^ n1138 ;
  assign n5200 = n2778 ^ n1839 ^ 1'b0 ;
  assign n5201 = n4801 & ~n5200 ;
  assign n5198 = ( n1114 & ~n2402 ) | ( n1114 & n2834 ) | ( ~n2402 & n2834 ) ;
  assign n5199 = n5198 ^ n3951 ^ n1779 ;
  assign n5202 = n5201 ^ n5199 ^ n2583 ;
  assign n5203 = n5202 ^ n5187 ^ 1'b0 ;
  assign n5204 = n1312 & ~n5203 ;
  assign n5205 = n1769 & ~n2520 ;
  assign n5206 = ( n1932 & ~n3103 ) | ( n1932 & n5205 ) | ( ~n3103 & n5205 ) ;
  assign n5207 = ( n992 & n4654 ) | ( n992 & ~n5206 ) | ( n4654 & ~n5206 ) ;
  assign n5208 = n582 & ~n4037 ;
  assign n5209 = n5208 ^ n1043 ^ 1'b0 ;
  assign n5210 = ( ~n728 & n1304 ) | ( ~n728 & n5209 ) | ( n1304 & n5209 ) ;
  assign n5211 = n600 ^ n551 ^ 1'b0 ;
  assign n5212 = ~n1451 & n5211 ;
  assign n5213 = n3120 | n5212 ;
  assign n5214 = ( n3055 & n3093 ) | ( n3055 & n5213 ) | ( n3093 & n5213 ) ;
  assign n5215 = n5214 ^ n5069 ^ n3131 ;
  assign n5216 = n5215 ^ n3672 ^ x126 ;
  assign n5217 = n5216 ^ n2674 ^ 1'b0 ;
  assign n5218 = n227 & ~n5217 ;
  assign n5219 = x43 & ~n5218 ;
  assign n5220 = ( ~n1842 & n3065 ) | ( ~n1842 & n4115 ) | ( n3065 & n4115 ) ;
  assign n5221 = ~n3884 & n5220 ;
  assign n5222 = n5221 ^ n2677 ^ 1'b0 ;
  assign n5223 = ( n1740 & n3816 ) | ( n1740 & ~n5222 ) | ( n3816 & ~n5222 ) ;
  assign n5224 = n1050 & n3653 ;
  assign n5225 = n3737 & n5224 ;
  assign n5226 = n5225 ^ n1020 ^ x4 ;
  assign n5227 = n1854 | n3957 ;
  assign n5228 = n1687 & ~n5227 ;
  assign n5229 = n1643 ^ n642 ^ 1'b0 ;
  assign n5230 = n5228 | n5229 ;
  assign n5231 = n2353 & ~n5230 ;
  assign n5232 = n5231 ^ n1021 ^ 1'b0 ;
  assign n5233 = ~n2932 & n5232 ;
  assign n5234 = ~n5226 & n5233 ;
  assign n5235 = n2769 ^ n826 ^ n203 ;
  assign n5236 = n5235 ^ n5023 ^ n1479 ;
  assign n5237 = ( n1444 & ~n3857 ) | ( n1444 & n4264 ) | ( ~n3857 & n4264 ) ;
  assign n5238 = ( n4951 & n5236 ) | ( n4951 & ~n5237 ) | ( n5236 & ~n5237 ) ;
  assign n5244 = n2198 ^ n1828 ^ n767 ;
  assign n5245 = n5244 ^ n1828 ^ 1'b0 ;
  assign n5243 = n2536 ^ n905 ^ n738 ;
  assign n5240 = n2405 ^ n1187 ^ n1090 ;
  assign n5241 = n5240 ^ n3321 ^ n602 ;
  assign n5239 = n1483 & ~n3596 ;
  assign n5242 = n5241 ^ n5239 ^ 1'b0 ;
  assign n5246 = n5245 ^ n5243 ^ n5242 ;
  assign n5247 = ~n577 & n899 ;
  assign n5248 = n5247 ^ n1201 ^ 1'b0 ;
  assign n5249 = n3167 ^ n479 ^ 1'b0 ;
  assign n5250 = ( n3075 & n5248 ) | ( n3075 & ~n5249 ) | ( n5248 & ~n5249 ) ;
  assign n5251 = n4485 ^ n571 ^ 1'b0 ;
  assign n5252 = n4971 | n5251 ;
  assign n5253 = n5252 ^ n3837 ^ n2650 ;
  assign n5254 = n4507 ^ n4213 ^ 1'b0 ;
  assign n5255 = n2041 | n5254 ;
  assign n5256 = n4622 | n5255 ;
  assign n5258 = n144 & n636 ;
  assign n5259 = ~n2098 & n5258 ;
  assign n5257 = x41 & ~n1540 ;
  assign n5260 = n5259 ^ n5257 ^ 1'b0 ;
  assign n5261 = n4901 ^ n1265 ^ 1'b0 ;
  assign n5262 = n5260 & ~n5261 ;
  assign n5263 = n5262 ^ n3950 ^ 1'b0 ;
  assign n5264 = n2653 ^ n1143 ^ 1'b0 ;
  assign n5265 = n2302 & ~n5264 ;
  assign n5266 = ~n809 & n5077 ;
  assign n5267 = n5266 ^ n3913 ^ n1037 ;
  assign n5268 = ( n1533 & ~n5265 ) | ( n1533 & n5267 ) | ( ~n5265 & n5267 ) ;
  assign n5269 = ( x7 & n1698 ) | ( x7 & ~n1767 ) | ( n1698 & ~n1767 ) ;
  assign n5270 = ( ~n313 & n4511 ) | ( ~n313 & n5269 ) | ( n4511 & n5269 ) ;
  assign n5271 = n5126 ^ n1578 ^ n1308 ;
  assign n5272 = n4971 ^ n3604 ^ x107 ;
  assign n5273 = n5272 ^ n3579 ^ n1064 ;
  assign n5295 = n3949 ^ n3337 ^ n2099 ;
  assign n5296 = ( n1205 & n1722 ) | ( n1205 & n5295 ) | ( n1722 & n5295 ) ;
  assign n5274 = ~n783 & n2036 ;
  assign n5275 = n339 & n5274 ;
  assign n5276 = ( n2664 & n4701 ) | ( n2664 & n5275 ) | ( n4701 & n5275 ) ;
  assign n5277 = n3269 ^ n1809 ^ x45 ;
  assign n5278 = n5277 ^ n2616 ^ n723 ;
  assign n5279 = n5278 ^ n2449 ^ n264 ;
  assign n5280 = n974 | n5279 ;
  assign n5281 = n785 & ~n5280 ;
  assign n5286 = n1671 ^ x125 ^ 1'b0 ;
  assign n5282 = n2329 ^ n1038 ^ 1'b0 ;
  assign n5283 = n5136 & n5282 ;
  assign n5284 = n1981 | n5283 ;
  assign n5285 = n5284 ^ n702 ^ 1'b0 ;
  assign n5287 = n5286 ^ n5285 ^ n1299 ;
  assign n5288 = n2194 ^ n744 ^ 1'b0 ;
  assign n5289 = n3710 | n5288 ;
  assign n5290 = n5289 ^ n2034 ^ 1'b0 ;
  assign n5291 = n5287 | n5290 ;
  assign n5292 = n5291 ^ n4228 ^ n1336 ;
  assign n5293 = ( n4376 & n5281 ) | ( n4376 & n5292 ) | ( n5281 & n5292 ) ;
  assign n5294 = ( n589 & ~n5276 ) | ( n589 & n5293 ) | ( ~n5276 & n5293 ) ;
  assign n5297 = n5296 ^ n5294 ^ n217 ;
  assign n5298 = n2665 ^ n721 ^ 1'b0 ;
  assign n5299 = n1306 & n4239 ;
  assign n5300 = ~n350 & n5299 ;
  assign n5307 = n897 | n3927 ;
  assign n5308 = n3396 ^ n2103 ^ x122 ;
  assign n5309 = ( n1744 & ~n5307 ) | ( n1744 & n5308 ) | ( ~n5307 & n5308 ) ;
  assign n5301 = n2121 ^ n195 ^ 1'b0 ;
  assign n5302 = n2328 & ~n5301 ;
  assign n5303 = ( ~x88 & n4285 ) | ( ~x88 & n5302 ) | ( n4285 & n5302 ) ;
  assign n5304 = n5303 ^ n271 ^ 1'b0 ;
  assign n5305 = n1720 | n5304 ;
  assign n5306 = ( n3789 & n4489 ) | ( n3789 & n5305 ) | ( n4489 & n5305 ) ;
  assign n5310 = n5309 ^ n5306 ^ n760 ;
  assign n5312 = n1839 ^ n1255 ^ n308 ;
  assign n5311 = n4925 ^ n1148 ^ 1'b0 ;
  assign n5313 = n5312 ^ n5311 ^ n4346 ;
  assign n5314 = n5310 & n5313 ;
  assign n5315 = ~n3217 & n5314 ;
  assign n5316 = n3220 ^ n2020 ^ 1'b0 ;
  assign n5317 = ( ~n2643 & n2961 ) | ( ~n2643 & n3536 ) | ( n2961 & n3536 ) ;
  assign n5318 = ( n3282 & n5316 ) | ( n3282 & ~n5317 ) | ( n5316 & ~n5317 ) ;
  assign n5319 = n5318 ^ n3946 ^ 1'b0 ;
  assign n5320 = ( n5300 & n5315 ) | ( n5300 & ~n5319 ) | ( n5315 & ~n5319 ) ;
  assign n5327 = ~n2467 & n4265 ;
  assign n5323 = ~n789 & n4212 ;
  assign n5324 = ( n2734 & ~n4078 ) | ( n2734 & n5323 ) | ( ~n4078 & n5323 ) ;
  assign n5321 = n2611 ^ n1352 ^ n521 ;
  assign n5322 = ( ~n189 & n2953 ) | ( ~n189 & n5321 ) | ( n2953 & n5321 ) ;
  assign n5325 = n5324 ^ n5322 ^ n1244 ;
  assign n5326 = n4317 & n5325 ;
  assign n5328 = n5327 ^ n5326 ^ 1'b0 ;
  assign n5329 = n1067 ^ n468 ^ n416 ;
  assign n5330 = n5329 ^ n1904 ^ n442 ;
  assign n5331 = ~n433 & n5330 ;
  assign n5348 = n5312 ^ n3849 ^ 1'b0 ;
  assign n5349 = n4866 & n5348 ;
  assign n5350 = n5245 ^ n1632 ^ 1'b0 ;
  assign n5351 = ~n2089 & n5350 ;
  assign n5352 = n5351 ^ n2070 ^ 1'b0 ;
  assign n5353 = n5349 & ~n5352 ;
  assign n5354 = ( n516 & n658 ) | ( n516 & n1363 ) | ( n658 & n1363 ) ;
  assign n5355 = n217 & n935 ;
  assign n5356 = n5355 ^ n326 ^ 1'b0 ;
  assign n5357 = n5354 | n5356 ;
  assign n5358 = n5353 | n5357 ;
  assign n5359 = n4179 ^ n4061 ^ n2317 ;
  assign n5360 = ( n3573 & ~n5358 ) | ( n3573 & n5359 ) | ( ~n5358 & n5359 ) ;
  assign n5361 = ( n175 & ~n1047 ) | ( n175 & n5360 ) | ( ~n1047 & n5360 ) ;
  assign n5346 = n4894 ^ n471 ^ n180 ;
  assign n5342 = n4782 ^ n4147 ^ 1'b0 ;
  assign n5343 = n395 & ~n5342 ;
  assign n5340 = n1457 ^ n1278 ^ 1'b0 ;
  assign n5341 = n5340 ^ n5027 ^ n1459 ;
  assign n5344 = n5343 ^ n5341 ^ n1945 ;
  assign n5336 = n172 & n2279 ;
  assign n5337 = n5336 ^ n1877 ^ n1116 ;
  assign n5332 = n3947 ^ n3277 ^ n1603 ;
  assign n5333 = n3825 ^ n462 ^ 1'b0 ;
  assign n5334 = n5332 | n5333 ;
  assign n5335 = ( ~n1665 & n3270 ) | ( ~n1665 & n5334 ) | ( n3270 & n5334 ) ;
  assign n5338 = n5337 ^ n5335 ^ 1'b0 ;
  assign n5339 = n4256 & n5338 ;
  assign n5345 = n5344 ^ n5339 ^ n559 ;
  assign n5347 = n5346 ^ n5345 ^ 1'b0 ;
  assign n5362 = n5361 ^ n5347 ^ n499 ;
  assign n5363 = n2729 & ~n3250 ;
  assign n5364 = ~n1236 & n5363 ;
  assign n5365 = n5364 ^ n2424 ^ 1'b0 ;
  assign n5366 = n2276 & n2853 ;
  assign n5367 = n170 & n5366 ;
  assign n5368 = ( n898 & n3820 ) | ( n898 & n5367 ) | ( n3820 & n5367 ) ;
  assign n5369 = ( n328 & ~n2218 ) | ( n328 & n3284 ) | ( ~n2218 & n3284 ) ;
  assign n5370 = n424 | n2679 ;
  assign n5371 = n655 & ~n5370 ;
  assign n5372 = ( n2738 & n4819 ) | ( n2738 & n5371 ) | ( n4819 & n5371 ) ;
  assign n5373 = n963 | n1151 ;
  assign n5374 = n5373 ^ n628 ^ 1'b0 ;
  assign n5375 = n5374 ^ n2157 ^ 1'b0 ;
  assign n5376 = n5375 ^ n2208 ^ n1311 ;
  assign n5377 = n5376 ^ n3900 ^ n140 ;
  assign n5378 = n1066 | n5377 ;
  assign n5379 = n5372 | n5378 ;
  assign n5380 = n4061 ^ n4046 ^ n2350 ;
  assign n5381 = n683 | n1301 ;
  assign n5382 = n5380 & n5381 ;
  assign n5383 = n5382 ^ n3446 ^ 1'b0 ;
  assign n5385 = n213 ^ n151 ^ x28 ;
  assign n5384 = n2973 ^ n1642 ^ 1'b0 ;
  assign n5386 = n5385 ^ n5384 ^ n1878 ;
  assign n5390 = ( ~n388 & n1514 ) | ( ~n388 & n5243 ) | ( n1514 & n5243 ) ;
  assign n5388 = n3688 ^ n347 ^ 1'b0 ;
  assign n5389 = n5114 | n5388 ;
  assign n5391 = n5390 ^ n5389 ^ 1'b0 ;
  assign n5387 = n4024 ^ n1978 ^ n165 ;
  assign n5392 = n5391 ^ n5387 ^ n2170 ;
  assign n5393 = n1250 | n3068 ;
  assign n5394 = n4973 ^ n3431 ^ n321 ;
  assign n5395 = ( ~n1785 & n2747 ) | ( ~n1785 & n5394 ) | ( n2747 & n5394 ) ;
  assign n5396 = n5308 & ~n5395 ;
  assign n5397 = n5396 ^ n2210 ^ 1'b0 ;
  assign n5407 = ( x78 & n1009 ) | ( x78 & n4305 ) | ( n1009 & n4305 ) ;
  assign n5408 = ( ~n1052 & n1503 ) | ( ~n1052 & n5407 ) | ( n1503 & n5407 ) ;
  assign n5406 = n2357 ^ n2109 ^ x33 ;
  assign n5403 = n2136 & n4164 ;
  assign n5404 = ~n1721 & n5403 ;
  assign n5398 = n1804 ^ n1335 ^ n1206 ;
  assign n5399 = n1092 | n5398 ;
  assign n5400 = n2983 | n5399 ;
  assign n5401 = ~n336 & n5400 ;
  assign n5402 = n5401 ^ n633 ^ 1'b0 ;
  assign n5405 = n5404 ^ n5402 ^ x49 ;
  assign n5409 = n5408 ^ n5406 ^ n5405 ;
  assign n5410 = n2667 & n2736 ;
  assign n5411 = n573 & n5410 ;
  assign n5412 = ( n1744 & n3946 ) | ( n1744 & ~n5411 ) | ( n3946 & ~n5411 ) ;
  assign n5413 = ( ~n2320 & n4614 ) | ( ~n2320 & n5412 ) | ( n4614 & n5412 ) ;
  assign n5414 = n1376 | n3198 ;
  assign n5415 = ( ~n3035 & n3934 ) | ( ~n3035 & n5414 ) | ( n3934 & n5414 ) ;
  assign n5416 = n1494 ^ n697 ^ n353 ;
  assign n5417 = n3898 | n5416 ;
  assign n5418 = n5415 & ~n5417 ;
  assign n5419 = n3250 ^ n1618 ^ n691 ;
  assign n5420 = n5027 ^ n1778 ^ 1'b0 ;
  assign n5421 = n5419 & ~n5420 ;
  assign n5422 = n5421 ^ n4640 ^ n3902 ;
  assign n5423 = ~n478 & n1608 ;
  assign n5425 = ~n1421 & n2164 ;
  assign n5426 = ~n1060 & n5425 ;
  assign n5427 = n971 & ~n1141 ;
  assign n5428 = ~n3790 & n5427 ;
  assign n5429 = n5428 ^ n2942 ^ 1'b0 ;
  assign n5430 = ( n955 & n5426 ) | ( n955 & ~n5429 ) | ( n5426 & ~n5429 ) ;
  assign n5424 = n1729 ^ n1516 ^ n1480 ;
  assign n5431 = n5430 ^ n5424 ^ 1'b0 ;
  assign n5432 = n2087 & ~n5431 ;
  assign n5433 = n768 ^ n268 ^ 1'b0 ;
  assign n5434 = ( ~n566 & n1528 ) | ( ~n566 & n5433 ) | ( n1528 & n5433 ) ;
  assign n5435 = ( ~n688 & n1441 ) | ( ~n688 & n5340 ) | ( n1441 & n5340 ) ;
  assign n5436 = ( n1254 & n3847 ) | ( n1254 & ~n5435 ) | ( n3847 & ~n5435 ) ;
  assign n5437 = ~n5434 & n5436 ;
  assign n5441 = n238 & n604 ;
  assign n5442 = n1027 & n5441 ;
  assign n5443 = n5442 ^ n3619 ^ 1'b0 ;
  assign n5444 = n1508 ^ n981 ^ 1'b0 ;
  assign n5445 = ( n1648 & n1947 ) | ( n1648 & ~n5444 ) | ( n1947 & ~n5444 ) ;
  assign n5446 = n5443 | n5445 ;
  assign n5447 = n4619 & ~n5446 ;
  assign n5448 = ( x65 & x115 ) | ( x65 & n5447 ) | ( x115 & n5447 ) ;
  assign n5449 = n5448 ^ n2919 ^ 1'b0 ;
  assign n5438 = ( n614 & n1289 ) | ( n614 & n1900 ) | ( n1289 & n1900 ) ;
  assign n5439 = ( n783 & n814 ) | ( n783 & ~n5438 ) | ( n814 & ~n5438 ) ;
  assign n5440 = n3104 & n5439 ;
  assign n5450 = n5449 ^ n5440 ^ 1'b0 ;
  assign n5451 = n4006 ^ n3684 ^ n1619 ;
  assign n5452 = n5451 ^ n617 ^ 1'b0 ;
  assign n5453 = n4608 & n5452 ;
  assign n5454 = n497 ^ n232 ^ 1'b0 ;
  assign n5455 = x30 & n5454 ;
  assign n5456 = ~n992 & n5455 ;
  assign n5457 = n5456 ^ n1020 ^ 1'b0 ;
  assign n5458 = n4148 & ~n4622 ;
  assign n5459 = ( ~n2852 & n3520 ) | ( ~n2852 & n5004 ) | ( n3520 & n5004 ) ;
  assign n5460 = n2713 ^ n2430 ^ x125 ;
  assign n5461 = ~n434 & n5307 ;
  assign n5462 = n5461 ^ x62 ^ 1'b0 ;
  assign n5469 = ~n1850 & n4287 ;
  assign n5466 = n1643 ^ n544 ^ n384 ;
  assign n5465 = n1148 ^ n627 ^ n464 ;
  assign n5467 = n5466 ^ n5465 ^ n3887 ;
  assign n5468 = n5467 ^ n5424 ^ n4236 ;
  assign n5463 = n3226 ^ n962 ^ 1'b0 ;
  assign n5464 = n3643 & ~n5463 ;
  assign n5470 = n5469 ^ n5468 ^ n5464 ;
  assign n5471 = ( ~n4790 & n5462 ) | ( ~n4790 & n5470 ) | ( n5462 & n5470 ) ;
  assign n5472 = ( x114 & n639 ) | ( x114 & ~n1280 ) | ( n639 & ~n1280 ) ;
  assign n5473 = n3361 ^ n2963 ^ 1'b0 ;
  assign n5474 = n1921 & n5473 ;
  assign n5475 = n4505 ^ n1363 ^ 1'b0 ;
  assign n5476 = n5474 & n5475 ;
  assign n5477 = ( n2430 & n5472 ) | ( n2430 & n5476 ) | ( n5472 & n5476 ) ;
  assign n5478 = n750 & ~n5477 ;
  assign n5479 = ( ~n861 & n2896 ) | ( ~n861 & n5478 ) | ( n2896 & n5478 ) ;
  assign n5480 = ~n902 & n2269 ;
  assign n5481 = ~n1709 & n4067 ;
  assign n5497 = n2828 ^ n2262 ^ n369 ;
  assign n5483 = x120 & ~n242 ;
  assign n5484 = n5483 ^ x75 ^ 1'b0 ;
  assign n5485 = n3387 | n5484 ;
  assign n5486 = n1547 ^ n1120 ^ n780 ;
  assign n5487 = n5486 ^ n1399 ^ n442 ;
  assign n5488 = ( n870 & n1085 ) | ( n870 & n1359 ) | ( n1085 & n1359 ) ;
  assign n5489 = ( n229 & ~n825 ) | ( n229 & n1750 ) | ( ~n825 & n1750 ) ;
  assign n5490 = n731 & ~n5489 ;
  assign n5491 = ( ~x62 & n1130 ) | ( ~x62 & n5490 ) | ( n1130 & n5490 ) ;
  assign n5492 = n2897 & ~n5491 ;
  assign n5493 = n1747 & n5492 ;
  assign n5494 = n5488 & ~n5493 ;
  assign n5495 = n5487 & ~n5494 ;
  assign n5496 = ~n5485 & n5495 ;
  assign n5498 = n5497 ^ n5496 ^ 1'b0 ;
  assign n5499 = n927 & n5498 ;
  assign n5482 = n490 | n4602 ;
  assign n5500 = n5499 ^ n5482 ^ 1'b0 ;
  assign n5501 = ( ~n1517 & n3298 ) | ( ~n1517 & n3589 ) | ( n3298 & n3589 ) ;
  assign n5502 = n2201 | n5031 ;
  assign n5503 = n1311 & n3200 ;
  assign n5504 = ( n1910 & n2194 ) | ( n1910 & n3450 ) | ( n2194 & n3450 ) ;
  assign n5505 = n833 | n5504 ;
  assign n5506 = n1067 & ~n5505 ;
  assign n5507 = n5506 ^ n2877 ^ n1998 ;
  assign n5508 = n5507 ^ n4946 ^ n1336 ;
  assign n5509 = ( ~n2141 & n2870 ) | ( ~n2141 & n4271 ) | ( n2870 & n4271 ) ;
  assign n5510 = n1277 & ~n5509 ;
  assign n5511 = ~n255 & n799 ;
  assign n5512 = n5511 ^ n2168 ^ 1'b0 ;
  assign n5513 = n5512 ^ n4085 ^ n1568 ;
  assign n5514 = n1878 ^ n1485 ^ 1'b0 ;
  assign n5515 = n5514 ^ n4079 ^ n643 ;
  assign n5516 = ( n1230 & n2072 ) | ( n1230 & n5515 ) | ( n2072 & n5515 ) ;
  assign n5517 = n5516 ^ n5321 ^ 1'b0 ;
  assign n5518 = n1984 & n5517 ;
  assign n5521 = n2998 ^ n1559 ^ n1375 ;
  assign n5522 = n1377 & ~n2190 ;
  assign n5523 = ( n2221 & n5521 ) | ( n2221 & ~n5522 ) | ( n5521 & ~n5522 ) ;
  assign n5519 = ~n1789 & n5265 ;
  assign n5520 = n4935 & n5519 ;
  assign n5524 = n5523 ^ n5520 ^ n3215 ;
  assign n5525 = n1123 ^ n192 ^ 1'b0 ;
  assign n5526 = n1810 ^ n205 ^ x70 ;
  assign n5527 = n1359 | n3854 ;
  assign n5528 = n5527 ^ n3357 ^ 1'b0 ;
  assign n5529 = n5526 & n5528 ;
  assign n5530 = ( n463 & n1161 ) | ( n463 & ~n3725 ) | ( n1161 & ~n3725 ) ;
  assign n5531 = ( n1179 & ~n2804 ) | ( n1179 & n5530 ) | ( ~n2804 & n5530 ) ;
  assign n5534 = ( n333 & n1042 ) | ( n333 & ~n1972 ) | ( n1042 & ~n1972 ) ;
  assign n5535 = n4962 & ~n5534 ;
  assign n5532 = n3324 & ~n3962 ;
  assign n5533 = ~n860 & n5532 ;
  assign n5536 = n5535 ^ n5533 ^ n2751 ;
  assign n5541 = n195 & n289 ;
  assign n5542 = n3986 & n5541 ;
  assign n5543 = ~n2823 & n5542 ;
  assign n5537 = n1529 | n2335 ;
  assign n5538 = n5537 ^ n2644 ^ 1'b0 ;
  assign n5539 = n3431 & ~n5538 ;
  assign n5540 = n5032 & n5539 ;
  assign n5544 = n5543 ^ n5540 ^ 1'b0 ;
  assign n5545 = ( x32 & n2742 ) | ( x32 & ~n5544 ) | ( n2742 & ~n5544 ) ;
  assign n5546 = n4952 ^ n2312 ^ n1173 ;
  assign n5547 = ( n3853 & n4632 ) | ( n3853 & ~n5546 ) | ( n4632 & ~n5546 ) ;
  assign n5548 = ( x94 & n5545 ) | ( x94 & ~n5547 ) | ( n5545 & ~n5547 ) ;
  assign n5557 = n1575 ^ n182 ^ n156 ;
  assign n5556 = ( n2115 & n2502 ) | ( n2115 & ~n2872 ) | ( n2502 & ~n2872 ) ;
  assign n5549 = n2739 & ~n5142 ;
  assign n5550 = n3684 ^ n3097 ^ 1'b0 ;
  assign n5551 = n5550 ^ x49 ^ 1'b0 ;
  assign n5552 = ( n3450 & n5549 ) | ( n3450 & n5551 ) | ( n5549 & n5551 ) ;
  assign n5553 = ( n458 & ~n3704 ) | ( n458 & n5552 ) | ( ~n3704 & n5552 ) ;
  assign n5554 = n4600 ^ n1125 ^ 1'b0 ;
  assign n5555 = ( n1428 & n5553 ) | ( n1428 & ~n5554 ) | ( n5553 & ~n5554 ) ;
  assign n5558 = n5557 ^ n5556 ^ n5555 ;
  assign n5559 = n2840 ^ n349 ^ 1'b0 ;
  assign n5560 = n5559 ^ n2140 ^ n1804 ;
  assign n5561 = n559 & ~n5560 ;
  assign n5562 = n1969 & n5561 ;
  assign n5563 = n3503 | n5562 ;
  assign n5564 = n5563 ^ n2353 ^ 1'b0 ;
  assign n5568 = ( x107 & n2377 ) | ( x107 & n3814 ) | ( n2377 & n3814 ) ;
  assign n5567 = n2805 & ~n3904 ;
  assign n5569 = n5568 ^ n5567 ^ 1'b0 ;
  assign n5566 = n3552 ^ n2720 ^ n2648 ;
  assign n5565 = n2635 ^ n294 ^ 1'b0 ;
  assign n5570 = n5569 ^ n5566 ^ n5565 ;
  assign n5571 = n823 & n3092 ;
  assign n5572 = n2936 & n5571 ;
  assign n5573 = ( n1086 & n5433 ) | ( n1086 & n5572 ) | ( n5433 & n5572 ) ;
  assign n5574 = ( n1763 & n2877 ) | ( n1763 & ~n5573 ) | ( n2877 & ~n5573 ) ;
  assign n5575 = ~n2113 & n2530 ;
  assign n5576 = n5575 ^ n3082 ^ 1'b0 ;
  assign n5577 = n4819 & ~n5576 ;
  assign n5578 = n5577 ^ n4841 ^ 1'b0 ;
  assign n5579 = n3106 ^ n655 ^ 1'b0 ;
  assign n5580 = ~n5578 & n5579 ;
  assign n5581 = n3871 ^ n2717 ^ 1'b0 ;
  assign n5582 = ( ~x104 & n502 ) | ( ~x104 & n718 ) | ( n502 & n718 ) ;
  assign n5583 = n5582 ^ n2551 ^ n701 ;
  assign n5584 = n1899 | n4128 ;
  assign n5585 = n5584 ^ x68 ^ 1'b0 ;
  assign n5588 = n5467 ^ n3860 ^ 1'b0 ;
  assign n5589 = n478 | n5588 ;
  assign n5586 = ( ~n604 & n1074 ) | ( ~n604 & n2585 ) | ( n1074 & n2585 ) ;
  assign n5587 = n1158 | n5586 ;
  assign n5590 = n5589 ^ n5587 ^ 1'b0 ;
  assign n5594 = n2709 ^ n1692 ^ 1'b0 ;
  assign n5595 = n5594 ^ n1772 ^ n701 ;
  assign n5596 = n1400 ^ n774 ^ 1'b0 ;
  assign n5597 = n5341 ^ n1573 ^ 1'b0 ;
  assign n5598 = n5596 & ~n5597 ;
  assign n5599 = ( n2380 & n5595 ) | ( n2380 & n5598 ) | ( n5595 & n5598 ) ;
  assign n5600 = ~n1600 & n5599 ;
  assign n5601 = ~n3790 & n5600 ;
  assign n5591 = ( n494 & n2376 ) | ( n494 & n3184 ) | ( n2376 & n3184 ) ;
  assign n5592 = n2283 & n5591 ;
  assign n5593 = n5592 ^ n2917 ^ 1'b0 ;
  assign n5602 = n5601 ^ n5593 ^ n2319 ;
  assign n5603 = ( n1934 & ~n2070 ) | ( n1934 & n5602 ) | ( ~n2070 & n5602 ) ;
  assign n5604 = ( n689 & n1953 ) | ( n689 & n3952 ) | ( n1953 & n3952 ) ;
  assign n5605 = n5604 ^ n1767 ^ 1'b0 ;
  assign n5608 = n944 & n2941 ;
  assign n5609 = n5608 ^ n3456 ^ 1'b0 ;
  assign n5607 = n3035 & ~n3597 ;
  assign n5610 = n5609 ^ n5607 ^ 1'b0 ;
  assign n5606 = n494 & n1543 ;
  assign n5611 = n5610 ^ n5606 ^ 1'b0 ;
  assign n5612 = n5244 ^ n3323 ^ n3321 ;
  assign n5613 = ( n1320 & n2894 ) | ( n1320 & n3034 ) | ( n2894 & n3034 ) ;
  assign n5614 = n2238 & ~n4302 ;
  assign n5615 = n2405 & n5614 ;
  assign n5616 = ( n2448 & n2611 ) | ( n2448 & ~n5615 ) | ( n2611 & ~n5615 ) ;
  assign n5617 = ~n5613 & n5616 ;
  assign n5618 = n5617 ^ n4008 ^ 1'b0 ;
  assign n5619 = n5618 ^ n1031 ^ 1'b0 ;
  assign n5620 = ~n5612 & n5619 ;
  assign n5621 = ( n5605 & ~n5611 ) | ( n5605 & n5620 ) | ( ~n5611 & n5620 ) ;
  assign n5622 = n5312 ^ n1508 ^ 1'b0 ;
  assign n5623 = n4034 ^ n2600 ^ 1'b0 ;
  assign n5624 = n2464 ^ n1713 ^ n910 ;
  assign n5625 = n1572 & ~n5624 ;
  assign n5626 = ~n5623 & n5625 ;
  assign n5627 = ( ~n3647 & n5622 ) | ( ~n3647 & n5626 ) | ( n5622 & n5626 ) ;
  assign n5628 = n5594 ^ n1269 ^ n1074 ;
  assign n5629 = n5628 ^ n1718 ^ 1'b0 ;
  assign n5630 = n4629 ^ n1822 ^ n862 ;
  assign n5639 = n3887 ^ n3430 ^ n1306 ;
  assign n5631 = ~n1512 & n1643 ;
  assign n5632 = n5631 ^ n3941 ^ 1'b0 ;
  assign n5633 = n901 | n5632 ;
  assign n5634 = n5633 ^ n4859 ^ n2872 ;
  assign n5635 = n4739 ^ n2162 ^ n1896 ;
  assign n5636 = ~n2800 & n5635 ;
  assign n5637 = n5636 ^ n1177 ^ 1'b0 ;
  assign n5638 = ( n3022 & ~n5634 ) | ( n3022 & n5637 ) | ( ~n5634 & n5637 ) ;
  assign n5640 = n5639 ^ n5638 ^ 1'b0 ;
  assign n5641 = n5630 & n5640 ;
  assign n5644 = ( n721 & n1939 ) | ( n721 & n2264 ) | ( n1939 & n2264 ) ;
  assign n5645 = n1629 ^ n1627 ^ 1'b0 ;
  assign n5646 = ~n5644 & n5645 ;
  assign n5643 = n1068 | n5433 ;
  assign n5642 = n5168 ^ n3843 ^ n1155 ;
  assign n5647 = n5646 ^ n5643 ^ n5642 ;
  assign n5658 = ( n258 & n1215 ) | ( n258 & n2124 ) | ( n1215 & n2124 ) ;
  assign n5659 = ~x86 & n5658 ;
  assign n5650 = n3595 ^ n2060 ^ n453 ;
  assign n5651 = n5650 ^ n3125 ^ n2049 ;
  assign n5652 = n5651 ^ n2349 ^ n1589 ;
  assign n5653 = n2184 ^ n1246 ^ 1'b0 ;
  assign n5654 = ~n3226 & n5653 ;
  assign n5655 = n5654 ^ n5389 ^ x83 ;
  assign n5656 = n5655 ^ n2239 ^ n1494 ;
  assign n5657 = n5652 | n5656 ;
  assign n5648 = n4547 ^ n3887 ^ n2179 ;
  assign n5649 = n5648 ^ n3040 ^ n1394 ;
  assign n5660 = n5659 ^ n5657 ^ n5649 ;
  assign n5662 = n5025 ^ n4602 ^ n1757 ;
  assign n5663 = n2362 & n5662 ;
  assign n5661 = ( n1384 & ~n3173 ) | ( n1384 & n4882 ) | ( ~n3173 & n4882 ) ;
  assign n5664 = n5663 ^ n5661 ^ n5223 ;
  assign n5665 = ( n2026 & n3583 ) | ( n2026 & n4503 ) | ( n3583 & n4503 ) ;
  assign n5667 = n3591 & ~n5036 ;
  assign n5666 = n1072 | n3147 ;
  assign n5668 = n5667 ^ n5666 ^ 1'b0 ;
  assign n5669 = n2238 ^ n1228 ^ n1133 ;
  assign n5670 = ~x115 & n260 ;
  assign n5671 = ( n2040 & n5669 ) | ( n2040 & n5670 ) | ( n5669 & n5670 ) ;
  assign n5672 = ( n1207 & n5668 ) | ( n1207 & ~n5671 ) | ( n5668 & ~n5671 ) ;
  assign n5673 = n5672 ^ n2529 ^ 1'b0 ;
  assign n5674 = n5581 & n5673 ;
  assign n5675 = ( n499 & n1171 ) | ( n499 & ~n2518 ) | ( n1171 & ~n2518 ) ;
  assign n5676 = n1349 ^ n393 ^ 1'b0 ;
  assign n5677 = n5675 & ~n5676 ;
  assign n5678 = n3005 & n5341 ;
  assign n5679 = n1459 & ~n2668 ;
  assign n5680 = ( x75 & ~n5678 ) | ( x75 & n5679 ) | ( ~n5678 & n5679 ) ;
  assign n5681 = ( ~n2840 & n5677 ) | ( ~n2840 & n5680 ) | ( n5677 & n5680 ) ;
  assign n5682 = n5525 ^ n3195 ^ n1857 ;
  assign n5683 = n5682 ^ n4304 ^ n1340 ;
  assign n5684 = ( n2098 & n4388 ) | ( n2098 & n5683 ) | ( n4388 & n5683 ) ;
  assign n5687 = n1834 ^ n984 ^ n275 ;
  assign n5685 = ( n3108 & n3473 ) | ( n3108 & ~n4333 ) | ( n3473 & ~n4333 ) ;
  assign n5686 = n5685 ^ n4459 ^ n1282 ;
  assign n5688 = n5687 ^ n5686 ^ n4037 ;
  assign n5693 = n2903 ^ x78 ^ 1'b0 ;
  assign n5694 = n4563 | n5693 ;
  assign n5690 = ( n296 & ~n440 ) | ( n296 & n3081 ) | ( ~n440 & n3081 ) ;
  assign n5691 = n3173 & ~n5690 ;
  assign n5692 = n3413 & n5691 ;
  assign n5689 = n3872 ^ n2140 ^ n273 ;
  assign n5695 = n5694 ^ n5692 ^ n5689 ;
  assign n5696 = n5695 ^ n4706 ^ n2919 ;
  assign n5697 = n3242 | n5426 ;
  assign n5702 = n1322 ^ n1162 ^ 1'b0 ;
  assign n5698 = n2024 ^ n835 ^ n605 ;
  assign n5699 = n4761 ^ n2405 ^ 1'b0 ;
  assign n5700 = n5698 & n5699 ;
  assign n5701 = n5700 ^ n3136 ^ 1'b0 ;
  assign n5703 = n5702 ^ n5701 ^ 1'b0 ;
  assign n5704 = ( n743 & n2960 ) | ( n743 & n5286 ) | ( n2960 & n5286 ) ;
  assign n5705 = ( n616 & n4294 ) | ( n616 & n5704 ) | ( n4294 & n5704 ) ;
  assign n5706 = n2339 & ~n5705 ;
  assign n5712 = x13 & n261 ;
  assign n5713 = n5712 ^ n493 ^ 1'b0 ;
  assign n5710 = n1635 ^ n905 ^ 1'b0 ;
  assign n5711 = n5710 ^ n5149 ^ n4673 ;
  assign n5708 = x115 & ~n2047 ;
  assign n5709 = n5708 ^ n1220 ^ 1'b0 ;
  assign n5714 = n5713 ^ n5711 ^ n5709 ;
  assign n5707 = n2707 ^ x85 ^ 1'b0 ;
  assign n5715 = n5714 ^ n5707 ^ n2085 ;
  assign n5717 = n4815 ^ n2239 ^ n562 ;
  assign n5716 = ( ~n760 & n1703 ) | ( ~n760 & n3579 ) | ( n1703 & n3579 ) ;
  assign n5718 = n5717 ^ n5716 ^ n1657 ;
  assign n5719 = ( n4205 & ~n4273 ) | ( n4205 & n5718 ) | ( ~n4273 & n5718 ) ;
  assign n5720 = n640 & n5719 ;
  assign n5721 = n5328 & n5720 ;
  assign n5722 = n387 & ~n5100 ;
  assign n5723 = n2588 | n3664 ;
  assign n5724 = ( n511 & n934 ) | ( n511 & ~n2031 ) | ( n934 & ~n2031 ) ;
  assign n5725 = n5724 ^ n3197 ^ 1'b0 ;
  assign n5726 = ( n2732 & n5381 ) | ( n2732 & n5725 ) | ( n5381 & n5725 ) ;
  assign n5727 = n4342 & n5726 ;
  assign n5728 = ( ~n5722 & n5723 ) | ( ~n5722 & n5727 ) | ( n5723 & n5727 ) ;
  assign n5729 = n4586 ^ n2002 ^ 1'b0 ;
  assign n5730 = x99 & ~n793 ;
  assign n5731 = ( n623 & ~n4294 ) | ( n623 & n5730 ) | ( ~n4294 & n5730 ) ;
  assign n5732 = n5731 ^ n5305 ^ n1986 ;
  assign n5733 = ~n5646 & n5732 ;
  assign n5737 = n4111 ^ n3070 ^ n1661 ;
  assign n5738 = n5737 ^ n231 ^ 1'b0 ;
  assign n5735 = ( n1759 & n2688 ) | ( n1759 & n3315 ) | ( n2688 & n3315 ) ;
  assign n5734 = n4796 ^ n4746 ^ n1646 ;
  assign n5736 = n5735 ^ n5734 ^ n2491 ;
  assign n5739 = n5738 ^ n5736 ^ n5007 ;
  assign n5743 = n258 & n4175 ;
  assign n5744 = n5743 ^ n724 ^ 1'b0 ;
  assign n5741 = ( x93 & n3494 ) | ( x93 & ~n3682 ) | ( n3494 & ~n3682 ) ;
  assign n5740 = ( ~n202 & n247 ) | ( ~n202 & n1148 ) | ( n247 & n1148 ) ;
  assign n5742 = n5741 ^ n5740 ^ n1761 ;
  assign n5745 = n5744 ^ n5742 ^ 1'b0 ;
  assign n5746 = n336 | n5745 ;
  assign n5752 = x100 & n378 ;
  assign n5753 = n2147 & n5752 ;
  assign n5747 = n214 & n3102 ;
  assign n5748 = n1705 & n5747 ;
  assign n5749 = n2919 | n5748 ;
  assign n5750 = n1463 | n5749 ;
  assign n5751 = n5750 ^ n1647 ^ n1416 ;
  assign n5754 = n5753 ^ n5751 ^ 1'b0 ;
  assign n5755 = n5754 ^ n5053 ^ 1'b0 ;
  assign n5756 = n5746 | n5755 ;
  assign n5758 = ( n1632 & n3275 ) | ( n1632 & n5279 ) | ( n3275 & n5279 ) ;
  assign n5757 = n3576 ^ n2087 ^ n163 ;
  assign n5759 = n5758 ^ n5757 ^ n734 ;
  assign n5760 = ( n2903 & ~n3941 ) | ( n2903 & n5037 ) | ( ~n3941 & n5037 ) ;
  assign n5761 = n955 & ~n2784 ;
  assign n5762 = n5761 ^ n4366 ^ 1'b0 ;
  assign n5763 = ( n2302 & n2894 ) | ( n2302 & n5359 ) | ( n2894 & n5359 ) ;
  assign n5764 = n4191 ^ n2579 ^ 1'b0 ;
  assign n5765 = n1787 & n5764 ;
  assign n5766 = ( n509 & ~n862 ) | ( n509 & n5765 ) | ( ~n862 & n5765 ) ;
  assign n5767 = ( n1343 & n2330 ) | ( n1343 & n3169 ) | ( n2330 & n3169 ) ;
  assign n5768 = x72 & ~n1877 ;
  assign n5769 = n5768 ^ n1971 ^ 1'b0 ;
  assign n5770 = n5767 & n5769 ;
  assign n5771 = n5770 ^ n3822 ^ 1'b0 ;
  assign n5772 = n4878 ^ n340 ^ 1'b0 ;
  assign n5773 = n636 & ~n5772 ;
  assign n5774 = n3311 ^ x121 ^ 1'b0 ;
  assign n5775 = ( n3165 & n3215 ) | ( n3165 & ~n4925 ) | ( n3215 & ~n4925 ) ;
  assign n5776 = n5775 ^ n4341 ^ 1'b0 ;
  assign n5777 = n4097 ^ n352 ^ 1'b0 ;
  assign n5778 = n5777 ^ n4740 ^ n200 ;
  assign n5783 = ( n547 & n3641 ) | ( n547 & ~n5241 ) | ( n3641 & ~n5241 ) ;
  assign n5779 = n2028 ^ n695 ^ 1'b0 ;
  assign n5780 = n4341 | n5779 ;
  assign n5781 = n1347 & ~n5780 ;
  assign n5782 = n5781 ^ n668 ^ 1'b0 ;
  assign n5784 = n5783 ^ n5782 ^ 1'b0 ;
  assign n5785 = n2798 & ~n5784 ;
  assign n5786 = n5778 & n5785 ;
  assign n5787 = n1482 & ~n4597 ;
  assign n5788 = ( ~n214 & n4934 ) | ( ~n214 & n5787 ) | ( n4934 & n5787 ) ;
  assign n5789 = n3934 ^ n3623 ^ n3190 ;
  assign n5790 = n3883 ^ n3055 ^ n2561 ;
  assign n5791 = ~n573 & n5790 ;
  assign n5792 = n5791 ^ n755 ^ 1'b0 ;
  assign n5793 = n4492 ^ n2712 ^ n605 ;
  assign n5794 = n5793 ^ n2771 ^ n2667 ;
  assign n5795 = n482 & n3885 ;
  assign n5796 = ~n524 & n5795 ;
  assign n5797 = ( n2688 & ~n4830 ) | ( n2688 & n5796 ) | ( ~n4830 & n5796 ) ;
  assign n5799 = n1421 ^ n820 ^ 1'b0 ;
  assign n5800 = n5710 | n5799 ;
  assign n5801 = n5800 ^ n3613 ^ 1'b0 ;
  assign n5798 = ( n963 & n1862 ) | ( n963 & n3458 ) | ( n1862 & n3458 ) ;
  assign n5802 = n5801 ^ n5798 ^ n3251 ;
  assign n5803 = n2570 & ~n5802 ;
  assign n5804 = n5803 ^ n583 ^ 1'b0 ;
  assign n5805 = ( n5106 & n5797 ) | ( n5106 & ~n5804 ) | ( n5797 & ~n5804 ) ;
  assign n5806 = x74 & ~n1228 ;
  assign n5807 = ~n341 & n5806 ;
  assign n5808 = n5807 ^ n739 ^ x62 ;
  assign n5809 = n1959 & ~n5808 ;
  assign n5810 = n5809 ^ n2823 ^ 1'b0 ;
  assign n5811 = n2482 & ~n5810 ;
  assign n5812 = ~n2955 & n5811 ;
  assign n5821 = ( ~n808 & n1863 ) | ( ~n808 & n3509 ) | ( n1863 & n3509 ) ;
  assign n5822 = x76 & ~n5821 ;
  assign n5823 = n5822 ^ n2375 ^ 1'b0 ;
  assign n5824 = n5199 | n5823 ;
  assign n5817 = n4610 ^ n3053 ^ 1'b0 ;
  assign n5818 = ( ~n2380 & n3799 ) | ( ~n2380 & n5817 ) | ( n3799 & n5817 ) ;
  assign n5813 = n2309 | n3603 ;
  assign n5814 = n277 & n5813 ;
  assign n5815 = n5814 ^ n647 ^ 1'b0 ;
  assign n5816 = n923 | n5815 ;
  assign n5819 = n5818 ^ n5816 ^ n2685 ;
  assign n5820 = n5819 ^ n2479 ^ n1511 ;
  assign n5825 = n5824 ^ n5820 ^ n526 ;
  assign n5826 = n1388 ^ n347 ^ 1'b0 ;
  assign n5827 = n4834 ^ n2430 ^ n2146 ;
  assign n5828 = ( ~n1047 & n1877 ) | ( ~n1047 & n5827 ) | ( n1877 & n5827 ) ;
  assign n5829 = ( n161 & n991 ) | ( n161 & ~n5828 ) | ( n991 & ~n5828 ) ;
  assign n5830 = ( n1517 & ~n4318 ) | ( n1517 & n5829 ) | ( ~n4318 & n5829 ) ;
  assign n5831 = n5491 ^ n1601 ^ 1'b0 ;
  assign n5832 = n4967 | n5831 ;
  assign n5833 = n2377 ^ n780 ^ n762 ;
  assign n5834 = ( n4789 & n5167 ) | ( n4789 & ~n5833 ) | ( n5167 & ~n5833 ) ;
  assign n5836 = ( ~n3869 & n4152 ) | ( ~n3869 & n4690 ) | ( n4152 & n4690 ) ;
  assign n5835 = ( ~n1356 & n2219 ) | ( ~n1356 & n2235 ) | ( n2219 & n2235 ) ;
  assign n5837 = n5836 ^ n5835 ^ 1'b0 ;
  assign n5838 = n5706 & ~n5837 ;
  assign n5839 = n423 & ~n5559 ;
  assign n5840 = n5839 ^ n4699 ^ 1'b0 ;
  assign n5841 = ( x38 & ~n4139 ) | ( x38 & n4746 ) | ( ~n4139 & n4746 ) ;
  assign n5842 = ~n4006 & n5841 ;
  assign n5843 = ( n4735 & n5840 ) | ( n4735 & n5842 ) | ( n5840 & n5842 ) ;
  assign n5844 = n5843 ^ n3176 ^ n1904 ;
  assign n5845 = ( n4461 & ~n4574 ) | ( n4461 & n5062 ) | ( ~n4574 & n5062 ) ;
  assign n5846 = n1673 ^ n1203 ^ 1'b0 ;
  assign n5847 = n5149 & n5846 ;
  assign n5848 = n5847 ^ n488 ^ 1'b0 ;
  assign n5849 = ( n1346 & n2102 ) | ( n1346 & ~n5848 ) | ( n2102 & ~n5848 ) ;
  assign n5850 = ~n553 & n973 ;
  assign n5851 = n5850 ^ n5414 ^ 1'b0 ;
  assign n5852 = ~n1716 & n5851 ;
  assign n5853 = n5852 ^ n4186 ^ 1'b0 ;
  assign n5854 = ~n5849 & n5853 ;
  assign n5855 = n2827 ^ n213 ^ 1'b0 ;
  assign n5856 = n1808 & n5855 ;
  assign n5857 = ~n1189 & n5856 ;
  assign n5858 = ( ~x82 & n1373 ) | ( ~x82 & n4739 ) | ( n1373 & n4739 ) ;
  assign n5859 = ( n5854 & n5857 ) | ( n5854 & ~n5858 ) | ( n5857 & ~n5858 ) ;
  assign n5860 = n5197 ^ n1663 ^ 1'b0 ;
  assign n5861 = n4878 ^ n3717 ^ n1525 ;
  assign n5863 = ( n509 & n2401 ) | ( n509 & n5121 ) | ( n2401 & n5121 ) ;
  assign n5862 = n1966 ^ n1188 ^ 1'b0 ;
  assign n5864 = n5863 ^ n5862 ^ n516 ;
  assign n5865 = n4806 & ~n5864 ;
  assign n5867 = x41 & ~n3416 ;
  assign n5868 = n5867 ^ n1713 ^ 1'b0 ;
  assign n5866 = n2762 | n4785 ;
  assign n5869 = n5868 ^ n5866 ^ 1'b0 ;
  assign n5870 = n5865 | n5869 ;
  assign n5871 = n894 ^ n577 ^ x60 ;
  assign n5872 = ( ~n1882 & n2485 ) | ( ~n1882 & n5871 ) | ( n2485 & n5871 ) ;
  assign n5873 = n5391 ^ n1588 ^ 1'b0 ;
  assign n5876 = n2957 ^ n2622 ^ n1721 ;
  assign n5874 = ( n912 & ~n2847 ) | ( n912 & n4911 ) | ( ~n2847 & n4911 ) ;
  assign n5875 = n2002 | n5874 ;
  assign n5877 = n5876 ^ n5875 ^ n4508 ;
  assign n5878 = n2602 ^ n2228 ^ 1'b0 ;
  assign n5879 = n5022 | n5878 ;
  assign n5880 = n5877 | n5879 ;
  assign n5881 = ~n1924 & n2165 ;
  assign n5882 = n5881 ^ x110 ^ 1'b0 ;
  assign n5883 = n1190 ^ n843 ^ n190 ;
  assign n5884 = n5883 ^ n665 ^ 1'b0 ;
  assign n5885 = n5882 | n5884 ;
  assign n5886 = n5885 ^ n4356 ^ n386 ;
  assign n5889 = n3833 ^ n1354 ^ 1'b0 ;
  assign n5890 = ( n2212 & n4034 ) | ( n2212 & ~n5889 ) | ( n4034 & ~n5889 ) ;
  assign n5887 = ( n1919 & n2486 ) | ( n1919 & ~n4764 ) | ( n2486 & ~n4764 ) ;
  assign n5888 = n5836 | n5887 ;
  assign n5891 = n5890 ^ n5888 ^ 1'b0 ;
  assign n5892 = ( ~n132 & n2145 ) | ( ~n132 & n2702 ) | ( n2145 & n2702 ) ;
  assign n5893 = ~n386 & n2165 ;
  assign n5894 = n5893 ^ n1121 ^ 1'b0 ;
  assign n5895 = n5894 ^ n1343 ^ 1'b0 ;
  assign n5896 = n1945 & n5895 ;
  assign n5897 = ( n1051 & n5892 ) | ( n1051 & n5896 ) | ( n5892 & n5896 ) ;
  assign n5898 = n840 & ~n5897 ;
  assign n5899 = n3580 & ~n3801 ;
  assign n5900 = ( x32 & n3188 ) | ( x32 & ~n3278 ) | ( n3188 & ~n3278 ) ;
  assign n5901 = ~n1376 & n5900 ;
  assign n5902 = n5734 & n5901 ;
  assign n5903 = n1123 ^ n820 ^ 1'b0 ;
  assign n5904 = n5594 & ~n5903 ;
  assign n5905 = n2953 ^ n738 ^ n333 ;
  assign n5914 = n305 ^ x24 ^ 1'b0 ;
  assign n5915 = n408 & n5914 ;
  assign n5916 = n5915 ^ n3776 ^ n1308 ;
  assign n5906 = ( ~n329 & n1240 ) | ( ~n329 & n3141 ) | ( n1240 & n3141 ) ;
  assign n5910 = ( n1680 & ~n1833 ) | ( n1680 & n4649 ) | ( ~n1833 & n4649 ) ;
  assign n5907 = n695 & n2220 ;
  assign n5908 = ~n218 & n5907 ;
  assign n5909 = ( ~n897 & n3546 ) | ( ~n897 & n5908 ) | ( n3546 & n5908 ) ;
  assign n5911 = n5910 ^ n5909 ^ 1'b0 ;
  assign n5912 = n5906 & n5911 ;
  assign n5913 = ( n352 & ~n5106 ) | ( n352 & n5912 ) | ( ~n5106 & n5912 ) ;
  assign n5917 = n5916 ^ n5913 ^ n4919 ;
  assign n5918 = n3962 ^ n3319 ^ 1'b0 ;
  assign n5919 = n349 & ~n2779 ;
  assign n5920 = x10 & ~n5919 ;
  assign n5921 = n5920 ^ n4134 ^ 1'b0 ;
  assign n5922 = n5921 ^ n4994 ^ n1417 ;
  assign n5923 = n355 & n488 ;
  assign n5924 = n5923 ^ n1893 ^ 1'b0 ;
  assign n5925 = n5924 ^ n1973 ^ n529 ;
  assign n5926 = n4734 ^ n1914 ^ x116 ;
  assign n5927 = n5926 ^ n4557 ^ x1 ;
  assign n5928 = ( n414 & n4269 ) | ( n414 & ~n4878 ) | ( n4269 & ~n4878 ) ;
  assign n5929 = n941 & ~n5928 ;
  assign n5930 = n418 ^ n157 ^ 1'b0 ;
  assign n5932 = n2389 | n4604 ;
  assign n5931 = n3192 ^ n131 ^ x37 ;
  assign n5933 = n5932 ^ n5931 ^ n4768 ;
  assign n5934 = n2994 ^ n2058 ^ 1'b0 ;
  assign n5935 = n4092 & n5934 ;
  assign n5936 = n292 & ~n1815 ;
  assign n5937 = ~n5935 & n5936 ;
  assign n5938 = ~n199 & n5451 ;
  assign n5939 = n5938 ^ n1350 ^ 1'b0 ;
  assign n5940 = n5939 ^ n5007 ^ n1575 ;
  assign n5944 = n1260 ^ n1199 ^ 1'b0 ;
  assign n5945 = n2283 & ~n5944 ;
  assign n5941 = n2380 | n3553 ;
  assign n5942 = n4918 & ~n5941 ;
  assign n5943 = n689 & n5942 ;
  assign n5946 = n5945 ^ n5943 ^ n319 ;
  assign n5947 = ( n2020 & n2306 ) | ( n2020 & n4366 ) | ( n2306 & n4366 ) ;
  assign n5948 = ( ~n2873 & n2983 ) | ( ~n2873 & n5089 ) | ( n2983 & n5089 ) ;
  assign n5949 = ~n5947 & n5948 ;
  assign n5950 = n5949 ^ n3687 ^ n1745 ;
  assign n5951 = n5950 ^ n5138 ^ 1'b0 ;
  assign n5952 = ~n2878 & n5951 ;
  assign n5953 = n335 | n505 ;
  assign n5954 = n613 & ~n5953 ;
  assign n5955 = n5954 ^ n3613 ^ n1659 ;
  assign n5956 = n5955 ^ n4202 ^ n1397 ;
  assign n5957 = ( n598 & n2252 ) | ( n598 & ~n3098 ) | ( n2252 & ~n3098 ) ;
  assign n5958 = ( n2144 & ~n3937 ) | ( n2144 & n5957 ) | ( ~n3937 & n5957 ) ;
  assign n5959 = ( n4282 & ~n5956 ) | ( n4282 & n5958 ) | ( ~n5956 & n5958 ) ;
  assign n5960 = n1720 ^ n753 ^ 1'b0 ;
  assign n5961 = n1574 | n3430 ;
  assign n5962 = n5945 | n5961 ;
  assign n5963 = n1640 ^ n1632 ^ n731 ;
  assign n5964 = n5962 & n5963 ;
  assign n5965 = n5964 ^ n5714 ^ 1'b0 ;
  assign n5966 = n5530 & n5534 ;
  assign n5967 = n5966 ^ n2265 ^ 1'b0 ;
  assign n5968 = ( n5960 & n5965 ) | ( n5960 & n5967 ) | ( n5965 & n5967 ) ;
  assign n5969 = ( n899 & ~n1213 ) | ( n899 & n5411 ) | ( ~n1213 & n5411 ) ;
  assign n5970 = ~n5968 & n5969 ;
  assign n5971 = ~n1632 & n5970 ;
  assign n5973 = ( n1329 & n1628 ) | ( n1329 & ~n3887 ) | ( n1628 & ~n3887 ) ;
  assign n5972 = ~n1723 & n4804 ;
  assign n5974 = n5973 ^ n5972 ^ x35 ;
  assign n5977 = n2421 ^ n1421 ^ 1'b0 ;
  assign n5978 = n1518 | n5977 ;
  assign n5979 = ( n2002 & n2902 ) | ( n2002 & ~n5978 ) | ( n2902 & ~n5978 ) ;
  assign n5975 = n359 | n3254 ;
  assign n5976 = n5975 ^ n5276 ^ n3785 ;
  assign n5980 = n5979 ^ n5976 ^ n2152 ;
  assign n5981 = ( n2338 & n5149 ) | ( n2338 & ~n5201 ) | ( n5149 & ~n5201 ) ;
  assign n5982 = n5981 ^ n1990 ^ 1'b0 ;
  assign n5983 = n5982 ^ n3316 ^ 1'b0 ;
  assign n5984 = n4979 | n5983 ;
  assign n5985 = n5650 ^ n1932 ^ n237 ;
  assign n5986 = n5985 ^ n3102 ^ n457 ;
  assign n5987 = n5986 ^ n1864 ^ n861 ;
  assign n5988 = ( n2813 & n5984 ) | ( n2813 & ~n5987 ) | ( n5984 & ~n5987 ) ;
  assign n5989 = ~n1920 & n5650 ;
  assign n5990 = n5989 ^ n1411 ^ 1'b0 ;
  assign n5991 = n2045 | n5990 ;
  assign n5992 = n498 & ~n5753 ;
  assign n5993 = ~n2267 & n5992 ;
  assign n5994 = n5993 ^ n4508 ^ n3409 ;
  assign n5995 = x24 & ~x122 ;
  assign n5998 = ~n393 & n5100 ;
  assign n5996 = n1304 ^ n382 ^ x124 ;
  assign n5997 = ~n1982 & n5996 ;
  assign n5999 = n5998 ^ n5997 ^ n3486 ;
  assign n6000 = n5445 ^ n2118 ^ 1'b0 ;
  assign n6001 = ( n408 & n1537 ) | ( n408 & n2639 ) | ( n1537 & n2639 ) ;
  assign n6002 = ( ~x15 & n3147 ) | ( ~x15 & n6001 ) | ( n3147 & n6001 ) ;
  assign n6003 = n6002 ^ n4087 ^ 1'b0 ;
  assign n6004 = n6000 & n6003 ;
  assign n6005 = ~n5999 & n6004 ;
  assign n6006 = n6005 ^ n4437 ^ 1'b0 ;
  assign n6013 = n5277 ^ n2237 ^ n1444 ;
  assign n6007 = n2754 ^ n367 ^ 1'b0 ;
  assign n6008 = n424 | n6007 ;
  assign n6009 = n224 | n1158 ;
  assign n6010 = n6008 & ~n6009 ;
  assign n6011 = n6010 ^ n3099 ^ n223 ;
  assign n6012 = n6011 ^ n1889 ^ n1754 ;
  assign n6014 = n6013 ^ n6012 ^ n4760 ;
  assign n6015 = ~n2779 & n4179 ;
  assign n6016 = n5142 ^ n317 ^ n306 ;
  assign n6017 = ( n710 & ~n4797 ) | ( n710 & n6016 ) | ( ~n4797 & n6016 ) ;
  assign n6018 = n5394 ^ n3546 ^ n2375 ;
  assign n6019 = ( ~n3600 & n6017 ) | ( ~n3600 & n6018 ) | ( n6017 & n6018 ) ;
  assign n6020 = n6019 ^ n473 ^ 1'b0 ;
  assign n6021 = n2800 & ~n6020 ;
  assign n6029 = ( x82 & n1414 ) | ( x82 & n1675 ) | ( n1414 & n1675 ) ;
  assign n6027 = ( n2174 & ~n2716 ) | ( n2174 & n3601 ) | ( ~n2716 & n3601 ) ;
  assign n6028 = n6027 ^ n3466 ^ n1513 ;
  assign n6022 = ~n393 & n2630 ;
  assign n6023 = n6022 ^ n1780 ^ 1'b0 ;
  assign n6024 = n6023 ^ n2213 ^ x3 ;
  assign n6025 = ~n4676 & n6024 ;
  assign n6026 = n6025 ^ n308 ^ 1'b0 ;
  assign n6030 = n6029 ^ n6028 ^ n6026 ;
  assign n6031 = n3989 & ~n4962 ;
  assign n6036 = n2790 ^ n1379 ^ 1'b0 ;
  assign n6037 = n2434 & ~n6036 ;
  assign n6032 = n2330 ^ n2253 ^ 1'b0 ;
  assign n6033 = n426 | n3673 ;
  assign n6034 = n6032 & ~n6033 ;
  assign n6035 = ~n2927 & n6034 ;
  assign n6038 = n6037 ^ n6035 ^ 1'b0 ;
  assign n6039 = n4677 ^ n1184 ^ 1'b0 ;
  assign n6040 = n6039 ^ n4176 ^ n2920 ;
  assign n6041 = n3856 ^ n2980 ^ n2211 ;
  assign n6042 = ( n2020 & n2860 ) | ( n2020 & n4730 ) | ( n2860 & n4730 ) ;
  assign n6043 = n6042 ^ n3592 ^ n757 ;
  assign n6044 = ( n2281 & n5133 ) | ( n2281 & n6043 ) | ( n5133 & n6043 ) ;
  assign n6045 = ( n2308 & ~n3540 ) | ( n2308 & n6044 ) | ( ~n3540 & n6044 ) ;
  assign n6046 = n5621 & n6045 ;
  assign n6047 = n6046 ^ n5826 ^ 1'b0 ;
  assign n6048 = n3103 & ~n6047 ;
  assign n6049 = n5506 ^ n3505 ^ n2141 ;
  assign n6050 = n4220 ^ x4 ^ 1'b0 ;
  assign n6051 = n6049 & ~n6050 ;
  assign n6052 = n3998 ^ n2036 ^ n950 ;
  assign n6053 = n6052 ^ n5206 ^ 1'b0 ;
  assign n6054 = n6051 & ~n6053 ;
  assign n6055 = x96 & ~n3849 ;
  assign n6056 = n6055 ^ n3801 ^ 1'b0 ;
  assign n6057 = n4384 ^ n2173 ^ n2092 ;
  assign n6058 = n6057 ^ n1589 ^ n1463 ;
  assign n6059 = n5734 ^ n594 ^ 1'b0 ;
  assign n6060 = n5206 | n6059 ;
  assign n6061 = n3761 | n6060 ;
  assign n6062 = n518 | n6061 ;
  assign n6065 = ( n423 & n4492 ) | ( n423 & ~n5048 ) | ( n4492 & ~n5048 ) ;
  assign n6063 = n3772 ^ n2750 ^ 1'b0 ;
  assign n6064 = n5276 & n6063 ;
  assign n6066 = n6065 ^ n6064 ^ n2457 ;
  assign n6067 = n4189 ^ n2314 ^ 1'b0 ;
  assign n6068 = ~n1312 & n3711 ;
  assign n6073 = ( ~n443 & n1152 ) | ( ~n443 & n1409 ) | ( n1152 & n1409 ) ;
  assign n6071 = n1247 & ~n1542 ;
  assign n6069 = n3238 ^ n2970 ^ n463 ;
  assign n6070 = n2228 & n6069 ;
  assign n6072 = n6071 ^ n6070 ^ 1'b0 ;
  assign n6074 = n6073 ^ n6072 ^ n392 ;
  assign n6075 = n6074 ^ n4860 ^ n259 ;
  assign n6076 = ~n1255 & n3277 ;
  assign n6077 = n6076 ^ n3237 ^ 1'b0 ;
  assign n6078 = ( n1465 & ~n3885 ) | ( n1465 & n6077 ) | ( ~n3885 & n6077 ) ;
  assign n6079 = ~n913 & n6078 ;
  assign n6083 = n3684 ^ n761 ^ n484 ;
  assign n6084 = n6083 ^ n350 ^ 1'b0 ;
  assign n6080 = ( x30 & n340 ) | ( x30 & ~n5465 ) | ( n340 & ~n5465 ) ;
  assign n6081 = ( n406 & n1612 ) | ( n406 & n3309 ) | ( n1612 & n3309 ) ;
  assign n6082 = ( ~n2257 & n6080 ) | ( ~n2257 & n6081 ) | ( n6080 & n6081 ) ;
  assign n6085 = n6084 ^ n6082 ^ 1'b0 ;
  assign n6086 = n175 | n2632 ;
  assign n6087 = n2293 ^ n1796 ^ n486 ;
  assign n6091 = n4645 ^ n3652 ^ n1893 ;
  assign n6092 = n1213 ^ n326 ^ 1'b0 ;
  assign n6093 = n6024 & n6092 ;
  assign n6094 = ~n6091 & n6093 ;
  assign n6088 = n5075 ^ n4223 ^ n1951 ;
  assign n6089 = n5296 & n6088 ;
  assign n6090 = n6089 ^ n2792 ^ 1'b0 ;
  assign n6095 = n6094 ^ n6090 ^ 1'b0 ;
  assign n6096 = n6087 | n6095 ;
  assign n6099 = n1184 | n2586 ;
  assign n6097 = n3714 ^ n497 ^ 1'b0 ;
  assign n6098 = n5892 | n6097 ;
  assign n6100 = n6099 ^ n6098 ^ 1'b0 ;
  assign n6106 = n424 | n2302 ;
  assign n6107 = n6106 ^ n4024 ^ n3393 ;
  assign n6104 = n4577 ^ n1609 ^ 1'b0 ;
  assign n6105 = n6104 ^ n3874 ^ n2312 ;
  assign n6108 = n6107 ^ n6105 ^ x61 ;
  assign n6101 = n809 ^ n315 ^ 1'b0 ;
  assign n6102 = n3698 & ~n6101 ;
  assign n6103 = n6102 ^ n4617 ^ 1'b0 ;
  assign n6109 = n6108 ^ n6103 ^ n6055 ;
  assign n6110 = n6109 ^ n4136 ^ 1'b0 ;
  assign n6111 = n4424 & n6110 ;
  assign n6112 = n894 & ~n2190 ;
  assign n6113 = ~n711 & n6112 ;
  assign n6114 = n2328 | n6113 ;
  assign n6115 = n6114 ^ n4640 ^ n3402 ;
  assign n6119 = x59 & n1947 ;
  assign n6120 = n1719 & n6119 ;
  assign n6116 = n1514 ^ n1494 ^ n802 ;
  assign n6117 = n6116 ^ n2070 ^ 1'b0 ;
  assign n6118 = x118 & n6117 ;
  assign n6121 = n6120 ^ n6118 ^ n359 ;
  assign n6122 = n2578 ^ n2000 ^ n1438 ;
  assign n6123 = n3615 ^ n1386 ^ n1119 ;
  assign n6124 = n3049 & ~n6123 ;
  assign n6125 = ( n400 & n424 ) | ( n400 & ~n4452 ) | ( n424 & ~n4452 ) ;
  assign n6126 = n6125 ^ n2198 ^ n2075 ;
  assign n6135 = n425 & n2126 ;
  assign n6136 = ( x97 & ~n2237 ) | ( x97 & n6135 ) | ( ~n2237 & n6135 ) ;
  assign n6137 = ~n4543 & n6136 ;
  assign n6138 = n3486 & n6137 ;
  assign n6127 = n583 ^ n490 ^ 1'b0 ;
  assign n6128 = ~n1755 & n6127 ;
  assign n6129 = n1116 ^ n588 ^ n287 ;
  assign n6130 = n6129 ^ n4314 ^ 1'b0 ;
  assign n6131 = n6128 & ~n6130 ;
  assign n6132 = n6131 ^ x30 ^ 1'b0 ;
  assign n6133 = n5404 ^ n683 ^ 1'b0 ;
  assign n6134 = ( n525 & n6132 ) | ( n525 & n6133 ) | ( n6132 & n6133 ) ;
  assign n6139 = n6138 ^ n6134 ^ x6 ;
  assign n6140 = ~n1265 & n6139 ;
  assign n6141 = n5562 ^ n1953 ^ 1'b0 ;
  assign n6142 = n4366 ^ n2172 ^ n1127 ;
  assign n6143 = n6142 ^ n2215 ^ n605 ;
  assign n6144 = n1204 | n3454 ;
  assign n6145 = n3686 & ~n6144 ;
  assign n6146 = ( n4015 & n6143 ) | ( n4015 & n6145 ) | ( n6143 & n6145 ) ;
  assign n6147 = n6146 ^ n3852 ^ 1'b0 ;
  assign n6148 = n6141 & ~n6147 ;
  assign n6149 = ( n604 & ~n2285 ) | ( n604 & n3237 ) | ( ~n2285 & n3237 ) ;
  assign n6150 = n6149 ^ n2915 ^ n1620 ;
  assign n6151 = n6150 ^ n1708 ^ 1'b0 ;
  assign n6152 = ~n1562 & n6151 ;
  assign n6153 = n6142 ^ n3467 ^ n200 ;
  assign n6154 = ( ~n1290 & n5642 ) | ( ~n1290 & n6153 ) | ( n5642 & n6153 ) ;
  assign n6155 = n1573 & ~n2305 ;
  assign n6156 = n3319 & n6155 ;
  assign n6157 = n6156 ^ n2643 ^ n465 ;
  assign n6158 = n2624 ^ n669 ^ n270 ;
  assign n6159 = n6158 ^ n4945 ^ 1'b0 ;
  assign n6160 = n1490 & ~n4143 ;
  assign n6161 = n6160 ^ n2109 ^ 1'b0 ;
  assign n6162 = n6161 ^ n365 ^ n266 ;
  assign n6165 = n2607 ^ n2392 ^ 1'b0 ;
  assign n6166 = ~n2047 & n6165 ;
  assign n6167 = ~n5724 & n6166 ;
  assign n6163 = n686 | n4186 ;
  assign n6164 = n6163 ^ n4645 ^ 1'b0 ;
  assign n6168 = n6167 ^ n6164 ^ n3120 ;
  assign n6169 = ~n6162 & n6168 ;
  assign n6170 = n6169 ^ x75 ^ 1'b0 ;
  assign n6171 = ~n2392 & n6135 ;
  assign n6172 = n4375 & n6171 ;
  assign n6173 = ( n944 & ~n1594 ) | ( n944 & n6172 ) | ( ~n1594 & n6172 ) ;
  assign n6174 = n6173 ^ n2802 ^ 1'b0 ;
  assign n6175 = n2151 ^ n1021 ^ 1'b0 ;
  assign n6176 = n3085 | n6175 ;
  assign n6177 = n6176 ^ n4139 ^ 1'b0 ;
  assign n6178 = n1402 & ~n4405 ;
  assign n6179 = n6178 ^ n2854 ^ n1299 ;
  assign n6180 = n1949 & ~n1962 ;
  assign n6195 = n2248 ^ n1961 ^ n1796 ;
  assign n6196 = n406 | n1114 ;
  assign n6197 = n6196 ^ n3580 ^ 1'b0 ;
  assign n6198 = ~n4972 & n6197 ;
  assign n6199 = ( n2379 & n6195 ) | ( n2379 & n6198 ) | ( n6195 & n6198 ) ;
  assign n6203 = n575 | n3703 ;
  assign n6200 = n5074 ^ n2930 ^ 1'b0 ;
  assign n6201 = ~n4624 & n6200 ;
  assign n6202 = n6201 ^ n1863 ^ n232 ;
  assign n6204 = n6203 ^ n6202 ^ 1'b0 ;
  assign n6205 = n6204 ^ n1136 ^ 1'b0 ;
  assign n6206 = ~n6199 & n6205 ;
  assign n6181 = n3710 ^ n1695 ^ n259 ;
  assign n6191 = ( ~n1353 & n5376 ) | ( ~n1353 & n6130 ) | ( n5376 & n6130 ) ;
  assign n6182 = ( ~n1862 & n1930 ) | ( ~n1862 & n1994 ) | ( n1930 & n1994 ) ;
  assign n6183 = n1708 | n2081 ;
  assign n6184 = n1862 ^ n241 ^ x23 ;
  assign n6185 = n4349 ^ n3587 ^ n865 ;
  assign n6186 = ( ~n995 & n1566 ) | ( ~n995 & n2247 ) | ( n1566 & n2247 ) ;
  assign n6187 = ( ~n1781 & n6185 ) | ( ~n1781 & n6186 ) | ( n6185 & n6186 ) ;
  assign n6188 = n6184 & ~n6187 ;
  assign n6189 = ~n6183 & n6188 ;
  assign n6190 = n6182 & ~n6189 ;
  assign n6192 = n6191 ^ n6190 ^ 1'b0 ;
  assign n6193 = n6192 ^ n1238 ^ 1'b0 ;
  assign n6194 = ~n6181 & n6193 ;
  assign n6207 = n6206 ^ n6194 ^ n2054 ;
  assign n6208 = n4435 ^ n3949 ^ n661 ;
  assign n6211 = n4151 ^ n1652 ^ 1'b0 ;
  assign n6212 = n4111 & n6211 ;
  assign n6213 = n6212 ^ n2665 ^ n2121 ;
  assign n6209 = n2750 ^ n1145 ^ n1074 ;
  assign n6210 = n5885 | n6209 ;
  assign n6214 = n6213 ^ n6210 ^ n4660 ;
  assign n6215 = n4794 ^ n2802 ^ n1874 ;
  assign n6216 = n6215 ^ n4846 ^ n2965 ;
  assign n6217 = ~n741 & n3910 ;
  assign n6218 = n6217 ^ n2108 ^ 1'b0 ;
  assign n6219 = ( n5150 & ~n6091 ) | ( n5150 & n6218 ) | ( ~n6091 & n6218 ) ;
  assign n6220 = n6219 ^ n4750 ^ 1'b0 ;
  assign n6221 = ~n2335 & n6220 ;
  assign n6222 = ( x9 & n591 ) | ( x9 & ~n6221 ) | ( n591 & ~n6221 ) ;
  assign n6223 = n1410 & ~n6222 ;
  assign n6224 = n591 & ~n1642 ;
  assign n6225 = n3877 & n6224 ;
  assign n6226 = n6225 ^ n293 ^ 1'b0 ;
  assign n6227 = ( n3119 & n4567 ) | ( n3119 & n6226 ) | ( n4567 & n6226 ) ;
  assign n6228 = ( n393 & n3851 ) | ( n393 & n6227 ) | ( n3851 & n6227 ) ;
  assign n6233 = n2436 & n3409 ;
  assign n6234 = ( n1494 & ~n3691 ) | ( n1494 & n5201 ) | ( ~n3691 & n5201 ) ;
  assign n6235 = n6233 | n6234 ;
  assign n6230 = n2149 & ~n2486 ;
  assign n6229 = x2 | n317 ;
  assign n6231 = n6230 ^ n6229 ^ n2612 ;
  assign n6232 = n6231 ^ n4513 ^ n4428 ;
  assign n6236 = n6235 ^ n6232 ^ n1529 ;
  assign n6237 = ( x75 & n1482 ) | ( x75 & n3687 ) | ( n1482 & n3687 ) ;
  assign n6239 = ( ~n991 & n1884 ) | ( ~n991 & n3592 ) | ( n1884 & n3592 ) ;
  assign n6240 = ( n745 & n914 ) | ( n745 & n6239 ) | ( n914 & n6239 ) ;
  assign n6238 = ( ~n200 & n389 ) | ( ~n200 & n2531 ) | ( n389 & n2531 ) ;
  assign n6241 = n6240 ^ n6238 ^ 1'b0 ;
  assign n6242 = n6237 & n6241 ;
  assign n6243 = ( n2969 & n4320 ) | ( n2969 & n6242 ) | ( n4320 & n6242 ) ;
  assign n6244 = ( n4881 & ~n6236 ) | ( n4881 & n6243 ) | ( ~n6236 & n6243 ) ;
  assign n6251 = n627 & ~n802 ;
  assign n6245 = ~n763 & n775 ;
  assign n6246 = ~n2672 & n6245 ;
  assign n6247 = n1868 & n6246 ;
  assign n6248 = x13 | n6247 ;
  assign n6249 = n3377 & n6248 ;
  assign n6250 = n6249 ^ n2311 ^ 1'b0 ;
  assign n6252 = n6251 ^ n6250 ^ n2750 ;
  assign n6253 = n1042 & ~n3062 ;
  assign n6254 = ( n1644 & ~n4003 ) | ( n1644 & n4907 ) | ( ~n4003 & n4907 ) ;
  assign n6261 = n3772 ^ n2552 ^ n1023 ;
  assign n6262 = n1842 | n6261 ;
  assign n6263 = n2031 & ~n6262 ;
  assign n6258 = n2646 ^ n1887 ^ 1'b0 ;
  assign n6259 = n4313 ^ n2262 ^ 1'b0 ;
  assign n6260 = ~n6258 & n6259 ;
  assign n6256 = n2070 ^ n1887 ^ n335 ;
  assign n6255 = n2702 | n4919 ;
  assign n6257 = n6256 ^ n6255 ^ 1'b0 ;
  assign n6264 = n6263 ^ n6260 ^ n6257 ;
  assign n6267 = ( ~n451 & n1982 ) | ( ~n451 & n2262 ) | ( n1982 & n2262 ) ;
  assign n6268 = n1527 & n6267 ;
  assign n6265 = n1572 & ~n1753 ;
  assign n6266 = n3031 & n6265 ;
  assign n6269 = n6268 ^ n6266 ^ 1'b0 ;
  assign n6270 = n1377 ^ n406 ^ 1'b0 ;
  assign n6271 = n5530 ^ n4496 ^ 1'b0 ;
  assign n6272 = n4343 & n6271 ;
  assign n6273 = n2972 ^ n2912 ^ n820 ;
  assign n6274 = n6101 ^ n2507 ^ 1'b0 ;
  assign n6275 = ( n203 & ~n953 ) | ( n203 & n4103 ) | ( ~n953 & n4103 ) ;
  assign n6276 = ( ~n581 & n3285 ) | ( ~n581 & n6275 ) | ( n3285 & n6275 ) ;
  assign n6277 = n6143 ^ n4743 ^ 1'b0 ;
  assign n6280 = n566 & ~n1189 ;
  assign n6279 = x85 & ~n3053 ;
  assign n6278 = ( n291 & ~n1493 ) | ( n291 & n3732 ) | ( ~n1493 & n3732 ) ;
  assign n6281 = n6280 ^ n6279 ^ n6278 ;
  assign n6282 = n6281 ^ n1231 ^ 1'b0 ;
  assign n6283 = n4629 ^ n1450 ^ 1'b0 ;
  assign n6284 = n5868 | n6283 ;
  assign n6286 = n4473 ^ n2357 ^ 1'b0 ;
  assign n6287 = n1330 | n6286 ;
  assign n6288 = n6287 ^ n1287 ^ n818 ;
  assign n6289 = n4645 ^ x38 ^ 1'b0 ;
  assign n6290 = n6289 ^ n762 ^ n659 ;
  assign n6291 = ( n2563 & n6288 ) | ( n2563 & n6290 ) | ( n6288 & n6290 ) ;
  assign n6285 = n2946 ^ n494 ^ n139 ;
  assign n6292 = n6291 ^ n6285 ^ 1'b0 ;
  assign n6293 = ~n6284 & n6292 ;
  assign n6294 = n4059 ^ n835 ^ 1'b0 ;
  assign n6295 = n6294 ^ n2375 ^ x22 ;
  assign n6297 = ( n205 & n1396 ) | ( n205 & ~n3912 ) | ( n1396 & ~n3912 ) ;
  assign n6296 = n1475 | n2464 ;
  assign n6298 = n6297 ^ n6296 ^ 1'b0 ;
  assign n6299 = ( ~n132 & n160 ) | ( ~n132 & n6298 ) | ( n160 & n6298 ) ;
  assign n6300 = n4595 ^ n1578 ^ 1'b0 ;
  assign n6301 = n2137 ^ n1601 ^ 1'b0 ;
  assign n6302 = n1785 & n6301 ;
  assign n6303 = n6288 & n6302 ;
  assign n6304 = n6303 ^ n240 ^ 1'b0 ;
  assign n6305 = n5430 ^ n4168 ^ n1961 ;
  assign n6306 = n6305 ^ n6018 ^ 1'b0 ;
  assign n6307 = n6306 ^ n4624 ^ n2669 ;
  assign n6308 = n4288 ^ n1500 ^ 1'b0 ;
  assign n6309 = n1996 | n6034 ;
  assign n6310 = n6309 ^ n5325 ^ x103 ;
  assign n6311 = n3160 ^ n2775 ^ n1638 ;
  assign n6312 = n6311 ^ n5337 ^ n3685 ;
  assign n6321 = n3714 ^ n3279 ^ 1'b0 ;
  assign n6313 = n5027 ^ n3413 ^ n1155 ;
  assign n6314 = ( n908 & ~n1489 ) | ( n908 & n3579 ) | ( ~n1489 & n3579 ) ;
  assign n6315 = n2859 ^ n2083 ^ 1'b0 ;
  assign n6316 = n6314 & n6315 ;
  assign n6317 = x75 & n3713 ;
  assign n6318 = ~n6000 & n6317 ;
  assign n6319 = n6316 & ~n6318 ;
  assign n6320 = n6313 & n6319 ;
  assign n6322 = n6321 ^ n6320 ^ x85 ;
  assign n6323 = n4886 ^ n1902 ^ 1'b0 ;
  assign n6324 = ~n3648 & n6323 ;
  assign n6325 = n1743 ^ x12 ^ 1'b0 ;
  assign n6326 = n3684 & n6325 ;
  assign n6327 = n6326 ^ n2844 ^ 1'b0 ;
  assign n6328 = ( n4192 & n6324 ) | ( n4192 & n6327 ) | ( n6324 & n6327 ) ;
  assign n6329 = n6328 ^ n2321 ^ 1'b0 ;
  assign n6330 = ( n535 & n2420 ) | ( n535 & n3092 ) | ( n2420 & n3092 ) ;
  assign n6331 = n2026 & n6330 ;
  assign n6332 = n969 & n6331 ;
  assign n6333 = n937 & ~n1337 ;
  assign n6334 = ( ~n2470 & n6099 ) | ( ~n2470 & n6333 ) | ( n6099 & n6333 ) ;
  assign n6335 = ( n4292 & ~n4574 ) | ( n4292 & n5702 ) | ( ~n4574 & n5702 ) ;
  assign n6336 = ( n933 & ~n6297 ) | ( n933 & n6335 ) | ( ~n6297 & n6335 ) ;
  assign n6337 = n1529 & n4365 ;
  assign n6338 = n2857 ^ n1581 ^ n668 ;
  assign n6339 = ( ~n3123 & n6337 ) | ( ~n3123 & n6338 ) | ( n6337 & n6338 ) ;
  assign n6340 = n758 & n6339 ;
  assign n6341 = n1341 & n6340 ;
  assign n6342 = ( ~n2028 & n4983 ) | ( ~n2028 & n6341 ) | ( n4983 & n6341 ) ;
  assign n6347 = ~n2311 & n4329 ;
  assign n6348 = n500 ^ n275 ^ 1'b0 ;
  assign n6349 = n3464 | n6348 ;
  assign n6350 = n1685 & ~n6349 ;
  assign n6351 = n1851 & ~n5687 ;
  assign n6352 = n4519 ^ n4217 ^ n243 ;
  assign n6353 = n6352 ^ n6016 ^ n4092 ;
  assign n6354 = ( n3890 & n6351 ) | ( n3890 & ~n6353 ) | ( n6351 & ~n6353 ) ;
  assign n6355 = ( n6347 & n6350 ) | ( n6347 & ~n6354 ) | ( n6350 & ~n6354 ) ;
  assign n6343 = n1166 & n4520 ;
  assign n6344 = ( n553 & n2884 ) | ( n553 & ~n6343 ) | ( n2884 & ~n6343 ) ;
  assign n6345 = n3317 | n6344 ;
  assign n6346 = n6345 ^ n1352 ^ 1'b0 ;
  assign n6356 = n6355 ^ n6346 ^ 1'b0 ;
  assign n6357 = ( x97 & ~n140 ) | ( x97 & n1839 ) | ( ~n140 & n1839 ) ;
  assign n6358 = ( n201 & n2708 ) | ( n201 & n6357 ) | ( n2708 & n6357 ) ;
  assign n6363 = ( n605 & n1254 ) | ( n605 & n5710 ) | ( n1254 & n5710 ) ;
  assign n6361 = n5451 ^ n2801 ^ n488 ;
  assign n6362 = n6361 ^ n2653 ^ n578 ;
  assign n6364 = n6363 ^ n6362 ^ n3941 ;
  assign n6359 = n643 | n4690 ;
  assign n6360 = n350 | n6359 ;
  assign n6365 = n6364 ^ n6360 ^ n3491 ;
  assign n6366 = n1466 ^ n988 ^ 1'b0 ;
  assign n6367 = n6366 ^ n3738 ^ n2028 ;
  assign n6368 = n5407 ^ n1062 ^ 1'b0 ;
  assign n6369 = n3275 ^ n2658 ^ 1'b0 ;
  assign n6370 = n3609 & ~n6369 ;
  assign n6371 = ( ~n3443 & n6368 ) | ( ~n3443 & n6370 ) | ( n6368 & n6370 ) ;
  assign n6372 = n912 & ~n1910 ;
  assign n6373 = ~n3967 & n6372 ;
  assign n6374 = ( n269 & n528 ) | ( n269 & n1020 ) | ( n528 & n1020 ) ;
  assign n6375 = n6374 ^ n325 ^ 1'b0 ;
  assign n6376 = n5349 ^ n1108 ^ 1'b0 ;
  assign n6377 = n2858 ^ n2488 ^ n206 ;
  assign n6378 = n3060 & ~n6377 ;
  assign n6379 = n4870 & n6378 ;
  assign n6380 = n2813 ^ n2292 ^ n1119 ;
  assign n6384 = ( n2885 & n3271 ) | ( n2885 & ~n4361 ) | ( n3271 & ~n4361 ) ;
  assign n6381 = n6145 ^ n4213 ^ n4019 ;
  assign n6382 = n6381 ^ n3556 ^ 1'b0 ;
  assign n6383 = ~n1264 & n6382 ;
  assign n6385 = n6384 ^ n6383 ^ 1'b0 ;
  assign n6386 = n2789 ^ n1015 ^ n589 ;
  assign n6388 = n5569 ^ n2130 ^ n332 ;
  assign n6387 = n3934 & ~n4926 ;
  assign n6389 = n6388 ^ n6387 ^ 1'b0 ;
  assign n6390 = ( n1221 & n6386 ) | ( n1221 & n6389 ) | ( n6386 & n6389 ) ;
  assign n6391 = ~n6385 & n6390 ;
  assign n6392 = n6380 & n6391 ;
  assign n6396 = n5765 ^ n663 ^ 1'b0 ;
  assign n6393 = n6128 ^ n2473 ^ n1430 ;
  assign n6394 = ( ~n3835 & n4341 ) | ( ~n3835 & n6393 ) | ( n4341 & n6393 ) ;
  assign n6395 = n6394 ^ n3063 ^ n1228 ;
  assign n6397 = n6396 ^ n6395 ^ n586 ;
  assign n6403 = ( ~x46 & n2210 ) | ( ~x46 & n3558 ) | ( n2210 & n3558 ) ;
  assign n6412 = n1859 ^ x43 ^ 1'b0 ;
  assign n6413 = n5048 | n6412 ;
  assign n6414 = ( ~n238 & n3077 ) | ( ~n238 & n6413 ) | ( n3077 & n6413 ) ;
  assign n6404 = n1170 ^ n1081 ^ n902 ;
  assign n6405 = ~n2039 & n2847 ;
  assign n6406 = ~n2585 & n6405 ;
  assign n6407 = n6406 ^ n1901 ^ n1896 ;
  assign n6408 = n6407 ^ n2065 ^ n1949 ;
  assign n6409 = ( ~n3353 & n6404 ) | ( ~n3353 & n6408 ) | ( n6404 & n6408 ) ;
  assign n6410 = n1646 & ~n6409 ;
  assign n6411 = n6410 ^ n4976 ^ 1'b0 ;
  assign n6415 = n6414 ^ n6411 ^ 1'b0 ;
  assign n6416 = n6403 & ~n6415 ;
  assign n6398 = n716 & ~n3207 ;
  assign n6399 = ~n1759 & n6398 ;
  assign n6400 = ~n1322 & n5851 ;
  assign n6401 = n6399 & n6400 ;
  assign n6402 = n1969 | n6401 ;
  assign n6417 = n6416 ^ n6402 ^ 1'b0 ;
  assign n6418 = n1037 & ~n6417 ;
  assign n6419 = ( ~n4637 & n4925 ) | ( ~n4637 & n6178 ) | ( n4925 & n6178 ) ;
  assign n6420 = ( ~n2573 & n2846 ) | ( ~n2573 & n3784 ) | ( n2846 & n3784 ) ;
  assign n6421 = n2247 ^ n1681 ^ n759 ;
  assign n6422 = ( ~n1592 & n1703 ) | ( ~n1592 & n6421 ) | ( n1703 & n6421 ) ;
  assign n6423 = ( ~n5107 & n6420 ) | ( ~n5107 & n6422 ) | ( n6420 & n6422 ) ;
  assign n6425 = ( n516 & ~n576 ) | ( n516 & n4762 ) | ( ~n576 & n4762 ) ;
  assign n6424 = n6150 ^ n5932 ^ n2312 ;
  assign n6426 = n6425 ^ n6424 ^ n2903 ;
  assign n6427 = ( ~n1433 & n5152 ) | ( ~n1433 & n6426 ) | ( n5152 & n6426 ) ;
  assign n6428 = n6427 ^ n1714 ^ 1'b0 ;
  assign n6432 = n2854 ^ n2769 ^ x71 ;
  assign n6429 = n2669 | n5091 ;
  assign n6430 = n6429 ^ n2349 ^ 1'b0 ;
  assign n6431 = n6430 ^ n704 ^ n245 ;
  assign n6433 = n6432 ^ n6431 ^ n4735 ;
  assign n6434 = n4926 | n6038 ;
  assign n6435 = ( ~n4457 & n5320 ) | ( ~n4457 & n5391 ) | ( n5320 & n5391 ) ;
  assign n6436 = n6435 ^ n2751 ^ 1'b0 ;
  assign n6437 = n5894 ^ n2529 ^ n143 ;
  assign n6438 = ( n1513 & ~n1801 ) | ( n1513 & n5582 ) | ( ~n1801 & n5582 ) ;
  assign n6439 = n4990 & n6438 ;
  assign n6440 = ~n6437 & n6439 ;
  assign n6441 = n6440 ^ n4855 ^ n4164 ;
  assign n6442 = n4804 ^ n3006 ^ n1033 ;
  assign n6443 = n6442 ^ n5753 ^ n3401 ;
  assign n6444 = n3294 | n6443 ;
  assign n6445 = n3721 ^ n2844 ^ n353 ;
  assign n6446 = n2858 ^ n466 ^ n429 ;
  assign n6447 = n6446 ^ n2917 ^ n132 ;
  assign n6448 = n1125 ^ n703 ^ 1'b0 ;
  assign n6449 = ~n6447 & n6448 ;
  assign n6450 = n1255 | n3132 ;
  assign n6451 = n6450 ^ n6226 ^ 1'b0 ;
  assign n6452 = n5152 ^ n567 ^ n326 ;
  assign n6463 = n1676 & n4282 ;
  assign n6464 = ~n2579 & n6463 ;
  assign n6460 = ( x89 & ~n471 ) | ( x89 & n1606 ) | ( ~n471 & n1606 ) ;
  assign n6458 = n6363 ^ n1719 ^ x61 ;
  assign n6459 = n353 | n6458 ;
  assign n6461 = n6460 ^ n6459 ^ 1'b0 ;
  assign n6456 = n3146 ^ n2716 ^ 1'b0 ;
  assign n6453 = n3951 ^ n728 ^ 1'b0 ;
  assign n6454 = ~n3766 & n6453 ;
  assign n6455 = n4945 & n6454 ;
  assign n6457 = n6456 ^ n6455 ^ 1'b0 ;
  assign n6462 = n6461 ^ n6457 ^ x102 ;
  assign n6465 = n6464 ^ n6462 ^ n3185 ;
  assign n6466 = ( ~n382 & n805 ) | ( ~n382 & n3278 ) | ( n805 & n3278 ) ;
  assign n6467 = n6466 ^ n4561 ^ 1'b0 ;
  assign n6468 = n6467 ^ n4666 ^ 1'b0 ;
  assign n6469 = ~n2609 & n6468 ;
  assign n6470 = n563 & n2819 ;
  assign n6471 = n4046 & ~n6341 ;
  assign n6472 = n3588 & n6471 ;
  assign n6473 = n6470 & n6472 ;
  assign n6474 = n3792 & n6473 ;
  assign n6475 = n4062 & ~n5818 ;
  assign n6482 = n4365 | n4670 ;
  assign n6483 = n6482 ^ n581 ^ 1'b0 ;
  assign n6480 = n725 ^ n655 ^ n288 ;
  assign n6481 = n6480 ^ n3823 ^ n3226 ;
  assign n6476 = ( n502 & ~n3078 ) | ( n502 & n3093 ) | ( ~n3078 & n3093 ) ;
  assign n6477 = n953 | n6476 ;
  assign n6478 = n524 & n2851 ;
  assign n6479 = ( n2877 & n6477 ) | ( n2877 & n6478 ) | ( n6477 & n6478 ) ;
  assign n6484 = n6483 ^ n6481 ^ n6479 ;
  assign n6485 = n6182 ^ n2565 ^ n1377 ;
  assign n6486 = n4555 ^ n1045 ^ 1'b0 ;
  assign n6487 = n503 | n6486 ;
  assign n6488 = ( ~n4505 & n6485 ) | ( ~n4505 & n6487 ) | ( n6485 & n6487 ) ;
  assign n6489 = n907 ^ n870 ^ 1'b0 ;
  assign n6490 = n6489 ^ n375 ^ 1'b0 ;
  assign n6491 = ~n6175 & n6490 ;
  assign n6492 = ~n6488 & n6491 ;
  assign n6498 = ( n441 & ~n2816 ) | ( n441 & n4785 ) | ( ~n2816 & n4785 ) ;
  assign n6499 = ( n1992 & n5385 ) | ( n1992 & ~n6498 ) | ( n5385 & ~n6498 ) ;
  assign n6493 = n322 & n5504 ;
  assign n6494 = n2092 ^ n1126 ^ 1'b0 ;
  assign n6495 = ~n5753 & n6494 ;
  assign n6496 = n6495 ^ n1106 ^ 1'b0 ;
  assign n6497 = ~n6493 & n6496 ;
  assign n6500 = n6499 ^ n6497 ^ n5400 ;
  assign n6501 = n6492 | n6500 ;
  assign n6502 = n5031 & ~n6501 ;
  assign n6503 = n2706 ^ n801 ^ n509 ;
  assign n6504 = ( n1086 & n5286 ) | ( n1086 & ~n6503 ) | ( n5286 & ~n6503 ) ;
  assign n6505 = ( n1096 & ~n3320 ) | ( n1096 & n3552 ) | ( ~n3320 & n3552 ) ;
  assign n6506 = n6505 ^ n4440 ^ 1'b0 ;
  assign n6507 = ~n6246 & n6506 ;
  assign n6508 = n3019 ^ n2788 ^ n1213 ;
  assign n6509 = n6508 ^ n3801 ^ 1'b0 ;
  assign n6510 = n1795 ^ n413 ^ n334 ;
  assign n6511 = ( n1921 & n4371 ) | ( n1921 & n6510 ) | ( n4371 & n6510 ) ;
  assign n6512 = n6511 ^ n2594 ^ 1'b0 ;
  assign n6513 = n6509 & ~n6512 ;
  assign n6518 = n178 & n513 ;
  assign n6517 = n2112 | n2269 ;
  assign n6519 = n6518 ^ n6517 ^ 1'b0 ;
  assign n6523 = n1467 | n5147 ;
  assign n6524 = n6523 ^ n209 ^ 1'b0 ;
  assign n6522 = n3700 ^ n1912 ^ 1'b0 ;
  assign n6525 = n6524 ^ n6522 ^ n5191 ;
  assign n6520 = n1219 & ~n1991 ;
  assign n6521 = n6520 ^ n405 ^ n285 ;
  assign n6526 = n6525 ^ n6521 ^ 1'b0 ;
  assign n6527 = n6519 & ~n6526 ;
  assign n6514 = n459 & n5004 ;
  assign n6515 = n1780 | n6514 ;
  assign n6516 = n3817 | n6515 ;
  assign n6528 = n6527 ^ n6516 ^ n2520 ;
  assign n6529 = n4375 ^ n468 ^ x96 ;
  assign n6530 = n6529 ^ n6150 ^ n1623 ;
  assign n6531 = ( n2152 & ~n3022 ) | ( n2152 & n6530 ) | ( ~n3022 & n6530 ) ;
  assign n6532 = ( n865 & ~n2252 ) | ( n865 & n2320 ) | ( ~n2252 & n2320 ) ;
  assign n6533 = ( n2336 & n2830 ) | ( n2336 & n3452 ) | ( n2830 & n3452 ) ;
  assign n6534 = ( ~n1327 & n6532 ) | ( ~n1327 & n6533 ) | ( n6532 & n6533 ) ;
  assign n6535 = n5306 ^ n5121 ^ n1312 ;
  assign n6536 = x94 & n1588 ;
  assign n6537 = n3322 & n6536 ;
  assign n6538 = ( n2167 & n2701 ) | ( n2167 & n6099 ) | ( n2701 & n6099 ) ;
  assign n6539 = n2901 & ~n6538 ;
  assign n6540 = ( n2978 & ~n6537 ) | ( n2978 & n6539 ) | ( ~n6537 & n6539 ) ;
  assign n6541 = n5246 ^ n4802 ^ n2321 ;
  assign n6542 = ( ~n1375 & n1484 ) | ( ~n1375 & n6448 ) | ( n1484 & n6448 ) ;
  assign n6543 = ( n4848 & n4971 ) | ( n4848 & ~n6542 ) | ( n4971 & ~n6542 ) ;
  assign n6544 = n5307 ^ n2489 ^ n2078 ;
  assign n6545 = n5024 ^ n2668 ^ 1'b0 ;
  assign n6546 = n5321 & ~n6545 ;
  assign n6547 = n4592 & n6546 ;
  assign n6548 = n3016 ^ n1263 ^ 1'b0 ;
  assign n6549 = n6548 ^ n3635 ^ n234 ;
  assign n6550 = ( ~n6544 & n6547 ) | ( ~n6544 & n6549 ) | ( n6547 & n6549 ) ;
  assign n6551 = n6550 ^ n5583 ^ n5169 ;
  assign n6552 = ~n3375 & n4141 ;
  assign n6553 = ( n459 & n5423 ) | ( n459 & ~n5672 ) | ( n5423 & ~n5672 ) ;
  assign n6554 = ( ~n1920 & n2988 ) | ( ~n1920 & n6553 ) | ( n2988 & n6553 ) ;
  assign n6558 = ( n1082 & n1757 ) | ( n1082 & n2211 ) | ( n1757 & n2211 ) ;
  assign n6555 = ( ~n2479 & n2569 ) | ( ~n2479 & n3423 ) | ( n2569 & n3423 ) ;
  assign n6556 = ( n1271 & n2702 ) | ( n1271 & n6555 ) | ( n2702 & n6555 ) ;
  assign n6557 = ( n558 & n2936 ) | ( n558 & n6556 ) | ( n2936 & n6556 ) ;
  assign n6559 = n6558 ^ n6557 ^ 1'b0 ;
  assign n6565 = n4223 ^ n2018 ^ 1'b0 ;
  assign n6566 = n6565 ^ n5808 ^ 1'b0 ;
  assign n6560 = x71 ^ x52 ^ 1'b0 ;
  assign n6561 = ~n1553 & n2605 ;
  assign n6562 = n6561 ^ n1991 ^ x34 ;
  assign n6563 = n4232 & n6562 ;
  assign n6564 = ~n6560 & n6563 ;
  assign n6567 = n6566 ^ n6564 ^ 1'b0 ;
  assign n6568 = n6567 ^ n4973 ^ 1'b0 ;
  assign n6569 = n6568 ^ n4291 ^ n1506 ;
  assign n6570 = n1589 & n3144 ;
  assign n6571 = n1493 & n2270 ;
  assign n6572 = n6571 ^ n4624 ^ 1'b0 ;
  assign n6573 = ( n630 & n3360 ) | ( n630 & n6572 ) | ( n3360 & n6572 ) ;
  assign n6574 = n169 & n2151 ;
  assign n6575 = n2788 & n3766 ;
  assign n6576 = n6574 & n6575 ;
  assign n6577 = ~n6107 & n6576 ;
  assign n6583 = n1127 | n2117 ;
  assign n6584 = n6583 ^ n2547 ^ 1'b0 ;
  assign n6582 = ( n192 & n1876 ) | ( n192 & ~n6302 ) | ( n1876 & ~n6302 ) ;
  assign n6578 = n5512 ^ n3934 ^ 1'b0 ;
  assign n6579 = n5275 ^ n1772 ^ 1'b0 ;
  assign n6580 = n3191 | n6579 ;
  assign n6581 = ( n1858 & n6578 ) | ( n1858 & ~n6580 ) | ( n6578 & ~n6580 ) ;
  assign n6585 = n6584 ^ n6582 ^ n6581 ;
  assign n6588 = x100 & n2539 ;
  assign n6589 = ~n2145 & n6588 ;
  assign n6590 = ( ~n850 & n4205 ) | ( ~n850 & n6589 ) | ( n4205 & n6589 ) ;
  assign n6586 = ( n2113 & n3139 ) | ( n2113 & ~n3296 ) | ( n3139 & ~n3296 ) ;
  assign n6587 = n870 & ~n6586 ;
  assign n6591 = n6590 ^ n6587 ^ 1'b0 ;
  assign n6592 = ( n2943 & n3095 ) | ( n2943 & n6591 ) | ( n3095 & n6591 ) ;
  assign n6593 = n2511 | n6592 ;
  assign n6594 = ( n3557 & ~n6585 ) | ( n3557 & n6593 ) | ( ~n6585 & n6593 ) ;
  assign n6595 = n1212 ^ n342 ^ 1'b0 ;
  assign n6596 = n830 | n6595 ;
  assign n6597 = n1155 | n6596 ;
  assign n6598 = n4109 & ~n6597 ;
  assign n6599 = n6598 ^ n4241 ^ 1'b0 ;
  assign n6600 = n6599 ^ n4461 ^ n3522 ;
  assign n6603 = n4342 ^ n1761 ^ n979 ;
  assign n6601 = n5050 ^ n4564 ^ 1'b0 ;
  assign n6602 = n6601 ^ n5491 ^ n329 ;
  assign n6604 = n6603 ^ n6602 ^ n1863 ;
  assign n6605 = n2061 | n6604 ;
  assign n6607 = ( ~n1978 & n4405 ) | ( ~n1978 & n4622 ) | ( n4405 & n4622 ) ;
  assign n6606 = ( n1282 & ~n2130 ) | ( n1282 & n5491 ) | ( ~n2130 & n5491 ) ;
  assign n6608 = n6607 ^ n6606 ^ 1'b0 ;
  assign n6616 = n1878 & n5390 ;
  assign n6617 = ~n1192 & n6616 ;
  assign n6618 = ( x26 & n2636 ) | ( x26 & n6617 ) | ( n2636 & n6617 ) ;
  assign n6609 = n226 | n5783 ;
  assign n6610 = n6609 ^ n2605 ^ 1'b0 ;
  assign n6611 = x74 & n6610 ;
  assign n6612 = n5212 & ~n6611 ;
  assign n6613 = n3437 | n6099 ;
  assign n6614 = n6612 | n6613 ;
  assign n6615 = ~n5852 & n6614 ;
  assign n6619 = n6618 ^ n6615 ^ 1'b0 ;
  assign n6620 = ~n159 & n5336 ;
  assign n6621 = n475 & n6620 ;
  assign n6622 = n3856 | n6621 ;
  assign n6623 = ~n1027 & n6622 ;
  assign n6625 = ~n565 & n3721 ;
  assign n6626 = n6625 ^ n1241 ^ 1'b0 ;
  assign n6624 = ~n1264 & n3944 ;
  assign n6627 = n6626 ^ n6624 ^ 1'b0 ;
  assign n6628 = ( ~n662 & n2653 ) | ( ~n662 & n3335 ) | ( n2653 & n3335 ) ;
  assign n6629 = ( n489 & ~n6421 ) | ( n489 & n6628 ) | ( ~n6421 & n6628 ) ;
  assign n6630 = n6629 ^ n6042 ^ 1'b0 ;
  assign n6631 = n6462 ^ n4653 ^ 1'b0 ;
  assign n6632 = n719 & ~n2800 ;
  assign n6633 = n6632 ^ n5748 ^ 1'b0 ;
  assign n6634 = n6633 ^ n4701 ^ n1617 ;
  assign n6635 = ( ~x61 & n1056 ) | ( ~x61 & n1422 ) | ( n1056 & n1422 ) ;
  assign n6636 = n1834 | n6635 ;
  assign n6637 = ( n2178 & ~n2761 ) | ( n2178 & n6636 ) | ( ~n2761 & n6636 ) ;
  assign n6638 = n6637 ^ n2252 ^ 1'b0 ;
  assign n6639 = n838 ^ n420 ^ 1'b0 ;
  assign n6640 = n6639 ^ n6437 ^ n2665 ;
  assign n6641 = ~n1127 & n6640 ;
  assign n6642 = n5167 & n6641 ;
  assign n6643 = n2850 ^ n2248 ^ 1'b0 ;
  assign n6644 = ~n6642 & n6643 ;
  assign n6645 = ( n503 & n3439 ) | ( n503 & n4944 ) | ( n3439 & n4944 ) ;
  assign n6646 = n6645 ^ n5506 ^ n4514 ;
  assign n6647 = n1919 & n6646 ;
  assign n6656 = n3648 ^ n3582 ^ n2846 ;
  assign n6653 = n3232 ^ n2812 ^ n180 ;
  assign n6654 = ( ~n4624 & n6162 ) | ( ~n4624 & n6653 ) | ( n6162 & n6653 ) ;
  assign n6655 = ( n828 & ~n2041 ) | ( n828 & n6654 ) | ( ~n2041 & n6654 ) ;
  assign n6650 = n5272 ^ n4034 ^ n3238 ;
  assign n6651 = n6650 ^ n3885 ^ n3443 ;
  assign n6648 = ~n607 & n3658 ;
  assign n6649 = n6648 ^ n418 ^ 1'b0 ;
  assign n6652 = n6651 ^ n6649 ^ n332 ;
  assign n6657 = n6656 ^ n6655 ^ n6652 ;
  assign n6658 = n2768 | n4762 ;
  assign n6663 = n416 | n1199 ;
  assign n6664 = n4314 | n6663 ;
  assign n6661 = n5416 ^ n3387 ^ n395 ;
  assign n6659 = n4205 ^ n3713 ^ 1'b0 ;
  assign n6660 = n4445 & ~n6659 ;
  assign n6662 = n6661 ^ n6660 ^ n2777 ;
  assign n6665 = n6664 ^ n6662 ^ n491 ;
  assign n6666 = n2653 | n6665 ;
  assign n6667 = n1545 & ~n6666 ;
  assign n6668 = ( n1084 & n6658 ) | ( n1084 & ~n6667 ) | ( n6658 & ~n6667 ) ;
  assign n6669 = ~n357 & n2652 ;
  assign n6670 = n6669 ^ n3026 ^ 1'b0 ;
  assign n6671 = n1516 | n6670 ;
  assign n6672 = n6671 ^ n5048 ^ n3083 ;
  assign n6673 = ( n5295 & n6109 ) | ( n5295 & ~n6672 ) | ( n6109 & ~n6672 ) ;
  assign n6674 = ~n858 & n1370 ;
  assign n6675 = n6674 ^ n2974 ^ 1'b0 ;
  assign n6676 = n6099 ^ n3054 ^ 1'b0 ;
  assign n6677 = ( n668 & n1181 ) | ( n668 & ~n4619 ) | ( n1181 & ~n4619 ) ;
  assign n6678 = n6677 ^ n4656 ^ n1581 ;
  assign n6679 = ~n2296 & n6678 ;
  assign n6680 = ( n735 & n1004 ) | ( n735 & n1516 ) | ( n1004 & n1516 ) ;
  assign n6681 = ( n1640 & ~n4356 ) | ( n1640 & n6680 ) | ( ~n4356 & n6680 ) ;
  assign n6682 = ~n3188 & n4015 ;
  assign n6683 = n6682 ^ n6489 ^ n640 ;
  assign n6684 = ( ~n1334 & n3354 ) | ( ~n1334 & n3365 ) | ( n3354 & n3365 ) ;
  assign n6685 = n4367 & ~n6684 ;
  assign n6686 = n4143 ^ n2295 ^ n2011 ;
  assign n6687 = ~n5723 & n6686 ;
  assign n6688 = n6687 ^ n1278 ^ 1'b0 ;
  assign n6689 = n1762 & ~n6688 ;
  assign n6690 = ~n3944 & n6689 ;
  assign n6691 = n1375 ^ n1347 ^ 1'b0 ;
  assign n6692 = n1290 & ~n6691 ;
  assign n6693 = n6692 ^ n6073 ^ n2003 ;
  assign n6694 = n6693 ^ n2057 ^ 1'b0 ;
  assign n6695 = n705 & ~n6602 ;
  assign n6696 = n5634 & n6695 ;
  assign n6697 = n6694 | n6696 ;
  assign n6698 = n4483 & n5512 ;
  assign n6699 = n1011 & ~n6698 ;
  assign n6710 = n3603 ^ n1238 ^ 1'b0 ;
  assign n6711 = n4143 | n6710 ;
  assign n6712 = n6711 ^ n3267 ^ 1'b0 ;
  assign n6713 = n3443 | n6712 ;
  assign n6714 = n6713 ^ n3785 ^ n1267 ;
  assign n6707 = n2792 ^ n1254 ^ n588 ;
  assign n6708 = n3164 | n6707 ;
  assign n6709 = n6708 ^ n1356 ^ 1'b0 ;
  assign n6700 = ( n225 & n1625 ) | ( n225 & n4353 ) | ( n1625 & n4353 ) ;
  assign n6701 = n6700 ^ x73 ^ 1'b0 ;
  assign n6702 = n145 & ~n5589 ;
  assign n6703 = n477 & n6702 ;
  assign n6704 = n4441 | n6703 ;
  assign n6705 = n3931 | n6704 ;
  assign n6706 = n6701 & ~n6705 ;
  assign n6715 = n6714 ^ n6709 ^ n6706 ;
  assign n6716 = n6290 ^ n4310 ^ 1'b0 ;
  assign n6717 = n6185 & ~n6716 ;
  assign n6718 = n6717 ^ n211 ^ 1'b0 ;
  assign n6719 = ~n531 & n3557 ;
  assign n6720 = n1779 | n1810 ;
  assign n6721 = ~n6464 & n6720 ;
  assign n6722 = ( n2665 & n6719 ) | ( n2665 & ~n6721 ) | ( n6719 & ~n6721 ) ;
  assign n6723 = n6109 & n6722 ;
  assign n6724 = n4954 ^ n4630 ^ 1'b0 ;
  assign n6725 = n6724 ^ n2889 ^ 1'b0 ;
  assign n6726 = n173 & ~n6725 ;
  assign n6727 = n6726 ^ n4280 ^ 1'b0 ;
  assign n6728 = n3498 & n6727 ;
  assign n6729 = n6728 ^ n5568 ^ 1'b0 ;
  assign n6731 = ( ~n1250 & n2530 ) | ( ~n1250 & n3790 ) | ( n2530 & n3790 ) ;
  assign n6730 = n2884 ^ n578 ^ 1'b0 ;
  assign n6732 = n6731 ^ n6730 ^ 1'b0 ;
  assign n6733 = n6732 ^ n3122 ^ n1227 ;
  assign n6734 = ( n1334 & ~n3772 ) | ( n1334 & n4100 ) | ( ~n3772 & n4100 ) ;
  assign n6735 = n3655 & n4742 ;
  assign n6736 = n6735 ^ n4353 ^ 1'b0 ;
  assign n6737 = ( n1765 & n6734 ) | ( n1765 & n6736 ) | ( n6734 & n6736 ) ;
  assign n6738 = n6737 ^ n4331 ^ n143 ;
  assign n6739 = ( ~n1373 & n1650 ) | ( ~n1373 & n3250 ) | ( n1650 & n3250 ) ;
  assign n6740 = n6739 ^ n5753 ^ n3306 ;
  assign n6741 = n2126 | n6740 ;
  assign n6742 = n1042 & ~n6741 ;
  assign n6743 = n2273 & n6742 ;
  assign n6744 = n6743 ^ n3944 ^ 1'b0 ;
  assign n6745 = n488 & n6744 ;
  assign n6746 = n3293 ^ n1312 ^ 1'b0 ;
  assign n6747 = n372 | n3443 ;
  assign n6748 = n6747 ^ n328 ^ 1'b0 ;
  assign n6749 = ( n1998 & n6136 ) | ( n1998 & ~n6748 ) | ( n6136 & ~n6748 ) ;
  assign n6750 = ( n2208 & n6746 ) | ( n2208 & ~n6749 ) | ( n6746 & ~n6749 ) ;
  assign n6751 = ( ~n3948 & n5191 ) | ( ~n3948 & n6750 ) | ( n5191 & n6750 ) ;
  assign n6752 = n2113 & ~n5162 ;
  assign n6753 = n2228 & ~n2363 ;
  assign n6754 = n4967 & n6753 ;
  assign n6755 = n6752 | n6754 ;
  assign n6756 = n6755 ^ n130 ^ 1'b0 ;
  assign n6757 = n6756 ^ x1 ^ 1'b0 ;
  assign n6758 = n6518 & n6757 ;
  assign n6759 = n3990 ^ n975 ^ n645 ;
  assign n6760 = ( n535 & n2307 ) | ( n535 & ~n6759 ) | ( n2307 & ~n6759 ) ;
  assign n6761 = ~n443 & n984 ;
  assign n6762 = ~n6760 & n6761 ;
  assign n6763 = ( n1186 & n3115 ) | ( n1186 & n6762 ) | ( n3115 & n6762 ) ;
  assign n6764 = n1396 ^ n933 ^ 1'b0 ;
  assign n6765 = ~n526 & n4427 ;
  assign n6766 = n1524 ^ n1193 ^ n429 ;
  assign n6767 = ~n2486 & n6766 ;
  assign n6768 = n5259 & n6767 ;
  assign n6769 = n3692 & n4551 ;
  assign n6770 = n6769 ^ n5633 ^ 1'b0 ;
  assign n6771 = ~n774 & n1682 ;
  assign n6772 = ( n6768 & n6770 ) | ( n6768 & ~n6771 ) | ( n6770 & ~n6771 ) ;
  assign n6773 = ( n173 & n1276 ) | ( n173 & ~n6772 ) | ( n1276 & ~n6772 ) ;
  assign n6774 = n6773 ^ n2672 ^ 1'b0 ;
  assign n6775 = ~n6742 & n6774 ;
  assign n6776 = n2800 ^ x56 ^ 1'b0 ;
  assign n6777 = n6776 ^ n3712 ^ n3226 ;
  assign n6780 = n2619 | n5438 ;
  assign n6781 = n6780 ^ n6218 ^ 1'b0 ;
  assign n6778 = ( ~n2078 & n2141 ) | ( ~n2078 & n3093 ) | ( n2141 & n3093 ) ;
  assign n6779 = ( ~n2460 & n6658 ) | ( ~n2460 & n6778 ) | ( n6658 & n6778 ) ;
  assign n6782 = n6781 ^ n6779 ^ 1'b0 ;
  assign n6783 = ( ~n1617 & n2321 ) | ( ~n1617 & n4377 ) | ( n2321 & n4377 ) ;
  assign n6784 = x112 & ~n953 ;
  assign n6785 = n6784 ^ n2165 ^ 1'b0 ;
  assign n6786 = ( n600 & n5986 ) | ( n600 & n6785 ) | ( n5986 & n6785 ) ;
  assign n6787 = ( n3571 & n6783 ) | ( n3571 & n6786 ) | ( n6783 & n6786 ) ;
  assign n6788 = n4791 ^ n4285 ^ n841 ;
  assign n6796 = n1936 ^ x109 ^ 1'b0 ;
  assign n6791 = n507 | n6589 ;
  assign n6792 = n5332 & ~n6791 ;
  assign n6793 = n1920 | n6792 ;
  assign n6794 = x21 | n6793 ;
  assign n6795 = n6794 ^ n6199 ^ n2501 ;
  assign n6789 = n4107 & ~n5206 ;
  assign n6790 = ~n705 & n6789 ;
  assign n6797 = n6796 ^ n6795 ^ n6790 ;
  assign n6798 = n3654 ^ n1323 ^ n1019 ;
  assign n6799 = ~n3581 & n6798 ;
  assign n6800 = n6161 ^ n2316 ^ n1225 ;
  assign n6801 = n1945 & ~n5291 ;
  assign n6802 = n6801 ^ n6113 ^ 1'b0 ;
  assign n6803 = n4746 & n6802 ;
  assign n6804 = ~n4693 & n6803 ;
  assign n6805 = ( n4259 & ~n5009 ) | ( n4259 & n6802 ) | ( ~n5009 & n6802 ) ;
  assign n6806 = ~n6804 & n6805 ;
  assign n6809 = n881 & n981 ;
  assign n6810 = ( ~n5416 & n5882 ) | ( ~n5416 & n6809 ) | ( n5882 & n6809 ) ;
  assign n6807 = n877 & ~n1301 ;
  assign n6808 = ( n2491 & n4284 ) | ( n2491 & n6807 ) | ( n4284 & n6807 ) ;
  assign n6811 = n6810 ^ n6808 ^ n1754 ;
  assign n6815 = n5248 ^ n726 ^ n357 ;
  assign n6816 = n6815 ^ n4459 ^ n2032 ;
  assign n6817 = n4914 & ~n6816 ;
  assign n6818 = n2381 & n6817 ;
  assign n6812 = n2701 ^ n1414 ^ n1081 ;
  assign n6813 = ( n1690 & n3271 ) | ( n1690 & ~n6812 ) | ( n3271 & ~n6812 ) ;
  assign n6814 = ( n1878 & ~n5449 ) | ( n1878 & n6813 ) | ( ~n5449 & n6813 ) ;
  assign n6819 = n6818 ^ n6814 ^ 1'b0 ;
  assign n6821 = n4514 ^ n994 ^ n573 ;
  assign n6820 = n556 & ~n1051 ;
  assign n6822 = n6821 ^ n6820 ^ n1891 ;
  assign n6823 = ( n2026 & n3168 ) | ( n2026 & ~n5310 ) | ( n3168 & ~n5310 ) ;
  assign n6824 = n6823 ^ n6077 ^ 1'b0 ;
  assign n6825 = ~n995 & n6824 ;
  assign n6827 = n1568 & ~n3355 ;
  assign n6828 = n643 & n6827 ;
  assign n6826 = n2443 ^ x62 ^ 1'b0 ;
  assign n6829 = n6828 ^ n6826 ^ n3066 ;
  assign n6830 = n1391 & n5077 ;
  assign n6831 = ( n3690 & n6829 ) | ( n3690 & n6830 ) | ( n6829 & n6830 ) ;
  assign n6832 = ( ~n1312 & n1738 ) | ( ~n1312 & n3712 ) | ( n1738 & n3712 ) ;
  assign n6833 = n6832 ^ n1713 ^ 1'b0 ;
  assign n6834 = n4113 & n4518 ;
  assign n6835 = n6834 ^ n6200 ^ 1'b0 ;
  assign n6836 = n847 | n3686 ;
  assign n6837 = n6586 & ~n6836 ;
  assign n6838 = n1271 & n6837 ;
  assign n6839 = n6838 ^ n3490 ^ 1'b0 ;
  assign n6840 = n6839 ^ n6040 ^ 1'b0 ;
  assign n6841 = n2184 & ~n3606 ;
  assign n6842 = ~n6328 & n6841 ;
  assign n6843 = n2366 ^ n1678 ^ 1'b0 ;
  assign n6844 = n1479 | n1769 ;
  assign n6845 = ( n2619 & ~n6843 ) | ( n2619 & n6844 ) | ( ~n6843 & n6844 ) ;
  assign n6846 = n1574 & n4521 ;
  assign n6847 = n6846 ^ n1263 ^ 1'b0 ;
  assign n6848 = n5394 ^ n3604 ^ 1'b0 ;
  assign n6849 = n6847 | n6848 ;
  assign n6850 = n312 | n3186 ;
  assign n6851 = n4683 | n6850 ;
  assign n6852 = ( n3464 & n4437 ) | ( n3464 & ~n6851 ) | ( n4437 & ~n6851 ) ;
  assign n6872 = n4882 ^ n2761 ^ 1'b0 ;
  assign n6871 = n2997 ^ n2366 ^ n2279 ;
  assign n6873 = n6872 ^ n6871 ^ n3333 ;
  assign n6874 = ( ~n2103 & n2674 ) | ( ~n2103 & n6873 ) | ( n2674 & n6873 ) ;
  assign n6868 = ~n2437 & n4768 ;
  assign n6869 = n6408 & ~n6868 ;
  assign n6867 = n2680 & n3122 ;
  assign n6870 = n6869 ^ n6867 ^ n4721 ;
  assign n6863 = n293 & ~n5488 ;
  assign n6864 = ~n548 & n6863 ;
  assign n6858 = ( n596 & n2238 ) | ( n596 & n5215 ) | ( n2238 & n5215 ) ;
  assign n6859 = n796 | n2961 ;
  assign n6860 = ( n4213 & n6858 ) | ( n4213 & n6859 ) | ( n6858 & n6859 ) ;
  assign n6853 = n5048 ^ n1869 ^ 1'b0 ;
  assign n6854 = ~n2493 & n6853 ;
  assign n6855 = n3319 ^ n213 ^ 1'b0 ;
  assign n6856 = n6854 & ~n6855 ;
  assign n6857 = ~n3851 & n6856 ;
  assign n6861 = n6860 ^ n6857 ^ 1'b0 ;
  assign n6862 = n2697 & n6861 ;
  assign n6865 = n6864 ^ n6862 ^ 1'b0 ;
  assign n6866 = ( n458 & n3782 ) | ( n458 & ~n6865 ) | ( n3782 & ~n6865 ) ;
  assign n6875 = n6874 ^ n6870 ^ n6866 ;
  assign n6876 = ( n456 & n3613 ) | ( n456 & n4749 ) | ( n3613 & n4749 ) ;
  assign n6877 = n3809 | n6876 ;
  assign n6878 = n2640 & ~n6877 ;
  assign n6883 = n4056 ^ n2429 ^ n1171 ;
  assign n6880 = n6077 ^ n1725 ^ x21 ;
  assign n6879 = ( ~n1501 & n2248 ) | ( ~n1501 & n5201 ) | ( n2248 & n5201 ) ;
  assign n6881 = n6880 ^ n6879 ^ x112 ;
  assign n6882 = ~n3333 & n6881 ;
  assign n6884 = n6883 ^ n6882 ^ n1171 ;
  assign n6888 = ( n1382 & n2007 ) | ( n1382 & n6470 ) | ( n2007 & n6470 ) ;
  assign n6889 = n1148 & ~n5713 ;
  assign n6890 = n6888 & n6889 ;
  assign n6885 = n2262 ^ n2167 ^ 1'b0 ;
  assign n6886 = ( n1107 & n5897 ) | ( n1107 & ~n6885 ) | ( n5897 & ~n6885 ) ;
  assign n6887 = ( ~n2386 & n4134 ) | ( ~n2386 & n6886 ) | ( n4134 & n6886 ) ;
  assign n6891 = n6890 ^ n6887 ^ n505 ;
  assign n6892 = ( n2928 & n5932 ) | ( n2928 & n6443 ) | ( n5932 & n6443 ) ;
  assign n6897 = ( n453 & ~n2524 ) | ( n453 & n3309 ) | ( ~n2524 & n3309 ) ;
  assign n6893 = n1186 ^ n284 ^ 1'b0 ;
  assign n6894 = n6893 ^ n2279 ^ 1'b0 ;
  assign n6895 = n1250 | n6894 ;
  assign n6896 = ( ~n2160 & n6489 ) | ( ~n2160 & n6895 ) | ( n6489 & n6895 ) ;
  assign n6898 = n6897 ^ n6896 ^ n4917 ;
  assign n6899 = n3622 ^ n1946 ^ n663 ;
  assign n6900 = ( n4117 & n6898 ) | ( n4117 & ~n6899 ) | ( n6898 & ~n6899 ) ;
  assign n6901 = ~n3157 & n6900 ;
  assign n6902 = n1168 ^ n352 ^ 1'b0 ;
  assign n6903 = n6901 & n6902 ;
  assign n6904 = ( n996 & n4878 ) | ( n996 & n5960 ) | ( n4878 & n5960 ) ;
  assign n6905 = n471 & ~n1546 ;
  assign n6906 = ( n4053 & ~n6904 ) | ( n4053 & n6905 ) | ( ~n6904 & n6905 ) ;
  assign n6907 = ( n2982 & n4629 ) | ( n2982 & ~n6483 ) | ( n4629 & ~n6483 ) ;
  assign n6908 = n2053 & n5750 ;
  assign n6909 = n4841 ^ n3918 ^ 1'b0 ;
  assign n6910 = n6908 & ~n6909 ;
  assign n6911 = ( n2317 & n6907 ) | ( n2317 & ~n6910 ) | ( n6907 & ~n6910 ) ;
  assign n6912 = n6911 ^ n2834 ^ n1955 ;
  assign n6913 = n2543 ^ n681 ^ 1'b0 ;
  assign n6918 = n1764 ^ n487 ^ 1'b0 ;
  assign n6919 = ( n1776 & ~n2065 ) | ( n1776 & n6918 ) | ( ~n2065 & n6918 ) ;
  assign n6917 = n5099 ^ n2507 ^ 1'b0 ;
  assign n6914 = n1666 | n1702 ;
  assign n6915 = n5534 ^ n4491 ^ n4169 ;
  assign n6916 = ( n329 & ~n6914 ) | ( n329 & n6915 ) | ( ~n6914 & n6915 ) ;
  assign n6920 = n6919 ^ n6917 ^ n6916 ;
  assign n6921 = n6322 ^ n5609 ^ n493 ;
  assign n6922 = n2848 ^ n2368 ^ 1'b0 ;
  assign n6923 = n1120 & n6922 ;
  assign n6924 = n6923 ^ n4815 ^ 1'b0 ;
  assign n6925 = n3828 & n6772 ;
  assign n6926 = n5854 ^ n1071 ^ 1'b0 ;
  assign n6927 = n1942 & ~n6926 ;
  assign n6928 = ( n4217 & n4415 ) | ( n4217 & ~n6927 ) | ( n4415 & ~n6927 ) ;
  assign n6929 = n5223 ^ n704 ^ n180 ;
  assign n6930 = ~n867 & n1661 ;
  assign n6931 = ~n5541 & n6930 ;
  assign n6932 = n1241 & ~n6931 ;
  assign n6933 = n6932 ^ n3193 ^ 1'b0 ;
  assign n6934 = n325 & ~n1700 ;
  assign n6935 = n6933 & n6934 ;
  assign n6936 = n310 | n4739 ;
  assign n6937 = n668 & ~n6936 ;
  assign n6938 = ( ~n1284 & n1339 ) | ( ~n1284 & n1480 ) | ( n1339 & n1480 ) ;
  assign n6939 = ( n1359 & n1659 ) | ( n1359 & n6938 ) | ( n1659 & n6938 ) ;
  assign n6940 = n6939 ^ n6369 ^ n918 ;
  assign n6941 = ( ~n5591 & n6937 ) | ( ~n5591 & n6940 ) | ( n6937 & n6940 ) ;
  assign n6942 = n4204 ^ n2592 ^ n1706 ;
  assign n6943 = ( n789 & n1721 ) | ( n789 & n3318 ) | ( n1721 & n3318 ) ;
  assign n6944 = n6943 ^ n386 ^ 1'b0 ;
  assign n6945 = n6942 & ~n6944 ;
  assign n6946 = n6291 ^ n5024 ^ n2281 ;
  assign n6947 = n6946 ^ n5187 ^ 1'b0 ;
  assign n6948 = ~n490 & n6947 ;
  assign n6949 = ( ~n245 & n3626 ) | ( ~n245 & n5504 ) | ( n3626 & n5504 ) ;
  assign n6950 = n1570 & n2973 ;
  assign n6951 = ( ~n866 & n2099 ) | ( ~n866 & n6950 ) | ( n2099 & n6950 ) ;
  assign n6952 = n6951 ^ n6469 ^ n4786 ;
  assign n6953 = ~n689 & n1242 ;
  assign n6954 = n6953 ^ n2695 ^ n1315 ;
  assign n6955 = ( n2794 & n6510 ) | ( n2794 & ~n6954 ) | ( n6510 & ~n6954 ) ;
  assign n6956 = ( n6546 & ~n6721 ) | ( n6546 & n6955 ) | ( ~n6721 & n6955 ) ;
  assign n6957 = ( n1264 & n1361 ) | ( n1264 & n2569 ) | ( n1361 & n2569 ) ;
  assign n6958 = ( n2141 & ~n6956 ) | ( n2141 & n6957 ) | ( ~n6956 & n6957 ) ;
  assign n6959 = n6478 | n6792 ;
  assign n6960 = n2339 ^ n1481 ^ 1'b0 ;
  assign n6961 = ( n331 & n1973 ) | ( n331 & ~n2621 ) | ( n1973 & ~n2621 ) ;
  assign n6962 = n2952 | n6961 ;
  assign n6963 = n6962 ^ n6090 ^ 1'b0 ;
  assign n6964 = n233 & ~n5599 ;
  assign n6965 = n6964 ^ n5379 ^ n5246 ;
  assign n6966 = ( n6960 & ~n6963 ) | ( n6960 & n6965 ) | ( ~n6963 & n6965 ) ;
  assign n6967 = ( ~n963 & n3102 ) | ( ~n963 & n3489 ) | ( n3102 & n3489 ) ;
  assign n6968 = n6967 ^ n1910 ^ n1230 ;
  assign n6969 = n1376 | n2212 ;
  assign n6970 = n6969 ^ n1682 ^ 1'b0 ;
  assign n6971 = ( n3561 & n6968 ) | ( n3561 & n6970 ) | ( n6968 & n6970 ) ;
  assign n6972 = ~n543 & n6971 ;
  assign n6973 = n4701 ^ n3421 ^ n1741 ;
  assign n6974 = n2578 ^ n1729 ^ 1'b0 ;
  assign n6975 = ( n760 & n1290 ) | ( n760 & n6974 ) | ( n1290 & n6974 ) ;
  assign n6976 = n6975 ^ n5818 ^ n4385 ;
  assign n6977 = ( n2524 & ~n6973 ) | ( n2524 & n6976 ) | ( ~n6973 & n6976 ) ;
  assign n6978 = n6972 & n6977 ;
  assign n6979 = ( n2552 & n3478 ) | ( n2552 & ~n6812 ) | ( n3478 & ~n6812 ) ;
  assign n6980 = n6979 ^ n2800 ^ 1'b0 ;
  assign n6981 = n3651 ^ n1912 ^ 1'b0 ;
  assign n6982 = n2434 & ~n6981 ;
  assign n6983 = n6982 ^ n6335 ^ n2568 ;
  assign n6984 = n6983 ^ n5935 ^ n2909 ;
  assign n6985 = n1738 ^ n820 ^ n360 ;
  assign n6986 = ~n766 & n6985 ;
  assign n6987 = ~n2989 & n6986 ;
  assign n6988 = ( n2729 & n4948 ) | ( n2729 & ~n6746 ) | ( n4948 & ~n6746 ) ;
  assign n6989 = n1220 ^ n411 ^ 1'b0 ;
  assign n6990 = x15 & n6989 ;
  assign n6991 = ( n1212 & n2225 ) | ( n1212 & n5241 ) | ( n2225 & n5241 ) ;
  assign n6992 = ( n3526 & n6990 ) | ( n3526 & ~n6991 ) | ( n6990 & ~n6991 ) ;
  assign n6993 = ( n6987 & n6988 ) | ( n6987 & n6992 ) | ( n6988 & n6992 ) ;
  assign n6994 = n6071 ^ n5646 ^ n2234 ;
  assign n6995 = n3016 ^ n1715 ^ x40 ;
  assign n6996 = n6886 ^ n719 ^ 1'b0 ;
  assign n6997 = ( n2032 & n6995 ) | ( n2032 & ~n6996 ) | ( n6995 & ~n6996 ) ;
  assign n6998 = ( n277 & n6994 ) | ( n277 & ~n6997 ) | ( n6994 & ~n6997 ) ;
  assign n6999 = ~n2178 & n2959 ;
  assign n7000 = ( ~n6187 & n6195 ) | ( ~n6187 & n6999 ) | ( n6195 & n6999 ) ;
  assign n7001 = n5033 ^ n1610 ^ 1'b0 ;
  assign n7002 = n7000 & n7001 ;
  assign n7003 = n2024 ^ n1640 ^ n1273 ;
  assign n7004 = ( n1430 & n6065 ) | ( n1430 & ~n7003 ) | ( n6065 & ~n7003 ) ;
  assign n7005 = ~n3066 & n7004 ;
  assign n7006 = n7005 ^ n4798 ^ 1'b0 ;
  assign n7007 = ~n6407 & n7006 ;
  assign n7008 = ~n7002 & n7007 ;
  assign n7009 = n4884 ^ n2079 ^ 1'b0 ;
  assign n7010 = n4333 & n7009 ;
  assign n7012 = n3900 ^ n3770 ^ n2305 ;
  assign n7013 = n2379 ^ n2258 ^ 1'b0 ;
  assign n7014 = ( n1148 & ~n7012 ) | ( n1148 & n7013 ) | ( ~n7012 & n7013 ) ;
  assign n7015 = n7014 ^ n1650 ^ 1'b0 ;
  assign n7011 = ~n4150 & n5657 ;
  assign n7016 = n7015 ^ n7011 ^ 1'b0 ;
  assign n7017 = n3917 ^ n1517 ^ n1021 ;
  assign n7018 = ~n2015 & n4632 ;
  assign n7020 = n2791 ^ n480 ^ 1'b0 ;
  assign n7021 = ~n998 & n7020 ;
  assign n7022 = ~n2141 & n7021 ;
  assign n7019 = n395 & ~n2185 ;
  assign n7023 = n7022 ^ n7019 ^ 1'b0 ;
  assign n7024 = n537 | n928 ;
  assign n7025 = n5547 & ~n7024 ;
  assign n7026 = n5293 ^ n699 ^ 1'b0 ;
  assign n7027 = n2811 & ~n7026 ;
  assign n7035 = ( n267 & n4090 ) | ( n267 & n4492 ) | ( n4090 & n4492 ) ;
  assign n7036 = n2417 ^ n1595 ^ n1130 ;
  assign n7037 = n445 & ~n7036 ;
  assign n7038 = ( n3049 & ~n7035 ) | ( n3049 & n7037 ) | ( ~n7035 & n7037 ) ;
  assign n7032 = n2495 ^ n1121 ^ 1'b0 ;
  assign n7033 = n2949 | n7032 ;
  assign n7028 = n3699 ^ n537 ^ x92 ;
  assign n7029 = n7028 ^ n3898 ^ n2129 ;
  assign n7030 = ( n991 & n1993 ) | ( n991 & n3191 ) | ( n1993 & n3191 ) ;
  assign n7031 = n7029 | n7030 ;
  assign n7034 = n7033 ^ n7031 ^ n6899 ;
  assign n7039 = n7038 ^ n7034 ^ n2377 ;
  assign n7040 = n2857 ^ x111 ^ 1'b0 ;
  assign n7041 = n7040 ^ n2660 ^ n1804 ;
  assign n7042 = ~n1425 & n7041 ;
  assign n7044 = n2562 & ~n5277 ;
  assign n7045 = n7044 ^ n277 ^ 1'b0 ;
  assign n7043 = n3385 ^ n2464 ^ n373 ;
  assign n7046 = n7045 ^ n7043 ^ n6805 ;
  assign n7047 = ( n3271 & n4996 ) | ( n3271 & n7046 ) | ( n4996 & n7046 ) ;
  assign n7048 = n5880 ^ n3127 ^ 1'b0 ;
  assign n7049 = ~n6544 & n7048 ;
  assign n7050 = ( ~n1819 & n1927 ) | ( ~n1819 & n5652 ) | ( n1927 & n5652 ) ;
  assign n7051 = ( n4977 & n6309 ) | ( n4977 & n7050 ) | ( n6309 & n7050 ) ;
  assign n7052 = ( n3187 & n4743 ) | ( n3187 & n5445 ) | ( n4743 & n5445 ) ;
  assign n7053 = n7052 ^ n4212 ^ n1367 ;
  assign n7054 = n2376 & n7053 ;
  assign n7055 = n7054 ^ n4130 ^ 1'b0 ;
  assign n7056 = n3714 ^ n2221 ^ n1287 ;
  assign n7057 = ( n271 & n3684 ) | ( n271 & ~n5184 ) | ( n3684 & ~n5184 ) ;
  assign n7058 = ( ~n4154 & n7056 ) | ( ~n4154 & n7057 ) | ( n7056 & n7057 ) ;
  assign n7066 = n3120 ^ n1925 ^ n1284 ;
  assign n7062 = n6589 ^ n4746 ^ n2918 ;
  assign n7063 = n7062 ^ n5296 ^ n4488 ;
  assign n7064 = ( ~n585 & n2071 ) | ( ~n585 & n7063 ) | ( n2071 & n7063 ) ;
  assign n7065 = n7064 ^ n6289 ^ n2115 ;
  assign n7059 = n1118 ^ n689 ^ n144 ;
  assign n7060 = n7059 ^ n3330 ^ n1537 ;
  assign n7061 = x57 & n7060 ;
  assign n7067 = n7066 ^ n7065 ^ n7061 ;
  assign n7068 = ( n2886 & n4261 ) | ( n2886 & n4966 ) | ( n4261 & n4966 ) ;
  assign n7069 = ~n3285 & n7068 ;
  assign n7070 = ~n2886 & n7069 ;
  assign n7075 = n3138 & n4485 ;
  assign n7076 = n239 & n7075 ;
  assign n7077 = n214 & ~n1125 ;
  assign n7078 = n3072 | n7077 ;
  assign n7079 = n7076 & ~n7078 ;
  assign n7080 = n7079 ^ n2296 ^ n1362 ;
  assign n7071 = n4751 ^ x42 ^ 1'b0 ;
  assign n7072 = n346 | n7071 ;
  assign n7073 = n7072 ^ n5424 ^ n4670 ;
  assign n7074 = n6123 & n7073 ;
  assign n7081 = n7080 ^ n7074 ^ 1'b0 ;
  assign n7082 = ~n767 & n2612 ;
  assign n7083 = ~n5589 & n7082 ;
  assign n7084 = n7083 ^ n2592 ^ n2488 ;
  assign n7085 = n7084 ^ n2112 ^ n541 ;
  assign n7086 = ( n1315 & ~n1411 ) | ( n1315 & n1480 ) | ( ~n1411 & n1480 ) ;
  assign n7087 = n4756 & ~n7086 ;
  assign n7088 = ( ~n1047 & n1449 ) | ( ~n1047 & n6029 ) | ( n1449 & n6029 ) ;
  assign n7089 = n7088 ^ n2965 ^ n1355 ;
  assign n7090 = n5509 ^ n1982 ^ n214 ;
  assign n7091 = n7090 ^ n4102 ^ 1'b0 ;
  assign n7092 = n7091 ^ n2805 ^ n748 ;
  assign n7093 = n6794 ^ n1235 ^ 1'b0 ;
  assign n7095 = ~n1266 & n4704 ;
  assign n7096 = n5793 & n7095 ;
  assign n7094 = n5931 ^ n5198 ^ 1'b0 ;
  assign n7097 = n7096 ^ n7094 ^ n2949 ;
  assign n7098 = n1569 ^ n1181 ^ n974 ;
  assign n7099 = n7098 ^ n3021 ^ 1'b0 ;
  assign n7100 = n2779 & ~n7099 ;
  assign n7101 = n3100 | n3408 ;
  assign n7102 = n6631 | n7101 ;
  assign n7103 = ( n2548 & n4646 ) | ( n2548 & n5414 ) | ( n4646 & n5414 ) ;
  assign n7104 = n6212 & ~n7103 ;
  assign n7105 = n7104 ^ n5525 ^ 1'b0 ;
  assign n7106 = n2697 ^ n1764 ^ x32 ;
  assign n7107 = n7106 ^ n6452 ^ n1809 ;
  assign n7108 = n5732 ^ n5202 ^ n3080 ;
  assign n7109 = n7108 ^ n4081 ^ 1'b0 ;
  assign n7110 = n258 & ~n5800 ;
  assign n7111 = n7110 ^ n1936 ^ n1485 ;
  assign n7112 = n3151 ^ n2931 ^ 1'b0 ;
  assign n7113 = ( n2754 & n3156 ) | ( n2754 & n7112 ) | ( n3156 & n7112 ) ;
  assign n7114 = ( n4174 & ~n7111 ) | ( n4174 & n7113 ) | ( ~n7111 & n7113 ) ;
  assign n7115 = n7114 ^ n5349 ^ n2873 ;
  assign n7116 = ~n2742 & n3379 ;
  assign n7117 = n7116 ^ n2210 ^ 1'b0 ;
  assign n7118 = ( ~n1517 & n6590 ) | ( ~n1517 & n7117 ) | ( n6590 & n7117 ) ;
  assign n7122 = n4033 ^ n3121 ^ x98 ;
  assign n7119 = n2698 & ~n4585 ;
  assign n7120 = n7119 ^ n6363 ^ 1'b0 ;
  assign n7121 = n7120 ^ n5833 ^ 1'b0 ;
  assign n7123 = n7122 ^ n7121 ^ n4684 ;
  assign n7124 = n1373 & ~n6150 ;
  assign n7125 = n7124 ^ n4798 ^ n3096 ;
  assign n7126 = ( ~n4307 & n5244 ) | ( ~n4307 & n7125 ) | ( n5244 & n7125 ) ;
  assign n7127 = n1722 | n2495 ;
  assign n7133 = n2243 ^ n743 ^ n290 ;
  assign n7134 = n4425 ^ n2214 ^ x66 ;
  assign n7135 = ( n3611 & n7133 ) | ( n3611 & n7134 ) | ( n7133 & n7134 ) ;
  assign n7136 = n5244 & n7135 ;
  assign n7128 = ~n839 & n1280 ;
  assign n7129 = ~n5336 & n7128 ;
  assign n7130 = n2596 & ~n7129 ;
  assign n7131 = n3495 & n7130 ;
  assign n7132 = n7131 ^ n3224 ^ 1'b0 ;
  assign n7137 = n7136 ^ n7132 ^ x24 ;
  assign n7138 = n1336 ^ n339 ^ n266 ;
  assign n7139 = ( ~n1261 & n5710 ) | ( ~n1261 & n7138 ) | ( n5710 & n7138 ) ;
  assign n7140 = n7139 ^ n954 ^ 1'b0 ;
  assign n7141 = n4083 & n7140 ;
  assign n7142 = n3021 ^ n2249 ^ 1'b0 ;
  assign n7143 = n7141 & ~n7142 ;
  assign n7144 = ( n192 & n303 ) | ( n192 & n1124 ) | ( n303 & n1124 ) ;
  assign n7145 = ( x36 & n505 ) | ( x36 & ~n2702 ) | ( n505 & ~n2702 ) ;
  assign n7146 = n7145 ^ n5687 ^ x127 ;
  assign n7147 = n7146 ^ n1713 ^ n1140 ;
  assign n7148 = ( ~n2668 & n2997 ) | ( ~n2668 & n7147 ) | ( n2997 & n7147 ) ;
  assign n7149 = ( n148 & n3518 ) | ( n148 & ~n4675 ) | ( n3518 & ~n4675 ) ;
  assign n7150 = ( n3528 & ~n3898 ) | ( n3528 & n7149 ) | ( ~n3898 & n7149 ) ;
  assign n7151 = n7148 & n7150 ;
  assign n7152 = n6555 & n7151 ;
  assign n7153 = n7152 ^ n3786 ^ n1904 ;
  assign n7155 = n2276 ^ n1222 ^ n827 ;
  assign n7154 = n2753 ^ n2608 ^ n2280 ;
  assign n7156 = n7155 ^ n7154 ^ 1'b0 ;
  assign n7157 = x113 & n7156 ;
  assign n7162 = n843 & ~n1079 ;
  assign n7163 = n7162 ^ n418 ^ 1'b0 ;
  assign n7164 = ( ~n1772 & n4241 ) | ( ~n1772 & n7163 ) | ( n4241 & n7163 ) ;
  assign n7159 = ( x82 & n369 ) | ( x82 & ~n6854 ) | ( n369 & ~n6854 ) ;
  assign n7160 = ( n313 & ~n1284 ) | ( n313 & n7159 ) | ( ~n1284 & n7159 ) ;
  assign n7158 = n3775 & n5372 ;
  assign n7161 = n7160 ^ n7158 ^ n728 ;
  assign n7165 = n7164 ^ n7161 ^ n3691 ;
  assign n7166 = n7165 ^ n7018 ^ n4155 ;
  assign n7168 = ( x75 & ~n1082 ) | ( x75 & n4205 ) | ( ~n1082 & n4205 ) ;
  assign n7167 = n3250 | n5398 ;
  assign n7169 = n7168 ^ n7167 ^ 1'b0 ;
  assign n7170 = n5058 & n7169 ;
  assign n7171 = n261 & ~n2294 ;
  assign n7172 = n3969 | n7171 ;
  assign n7173 = n7172 ^ n596 ^ 1'b0 ;
  assign n7174 = ( n2175 & n6002 ) | ( n2175 & n7173 ) | ( n6002 & n7173 ) ;
  assign n7175 = ( n5550 & n7170 ) | ( n5550 & ~n7174 ) | ( n7170 & ~n7174 ) ;
  assign n7177 = ( n218 & ~n405 ) | ( n218 & n4519 ) | ( ~n405 & n4519 ) ;
  assign n7176 = ( n1313 & ~n3248 ) | ( n1313 & n6939 ) | ( ~n3248 & n6939 ) ;
  assign n7178 = n7177 ^ n7176 ^ n4103 ;
  assign n7179 = ( ~n1861 & n4029 ) | ( ~n1861 & n4947 ) | ( n4029 & n4947 ) ;
  assign n7180 = ( n190 & n2105 ) | ( n190 & n7179 ) | ( n2105 & n7179 ) ;
  assign n7181 = n4461 | n7180 ;
  assign n7182 = x7 | n7181 ;
  assign n7183 = n7182 ^ n1445 ^ 1'b0 ;
  assign n7184 = n5817 | n7183 ;
  assign n7188 = n1407 & ~n3175 ;
  assign n7189 = n7188 ^ x108 ^ 1'b0 ;
  assign n7185 = ( x63 & ~n231 ) | ( x63 & n3626 ) | ( ~n231 & n3626 ) ;
  assign n7186 = n3928 & n7185 ;
  assign n7187 = ~n1984 & n7186 ;
  assign n7190 = n7189 ^ n7187 ^ n3113 ;
  assign n7191 = n5726 | n7190 ;
  assign n7192 = ~n3055 & n6871 ;
  assign n7194 = ( ~n1880 & n1992 ) | ( ~n1880 & n4000 ) | ( n1992 & n4000 ) ;
  assign n7193 = ( n518 & ~n1176 ) | ( n518 & n5615 ) | ( ~n1176 & n5615 ) ;
  assign n7195 = n7194 ^ n7193 ^ 1'b0 ;
  assign n7196 = n7192 | n7195 ;
  assign n7197 = ( n1583 & n2803 ) | ( n1583 & ~n3693 ) | ( n2803 & ~n3693 ) ;
  assign n7198 = n2330 ^ n2117 ^ n1703 ;
  assign n7200 = n2015 ^ n628 ^ 1'b0 ;
  assign n7199 = n6185 ^ n2632 ^ n1541 ;
  assign n7201 = n7200 ^ n7199 ^ 1'b0 ;
  assign n7202 = n1370 ^ n413 ^ x65 ;
  assign n7203 = n2592 | n7202 ;
  assign n7204 = n7203 ^ n643 ^ 1'b0 ;
  assign n7205 = ( n1061 & ~n4530 ) | ( n1061 & n7204 ) | ( ~n4530 & n7204 ) ;
  assign n7206 = ( n7198 & ~n7201 ) | ( n7198 & n7205 ) | ( ~n7201 & n7205 ) ;
  assign n7209 = n2739 ^ n2237 ^ x8 ;
  assign n7210 = ( ~n1623 & n6933 ) | ( ~n1623 & n7209 ) | ( n6933 & n7209 ) ;
  assign n7211 = n7210 ^ n617 ^ n603 ;
  assign n7207 = n4104 ^ n2156 ^ 1'b0 ;
  assign n7208 = n3361 & n7207 ;
  assign n7212 = n7211 ^ n7208 ^ 1'b0 ;
  assign n7213 = n1205 ^ n627 ^ 1'b0 ;
  assign n7214 = n5957 & n7213 ;
  assign n7215 = ( x112 & n812 ) | ( x112 & ~n2094 ) | ( n812 & ~n2094 ) ;
  assign n7216 = n7215 ^ n3847 ^ n992 ;
  assign n7217 = ( ~n455 & n7214 ) | ( ~n455 & n7216 ) | ( n7214 & n7216 ) ;
  assign n7218 = ( n411 & ~n4311 ) | ( n411 & n7217 ) | ( ~n4311 & n7217 ) ;
  assign n7219 = n4952 ^ n4092 ^ 1'b0 ;
  assign n7220 = ~n4611 & n7219 ;
  assign n7221 = ~n4475 & n7220 ;
  assign n7222 = n7221 ^ n3131 ^ 1'b0 ;
  assign n7223 = n7218 & ~n7222 ;
  assign n7224 = n3690 ^ n1171 ^ n826 ;
  assign n7225 = ( n685 & ~n2630 ) | ( n685 & n7224 ) | ( ~n2630 & n7224 ) ;
  assign n7226 = n7225 ^ n6688 ^ 1'b0 ;
  assign n7228 = n418 | n3632 ;
  assign n7229 = n7228 ^ n4343 ^ 1'b0 ;
  assign n7227 = n2536 & n5724 ;
  assign n7230 = n7229 ^ n7227 ^ 1'b0 ;
  assign n7231 = n669 & ~n3336 ;
  assign n7232 = n7231 ^ x25 ^ 1'b0 ;
  assign n7233 = n2518 & ~n7232 ;
  assign n7234 = n5442 ^ n1371 ^ n708 ;
  assign n7235 = n7234 ^ n1183 ^ 1'b0 ;
  assign n7236 = ~n1228 & n7235 ;
  assign n7237 = ( n4950 & n7233 ) | ( n4950 & ~n7236 ) | ( n7233 & ~n7236 ) ;
  assign n7239 = n6087 ^ n5761 ^ n3187 ;
  assign n7238 = n1720 | n3901 ;
  assign n7240 = n7239 ^ n7238 ^ 1'b0 ;
  assign n7241 = n6612 ^ n2676 ^ 1'b0 ;
  assign n7242 = n2147 ^ n1114 ^ n433 ;
  assign n7243 = n2149 ^ x44 ^ 1'b0 ;
  assign n7244 = n938 | n7243 ;
  assign n7245 = n7244 ^ n3327 ^ n988 ;
  assign n7246 = n7245 ^ n5383 ^ n2185 ;
  assign n7247 = ( ~n4458 & n7242 ) | ( ~n4458 & n7246 ) | ( n7242 & n7246 ) ;
  assign n7248 = n2518 & n5149 ;
  assign n7249 = ~n5394 & n7248 ;
  assign n7250 = ~n4789 & n5032 ;
  assign n7251 = n7250 ^ n1927 ^ 1'b0 ;
  assign n7252 = ~n7249 & n7251 ;
  assign n7258 = x68 & n823 ;
  assign n7259 = n2610 & n7258 ;
  assign n7260 = n7259 ^ n4640 ^ n2276 ;
  assign n7253 = n520 | n2329 ;
  assign n7254 = n1824 & ~n7253 ;
  assign n7255 = n1301 | n7254 ;
  assign n7256 = n3075 | n7255 ;
  assign n7257 = n3202 & n7256 ;
  assign n7261 = n7260 ^ n7257 ^ 1'b0 ;
  assign n7262 = ( n2448 & n2952 ) | ( n2448 & ~n3543 ) | ( n2952 & ~n3543 ) ;
  assign n7263 = n2961 | n7262 ;
  assign n7264 = n7263 ^ n2775 ^ 1'b0 ;
  assign n7265 = ~n2125 & n3382 ;
  assign n7266 = n7264 | n7265 ;
  assign n7267 = n2099 & n7266 ;
  assign n7268 = ( n143 & ~n2465 ) | ( n143 & n6424 ) | ( ~n2465 & n6424 ) ;
  assign n7269 = n4989 & n7268 ;
  assign n7270 = n203 & n214 ;
  assign n7271 = n4346 ^ x40 ^ 1'b0 ;
  assign n7272 = n489 & ~n7271 ;
  assign n7273 = ~n2862 & n7272 ;
  assign n7274 = n7270 & n7273 ;
  assign n7275 = n7274 ^ n6487 ^ n3680 ;
  assign n7276 = ( n4574 & ~n5065 ) | ( n4574 & n7275 ) | ( ~n5065 & n7275 ) ;
  assign n7277 = n5634 ^ n5191 ^ n3001 ;
  assign n7278 = n7277 ^ n1516 ^ 1'b0 ;
  assign n7279 = ~n6332 & n7278 ;
  assign n7280 = ( ~n3462 & n3783 ) | ( ~n3462 & n5162 ) | ( n3783 & n5162 ) ;
  assign n7282 = n705 & n2792 ;
  assign n7281 = ( n153 & n1989 ) | ( n153 & n4497 ) | ( n1989 & n4497 ) ;
  assign n7283 = n7282 ^ n7281 ^ 1'b0 ;
  assign n7284 = ~n7280 & n7283 ;
  assign n7285 = n7284 ^ n2350 ^ n762 ;
  assign n7286 = n2541 & n3267 ;
  assign n7287 = n6001 ^ n5337 ^ n343 ;
  assign n7288 = n880 | n7287 ;
  assign n7296 = ( n1663 & n4575 ) | ( n1663 & n6414 ) | ( n4575 & n6414 ) ;
  assign n7297 = ( n667 & n3860 ) | ( n667 & n7296 ) | ( n3860 & n7296 ) ;
  assign n7289 = n840 ^ n408 ^ 1'b0 ;
  assign n7290 = n1297 | n1524 ;
  assign n7291 = n5865 | n7290 ;
  assign n7292 = n4575 | n7291 ;
  assign n7293 = ~n2015 & n7292 ;
  assign n7294 = n4527 & n7293 ;
  assign n7295 = ( n2283 & n7289 ) | ( n2283 & n7294 ) | ( n7289 & n7294 ) ;
  assign n7298 = n7297 ^ n7295 ^ n2946 ;
  assign n7299 = n2224 ^ n1442 ^ n704 ;
  assign n7300 = x37 & n7299 ;
  assign n7301 = ~x72 & n7300 ;
  assign n7302 = n5948 & ~n7301 ;
  assign n7303 = n7302 ^ n4275 ^ 1'b0 ;
  assign n7304 = ( ~n975 & n2248 ) | ( ~n975 & n5027 ) | ( n2248 & n5027 ) ;
  assign n7305 = n7179 & n7304 ;
  assign n7306 = ~n1268 & n7305 ;
  assign n7307 = n7303 & ~n7306 ;
  assign n7308 = n5405 & n7307 ;
  assign n7310 = n294 & ~n3851 ;
  assign n7311 = ~n1441 & n7310 ;
  assign n7309 = n6018 ^ n1544 ^ n572 ;
  assign n7312 = n7311 ^ n7309 ^ n3483 ;
  assign n7313 = ~n3796 & n7312 ;
  assign n7314 = n6294 ^ n5746 ^ 1'b0 ;
  assign n7315 = ( ~n485 & n5346 ) | ( ~n485 & n7314 ) | ( n5346 & n7314 ) ;
  assign n7316 = n4740 ^ n1399 ^ 1'b0 ;
  assign n7317 = n2324 ^ n1931 ^ n1800 ;
  assign n7318 = ~n916 & n5332 ;
  assign n7319 = ( n2581 & n7317 ) | ( n2581 & ~n7318 ) | ( n7317 & ~n7318 ) ;
  assign n7320 = n7316 & ~n7319 ;
  assign n7321 = ( ~n1698 & n3023 ) | ( ~n1698 & n5490 ) | ( n3023 & n5490 ) ;
  assign n7322 = n7321 ^ n4201 ^ n264 ;
  assign n7323 = ( n390 & n1349 ) | ( n390 & ~n2765 ) | ( n1349 & ~n2765 ) ;
  assign n7324 = n7323 ^ n6721 ^ n5982 ;
  assign n7326 = n3657 ^ n3101 ^ 1'b0 ;
  assign n7327 = n7043 & ~n7326 ;
  assign n7325 = n3652 | n6294 ;
  assign n7328 = n7327 ^ n7325 ^ 1'b0 ;
  assign n7331 = n1136 ^ n467 ^ 1'b0 ;
  assign n7332 = n4739 | n7331 ;
  assign n7329 = n6280 ^ n3503 ^ 1'b0 ;
  assign n7330 = ~n3825 & n7329 ;
  assign n7333 = n7332 ^ n7330 ^ n4030 ;
  assign n7334 = n7333 ^ n5985 ^ n1659 ;
  assign n7335 = n7334 ^ n3118 ^ n553 ;
  assign n7336 = ( n1792 & n2134 ) | ( n1792 & ~n3764 ) | ( n2134 & ~n3764 ) ;
  assign n7337 = n6938 ^ n2560 ^ x69 ;
  assign n7338 = n7336 | n7337 ;
  assign n7339 = n1765 & ~n1940 ;
  assign n7340 = n7339 ^ n6069 ^ n2360 ;
  assign n7341 = n7340 ^ n6288 ^ n810 ;
  assign n7342 = ( ~n2376 & n4008 ) | ( ~n2376 & n7341 ) | ( n4008 & n7341 ) ;
  assign n7343 = ( ~n6909 & n7338 ) | ( ~n6909 & n7342 ) | ( n7338 & n7342 ) ;
  assign n7344 = ( n1975 & n4896 ) | ( n1975 & n7343 ) | ( n4896 & n7343 ) ;
  assign n7345 = n4121 ^ n3944 ^ 1'b0 ;
  assign n7346 = n1703 | n7345 ;
  assign n7347 = n2053 ^ n2047 ^ 1'b0 ;
  assign n7348 = n7347 ^ n3840 ^ n908 ;
  assign n7349 = ( n2305 & n2372 ) | ( n2305 & ~n4677 ) | ( n2372 & ~n4677 ) ;
  assign n7356 = x59 & n3712 ;
  assign n7357 = n7356 ^ n1597 ^ 1'b0 ;
  assign n7350 = n4304 ^ n2805 ^ n1376 ;
  assign n7351 = ( x102 & n5241 ) | ( x102 & ~n6651 ) | ( n5241 & ~n6651 ) ;
  assign n7352 = ( n3752 & ~n4255 ) | ( n3752 & n7351 ) | ( ~n4255 & n7351 ) ;
  assign n7353 = ( n2982 & ~n7350 ) | ( n2982 & n7352 ) | ( ~n7350 & n7352 ) ;
  assign n7354 = n2778 & ~n7353 ;
  assign n7355 = n3543 & n7354 ;
  assign n7358 = n7357 ^ n7355 ^ 1'b0 ;
  assign n7359 = ( n1437 & n1751 ) | ( n1437 & n2140 ) | ( n1751 & n2140 ) ;
  assign n7360 = ( n2851 & ~n4815 ) | ( n2851 & n7359 ) | ( ~n4815 & n7359 ) ;
  assign n7361 = ( n1645 & n3381 ) | ( n1645 & n7360 ) | ( n3381 & n7360 ) ;
  assign n7362 = n4662 ^ n4332 ^ x16 ;
  assign n7366 = n6950 ^ n2624 ^ 1'b0 ;
  assign n7367 = ~n3583 & n7366 ;
  assign n7363 = n1260 & ~n2271 ;
  assign n7364 = n7363 ^ n1332 ^ 1'b0 ;
  assign n7365 = n7364 ^ n3515 ^ n2191 ;
  assign n7368 = n7367 ^ n7365 ^ n5228 ;
  assign n7369 = ( n1661 & n1699 ) | ( n1661 & n5908 ) | ( n1699 & n5908 ) ;
  assign n7370 = n7369 ^ n3621 ^ 1'b0 ;
  assign n7376 = ( ~n1653 & n2643 ) | ( ~n1653 & n2791 ) | ( n2643 & n2791 ) ;
  assign n7372 = ~n1472 & n5275 ;
  assign n7371 = n1391 | n5128 ;
  assign n7373 = n7372 ^ n7371 ^ n4650 ;
  assign n7374 = n4487 & ~n7373 ;
  assign n7375 = ~n2349 & n7374 ;
  assign n7377 = n7376 ^ n7375 ^ n4880 ;
  assign n7378 = ( ~n5464 & n7370 ) | ( ~n5464 & n7377 ) | ( n7370 & n7377 ) ;
  assign n7379 = ( n715 & ~n1775 ) | ( n715 & n1962 ) | ( ~n1775 & n1962 ) ;
  assign n7380 = ( n1012 & n2391 ) | ( n1012 & n7379 ) | ( n2391 & n7379 ) ;
  assign n7381 = n4951 ^ n3353 ^ n2927 ;
  assign n7382 = n3842 ^ n2101 ^ 1'b0 ;
  assign n7383 = n6938 ^ n6617 ^ n197 ;
  assign n7384 = n5400 ^ n2158 ^ n553 ;
  assign n7385 = ( n807 & ~n823 ) | ( n807 & n3783 ) | ( ~n823 & n3783 ) ;
  assign n7386 = n7385 ^ n4878 ^ 1'b0 ;
  assign n7387 = n7386 ^ n1424 ^ 1'b0 ;
  assign n7388 = ~n7384 & n7387 ;
  assign n7389 = ( n4105 & n7383 ) | ( n4105 & ~n7388 ) | ( n7383 & ~n7388 ) ;
  assign n7390 = ( ~n170 & n7382 ) | ( ~n170 & n7389 ) | ( n7382 & n7389 ) ;
  assign n7397 = x84 & n2429 ;
  assign n7398 = n1607 & n7397 ;
  assign n7395 = n2885 ^ n2072 ^ n364 ;
  assign n7396 = n7395 ^ n5984 ^ 1'b0 ;
  assign n7391 = n440 & ~n5187 ;
  assign n7392 = n7391 ^ n2246 ^ 1'b0 ;
  assign n7393 = n7392 ^ n1551 ^ 1'b0 ;
  assign n7394 = n4523 & ~n7393 ;
  assign n7399 = n7398 ^ n7396 ^ n7394 ;
  assign n7400 = n1877 ^ n1302 ^ n816 ;
  assign n7401 = n373 & n996 ;
  assign n7402 = ( n1256 & ~n7400 ) | ( n1256 & n7401 ) | ( ~n7400 & n7401 ) ;
  assign n7403 = n5313 ^ n4143 ^ 1'b0 ;
  assign n7404 = n4285 ^ n451 ^ 1'b0 ;
  assign n7405 = n7404 ^ n1829 ^ 1'b0 ;
  assign n7406 = n2779 ^ n1854 ^ n408 ;
  assign n7407 = n3575 ^ n852 ^ 1'b0 ;
  assign n7408 = ( n850 & ~n4399 ) | ( n850 & n7407 ) | ( ~n4399 & n7407 ) ;
  assign n7409 = ( n1714 & n1849 ) | ( n1714 & n7408 ) | ( n1849 & n7408 ) ;
  assign n7410 = ( n1494 & ~n7406 ) | ( n1494 & n7409 ) | ( ~n7406 & n7409 ) ;
  assign n7411 = n6238 ^ n3044 ^ n1015 ;
  assign n7412 = ( n724 & ~n3730 ) | ( n724 & n4000 ) | ( ~n3730 & n4000 ) ;
  assign n7413 = ( n1407 & n3147 ) | ( n1407 & n7412 ) | ( n3147 & n7412 ) ;
  assign n7414 = n2446 ^ n1966 ^ n1167 ;
  assign n7415 = n4551 ^ n4274 ^ n3879 ;
  assign n7416 = ( n777 & n4434 ) | ( n777 & ~n7415 ) | ( n4434 & ~n7415 ) ;
  assign n7417 = n7416 ^ n5993 ^ n3308 ;
  assign n7421 = n3906 | n6401 ;
  assign n7418 = ~n2721 & n3265 ;
  assign n7419 = n3967 ^ n2191 ^ n2120 ;
  assign n7420 = n7418 & ~n7419 ;
  assign n7422 = n7421 ^ n7420 ^ 1'b0 ;
  assign n7423 = n6328 & n7422 ;
  assign n7424 = ~n7018 & n7423 ;
  assign n7425 = ( n447 & n478 ) | ( n447 & ~n7378 ) | ( n478 & ~n7378 ) ;
  assign n7426 = n6499 ^ n4041 ^ 1'b0 ;
  assign n7427 = n4100 & n7426 ;
  assign n7428 = ~n912 & n1738 ;
  assign n7429 = ( n214 & n673 ) | ( n214 & ~n3103 ) | ( n673 & ~n3103 ) ;
  assign n7430 = ( n3789 & ~n7428 ) | ( n3789 & n7429 ) | ( ~n7428 & n7429 ) ;
  assign n7431 = n3657 | n7430 ;
  assign n7432 = ( n4934 & n7427 ) | ( n4934 & ~n7431 ) | ( n7427 & ~n7431 ) ;
  assign n7443 = n2497 ^ n1048 ^ 1'b0 ;
  assign n7436 = ~n4782 & n6908 ;
  assign n7437 = n7436 ^ n5710 ^ 1'b0 ;
  assign n7438 = n1366 & n7437 ;
  assign n7439 = n6671 & n7438 ;
  assign n7440 = n5241 ^ n4749 ^ 1'b0 ;
  assign n7441 = n7439 | n7440 ;
  assign n7442 = n6297 | n7441 ;
  assign n7434 = ( n2516 & n5813 ) | ( n2516 & ~n6218 ) | ( n5813 & ~n6218 ) ;
  assign n7433 = ~n1116 & n1762 ;
  assign n7435 = n7434 ^ n7433 ^ 1'b0 ;
  assign n7444 = n7443 ^ n7442 ^ n7435 ;
  assign n7445 = n7444 ^ n5681 ^ n916 ;
  assign n7446 = ( n3690 & n7432 ) | ( n3690 & n7445 ) | ( n7432 & n7445 ) ;
  assign n7447 = ( n1047 & ~n4345 ) | ( n1047 & n7446 ) | ( ~n4345 & n7446 ) ;
  assign n7448 = n1843 & ~n5004 ;
  assign n7449 = n6107 ^ n5070 ^ 1'b0 ;
  assign n7450 = ~n4425 & n7449 ;
  assign n7451 = n7448 & n7450 ;
  assign n7452 = n5058 ^ n3917 ^ 1'b0 ;
  assign n7453 = n1493 & n7452 ;
  assign n7454 = n7453 ^ n6360 ^ 1'b0 ;
  assign n7455 = ( n1629 & n2249 ) | ( n1629 & ~n7454 ) | ( n2249 & ~n7454 ) ;
  assign n7471 = n5698 ^ n2757 ^ 1'b0 ;
  assign n7468 = n1867 ^ n1265 ^ n445 ;
  assign n7469 = n3762 ^ n1455 ^ n471 ;
  assign n7470 = ~n7468 & n7469 ;
  assign n7472 = n7471 ^ n7470 ^ 1'b0 ;
  assign n7464 = n1559 & n1932 ;
  assign n7465 = n7464 ^ n2258 ^ 1'b0 ;
  assign n7466 = n7465 ^ n1256 ^ n375 ;
  assign n7467 = n7466 ^ n4782 ^ n357 ;
  assign n7462 = n1573 ^ n1413 ^ 1'b0 ;
  assign n7459 = n2465 ^ n380 ^ x18 ;
  assign n7460 = n1840 & ~n7459 ;
  assign n7456 = n3985 ^ n593 ^ 1'b0 ;
  assign n7457 = n3889 | n7456 ;
  assign n7458 = n3912 | n7457 ;
  assign n7461 = n7460 ^ n7458 ^ n4044 ;
  assign n7463 = n7462 ^ n7461 ^ n3830 ;
  assign n7473 = n7472 ^ n7467 ^ n7463 ;
  assign n7476 = ( ~x109 & n1650 ) | ( ~x109 & n5644 ) | ( n1650 & n5644 ) ;
  assign n7474 = n6532 ^ n5321 ^ n4406 ;
  assign n7475 = ( n3000 & n5507 ) | ( n3000 & n7474 ) | ( n5507 & n7474 ) ;
  assign n7477 = n7476 ^ n7475 ^ n226 ;
  assign n7479 = n890 ^ x88 ^ 1'b0 ;
  assign n7478 = n420 & ~n3446 ;
  assign n7480 = n7479 ^ n7478 ^ 1'b0 ;
  assign n7481 = n2454 & ~n3507 ;
  assign n7482 = n5124 & n5681 ;
  assign n7483 = ~n293 & n1828 ;
  assign n7484 = n2920 & ~n7483 ;
  assign n7485 = n7484 ^ n6954 ^ 1'b0 ;
  assign n7486 = n238 & n7485 ;
  assign n7487 = ~n1425 & n7486 ;
  assign n7488 = n2930 ^ n1699 ^ n1531 ;
  assign n7489 = ~n4507 & n7488 ;
  assign n7490 = n7489 ^ n4020 ^ n1221 ;
  assign n7491 = n1130 ^ n556 ^ 1'b0 ;
  assign n7492 = n5131 ^ n4190 ^ n2114 ;
  assign n7493 = n4762 ^ n4551 ^ n2069 ;
  assign n7494 = n4190 ^ n3115 ^ n1285 ;
  assign n7495 = ( n6823 & n7493 ) | ( n6823 & n7494 ) | ( n7493 & n7494 ) ;
  assign n7496 = n2256 & n2729 ;
  assign n7497 = n7496 ^ n3347 ^ 1'b0 ;
  assign n7498 = n2908 ^ n1716 ^ n362 ;
  assign n7499 = n2982 ^ n2558 ^ 1'b0 ;
  assign n7500 = ~n4034 & n7499 ;
  assign n7501 = ~n7498 & n7500 ;
  assign n7502 = n7497 & ~n7501 ;
  assign n7503 = ~n7495 & n7502 ;
  assign n7504 = n4979 ^ n3431 ^ 1'b0 ;
  assign n7505 = n2059 & ~n7504 ;
  assign n7506 = ( n1818 & n4077 ) | ( n1818 & ~n7505 ) | ( n4077 & ~n7505 ) ;
  assign n7507 = n4670 ^ n1301 ^ 1'b0 ;
  assign n7508 = n7507 ^ n4880 ^ 1'b0 ;
  assign n7509 = n5294 | n7508 ;
  assign n7510 = n7083 ^ n3953 ^ 1'b0 ;
  assign n7511 = n7510 ^ n6897 ^ n1028 ;
  assign n7512 = n212 | n4014 ;
  assign n7513 = n6230 | n7512 ;
  assign n7514 = ( n671 & ~n1304 ) | ( n671 & n4326 ) | ( ~n1304 & n4326 ) ;
  assign n7515 = ( n7511 & n7513 ) | ( n7511 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7516 = n4670 ^ n2311 ^ 1'b0 ;
  assign n7517 = n4730 & n7516 ;
  assign n7518 = n3917 | n7517 ;
  assign n7519 = n7518 ^ x17 ^ 1'b0 ;
  assign n7520 = ( n2041 & n7515 ) | ( n2041 & ~n7519 ) | ( n7515 & ~n7519 ) ;
  assign n7521 = ( n568 & n2747 ) | ( n568 & ~n5228 ) | ( n2747 & ~n5228 ) ;
  assign n7522 = ( ~n2058 & n6099 ) | ( ~n2058 & n7521 ) | ( n6099 & n7521 ) ;
  assign n7523 = ( ~n7509 & n7520 ) | ( ~n7509 & n7522 ) | ( n7520 & n7522 ) ;
  assign n7524 = n7523 ^ n3247 ^ 1'b0 ;
  assign n7525 = n5101 ^ n4966 ^ 1'b0 ;
  assign n7526 = n5081 | n7525 ;
  assign n7527 = ( n1042 & n2582 ) | ( n1042 & ~n4947 ) | ( n2582 & ~n4947 ) ;
  assign n7528 = n7527 ^ n6893 ^ n6752 ;
  assign n7529 = n953 ^ x79 ^ 1'b0 ;
  assign n7530 = n1964 & ~n7529 ;
  assign n7531 = n5321 ^ n3963 ^ n3024 ;
  assign n7532 = ~n6347 & n7531 ;
  assign n7533 = n7532 ^ n3263 ^ 1'b0 ;
  assign n7534 = n7530 & n7533 ;
  assign n7535 = n7534 ^ n5298 ^ 1'b0 ;
  assign n7536 = n7535 ^ n1895 ^ 1'b0 ;
  assign n7537 = n2563 & n7536 ;
  assign n7538 = ( ~n2933 & n4454 ) | ( ~n2933 & n5086 ) | ( n4454 & n5086 ) ;
  assign n7539 = n1481 & ~n7538 ;
  assign n7540 = n7539 ^ x88 ^ 1'b0 ;
  assign n7541 = n6660 & ~n6868 ;
  assign n7542 = ~n1485 & n7541 ;
  assign n7543 = ( ~n1015 & n2493 ) | ( ~n1015 & n7542 ) | ( n2493 & n7542 ) ;
  assign n7544 = ( x7 & n484 ) | ( x7 & ~n1698 ) | ( n484 & ~n1698 ) ;
  assign n7545 = ( ~n2528 & n2988 ) | ( ~n2528 & n3364 ) | ( n2988 & n3364 ) ;
  assign n7546 = ( ~n1254 & n7544 ) | ( ~n1254 & n7545 ) | ( n7544 & n7545 ) ;
  assign n7547 = n2085 ^ n2070 ^ n1411 ;
  assign n7548 = n7547 ^ n2265 ^ n1519 ;
  assign n7549 = ( n1808 & ~n6586 ) | ( n1808 & n7548 ) | ( ~n6586 & n7548 ) ;
  assign n7550 = n7546 & n7549 ;
  assign n7551 = n7543 & n7550 ;
  assign n7558 = n2036 & n4531 ;
  assign n7559 = ~n3257 & n7558 ;
  assign n7560 = n1519 ^ n1038 ^ x117 ;
  assign n7561 = ( n6830 & n7559 ) | ( n6830 & ~n7560 ) | ( n7559 & ~n7560 ) ;
  assign n7562 = n7561 ^ n2635 ^ 1'b0 ;
  assign n7563 = n7295 | n7562 ;
  assign n7552 = n466 | n5521 ;
  assign n7553 = n1640 & n5998 ;
  assign n7554 = n7553 ^ n4988 ^ 1'b0 ;
  assign n7555 = n7552 | n7554 ;
  assign n7556 = ( x99 & ~n3169 ) | ( x99 & n7555 ) | ( ~n3169 & n7555 ) ;
  assign n7557 = ~n6239 & n7556 ;
  assign n7564 = n7563 ^ n7557 ^ 1'b0 ;
  assign n7565 = n2694 ^ n1037 ^ n398 ;
  assign n7566 = n1397 & n7060 ;
  assign n7567 = n2485 & n7566 ;
  assign n7568 = n6125 ^ n5655 ^ n2005 ;
  assign n7569 = ( n2405 & n7567 ) | ( n2405 & ~n7568 ) | ( n7567 & ~n7568 ) ;
  assign n7570 = ~n1971 & n7556 ;
  assign n7571 = n2510 & n7570 ;
  assign n7572 = n2375 ^ n214 ^ x74 ;
  assign n7573 = ( n2168 & n2865 ) | ( n2168 & ~n7572 ) | ( n2865 & ~n7572 ) ;
  assign n7577 = n7012 ^ n2375 ^ n1991 ;
  assign n7575 = n6967 ^ n6016 ^ n5259 ;
  assign n7574 = ~n462 & n3986 ;
  assign n7576 = n7575 ^ n7574 ^ 1'b0 ;
  assign n7578 = n7577 ^ n7576 ^ n7050 ;
  assign n7585 = n3034 ^ n2072 ^ 1'b0 ;
  assign n7581 = ~n1461 & n2902 ;
  assign n7582 = n3485 & n7581 ;
  assign n7583 = n7582 ^ n1494 ^ n700 ;
  assign n7580 = n7159 ^ n1513 ^ 1'b0 ;
  assign n7584 = n7583 ^ n7580 ^ n795 ;
  assign n7579 = ( n1948 & ~n2709 ) | ( n1948 & n6795 ) | ( ~n2709 & n6795 ) ;
  assign n7586 = n7585 ^ n7584 ^ n7579 ;
  assign n7587 = n2321 & ~n2625 ;
  assign n7588 = n7587 ^ n4058 ^ 1'b0 ;
  assign n7596 = n1942 | n6073 ;
  assign n7589 = ( n2000 & n2406 ) | ( n2000 & n3167 ) | ( n2406 & n3167 ) ;
  assign n7590 = n5827 & n7589 ;
  assign n7591 = ~n945 & n7590 ;
  assign n7592 = n1190 & ~n3285 ;
  assign n7593 = ( n252 & n1150 ) | ( n252 & n7592 ) | ( n1150 & n7592 ) ;
  assign n7594 = ( n1766 & n7591 ) | ( n1766 & ~n7593 ) | ( n7591 & ~n7593 ) ;
  assign n7595 = n7594 ^ n7542 ^ n1332 ;
  assign n7597 = n7596 ^ n7595 ^ 1'b0 ;
  assign n7598 = n7588 | n7597 ;
  assign n7599 = n622 & n5136 ;
  assign n7600 = ~n1887 & n7599 ;
  assign n7601 = ~n3380 & n7164 ;
  assign n7602 = ( n719 & ~n4144 ) | ( n719 & n7601 ) | ( ~n4144 & n7601 ) ;
  assign n7603 = ( n227 & n825 ) | ( n227 & ~n7602 ) | ( n825 & ~n7602 ) ;
  assign n7604 = n4541 | n7369 ;
  assign n7605 = n7603 & ~n7604 ;
  assign n7606 = n5643 ^ n3127 ^ 1'b0 ;
  assign n7607 = ( x121 & n130 ) | ( x121 & ~n2040 ) | ( n130 & ~n2040 ) ;
  assign n7608 = n1058 & n3952 ;
  assign n7609 = n7607 | n7608 ;
  assign n7610 = n1900 | n7609 ;
  assign n7611 = n7610 ^ n974 ^ n226 ;
  assign n7612 = ( n910 & n1024 ) | ( n910 & ~n5827 ) | ( n1024 & ~n5827 ) ;
  assign n7613 = ( n928 & n2510 ) | ( n928 & ~n3333 ) | ( n2510 & ~n3333 ) ;
  assign n7614 = n3259 & n7613 ;
  assign n7615 = n4213 & n7614 ;
  assign n7616 = n7615 ^ n6520 ^ 1'b0 ;
  assign n7617 = n5086 & n7616 ;
  assign n7618 = n5816 | n7617 ;
  assign n7620 = n3173 & n5632 ;
  assign n7621 = n1290 | n7620 ;
  assign n7619 = ~n4052 & n4314 ;
  assign n7622 = n7621 ^ n7619 ^ 1'b0 ;
  assign n7623 = ~n3237 & n3462 ;
  assign n7624 = ~n6519 & n7623 ;
  assign n7625 = ( n952 & ~n3474 ) | ( n952 & n4474 ) | ( ~n3474 & n4474 ) ;
  assign n7626 = n6883 & n7625 ;
  assign n7627 = ( ~n862 & n1199 ) | ( ~n862 & n1886 ) | ( n1199 & n1886 ) ;
  assign n7628 = n2003 ^ n294 ^ 1'b0 ;
  assign n7629 = n7628 ^ x52 ^ 1'b0 ;
  assign n7630 = ~n3815 & n7629 ;
  assign n7631 = ( ~n364 & n2672 ) | ( ~n364 & n6055 ) | ( n2672 & n6055 ) ;
  assign n7632 = ( n2476 & n3049 ) | ( n2476 & n7631 ) | ( n3049 & n7631 ) ;
  assign n7633 = ( n6225 & n7630 ) | ( n6225 & ~n7632 ) | ( n7630 & ~n7632 ) ;
  assign n7634 = ( n1679 & n7627 ) | ( n1679 & n7633 ) | ( n7627 & n7633 ) ;
  assign n7635 = n7634 ^ n3646 ^ 1'b0 ;
  assign n7636 = n7626 & n7635 ;
  assign n7637 = n2073 & n5632 ;
  assign n7638 = n7637 ^ n3847 ^ 1'b0 ;
  assign n7639 = ( ~n218 & n898 ) | ( ~n218 & n7638 ) | ( n898 & n7638 ) ;
  assign n7640 = n2627 & ~n6130 ;
  assign n7641 = n7640 ^ n1550 ^ 1'b0 ;
  assign n7642 = n1305 & ~n7641 ;
  assign n7643 = ( n526 & n1353 ) | ( n526 & ~n5163 ) | ( n1353 & ~n5163 ) ;
  assign n7644 = n5705 ^ n1571 ^ 1'b0 ;
  assign n7645 = n440 & n3500 ;
  assign n7646 = n2467 & n7645 ;
  assign n7647 = ( ~n697 & n7644 ) | ( ~n697 & n7646 ) | ( n7644 & n7646 ) ;
  assign n7648 = n4867 & n6685 ;
  assign n7649 = ~n6967 & n7136 ;
  assign n7652 = ( n699 & ~n1732 ) | ( n699 & n2624 ) | ( ~n1732 & n2624 ) ;
  assign n7653 = n6956 ^ n2346 ^ 1'b0 ;
  assign n7654 = n7652 & ~n7653 ;
  assign n7650 = n1715 | n7512 ;
  assign n7651 = n7650 ^ n403 ^ 1'b0 ;
  assign n7655 = n7654 ^ n7651 ^ 1'b0 ;
  assign n7656 = ~n3889 & n7655 ;
  assign n7657 = n1981 & ~n2885 ;
  assign n7658 = n4403 & n7617 ;
  assign n7659 = n7657 & n7658 ;
  assign n7660 = ~n5206 & n5650 ;
  assign n7661 = n3840 & n7660 ;
  assign n7662 = ( n2736 & n6011 ) | ( n2736 & n7661 ) | ( n6011 & n7661 ) ;
  assign n7663 = ( n1769 & n7144 ) | ( n1769 & n7662 ) | ( n7144 & n7662 ) ;
  assign n7664 = n5883 | n6240 ;
  assign n7665 = n1982 & ~n7664 ;
  assign n7666 = n6019 | n6954 ;
  assign n7667 = n589 & ~n7666 ;
  assign n7668 = n5362 & ~n7667 ;
  assign n7669 = n7588 & n7668 ;
  assign n7670 = ( n4568 & n5622 ) | ( n4568 & n7669 ) | ( n5622 & n7669 ) ;
  assign n7671 = n7041 ^ n4914 ^ 1'b0 ;
  assign n7672 = n2465 & n7671 ;
  assign n7673 = n6437 ^ n3007 ^ n1342 ;
  assign n7674 = ( n3127 & n5354 ) | ( n3127 & ~n7673 ) | ( n5354 & ~n7673 ) ;
  assign n7679 = n1839 | n1977 ;
  assign n7680 = n7679 ^ n3910 ^ 1'b0 ;
  assign n7676 = n3509 ^ n1739 ^ n739 ;
  assign n7675 = n3783 ^ n3354 ^ n1727 ;
  assign n7677 = n7676 ^ n7675 ^ 1'b0 ;
  assign n7678 = n7677 ^ n4195 ^ n3054 ;
  assign n7681 = n7680 ^ n7678 ^ 1'b0 ;
  assign n7682 = ( n2656 & n4473 ) | ( n2656 & n6408 ) | ( n4473 & n6408 ) ;
  assign n7683 = n1982 ^ n898 ^ 1'b0 ;
  assign n7684 = n1729 ^ n1557 ^ 1'b0 ;
  assign n7685 = n4474 & n7684 ;
  assign n7686 = ( n751 & ~n2019 ) | ( n751 & n7685 ) | ( ~n2019 & n7685 ) ;
  assign n7687 = n6083 ^ n4195 ^ 1'b0 ;
  assign n7688 = ~n3331 & n7687 ;
  assign n7689 = ( ~n7683 & n7686 ) | ( ~n7683 & n7688 ) | ( n7686 & n7688 ) ;
  assign n7690 = ( ~n1842 & n2030 ) | ( ~n1842 & n2889 ) | ( n2030 & n2889 ) ;
  assign n7691 = n7690 ^ n3642 ^ 1'b0 ;
  assign n7692 = n7691 ^ n7559 ^ n4325 ;
  assign n7693 = n7689 | n7692 ;
  assign n7694 = n7682 & ~n7693 ;
  assign n7699 = ~n4000 & n4502 ;
  assign n7700 = ~n1239 & n7699 ;
  assign n7701 = n7700 ^ n2611 ^ n1650 ;
  assign n7702 = n3778 & ~n7701 ;
  assign n7703 = n1353 & ~n7702 ;
  assign n7704 = n5090 & ~n6055 ;
  assign n7705 = n7704 ^ n7409 ^ n6008 ;
  assign n7706 = ( n509 & n7703 ) | ( n509 & ~n7705 ) | ( n7703 & ~n7705 ) ;
  assign n7697 = n3181 ^ n2092 ^ 1'b0 ;
  assign n7695 = n3103 & n4256 ;
  assign n7696 = ( n2527 & ~n5504 ) | ( n2527 & n7695 ) | ( ~n5504 & n7695 ) ;
  assign n7698 = n7697 ^ n7696 ^ n1861 ;
  assign n7707 = n7706 ^ n7698 ^ 1'b0 ;
  assign n7708 = n2842 & n6214 ;
  assign n7709 = n4288 & n5285 ;
  assign n7710 = n7709 ^ n3641 ^ 1'b0 ;
  assign n7711 = n2124 | n7710 ;
  assign n7712 = n7711 ^ n2077 ^ 1'b0 ;
  assign n7713 = ~n2201 & n5738 ;
  assign n7714 = ( n2605 & ~n4256 ) | ( n2605 & n4954 ) | ( ~n4256 & n4954 ) ;
  assign n7715 = ( n3130 & ~n3734 ) | ( n3130 & n6284 ) | ( ~n3734 & n6284 ) ;
  assign n7716 = ( n859 & n7714 ) | ( n859 & ~n7715 ) | ( n7714 & ~n7715 ) ;
  assign n7717 = n5364 ^ n4878 ^ n1434 ;
  assign n7718 = n7717 ^ n6745 ^ n4903 ;
  assign n7719 = n4102 ^ n1929 ^ 1'b0 ;
  assign n7720 = n972 | n7719 ;
  assign n7721 = ( ~n145 & n2975 ) | ( ~n145 & n6908 ) | ( n2975 & n6908 ) ;
  assign n7722 = n7721 ^ n1407 ^ n495 ;
  assign n7723 = ~n1100 & n2840 ;
  assign n7724 = n7723 ^ n1890 ^ 1'b0 ;
  assign n7725 = n1434 & n6684 ;
  assign n7726 = ( n1028 & n3238 ) | ( n1028 & n7725 ) | ( n3238 & n7725 ) ;
  assign n7727 = n5312 & ~n7726 ;
  assign n7728 = n7727 ^ n7505 ^ 1'b0 ;
  assign n7729 = ( n3654 & ~n7724 ) | ( n3654 & n7728 ) | ( ~n7724 & n7728 ) ;
  assign n7730 = n5123 ^ n2029 ^ n1441 ;
  assign n7731 = ~n3620 & n4168 ;
  assign n7732 = ~n5773 & n7731 ;
  assign n7749 = n2530 & ~n5490 ;
  assign n7733 = n1282 | n3699 ;
  assign n7734 = n7733 ^ x63 ^ 1'b0 ;
  assign n7735 = ( n1718 & n4202 ) | ( n1718 & ~n7489 ) | ( n4202 & ~n7489 ) ;
  assign n7736 = ( n1122 & n7734 ) | ( n1122 & n7735 ) | ( n7734 & n7735 ) ;
  assign n7737 = n3452 ^ n768 ^ 1'b0 ;
  assign n7738 = ~n7736 & n7737 ;
  assign n7739 = n7738 ^ n5972 ^ n5467 ;
  assign n7740 = n5724 ^ n3035 ^ 1'b0 ;
  assign n7741 = n7740 ^ n3557 ^ 1'b0 ;
  assign n7742 = n6939 ^ n3008 ^ 1'b0 ;
  assign n7743 = n7741 | n7742 ;
  assign n7744 = ( n4918 & ~n5604 ) | ( n4918 & n6200 ) | ( ~n5604 & n6200 ) ;
  assign n7745 = n7744 ^ n1532 ^ 1'b0 ;
  assign n7746 = n3008 & n7745 ;
  assign n7747 = ( n7739 & n7743 ) | ( n7739 & n7746 ) | ( n7743 & n7746 ) ;
  assign n7748 = n7747 ^ n5882 ^ n3833 ;
  assign n7750 = n7749 ^ n7748 ^ n810 ;
  assign n7762 = n841 | n2120 ;
  assign n7763 = n7762 ^ n3139 ^ 1'b0 ;
  assign n7764 = n7763 ^ n3142 ^ 1'b0 ;
  assign n7765 = n1220 & ~n7764 ;
  assign n7766 = n7765 ^ n3481 ^ 1'b0 ;
  assign n7760 = ( n1216 & n1251 ) | ( n1216 & ~n1998 ) | ( n1251 & ~n1998 ) ;
  assign n7761 = ( n5077 & ~n6677 ) | ( n5077 & n7760 ) | ( ~n6677 & n7760 ) ;
  assign n7767 = n7766 ^ n7761 ^ n2469 ;
  assign n7755 = n6430 ^ n3854 ^ 1'b0 ;
  assign n7756 = n6645 | n7755 ;
  assign n7757 = n7337 & n7756 ;
  assign n7758 = ( ~n1976 & n5196 ) | ( ~n1976 & n7757 ) | ( n5196 & n7757 ) ;
  assign n7752 = ( n271 & ~n1329 ) | ( n271 & n2476 ) | ( ~n1329 & n2476 ) ;
  assign n7753 = n1788 & ~n2785 ;
  assign n7754 = n7752 & n7753 ;
  assign n7759 = n7758 ^ n7754 ^ n7549 ;
  assign n7751 = ( ~n389 & n1216 ) | ( ~n389 & n5827 ) | ( n1216 & n5827 ) ;
  assign n7768 = n7767 ^ n7759 ^ n7751 ;
  assign n7769 = n5630 ^ n1335 ^ 1'b0 ;
  assign n7770 = n7769 ^ n6083 ^ n4633 ;
  assign n7771 = n275 | n4374 ;
  assign n7772 = ~n1884 & n7771 ;
  assign n7773 = n7772 ^ n5277 ^ 1'b0 ;
  assign n7774 = ( n2222 & n7173 ) | ( n2222 & n7773 ) | ( n7173 & n7773 ) ;
  assign n7775 = n3729 ^ n708 ^ x4 ;
  assign n7776 = n7775 ^ n6437 ^ n1900 ;
  assign n7779 = n6933 ^ n3548 ^ n2531 ;
  assign n7778 = n2695 & n4168 ;
  assign n7777 = n4683 ^ n3074 ^ n2269 ;
  assign n7780 = n7779 ^ n7778 ^ n7777 ;
  assign n7781 = ( n1805 & n4574 ) | ( n1805 & ~n7780 ) | ( n4574 & ~n7780 ) ;
  assign n7782 = n2274 ^ n665 ^ 1'b0 ;
  assign n7783 = x66 & ~n7782 ;
  assign n7784 = n6184 ^ n5295 ^ 1'b0 ;
  assign n7785 = ~n1949 & n7784 ;
  assign n7786 = n7783 & n7785 ;
  assign n7787 = x31 & n4502 ;
  assign n7788 = ( ~n1050 & n1374 ) | ( ~n1050 & n2265 ) | ( n1374 & n2265 ) ;
  assign n7789 = n7787 & n7788 ;
  assign n7790 = n7789 ^ n1834 ^ 1'b0 ;
  assign n7795 = n5277 ^ n1188 ^ n551 ;
  assign n7791 = n1457 ^ n777 ^ n753 ;
  assign n7792 = ( ~n2727 & n5651 ) | ( ~n2727 & n7791 ) | ( n5651 & n7791 ) ;
  assign n7793 = ~n3087 & n7792 ;
  assign n7794 = n2032 & n7793 ;
  assign n7796 = n7795 ^ n7794 ^ n1540 ;
  assign n7803 = n1874 ^ n465 ^ x46 ;
  assign n7804 = n3072 | n5928 ;
  assign n7805 = n7803 & ~n7804 ;
  assign n7812 = n7133 ^ n5404 ^ n1900 ;
  assign n7813 = ( n3388 & n6498 ) | ( n3388 & n7812 ) | ( n6498 & n7812 ) ;
  assign n7814 = n7813 ^ n1139 ^ 1'b0 ;
  assign n7811 = n1000 & n2616 ;
  assign n7806 = ( ~n1052 & n3404 ) | ( ~n1052 & n4420 ) | ( n3404 & n4420 ) ;
  assign n7807 = n7806 ^ n746 ^ n531 ;
  assign n7808 = n6574 ^ n3481 ^ 1'b0 ;
  assign n7809 = n7807 & n7808 ;
  assign n7810 = ( n3017 & ~n3106 ) | ( n3017 & n7809 ) | ( ~n3106 & n7809 ) ;
  assign n7815 = n7814 ^ n7811 ^ n7810 ;
  assign n7816 = ( ~n7408 & n7805 ) | ( ~n7408 & n7815 ) | ( n7805 & n7815 ) ;
  assign n7797 = n2316 & ~n4510 ;
  assign n7798 = ~n5465 & n7797 ;
  assign n7799 = n1880 & ~n2013 ;
  assign n7800 = n212 & n7799 ;
  assign n7801 = ( n2036 & ~n7204 ) | ( n2036 & n7800 ) | ( ~n7204 & n7800 ) ;
  assign n7802 = ~n7798 & n7801 ;
  assign n7817 = n7816 ^ n7802 ^ 1'b0 ;
  assign n7818 = ( n740 & ~n1575 ) | ( n740 & n4941 ) | ( ~n1575 & n4941 ) ;
  assign n7819 = ( x114 & n5186 ) | ( x114 & n7818 ) | ( n5186 & n7818 ) ;
  assign n7820 = n7819 ^ n3110 ^ n1436 ;
  assign n7821 = ~n218 & n4164 ;
  assign n7822 = ( n1306 & ~n7498 ) | ( n1306 & n7821 ) | ( ~n7498 & n7821 ) ;
  assign n7823 = n7822 ^ n1003 ^ x22 ;
  assign n7824 = n2011 ^ n1351 ^ n1289 ;
  assign n7825 = n7289 ^ n2543 ^ n623 ;
  assign n7826 = n7825 ^ n4239 ^ x84 ;
  assign n7827 = ( n350 & ~n746 ) | ( n350 & n1993 ) | ( ~n746 & n1993 ) ;
  assign n7828 = n3283 & n4779 ;
  assign n7829 = ~n7827 & n7828 ;
  assign n7830 = n3761 | n7829 ;
  assign n7831 = n7826 & ~n7830 ;
  assign n7832 = ( n2502 & n7824 ) | ( n2502 & ~n7831 ) | ( n7824 & ~n7831 ) ;
  assign n7842 = n7791 ^ n1804 ^ 1'b0 ;
  assign n7841 = n7734 ^ n467 ^ 1'b0 ;
  assign n7833 = n1954 & ~n4183 ;
  assign n7834 = n230 & n7833 ;
  assign n7835 = n3573 & ~n7834 ;
  assign n7836 = n6796 & n7835 ;
  assign n7837 = ( ~n6135 & n6330 ) | ( ~n6135 & n7836 ) | ( n6330 & n7836 ) ;
  assign n7838 = n1955 ^ n322 ^ 1'b0 ;
  assign n7839 = ~n7837 & n7838 ;
  assign n7840 = n7839 ^ n1475 ^ n1466 ;
  assign n7843 = n7842 ^ n7841 ^ n7840 ;
  assign n7849 = n2730 ^ n2144 ^ 1'b0 ;
  assign n7848 = n2614 | n2781 ;
  assign n7844 = ( ~n703 & n2218 ) | ( ~n703 & n2275 ) | ( n2218 & n2275 ) ;
  assign n7845 = ( n395 & n2117 ) | ( n395 & n6337 ) | ( n2117 & n6337 ) ;
  assign n7846 = n6850 ^ n3904 ^ n3869 ;
  assign n7847 = ( n7844 & ~n7845 ) | ( n7844 & n7846 ) | ( ~n7845 & n7846 ) ;
  assign n7850 = n7849 ^ n7848 ^ n7847 ;
  assign n7856 = ~n2335 & n4952 ;
  assign n7857 = n7856 ^ n2934 ^ 1'b0 ;
  assign n7858 = n7857 ^ n1470 ^ x85 ;
  assign n7859 = n7858 ^ n5034 ^ n3318 ;
  assign n7851 = n2061 ^ n1994 ^ 1'b0 ;
  assign n7852 = n234 & ~n7851 ;
  assign n7853 = n7852 ^ n3122 ^ n521 ;
  assign n7854 = ( n3995 & ~n5650 ) | ( n3995 & n7853 ) | ( ~n5650 & n7853 ) ;
  assign n7855 = ( n2151 & ~n2745 ) | ( n2151 & n7854 ) | ( ~n2745 & n7854 ) ;
  assign n7860 = n7859 ^ n7855 ^ n4473 ;
  assign n7861 = ~n3014 & n3382 ;
  assign n7862 = n7861 ^ n6522 ^ 1'b0 ;
  assign n7863 = n1190 & n1632 ;
  assign n7864 = ~n2228 & n7863 ;
  assign n7865 = n7862 | n7864 ;
  assign n7866 = n1738 & n2832 ;
  assign n7867 = n7866 ^ n1824 ^ 1'b0 ;
  assign n7868 = n4031 ^ n410 ^ n334 ;
  assign n7869 = ( n1996 & n7867 ) | ( n1996 & ~n7868 ) | ( n7867 & ~n7868 ) ;
  assign n7870 = n3130 & ~n7869 ;
  assign n7871 = n2539 & ~n3054 ;
  assign n7876 = n4565 & ~n6133 ;
  assign n7877 = n7876 ^ n7582 ^ 1'b0 ;
  assign n7878 = n7877 ^ n5930 ^ n270 ;
  assign n7875 = ( n4562 & n5897 ) | ( n4562 & ~n7150 ) | ( n5897 & ~n7150 ) ;
  assign n7872 = n4987 ^ n2826 ^ n1981 ;
  assign n7873 = n6976 | n7872 ;
  assign n7874 = n6823 | n7873 ;
  assign n7879 = n7878 ^ n7875 ^ n7874 ;
  assign n7880 = n7189 ^ n7014 ^ n867 ;
  assign n7881 = ( n664 & n4961 ) | ( n664 & n7880 ) | ( n4961 & n7880 ) ;
  assign n7882 = n2154 ^ n1793 ^ 1'b0 ;
  assign n7883 = n7882 ^ n4574 ^ 1'b0 ;
  assign n7884 = ~n3887 & n7883 ;
  assign n7885 = n5040 ^ n3981 ^ n3736 ;
  assign n7886 = ( n1580 & ~n2682 ) | ( n1580 & n4231 ) | ( ~n2682 & n4231 ) ;
  assign n7887 = n7886 ^ n4593 ^ 1'b0 ;
  assign n7888 = n619 & ~n1116 ;
  assign n7889 = ( n3376 & n5193 ) | ( n3376 & ~n7888 ) | ( n5193 & ~n7888 ) ;
  assign n7890 = n1550 & n7889 ;
  assign n7891 = n1217 ^ n583 ^ n329 ;
  assign n7892 = n2333 | n7891 ;
  assign n7893 = n4923 ^ n3544 ^ 1'b0 ;
  assign n7894 = n7892 | n7893 ;
  assign n7895 = ~n407 & n3971 ;
  assign n7896 = ~n7894 & n7895 ;
  assign n7897 = n7890 & n7896 ;
  assign n7898 = n2289 & ~n7669 ;
  assign n7899 = x66 & n1637 ;
  assign n7900 = n7899 ^ x28 ^ 1'b0 ;
  assign n7901 = ( n463 & ~n5551 ) | ( n463 & n7900 ) | ( ~n5551 & n7900 ) ;
  assign n7902 = ( n1428 & ~n2625 ) | ( n1428 & n3584 ) | ( ~n2625 & n3584 ) ;
  assign n7903 = ( ~n3746 & n7347 ) | ( ~n3746 & n7902 ) | ( n7347 & n7902 ) ;
  assign n7904 = ~n6520 & n7903 ;
  assign n7905 = n7904 ^ n3779 ^ 1'b0 ;
  assign n7906 = n7905 ^ n1332 ^ 1'b0 ;
  assign n7907 = n1312 & n4628 ;
  assign n7908 = n7907 ^ n3404 ^ 1'b0 ;
  assign n7909 = ( n7901 & n7906 ) | ( n7901 & n7908 ) | ( n7906 & n7908 ) ;
  assign n7913 = ~n2028 & n3200 ;
  assign n7912 = n2548 & ~n3690 ;
  assign n7910 = n2157 ^ n663 ^ x19 ;
  assign n7911 = ( n3664 & n5976 ) | ( n3664 & n7910 ) | ( n5976 & n7910 ) ;
  assign n7914 = n7913 ^ n7912 ^ n7911 ;
  assign n7915 = n3845 | n7914 ;
  assign n7917 = ( x93 & n702 ) | ( x93 & n1618 ) | ( n702 & n1618 ) ;
  assign n7916 = ( n1379 & ~n1679 ) | ( n1379 & n3376 ) | ( ~n1679 & n3376 ) ;
  assign n7918 = n7917 ^ n7916 ^ n5887 ;
  assign n7919 = n2069 & n5864 ;
  assign n7920 = n4934 ^ n2948 ^ 1'b0 ;
  assign n7921 = n2889 ^ n648 ^ 1'b0 ;
  assign n7922 = n7920 | n7921 ;
  assign n7923 = n5297 & n7922 ;
  assign n7924 = ( x75 & n3424 ) | ( x75 & n7923 ) | ( n3424 & n7923 ) ;
  assign n7925 = ~n3302 & n3573 ;
  assign n7926 = ~n7888 & n7925 ;
  assign n7927 = ( n357 & n1542 ) | ( n357 & ~n1870 ) | ( n1542 & ~n1870 ) ;
  assign n7928 = ( ~n4611 & n7270 ) | ( ~n4611 & n7927 ) | ( n7270 & n7927 ) ;
  assign n7929 = n7928 ^ n6532 ^ 1'b0 ;
  assign n7930 = n7929 ^ n6273 ^ n1062 ;
  assign n7931 = ( n2884 & ~n3553 ) | ( n2884 & n7383 ) | ( ~n3553 & n7383 ) ;
  assign n7932 = n7394 ^ n5383 ^ n270 ;
  assign n7933 = n4012 ^ n509 ^ 1'b0 ;
  assign n7934 = n3248 & n7933 ;
  assign n7936 = ~n1625 & n5005 ;
  assign n7937 = n1269 & n7936 ;
  assign n7935 = ( n921 & ~n1632 ) | ( n921 & n4010 ) | ( ~n1632 & n4010 ) ;
  assign n7938 = n7937 ^ n7935 ^ n562 ;
  assign n7939 = n7934 | n7938 ;
  assign n7940 = ( ~n3064 & n3862 ) | ( ~n3064 & n5593 ) | ( n3862 & n5593 ) ;
  assign n7944 = ~n4567 & n5871 ;
  assign n7941 = n3384 ^ n2761 ^ n1949 ;
  assign n7942 = n3026 & ~n7710 ;
  assign n7943 = ~n7941 & n7942 ;
  assign n7945 = n7944 ^ n7943 ^ n1256 ;
  assign n7946 = ( n313 & ~n7940 ) | ( n313 & n7945 ) | ( ~n7940 & n7945 ) ;
  assign n7947 = ( n763 & ~n2503 ) | ( n763 & n5908 ) | ( ~n2503 & n5908 ) ;
  assign n7948 = n7947 ^ n5037 ^ n498 ;
  assign n7949 = n7948 ^ n6401 ^ n1942 ;
  assign n7955 = ~n1924 & n3773 ;
  assign n7954 = n4973 ^ n2393 ^ 1'b0 ;
  assign n7956 = n7955 ^ n7954 ^ n1478 ;
  assign n7950 = n6796 ^ n4292 ^ 1'b0 ;
  assign n7951 = ( n926 & n1479 ) | ( n926 & ~n3683 ) | ( n1479 & ~n3683 ) ;
  assign n7952 = n7951 ^ n2473 ^ 1'b0 ;
  assign n7953 = ( ~n1376 & n7950 ) | ( ~n1376 & n7952 ) | ( n7950 & n7952 ) ;
  assign n7957 = n7956 ^ n7953 ^ n7037 ;
  assign n7958 = n4342 ^ n2725 ^ 1'b0 ;
  assign n7959 = n3119 | n7958 ;
  assign n7960 = ( n3247 & n7957 ) | ( n3247 & n7959 ) | ( n7957 & n7959 ) ;
  assign n7961 = ~n990 & n2206 ;
  assign n7962 = n7961 ^ n3986 ^ n553 ;
  assign n7963 = n7962 ^ n1176 ^ n569 ;
  assign n7964 = n7963 ^ n1863 ^ 1'b0 ;
  assign n7965 = n3916 & ~n7964 ;
  assign n7966 = x95 & ~n1759 ;
  assign n7967 = n6740 ^ n1999 ^ 1'b0 ;
  assign n7968 = ~n1326 & n7967 ;
  assign n7969 = n3790 & n7968 ;
  assign n7970 = n7966 & n7969 ;
  assign n7971 = n4214 | n5438 ;
  assign n7972 = n7971 ^ x25 ^ 1'b0 ;
  assign n7973 = n7970 & n7972 ;
  assign n7974 = n1506 | n4894 ;
  assign n7975 = n7613 ^ n5836 ^ n644 ;
  assign n7976 = ~n2005 & n2983 ;
  assign n7977 = n5851 ^ n4767 ^ n1035 ;
  assign n7978 = ( n1780 & ~n5927 ) | ( n1780 & n7977 ) | ( ~n5927 & n7977 ) ;
  assign n7979 = ~n2425 & n6709 ;
  assign n7980 = n7979 ^ n741 ^ 1'b0 ;
  assign n7983 = n6043 ^ n2474 ^ n1420 ;
  assign n7984 = n7983 ^ n7901 ^ n969 ;
  assign n7981 = ( n2211 & ~n3700 ) | ( n2211 & n6664 ) | ( ~n3700 & n6664 ) ;
  assign n7982 = n7981 ^ n3441 ^ n2531 ;
  assign n7985 = n7984 ^ n7982 ^ n7495 ;
  assign n7986 = n6212 ^ n5987 ^ n1660 ;
  assign n7989 = n378 & ~n1377 ;
  assign n7990 = ~n3800 & n7989 ;
  assign n7987 = n1222 | n4117 ;
  assign n7988 = n7824 | n7987 ;
  assign n7991 = n7990 ^ n7988 ^ n3766 ;
  assign n7992 = ( n3868 & n7437 ) | ( n3868 & ~n7991 ) | ( n7437 & ~n7991 ) ;
  assign n7993 = n6462 ^ n3600 ^ 1'b0 ;
  assign n7994 = n7992 & n7993 ;
  assign n7995 = n1544 | n2301 ;
  assign n7996 = n666 | n7995 ;
  assign n7997 = n7996 ^ n2321 ^ 1'b0 ;
  assign n7998 = n7994 & n7997 ;
  assign n7999 = ( n6974 & ~n7986 ) | ( n6974 & n7998 ) | ( ~n7986 & n7998 ) ;
  assign n8000 = n1168 | n4587 ;
  assign n8001 = n3016 & ~n8000 ;
  assign n8002 = x101 & n177 ;
  assign n8003 = n8002 ^ n873 ^ n272 ;
  assign n8004 = n306 & n4371 ;
  assign n8005 = n3347 & n8004 ;
  assign n8006 = n6840 & ~n8005 ;
  assign n8007 = n1573 & n8006 ;
  assign n8008 = n8007 ^ n3673 ^ n3333 ;
  assign n8009 = n4934 & ~n6510 ;
  assign n8010 = ~n4636 & n8009 ;
  assign n8011 = n2664 & ~n8010 ;
  assign n8012 = n3951 ^ n3395 ^ n1453 ;
  assign n8013 = n8012 ^ n653 ^ 1'b0 ;
  assign n8014 = n8011 & ~n8013 ;
  assign n8015 = n7661 ^ n4170 ^ n514 ;
  assign n8016 = ( n1517 & ~n3710 ) | ( n1517 & n4319 ) | ( ~n3710 & n4319 ) ;
  assign n8017 = n8015 | n8016 ;
  assign n8018 = n8017 ^ n4702 ^ 1'b0 ;
  assign n8019 = n2258 & n8018 ;
  assign n8022 = n4590 & n5846 ;
  assign n8023 = ~n1521 & n8022 ;
  assign n8024 = n8023 ^ n2842 ^ n2676 ;
  assign n8021 = ( n545 & n2163 ) | ( n545 & n5279 ) | ( n2163 & n5279 ) ;
  assign n8020 = n801 | n1139 ;
  assign n8025 = n8024 ^ n8021 ^ n8020 ;
  assign n8026 = ( n4102 & n8019 ) | ( n4102 & n8025 ) | ( n8019 & n8025 ) ;
  assign n8027 = n7059 ^ n4292 ^ n4095 ;
  assign n8033 = ( n182 & ~n1699 ) | ( n182 & n2998 ) | ( ~n1699 & n2998 ) ;
  assign n8035 = ( n206 & ~n1659 ) | ( n206 & n2545 ) | ( ~n1659 & n2545 ) ;
  assign n8034 = n3144 & ~n7430 ;
  assign n8036 = n8035 ^ n8034 ^ 1'b0 ;
  assign n8037 = ~n6626 & n8036 ;
  assign n8038 = ( n3320 & n8033 ) | ( n3320 & n8037 ) | ( n8033 & n8037 ) ;
  assign n8028 = n2729 ^ n1877 ^ n631 ;
  assign n8029 = n3333 | n8028 ;
  assign n8030 = n8029 ^ n5833 ^ 1'b0 ;
  assign n8031 = n6047 & ~n8030 ;
  assign n8032 = n8031 ^ n496 ^ 1'b0 ;
  assign n8039 = n8038 ^ n8032 ^ 1'b0 ;
  assign n8040 = ( ~n200 & n2545 ) | ( ~n200 & n3061 ) | ( n2545 & n3061 ) ;
  assign n8041 = n8040 ^ n1680 ^ 1'b0 ;
  assign n8042 = n6651 ^ n6233 ^ 1'b0 ;
  assign n8043 = ( n229 & ~n5787 ) | ( n229 & n8042 ) | ( ~n5787 & n8042 ) ;
  assign n8044 = n651 & ~n1567 ;
  assign n8045 = n8044 ^ n4264 ^ 1'b0 ;
  assign n8046 = ( n1610 & ~n7205 ) | ( n1610 & n8045 ) | ( ~n7205 & n8045 ) ;
  assign n8047 = ( n2521 & n2621 ) | ( n2521 & ~n4420 ) | ( n2621 & ~n4420 ) ;
  assign n8048 = n8047 ^ n666 ^ 1'b0 ;
  assign n8049 = n7187 ^ n6524 ^ n261 ;
  assign n8050 = n1609 | n3849 ;
  assign n8051 = n8050 ^ n164 ^ 1'b0 ;
  assign n8052 = n8049 | n8051 ;
  assign n8053 = ( n7825 & n8048 ) | ( n7825 & n8052 ) | ( n8048 & n8052 ) ;
  assign n8054 = n1947 ^ n1487 ^ 1'b0 ;
  assign n8055 = n8054 ^ n4015 ^ n236 ;
  assign n8056 = n8055 ^ n2238 ^ n206 ;
  assign n8057 = ( ~n555 & n2683 ) | ( ~n555 & n2701 ) | ( n2683 & n2701 ) ;
  assign n8058 = ( n841 & n1221 ) | ( n841 & ~n8057 ) | ( n1221 & ~n8057 ) ;
  assign n8059 = n543 & n8058 ;
  assign n8060 = n7507 ^ n7434 ^ n5979 ;
  assign n8061 = n2896 & ~n7582 ;
  assign n8062 = n8061 ^ n7984 ^ 1'b0 ;
  assign n8063 = n8060 | n8062 ;
  assign n8064 = n433 & ~n5863 ;
  assign n8065 = n8064 ^ n6476 ^ 1'b0 ;
  assign n8066 = n5384 & n6295 ;
  assign n8067 = n8066 ^ n2071 ^ 1'b0 ;
  assign n8068 = ( n310 & n4774 ) | ( n310 & n8067 ) | ( n4774 & n8067 ) ;
  assign n8069 = n2733 & ~n8068 ;
  assign n8070 = n3448 ^ n2269 ^ 1'b0 ;
  assign n8071 = n6511 & n8070 ;
  assign n8072 = ( n3310 & n4473 ) | ( n3310 & n6173 ) | ( n4473 & n6173 ) ;
  assign n8075 = n5833 ^ n1716 ^ n964 ;
  assign n8073 = n907 ^ n773 ^ 1'b0 ;
  assign n8074 = ( n2377 & n3741 ) | ( n2377 & n8073 ) | ( n3741 & n8073 ) ;
  assign n8076 = n8075 ^ n8074 ^ n3878 ;
  assign n8077 = ( n3526 & ~n3786 ) | ( n3526 & n4825 ) | ( ~n3786 & n4825 ) ;
  assign n8078 = n5008 ^ n4459 ^ n3857 ;
  assign n8079 = n2644 | n8078 ;
  assign n8080 = n8077 & ~n8079 ;
  assign n8081 = n1099 & ~n6864 ;
  assign n8082 = n1932 & n4455 ;
  assign n8083 = n255 | n8082 ;
  assign n8084 = n8081 | n8083 ;
  assign n8085 = n1269 & ~n1451 ;
  assign n8086 = n8085 ^ n7323 ^ 1'b0 ;
  assign n8087 = ~n8084 & n8086 ;
  assign n8088 = ( n8076 & n8080 ) | ( n8076 & n8087 ) | ( n8080 & n8087 ) ;
  assign n8089 = ( n8071 & n8072 ) | ( n8071 & ~n8088 ) | ( n8072 & ~n8088 ) ;
  assign n8095 = n6413 ^ n4361 ^ 1'b0 ;
  assign n8096 = ( n3058 & ~n4401 ) | ( n3058 & n8095 ) | ( ~n4401 & n8095 ) ;
  assign n8091 = n7935 ^ x46 ^ 1'b0 ;
  assign n8092 = ~n3788 & n8091 ;
  assign n8090 = n2570 & n7944 ;
  assign n8093 = n8092 ^ n8090 ^ 1'b0 ;
  assign n8094 = n1956 & ~n8093 ;
  assign n8097 = n8096 ^ n8094 ^ 1'b0 ;
  assign n8098 = n8097 ^ n4689 ^ n1075 ;
  assign n8099 = n5163 & ~n5176 ;
  assign n8100 = n8099 ^ n4625 ^ 1'b0 ;
  assign n8101 = ( n670 & ~n2299 ) | ( n670 & n4830 ) | ( ~n2299 & n4830 ) ;
  assign n8102 = ( n2899 & n7376 ) | ( n2899 & n8101 ) | ( n7376 & n8101 ) ;
  assign n8103 = n8102 ^ n7269 ^ n1556 ;
  assign n8104 = n3876 ^ n2646 ^ n2367 ;
  assign n8105 = ( ~n184 & n627 ) | ( ~n184 & n5049 ) | ( n627 & n5049 ) ;
  assign n8106 = n4555 & n8105 ;
  assign n8107 = n8104 & n8106 ;
  assign n8108 = n4077 | n4400 ;
  assign n8109 = ~n1050 & n4934 ;
  assign n8110 = n8109 ^ n1479 ^ 1'b0 ;
  assign n8111 = ~n4153 & n8110 ;
  assign n8112 = n1763 & n8111 ;
  assign n8113 = ~n2656 & n8112 ;
  assign n8114 = n1560 & ~n1893 ;
  assign n8116 = n7169 ^ n6759 ^ n2759 ;
  assign n8115 = n2322 | n5915 ;
  assign n8117 = n8116 ^ n8115 ^ 1'b0 ;
  assign n8118 = ( n3361 & ~n6182 ) | ( n3361 & n6804 ) | ( ~n6182 & n6804 ) ;
  assign n8124 = ( n4696 & n5780 ) | ( n4696 & n7096 ) | ( n5780 & n7096 ) ;
  assign n8125 = n6637 & ~n8124 ;
  assign n8126 = ~n4565 & n8125 ;
  assign n8119 = n6261 ^ n3324 ^ 1'b0 ;
  assign n8120 = n2427 | n8119 ;
  assign n8121 = ( n2287 & n7134 ) | ( n2287 & n8120 ) | ( n7134 & n8120 ) ;
  assign n8122 = n2961 | n8121 ;
  assign n8123 = n2322 & ~n8122 ;
  assign n8127 = n8126 ^ n8123 ^ n1519 ;
  assign n8128 = n8127 ^ n3423 ^ x47 ;
  assign n8129 = n7065 ^ n5466 ^ n2151 ;
  assign n8130 = n6916 ^ n6697 ^ n4781 ;
  assign n8132 = n6002 ^ n3911 ^ n1447 ;
  assign n8133 = ( n761 & n1351 ) | ( n761 & ~n5753 ) | ( n1351 & ~n5753 ) ;
  assign n8134 = n8132 & n8133 ;
  assign n8135 = n3752 & n8134 ;
  assign n8131 = ( n320 & n2817 ) | ( n320 & ~n7077 ) | ( n2817 & ~n7077 ) ;
  assign n8136 = n8135 ^ n8131 ^ n6688 ;
  assign n8137 = ~n3083 & n7613 ;
  assign n8138 = n8137 ^ n3125 ^ 1'b0 ;
  assign n8144 = ~n926 & n1576 ;
  assign n8139 = n6231 ^ n5191 ^ n1534 ;
  assign n8140 = n5487 ^ n2788 ^ n1562 ;
  assign n8141 = n5778 ^ n1421 ^ 1'b0 ;
  assign n8142 = n8140 & n8141 ;
  assign n8143 = n8139 & ~n8142 ;
  assign n8145 = n8144 ^ n8143 ^ n1538 ;
  assign n8146 = n1556 | n3210 ;
  assign n8147 = n3463 & n4330 ;
  assign n8148 = ( n7689 & n8146 ) | ( n7689 & ~n8147 ) | ( n8146 & ~n8147 ) ;
  assign n8151 = n4064 | n4330 ;
  assign n8152 = n2038 | n8151 ;
  assign n8153 = n8152 ^ n3123 ^ 1'b0 ;
  assign n8154 = ( ~n553 & n651 ) | ( ~n553 & n8153 ) | ( n651 & n8153 ) ;
  assign n8149 = n6479 ^ n1449 ^ 1'b0 ;
  assign n8150 = ~n742 & n8149 ;
  assign n8155 = n8154 ^ n8150 ^ 1'b0 ;
  assign n8156 = ~n1775 & n4794 ;
  assign n8157 = ( n2804 & n4859 ) | ( n2804 & ~n8156 ) | ( n4859 & ~n8156 ) ;
  assign n8158 = n699 & n7006 ;
  assign n8159 = n6454 ^ n1630 ^ 1'b0 ;
  assign n8160 = n8159 ^ n2396 ^ 1'b0 ;
  assign n8166 = n2206 ^ n909 ^ n598 ;
  assign n8165 = ~n207 & n2612 ;
  assign n8167 = n8166 ^ n8165 ^ 1'b0 ;
  assign n8161 = n5033 ^ n3145 ^ n3131 ;
  assign n8162 = n6258 ^ n2975 ^ n1113 ;
  assign n8163 = n8161 | n8162 ;
  assign n8164 = n8163 ^ n175 ^ 1'b0 ;
  assign n8168 = n8167 ^ n8164 ^ n7938 ;
  assign n8169 = ( n860 & n8160 ) | ( n860 & n8168 ) | ( n8160 & n8168 ) ;
  assign n8170 = ( n239 & n1042 ) | ( n239 & n1248 ) | ( n1042 & n1248 ) ;
  assign n8171 = n2140 & ~n8170 ;
  assign n8172 = n5277 & n8171 ;
  assign n8173 = n2515 | n3081 ;
  assign n8174 = n8173 ^ n1668 ^ 1'b0 ;
  assign n8175 = ( n1956 & n2384 ) | ( n1956 & ~n8174 ) | ( n2384 & ~n8174 ) ;
  assign n8176 = ~n998 & n2071 ;
  assign n8177 = ~n2167 & n8176 ;
  assign n8178 = n8177 ^ n1725 ^ 1'b0 ;
  assign n8179 = ( n2039 & n4010 ) | ( n2039 & n8178 ) | ( n4010 & n8178 ) ;
  assign n8180 = ( ~n3165 & n4980 ) | ( ~n3165 & n7880 ) | ( n4980 & n7880 ) ;
  assign n8182 = n3864 ^ n2366 ^ 1'b0 ;
  assign n8181 = ( n1525 & n3516 ) | ( n1525 & n3699 ) | ( n3516 & n3699 ) ;
  assign n8183 = n8182 ^ n8181 ^ n8071 ;
  assign n8184 = n8183 ^ n3640 ^ 1'b0 ;
  assign n8185 = n2520 & n8184 ;
  assign n8186 = n1992 & n7122 ;
  assign n8187 = ~n7365 & n8186 ;
  assign n8188 = n253 | n8187 ;
  assign n8189 = n8188 ^ n4886 ^ 1'b0 ;
  assign n8190 = n686 | n2329 ;
  assign n8191 = n8190 ^ n1442 ^ 1'b0 ;
  assign n8192 = n8191 ^ n3710 ^ n266 ;
  assign n8193 = ( n3524 & ~n6558 ) | ( n3524 & n8192 ) | ( ~n6558 & n8192 ) ;
  assign n8194 = ( n829 & ~n1114 ) | ( n829 & n6766 ) | ( ~n1114 & n6766 ) ;
  assign n8195 = n2918 ^ n1203 ^ n156 ;
  assign n8196 = n2359 & n8195 ;
  assign n8197 = n8196 ^ n5761 ^ 1'b0 ;
  assign n8198 = n8197 ^ n2990 ^ n918 ;
  assign n8199 = n8198 ^ n2061 ^ n1130 ;
  assign n8200 = ( n6732 & n8194 ) | ( n6732 & ~n8199 ) | ( n8194 & ~n8199 ) ;
  assign n8201 = n3075 & ~n6661 ;
  assign n8202 = ( n8193 & ~n8200 ) | ( n8193 & n8201 ) | ( ~n8200 & n8201 ) ;
  assign n8205 = n7882 ^ n3179 ^ n3026 ;
  assign n8206 = ~n1608 & n8205 ;
  assign n8210 = ~n2712 & n6664 ;
  assign n8207 = ( n1781 & n3165 ) | ( n1781 & ~n6001 ) | ( n3165 & ~n6001 ) ;
  assign n8208 = ( ~n1640 & n5056 ) | ( ~n1640 & n8207 ) | ( n5056 & n8207 ) ;
  assign n8209 = ~n3726 & n8208 ;
  assign n8211 = n8210 ^ n8209 ^ 1'b0 ;
  assign n8212 = n8211 ^ n3751 ^ 1'b0 ;
  assign n8213 = n8206 & ~n8212 ;
  assign n8203 = n4494 & n7352 ;
  assign n8204 = ~n7461 & n8203 ;
  assign n8214 = n8213 ^ n8204 ^ 1'b0 ;
  assign n8215 = n8214 ^ n2997 ^ n814 ;
  assign n8216 = n8215 ^ n5435 ^ 1'b0 ;
  assign n8217 = ( n984 & n2052 ) | ( n984 & ~n7600 ) | ( n2052 & ~n7600 ) ;
  assign n8218 = n6510 ^ n3358 ^ 1'b0 ;
  assign n8219 = n7739 ^ n2280 ^ 1'b0 ;
  assign n8220 = ~n8218 & n8219 ;
  assign n8221 = n2195 ^ n586 ^ x47 ;
  assign n8222 = n1038 ^ n695 ^ n350 ;
  assign n8223 = n8222 ^ n4862 ^ 1'b0 ;
  assign n8224 = ( n1967 & n8221 ) | ( n1967 & ~n8223 ) | ( n8221 & ~n8223 ) ;
  assign n8225 = n7280 ^ n3073 ^ 1'b0 ;
  assign n8226 = n585 & n8225 ;
  assign n8227 = ( n1226 & ~n3284 ) | ( n1226 & n8226 ) | ( ~n3284 & n8226 ) ;
  assign n8232 = ~n2828 & n3056 ;
  assign n8233 = n3736 & n8232 ;
  assign n8234 = n838 & ~n1489 ;
  assign n8235 = ( n3354 & n8233 ) | ( n3354 & ~n8234 ) | ( n8233 & ~n8234 ) ;
  assign n8230 = n1686 | n2386 ;
  assign n8228 = n1343 & ~n2521 ;
  assign n8229 = n8228 ^ n2072 ^ 1'b0 ;
  assign n8231 = n8230 ^ n8229 ^ n1628 ;
  assign n8236 = n8235 ^ n8231 ^ n8208 ;
  assign n8237 = n8236 ^ n6840 ^ 1'b0 ;
  assign n8238 = n2017 | n8237 ;
  assign n8239 = x36 & ~n275 ;
  assign n8240 = ~n4467 & n8239 ;
  assign n8241 = n214 | n673 ;
  assign n8242 = ( ~n770 & n4114 ) | ( ~n770 & n8116 ) | ( n4114 & n8116 ) ;
  assign n8243 = ( n588 & n3918 ) | ( n588 & n8242 ) | ( n3918 & n8242 ) ;
  assign n8244 = ( n8240 & n8241 ) | ( n8240 & ~n8243 ) | ( n8241 & ~n8243 ) ;
  assign n8245 = n2592 | n3187 ;
  assign n8246 = n5471 | n8245 ;
  assign n8247 = n8246 ^ n2454 ^ 1'b0 ;
  assign n8248 = n8244 & n8247 ;
  assign n8251 = n2707 ^ n2202 ^ n1205 ;
  assign n8252 = ( n4580 & ~n6770 ) | ( n4580 & n8251 ) | ( ~n6770 & n8251 ) ;
  assign n8249 = n4385 ^ n2926 ^ n2485 ;
  assign n8250 = ~n1002 & n8249 ;
  assign n8253 = n8252 ^ n8250 ^ 1'b0 ;
  assign n8254 = n8253 ^ n7896 ^ n2997 ;
  assign n8255 = ( ~n811 & n2375 ) | ( ~n811 & n6575 ) | ( n2375 & n6575 ) ;
  assign n8256 = n5341 ^ n816 ^ 1'b0 ;
  assign n8257 = ( n2020 & n3461 ) | ( n2020 & ~n8256 ) | ( n3461 & ~n8256 ) ;
  assign n8258 = n8257 ^ n2280 ^ n1269 ;
  assign n8259 = n8258 ^ n2086 ^ 1'b0 ;
  assign n8260 = ~n1110 & n8259 ;
  assign n8261 = n1677 & ~n8260 ;
  assign n8262 = ( n3226 & n8255 ) | ( n3226 & n8261 ) | ( n8255 & n8261 ) ;
  assign n8263 = n6843 ^ n6669 ^ 1'b0 ;
  assign n8264 = n4453 ^ n1868 ^ 1'b0 ;
  assign n8265 = n8263 & n8264 ;
  assign n8266 = n3395 ^ n1522 ^ 1'b0 ;
  assign n8270 = ( n1239 & ~n1882 ) | ( n1239 & n2368 ) | ( ~n1882 & n2368 ) ;
  assign n8271 = n8270 ^ n7350 ^ 1'b0 ;
  assign n8272 = ~n697 & n8271 ;
  assign n8267 = ~n5315 & n6576 ;
  assign n8268 = ~n2253 & n8267 ;
  assign n8269 = n2701 | n8268 ;
  assign n8273 = n8272 ^ n8269 ^ 1'b0 ;
  assign n8274 = ( n2464 & ~n8266 ) | ( n2464 & n8273 ) | ( ~n8266 & n8273 ) ;
  assign n8275 = n6636 ^ n3032 ^ 1'b0 ;
  assign n8276 = ~n1062 & n8057 ;
  assign n8277 = ( ~n1007 & n1113 ) | ( ~n1007 & n5068 ) | ( n1113 & n5068 ) ;
  assign n8278 = n8277 ^ n6669 ^ n324 ;
  assign n8279 = ( n2524 & ~n3937 ) | ( n2524 & n8278 ) | ( ~n3937 & n8278 ) ;
  assign n8280 = n4112 & ~n6720 ;
  assign n8281 = ( ~n1042 & n1266 ) | ( ~n1042 & n3651 ) | ( n1266 & n3651 ) ;
  assign n8282 = ( ~n2712 & n8280 ) | ( ~n2712 & n8281 ) | ( n8280 & n8281 ) ;
  assign n8283 = n4442 ^ n2566 ^ 1'b0 ;
  assign n8284 = n8283 ^ n6662 ^ 1'b0 ;
  assign n8285 = ( n8101 & n8282 ) | ( n8101 & ~n8284 ) | ( n8282 & ~n8284 ) ;
  assign n8286 = n6872 ^ n139 ^ 1'b0 ;
  assign n8287 = ( n5735 & n7431 ) | ( n5735 & n8286 ) | ( n7431 & n8286 ) ;
  assign n8292 = ( ~n506 & n1247 ) | ( ~n506 & n3675 ) | ( n1247 & n3675 ) ;
  assign n8288 = n1388 | n2678 ;
  assign n8289 = n508 & ~n8288 ;
  assign n8290 = n8289 ^ n7294 ^ n1500 ;
  assign n8291 = n8290 ^ n2178 ^ 1'b0 ;
  assign n8293 = n8292 ^ n8291 ^ n2790 ;
  assign n8294 = n2796 ^ n1315 ^ 1'b0 ;
  assign n8295 = n3584 & n8294 ;
  assign n8296 = n4135 & n8295 ;
  assign n8297 = n1608 & n8296 ;
  assign n8298 = ( n2393 & n3568 ) | ( n2393 & ~n5245 ) | ( n3568 & ~n5245 ) ;
  assign n8299 = n680 ^ n397 ^ 1'b0 ;
  assign n8300 = ( n2554 & ~n6288 ) | ( n2554 & n8299 ) | ( ~n6288 & n8299 ) ;
  assign n8301 = n8300 ^ n7583 ^ 1'b0 ;
  assign n8302 = n8298 | n8301 ;
  assign n8303 = ( n3580 & ~n3672 ) | ( n3580 & n8302 ) | ( ~n3672 & n8302 ) ;
  assign n8304 = n8303 ^ n6921 ^ n2568 ;
  assign n8305 = n4049 ^ n3833 ^ n1767 ;
  assign n8306 = n8305 ^ n4721 ^ n1686 ;
  assign n8318 = ( ~x33 & n1377 ) | ( ~x33 & n3617 ) | ( n1377 & n3617 ) ;
  assign n8319 = ( n2058 & n3379 ) | ( n2058 & n8318 ) | ( n3379 & n8318 ) ;
  assign n8316 = n5737 ^ n977 ^ n555 ;
  assign n8314 = n3069 ^ n2128 ^ n424 ;
  assign n8315 = n8314 ^ n3712 ^ n2092 ;
  assign n8311 = x65 & ~n1578 ;
  assign n8312 = ~n2506 & n8311 ;
  assign n8310 = n2844 & ~n6102 ;
  assign n8313 = n8312 ^ n8310 ^ 1'b0 ;
  assign n8317 = n8316 ^ n8315 ^ n8313 ;
  assign n8307 = n4006 ^ n1967 ^ n1252 ;
  assign n8308 = n1840 | n8307 ;
  assign n8309 = n8308 ^ n7583 ^ n6721 ;
  assign n8320 = n8319 ^ n8317 ^ n8309 ;
  assign n8321 = ( n1127 & ~n1260 ) | ( n1127 & n5537 ) | ( ~n1260 & n5537 ) ;
  assign n8322 = ( ~n1373 & n2646 ) | ( ~n1373 & n3229 ) | ( n2646 & n3229 ) ;
  assign n8323 = n8322 ^ n2801 ^ n2520 ;
  assign n8324 = n4961 ^ n4247 ^ n2727 ;
  assign n8325 = n8324 ^ n6885 ^ 1'b0 ;
  assign n8326 = n8323 & n8325 ;
  assign n8327 = n4373 ^ n3835 ^ x62 ;
  assign n8328 = ( n3626 & ~n4363 ) | ( n3626 & n5436 ) | ( ~n4363 & n5436 ) ;
  assign n8329 = n1362 & ~n6558 ;
  assign n8330 = ~n3324 & n8329 ;
  assign n8331 = n1538 & ~n4946 ;
  assign n8332 = n8330 & n8331 ;
  assign n8333 = n3044 ^ n1321 ^ x25 ;
  assign n8334 = n8333 ^ n7121 ^ n2132 ;
  assign n8335 = n5032 | n8221 ;
  assign n8336 = n8335 ^ n4784 ^ 1'b0 ;
  assign n8337 = ( n354 & ~n1450 ) | ( n354 & n8336 ) | ( ~n1450 & n8336 ) ;
  assign n8347 = n6807 ^ n1776 ^ 1'b0 ;
  assign n8340 = n4996 ^ n3261 ^ n1359 ;
  assign n8341 = n8340 ^ n1992 ^ n855 ;
  assign n8342 = ( n1601 & ~n4577 ) | ( n1601 & n8341 ) | ( ~n4577 & n8341 ) ;
  assign n8343 = ( n6271 & ~n6440 ) | ( n6271 & n8342 ) | ( ~n6440 & n8342 ) ;
  assign n8344 = n8343 ^ n2029 ^ x46 ;
  assign n8338 = n555 | n3897 ;
  assign n8339 = n8338 ^ n7224 ^ x101 ;
  assign n8345 = n8344 ^ n8339 ^ n5963 ;
  assign n8346 = n8345 ^ n1315 ^ 1'b0 ;
  assign n8348 = n8347 ^ n8346 ^ 1'b0 ;
  assign n8349 = n8337 & ~n8348 ;
  assign n8350 = n6494 ^ n5526 ^ n1220 ;
  assign n8351 = n8350 ^ n1172 ^ n663 ;
  assign n8352 = n2018 ^ n1261 ^ 1'b0 ;
  assign n8353 = n4782 | n8352 ;
  assign n8354 = n2116 | n8353 ;
  assign n8355 = n5183 & n8354 ;
  assign n8356 = n5711 | n8355 ;
  assign n8357 = n6900 ^ n4652 ^ n1703 ;
  assign n8358 = ( n1862 & n3834 ) | ( n1862 & ~n7749 ) | ( n3834 & ~n7749 ) ;
  assign n8359 = ( n2281 & n6534 ) | ( n2281 & n8358 ) | ( n6534 & n8358 ) ;
  assign n8360 = n5321 & ~n8359 ;
  assign n8361 = n5766 & n8360 ;
  assign n8363 = ( ~n1738 & n2514 ) | ( ~n1738 & n6158 ) | ( n2514 & n6158 ) ;
  assign n8362 = n5669 ^ n1179 ^ n315 ;
  assign n8364 = n8363 ^ n8362 ^ 1'b0 ;
  assign n8365 = n400 | n3415 ;
  assign n8366 = n4901 & ~n8365 ;
  assign n8367 = n3817 & ~n8345 ;
  assign n8368 = ~n8366 & n8367 ;
  assign n8369 = ( ~n1685 & n3894 ) | ( ~n1685 & n5121 ) | ( n3894 & n5121 ) ;
  assign n8370 = n8369 ^ n6525 ^ n6164 ;
  assign n8371 = ( n324 & ~n535 ) | ( n324 & n8365 ) | ( ~n535 & n8365 ) ;
  assign n8372 = ( n2142 & ~n4495 ) | ( n2142 & n8371 ) | ( ~n4495 & n8371 ) ;
  assign n8373 = ( n2654 & ~n6694 ) | ( n2654 & n8372 ) | ( ~n6694 & n8372 ) ;
  assign n8375 = n5484 ^ n991 ^ n608 ;
  assign n8374 = n3164 ^ n2125 ^ n1775 ;
  assign n8376 = n8375 ^ n8374 ^ n6240 ;
  assign n8377 = n8376 ^ n2869 ^ n1506 ;
  assign n8378 = n3217 ^ n1958 ^ 1'b0 ;
  assign n8379 = n1763 ^ n541 ^ 1'b0 ;
  assign n8380 = n7706 & n8379 ;
  assign n8381 = n4534 ^ n1340 ^ n1015 ;
  assign n8382 = n8381 ^ n1184 ^ n917 ;
  assign n8384 = ( ~n711 & n1751 ) | ( ~n711 & n2994 ) | ( n1751 & n2994 ) ;
  assign n8383 = n6198 ^ n529 ^ 1'b0 ;
  assign n8385 = n8384 ^ n8383 ^ n1066 ;
  assign n8386 = ~n3360 & n3522 ;
  assign n8387 = n8386 ^ n2999 ^ 1'b0 ;
  assign n8388 = n8387 ^ n2863 ^ 1'b0 ;
  assign n8389 = ( ~n8382 & n8385 ) | ( ~n8382 & n8388 ) | ( n8385 & n8388 ) ;
  assign n8390 = n1386 ^ n1180 ^ 1'b0 ;
  assign n8391 = ( n2244 & n3849 ) | ( n2244 & n5919 ) | ( n3849 & n5919 ) ;
  assign n8392 = n8391 ^ n5800 ^ 1'b0 ;
  assign n8393 = n8390 & n8392 ;
  assign n8394 = n3017 ^ n2780 ^ n1177 ;
  assign n8395 = n8394 ^ n5374 ^ n2733 ;
  assign n8396 = ( n1084 & n8393 ) | ( n1084 & n8395 ) | ( n8393 & n8395 ) ;
  assign n8402 = n8132 ^ n5916 ^ 1'b0 ;
  assign n8399 = n7749 ^ n945 ^ n653 ;
  assign n8400 = n8399 ^ n7429 ^ n2053 ;
  assign n8397 = n1843 | n8082 ;
  assign n8398 = n3488 & ~n8397 ;
  assign n8401 = n8400 ^ n8398 ^ n1440 ;
  assign n8403 = n8402 ^ n8401 ^ n3037 ;
  assign n8404 = n6199 ^ n1571 ^ 1'b0 ;
  assign n8405 = n1745 | n8404 ;
  assign n8406 = n6302 ^ n864 ^ 1'b0 ;
  assign n8414 = ( ~n757 & n1778 ) | ( ~n757 & n2195 ) | ( n1778 & n2195 ) ;
  assign n8412 = n3365 ^ n1379 ^ n1201 ;
  assign n8409 = ( n1715 & n2741 ) | ( n1715 & ~n2828 ) | ( n2741 & ~n2828 ) ;
  assign n8407 = n5787 ^ n1606 ^ 1'b0 ;
  assign n8408 = n4157 | n8407 ;
  assign n8410 = n8409 ^ n8408 ^ 1'b0 ;
  assign n8411 = n3619 & ~n8410 ;
  assign n8413 = n8412 ^ n8411 ^ 1'b0 ;
  assign n8415 = n8414 ^ n8413 ^ n4867 ;
  assign n8416 = n3358 & ~n6389 ;
  assign n8417 = n8416 ^ n6801 ^ n856 ;
  assign n8418 = ( n507 & ~n828 ) | ( n507 & n4499 ) | ( ~n828 & n4499 ) ;
  assign n8419 = ( n1125 & ~n5612 ) | ( n1125 & n5908 ) | ( ~n5612 & n5908 ) ;
  assign n8421 = n2713 ^ n1860 ^ 1'b0 ;
  assign n8422 = n8421 ^ n5525 ^ 1'b0 ;
  assign n8420 = x83 & ~n1348 ;
  assign n8423 = n8422 ^ n8420 ^ 1'b0 ;
  assign n8424 = n3470 & ~n8423 ;
  assign n8433 = n1095 ^ n785 ^ n549 ;
  assign n8431 = n2153 & n2778 ;
  assign n8432 = ( ~n4868 & n6914 ) | ( ~n4868 & n8431 ) | ( n6914 & n8431 ) ;
  assign n8434 = n8433 ^ n8432 ^ 1'b0 ;
  assign n8430 = n425 & n4589 ;
  assign n8426 = n8174 ^ n1783 ^ n581 ;
  assign n8425 = ( n5168 & n6452 ) | ( n5168 & ~n7854 ) | ( n6452 & ~n7854 ) ;
  assign n8427 = n8426 ^ n8425 ^ 1'b0 ;
  assign n8428 = n726 & ~n8427 ;
  assign n8429 = ~n7321 & n8428 ;
  assign n8435 = n8434 ^ n8430 ^ n8429 ;
  assign n8436 = n3229 | n8283 ;
  assign n8437 = n8436 ^ n7043 ^ 1'b0 ;
  assign n8438 = ~n1051 & n1291 ;
  assign n8439 = n8438 ^ n2303 ^ 1'b0 ;
  assign n8440 = ( n957 & ~n7407 ) | ( n957 & n8439 ) | ( ~n7407 & n8439 ) ;
  assign n8441 = n8440 ^ n7184 ^ 1'b0 ;
  assign n8442 = n8437 & n8441 ;
  assign n8444 = ( x95 & n3108 ) | ( x95 & ~n3249 ) | ( n3108 & ~n3249 ) ;
  assign n8443 = n971 & n1426 ;
  assign n8445 = n8444 ^ n8443 ^ 1'b0 ;
  assign n8446 = n8445 ^ n6766 ^ n5367 ;
  assign n8447 = n1895 | n8446 ;
  assign n8448 = n1282 & ~n8447 ;
  assign n8449 = n6586 ^ n4667 ^ 1'b0 ;
  assign n8450 = n8449 ^ n6678 ^ n5650 ;
  assign n8451 = ( n8442 & ~n8448 ) | ( n8442 & n8450 ) | ( ~n8448 & n8450 ) ;
  assign n8452 = ( ~n775 & n3853 ) | ( ~n775 & n5880 ) | ( n3853 & n5880 ) ;
  assign n8453 = n5929 ^ n3309 ^ n1097 ;
  assign n8454 = ( n1698 & n2308 ) | ( n1698 & n8453 ) | ( n2308 & n8453 ) ;
  assign n8455 = ~n5443 & n8454 ;
  assign n8456 = n8455 ^ n7343 ^ 1'b0 ;
  assign n8457 = n8456 ^ n6537 ^ n5180 ;
  assign n8458 = n2914 ^ n1754 ^ 1'b0 ;
  assign n8459 = ~n3284 & n8458 ;
  assign n8460 = ~n2478 & n7149 ;
  assign n8461 = n3814 ^ n2448 ^ 1'b0 ;
  assign n8462 = n8461 ^ n4228 ^ n3666 ;
  assign n8463 = ( n1350 & n4107 ) | ( n1350 & ~n8462 ) | ( n4107 & ~n8462 ) ;
  assign n8464 = ( n4925 & n7571 ) | ( n4925 & n8463 ) | ( n7571 & n8463 ) ;
  assign n8466 = n2751 ^ n2672 ^ n754 ;
  assign n8465 = n614 & ~n3735 ;
  assign n8467 = n8466 ^ n8465 ^ 1'b0 ;
  assign n8471 = n3616 ^ n1957 ^ n1684 ;
  assign n8472 = n7209 & n8471 ;
  assign n8473 = n2372 & n8472 ;
  assign n8469 = n1092 | n1188 ;
  assign n8468 = n3842 ^ n3336 ^ n861 ;
  assign n8470 = n8469 ^ n8468 ^ 1'b0 ;
  assign n8474 = n8473 ^ n8470 ^ n6585 ;
  assign n8475 = n2340 ^ n1637 ^ n855 ;
  assign n8476 = ~n7717 & n8475 ;
  assign n8477 = n4040 & n8476 ;
  assign n8478 = n3432 ^ n2857 ^ 1'b0 ;
  assign n8479 = n8478 ^ n6021 ^ 1'b0 ;
  assign n8480 = n1207 | n7690 ;
  assign n8481 = n8480 ^ n2262 ^ 1'b0 ;
  assign n8482 = x69 & n8481 ;
  assign n8483 = n8482 ^ n6464 ^ n1061 ;
  assign n8484 = n7312 ^ n3291 ^ 1'b0 ;
  assign n8485 = n8483 & ~n8484 ;
  assign n8486 = n8485 ^ n1447 ^ 1'b0 ;
  assign n8487 = n3027 ^ n2976 ^ n1624 ;
  assign n8488 = n8487 ^ n5240 ^ n1680 ;
  assign n8489 = n8488 ^ n6655 ^ n1648 ;
  assign n8494 = n3358 ^ n2860 ^ n2784 ;
  assign n8495 = n8494 ^ n1609 ^ n549 ;
  assign n8496 = n1745 | n8495 ;
  assign n8497 = ( n2129 & n5632 ) | ( n2129 & n8496 ) | ( n5632 & n8496 ) ;
  assign n8498 = n8497 ^ n5022 ^ n4420 ;
  assign n8490 = n6290 ^ n2209 ^ n844 ;
  assign n8491 = ~n4039 & n8490 ;
  assign n8492 = ~n6897 & n8491 ;
  assign n8493 = n8492 ^ n5316 ^ 1'b0 ;
  assign n8499 = n8498 ^ n8493 ^ 1'b0 ;
  assign n8500 = n4874 ^ n1647 ^ n912 ;
  assign n8501 = n8500 ^ n7031 ^ 1'b0 ;
  assign n8502 = n4217 & ~n8501 ;
  assign n8503 = n4164 ^ n3029 ^ n2733 ;
  assign n8504 = n352 | n8503 ;
  assign n8505 = n8504 ^ n4825 ^ 1'b0 ;
  assign n8506 = n3022 ^ n701 ^ 1'b0 ;
  assign n8507 = ~n7834 & n8506 ;
  assign n8508 = ~n3183 & n8507 ;
  assign n8509 = n180 & n8508 ;
  assign n8510 = n8509 ^ n5855 ^ n1215 ;
  assign n8511 = n6422 ^ n4602 ^ n1090 ;
  assign n8512 = n2375 & n6052 ;
  assign n8513 = n8512 ^ n2542 ^ 1'b0 ;
  assign n8514 = ( n2384 & ~n2622 ) | ( n2384 & n8513 ) | ( ~n2622 & n8513 ) ;
  assign n8515 = ( n4134 & ~n8511 ) | ( n4134 & n8514 ) | ( ~n8511 & n8514 ) ;
  assign n8516 = n1633 & ~n5264 ;
  assign n8517 = n4231 & n8516 ;
  assign n8518 = n4527 & n8517 ;
  assign n8522 = ( n394 & n2376 ) | ( n394 & ~n3997 ) | ( n2376 & ~n3997 ) ;
  assign n8519 = ( n1633 & ~n2129 ) | ( n1633 & n4188 ) | ( ~n2129 & n4188 ) ;
  assign n8520 = x44 & ~n8519 ;
  assign n8521 = n8520 ^ n596 ^ 1'b0 ;
  assign n8523 = n8522 ^ n8521 ^ n8186 ;
  assign n8524 = n497 & ~n3072 ;
  assign n8525 = n3855 & n8524 ;
  assign n8526 = n810 | n4939 ;
  assign n8527 = n8152 ^ n2103 ^ 1'b0 ;
  assign n8528 = n8527 ^ n1257 ^ 1'b0 ;
  assign n8529 = n5910 ^ n704 ^ x24 ;
  assign n8530 = n6851 & ~n8529 ;
  assign n8531 = n380 & n8002 ;
  assign n8532 = n8235 ^ n5100 ^ 1'b0 ;
  assign n8533 = n3919 ^ n3522 ^ n916 ;
  assign n8534 = ( ~n2212 & n8532 ) | ( ~n2212 & n8533 ) | ( n8532 & n8533 ) ;
  assign n8535 = ( n4056 & n8531 ) | ( n4056 & n8534 ) | ( n8531 & n8534 ) ;
  assign n8536 = n2842 & ~n8535 ;
  assign n8537 = ~n8530 & n8536 ;
  assign n8541 = n2504 ^ n2194 ^ n1958 ;
  assign n8542 = n7383 ^ n2276 ^ 1'b0 ;
  assign n8543 = n2360 | n8542 ;
  assign n8544 = ( n7168 & ~n8541 ) | ( n7168 & n8543 ) | ( ~n8541 & n8543 ) ;
  assign n8538 = n1069 & n2697 ;
  assign n8539 = n8538 ^ n875 ^ 1'b0 ;
  assign n8540 = ( n5424 & n5537 ) | ( n5424 & ~n8539 ) | ( n5537 & ~n8539 ) ;
  assign n8545 = n8544 ^ n8540 ^ n8486 ;
  assign n8546 = ( n357 & ~n1377 ) | ( n357 & n6280 ) | ( ~n1377 & n6280 ) ;
  assign n8547 = n8546 ^ n3265 ^ n1269 ;
  assign n8548 = n8547 ^ n7902 ^ n738 ;
  assign n8549 = ~n4895 & n8230 ;
  assign n8550 = n1114 & n8549 ;
  assign n8551 = n766 | n8299 ;
  assign n8552 = n3848 | n8551 ;
  assign n8553 = n8552 ^ n245 ^ 1'b0 ;
  assign n8556 = n313 & ~n3929 ;
  assign n8554 = n4489 & n7323 ;
  assign n8555 = n5303 & n8554 ;
  assign n8557 = n8556 ^ n8555 ^ n2588 ;
  assign n8558 = n2519 ^ n2460 ^ 1'b0 ;
  assign n8559 = n1476 & ~n8558 ;
  assign n8561 = n5051 ^ n2640 ^ n844 ;
  assign n8560 = n7857 ^ n6446 ^ n1372 ;
  assign n8562 = n8561 ^ n8560 ^ 1'b0 ;
  assign n8563 = n8559 & n8562 ;
  assign n8564 = n1657 & ~n4153 ;
  assign n8565 = n8564 ^ n699 ^ 1'b0 ;
  assign n8566 = n1687 ^ n445 ^ 1'b0 ;
  assign n8567 = ( n2170 & n8565 ) | ( n2170 & ~n8566 ) | ( n8565 & ~n8566 ) ;
  assign n8568 = n6321 & ~n8567 ;
  assign n8569 = n6414 & n8568 ;
  assign n8570 = n3422 & ~n4606 ;
  assign n8571 = n8570 ^ n5910 ^ n4891 ;
  assign n8572 = n8449 ^ n2406 ^ 1'b0 ;
  assign n8573 = n8571 & n8572 ;
  assign n8574 = n8573 ^ n3935 ^ 1'b0 ;
  assign n8575 = n4768 & ~n5156 ;
  assign n8576 = n8575 ^ n6777 ^ 1'b0 ;
  assign n8577 = ( n1228 & ~n6790 ) | ( n1228 & n8576 ) | ( ~n6790 & n8576 ) ;
  assign n8578 = ( n8569 & ~n8574 ) | ( n8569 & n8577 ) | ( ~n8574 & n8577 ) ;
  assign n8579 = n5490 ^ n514 ^ 1'b0 ;
  assign n8580 = n6337 ^ n3679 ^ 1'b0 ;
  assign n8581 = n2779 & n8580 ;
  assign n8582 = ~n8579 & n8581 ;
  assign n8583 = ( n331 & n2029 ) | ( n331 & ~n7339 ) | ( n2029 & ~n7339 ) ;
  assign n8584 = ( ~n2026 & n3009 ) | ( ~n2026 & n4170 ) | ( n3009 & n4170 ) ;
  assign n8585 = ~n7901 & n8584 ;
  assign n8586 = ~n947 & n8585 ;
  assign n8587 = ~n8583 & n8586 ;
  assign n8589 = ( n170 & n1333 ) | ( n170 & ~n2325 ) | ( n1333 & ~n2325 ) ;
  assign n8590 = ( n2421 & n4934 ) | ( n2421 & n8589 ) | ( n4934 & n8589 ) ;
  assign n8591 = ( n3506 & ~n4677 ) | ( n3506 & n8590 ) | ( ~n4677 & n8590 ) ;
  assign n8596 = n8591 ^ n3125 ^ 1'b0 ;
  assign n8597 = ~n5899 & n8596 ;
  assign n8588 = n5178 ^ n4488 ^ n1299 ;
  assign n8592 = ( ~n816 & n3889 ) | ( ~n816 & n8591 ) | ( n3889 & n8591 ) ;
  assign n8593 = ~n1619 & n8592 ;
  assign n8594 = n8593 ^ n7174 ^ 1'b0 ;
  assign n8595 = ~n8588 & n8594 ;
  assign n8598 = n8597 ^ n8595 ^ 1'b0 ;
  assign n8599 = n4566 ^ n4551 ^ x102 ;
  assign n8600 = ~n4521 & n8599 ;
  assign n8601 = n8600 ^ n6692 ^ n4217 ;
  assign n8607 = x107 & n2357 ;
  assign n8608 = n2634 & n8607 ;
  assign n8606 = n1297 & ~n1336 ;
  assign n8609 = n8608 ^ n8606 ^ 1'b0 ;
  assign n8602 = n296 & ~n994 ;
  assign n8603 = n8602 ^ n3597 ^ n1620 ;
  assign n8604 = n5945 ^ n2036 ^ 1'b0 ;
  assign n8605 = n8603 & ~n8604 ;
  assign n8610 = n8609 ^ n8605 ^ n5419 ;
  assign n8611 = n4244 ^ n3113 ^ n566 ;
  assign n8612 = ( n902 & n1728 ) | ( n902 & n8611 ) | ( n1728 & n8611 ) ;
  assign n8613 = ( n1180 & ~n2846 ) | ( n1180 & n8612 ) | ( ~n2846 & n8612 ) ;
  assign n8614 = n3251 | n5259 ;
  assign n8615 = n8614 ^ n4701 ^ n2870 ;
  assign n8616 = ( n273 & ~n2685 ) | ( n273 & n8615 ) | ( ~n2685 & n8615 ) ;
  assign n8617 = n5011 & ~n8097 ;
  assign n8622 = n1017 & ~n1199 ;
  assign n8623 = n3671 & n8622 ;
  assign n8624 = n2996 | n8399 ;
  assign n8625 = ( n2701 & ~n8623 ) | ( n2701 & n8624 ) | ( ~n8623 & n8624 ) ;
  assign n8618 = n6113 ^ n4504 ^ n4441 ;
  assign n8619 = n8618 ^ n8111 ^ n4406 ;
  assign n8620 = n8619 ^ n8078 ^ n3242 ;
  assign n8621 = n7952 | n8620 ;
  assign n8626 = n8625 ^ n8621 ^ n5016 ;
  assign n8627 = n8431 ^ n5610 ^ n5530 ;
  assign n8628 = n8627 ^ n2486 ^ n839 ;
  assign n8629 = n3196 ^ n1680 ^ n912 ;
  assign n8630 = ( ~n243 & n3169 ) | ( ~n243 & n8162 ) | ( n3169 & n8162 ) ;
  assign n8631 = ( ~n1763 & n5385 ) | ( ~n1763 & n7882 ) | ( n5385 & n7882 ) ;
  assign n8632 = ( n4655 & ~n6103 ) | ( n4655 & n8631 ) | ( ~n6103 & n8631 ) ;
  assign n8633 = n6199 & n8632 ;
  assign n8634 = ( n8629 & n8630 ) | ( n8629 & ~n8633 ) | ( n8630 & ~n8633 ) ;
  assign n8635 = ~n8628 & n8634 ;
  assign n8636 = n3038 & n8635 ;
  assign n8637 = n1845 | n7336 ;
  assign n8639 = ( ~n2685 & n3101 ) | ( ~n2685 & n7812 ) | ( n3101 & n7812 ) ;
  assign n8638 = n2710 ^ n2560 ^ 1'b0 ;
  assign n8640 = n8639 ^ n8638 ^ n4987 ;
  assign n8641 = ( n315 & n1492 ) | ( n315 & n4010 ) | ( n1492 & n4010 ) ;
  assign n8642 = n8641 ^ n6084 ^ 1'b0 ;
  assign n8643 = ~n1009 & n1305 ;
  assign n8644 = ~n1886 & n8643 ;
  assign n8645 = n8644 ^ n7787 ^ n3026 ;
  assign n8646 = ( n3200 & n5725 ) | ( n3200 & n7674 ) | ( n5725 & n7674 ) ;
  assign n8647 = n6968 ^ n6416 ^ 1'b0 ;
  assign n8648 = n8365 ^ n5957 ^ 1'b0 ;
  assign n8649 = n6796 ^ n1890 ^ n1322 ;
  assign n8650 = ( ~n1034 & n6885 ) | ( ~n1034 & n8649 ) | ( n6885 & n8649 ) ;
  assign n8651 = n2429 & ~n4946 ;
  assign n8652 = ( ~n1993 & n3169 ) | ( ~n1993 & n8651 ) | ( n3169 & n8651 ) ;
  assign n8653 = ( ~n5080 & n8650 ) | ( ~n5080 & n8652 ) | ( n8650 & n8652 ) ;
  assign n8655 = n2483 & n4061 ;
  assign n8654 = n6821 ^ n6282 ^ n964 ;
  assign n8656 = n8655 ^ n8654 ^ 1'b0 ;
  assign n8657 = n1948 & n8656 ;
  assign n8660 = ( n237 & ~n1434 ) | ( n237 & n1884 ) | ( ~n1434 & n1884 ) ;
  assign n8658 = ~n2851 & n8527 ;
  assign n8659 = ( n3249 & ~n4201 ) | ( n3249 & n8658 ) | ( ~n4201 & n8658 ) ;
  assign n8661 = n8660 ^ n8659 ^ n5196 ;
  assign n8662 = ( n741 & n1391 ) | ( n741 & ~n6403 ) | ( n1391 & ~n6403 ) ;
  assign n8663 = n8662 ^ n3543 ^ n566 ;
  assign n8664 = ( ~n2582 & n7602 ) | ( ~n2582 & n8663 ) | ( n7602 & n8663 ) ;
  assign n8665 = n6201 ^ n5016 ^ 1'b0 ;
  assign n8666 = ~n6548 & n8665 ;
  assign n8667 = ( ~n4304 & n8019 ) | ( ~n4304 & n8666 ) | ( n8019 & n8666 ) ;
  assign n8668 = n7471 ^ n312 ^ 1'b0 ;
  assign n8669 = ~n2089 & n8668 ;
  assign n8670 = n8669 ^ n1309 ^ 1'b0 ;
  assign n8671 = ~n2486 & n8670 ;
  assign n8672 = ~n965 & n8671 ;
  assign n8673 = n6180 ^ n909 ^ 1'b0 ;
  assign n8674 = ~n8672 & n8673 ;
  assign n8675 = n7734 ^ n3257 ^ 1'b0 ;
  assign n8676 = ~n561 & n4002 ;
  assign n8677 = n5744 ^ n4781 ^ n1628 ;
  assign n8678 = n8676 & n8677 ;
  assign n8679 = n3431 ^ n3264 ^ 1'b0 ;
  assign n8680 = x24 & n8679 ;
  assign n8681 = n7231 & n8680 ;
  assign n8682 = n8681 ^ n5969 ^ n1947 ;
  assign n8683 = ( n1341 & n2025 ) | ( n1341 & n7238 ) | ( n2025 & n7238 ) ;
  assign n8684 = n6033 & n7427 ;
  assign n8685 = ( n1205 & n4303 ) | ( n1205 & n7175 ) | ( n4303 & n7175 ) ;
  assign n8686 = ( ~n1151 & n1973 ) | ( ~n1151 & n3117 ) | ( n1973 & n3117 ) ;
  assign n8687 = n8686 ^ n2482 ^ 1'b0 ;
  assign n8688 = ~n6347 & n7472 ;
  assign n8689 = n3188 | n4972 ;
  assign n8690 = n8688 | n8689 ;
  assign n8691 = n1195 ^ n513 ^ 1'b0 ;
  assign n8692 = ( n1865 & n2908 ) | ( n1865 & ~n8691 ) | ( n2908 & ~n8691 ) ;
  assign n8693 = ( ~n2996 & n3488 ) | ( ~n2996 & n8692 ) | ( n3488 & n8692 ) ;
  assign n8694 = n8693 ^ n2689 ^ n1348 ;
  assign n8695 = ( n1662 & n3871 ) | ( n1662 & n4357 ) | ( n3871 & n4357 ) ;
  assign n8696 = n252 & n4551 ;
  assign n8697 = ( n3145 & n4461 ) | ( n3145 & n8696 ) | ( n4461 & n8696 ) ;
  assign n8698 = ( n2431 & n5957 ) | ( n2431 & ~n8697 ) | ( n5957 & ~n8697 ) ;
  assign n8699 = ( n2191 & n8695 ) | ( n2191 & n8698 ) | ( n8695 & n8698 ) ;
  assign n8700 = ( n4002 & n8694 ) | ( n4002 & n8699 ) | ( n8694 & n8699 ) ;
  assign n8701 = ( n1457 & n4717 ) | ( n1457 & n7644 ) | ( n4717 & n7644 ) ;
  assign n8702 = ( n310 & ~n734 ) | ( n310 & n4931 ) | ( ~n734 & n4931 ) ;
  assign n8703 = n485 & n816 ;
  assign n8704 = n1501 | n8703 ;
  assign n8705 = ( n7917 & ~n8702 ) | ( n7917 & n8704 ) | ( ~n8702 & n8704 ) ;
  assign n8706 = ( n738 & n8701 ) | ( n738 & n8705 ) | ( n8701 & n8705 ) ;
  assign n8707 = n389 & ~n2673 ;
  assign n8708 = n2543 ^ n851 ^ n131 ;
  assign n8711 = ( n2663 & ~n6237 ) | ( n2663 & n8614 ) | ( ~n6237 & n8614 ) ;
  assign n8709 = n1870 | n3890 ;
  assign n8710 = n8709 ^ n7530 ^ 1'b0 ;
  assign n8712 = n8711 ^ n8710 ^ n6713 ;
  assign n8713 = n7947 ^ n7801 ^ 1'b0 ;
  assign n8714 = n3454 | n8713 ;
  assign n8715 = n6408 ^ n1038 ^ 1'b0 ;
  assign n8716 = n1093 | n7290 ;
  assign n8717 = n8715 | n8716 ;
  assign n8718 = n7311 ^ n7243 ^ n7006 ;
  assign n8719 = ( ~n967 & n8717 ) | ( ~n967 & n8718 ) | ( n8717 & n8718 ) ;
  assign n8720 = ~n3079 & n3096 ;
  assign n8721 = n8720 ^ n1332 ^ 1'b0 ;
  assign n8722 = ~n7710 & n8721 ;
  assign n8723 = n8722 ^ n2646 ^ 1'b0 ;
  assign n8724 = n7439 ^ n6064 ^ 1'b0 ;
  assign n8725 = n827 & ~n8724 ;
  assign n8726 = n6943 ^ n5822 ^ n1019 ;
  assign n8727 = n1136 ^ n195 ^ 1'b0 ;
  assign n8728 = n8727 ^ n3816 ^ 1'b0 ;
  assign n8729 = ( n2044 & n2583 ) | ( n2044 & n6287 ) | ( n2583 & n6287 ) ;
  assign n8730 = n8729 ^ n5949 ^ n3148 ;
  assign n8731 = n8730 ^ n6128 ^ n5157 ;
  assign n8732 = n8731 ^ n8430 ^ 1'b0 ;
  assign n8733 = n5808 ^ n3151 ^ 1'b0 ;
  assign n8734 = n1213 & n8733 ;
  assign n8735 = n8734 ^ n5063 ^ 1'b0 ;
  assign n8740 = n3620 ^ n2306 ^ n2059 ;
  assign n8741 = n2282 | n8740 ;
  assign n8742 = n8741 ^ n545 ^ 1'b0 ;
  assign n8737 = n2607 ^ n1906 ^ n890 ;
  assign n8738 = n8737 ^ n3410 ^ n2798 ;
  assign n8736 = ( x5 & n1072 ) | ( x5 & ~n7922 ) | ( n1072 & ~n7922 ) ;
  assign n8739 = n8738 ^ n8736 ^ n4212 ;
  assign n8743 = n8742 ^ n8739 ^ n7646 ;
  assign n8744 = ( n1677 & n1727 ) | ( n1677 & n4153 ) | ( n1727 & n4153 ) ;
  assign n8745 = n8744 ^ n1259 ^ 1'b0 ;
  assign n8746 = n3007 | n8745 ;
  assign n8747 = n6023 & ~n8746 ;
  assign n8748 = n8747 ^ n3705 ^ 1'b0 ;
  assign n8749 = ( n3874 & ~n6682 ) | ( n3874 & n8748 ) | ( ~n6682 & n8748 ) ;
  assign n8753 = n3197 ^ n2559 ^ n2260 ;
  assign n8754 = n8753 ^ n1250 ^ n433 ;
  assign n8755 = n1445 & ~n8754 ;
  assign n8750 = ~n3159 & n8566 ;
  assign n8751 = ~n6104 & n8750 ;
  assign n8752 = n2642 & ~n8751 ;
  assign n8756 = n8755 ^ n8752 ^ n6898 ;
  assign n8757 = ( ~n5733 & n8749 ) | ( ~n5733 & n8756 ) | ( n8749 & n8756 ) ;
  assign n8758 = n3990 ^ n1463 ^ n1131 ;
  assign n8759 = n5702 ^ n1646 ^ 1'b0 ;
  assign n8760 = ( n2236 & ~n3192 ) | ( n2236 & n8759 ) | ( ~n3192 & n8759 ) ;
  assign n8761 = ~n8758 & n8760 ;
  assign n8762 = n2821 & n8761 ;
  assign n8763 = n1905 ^ n1486 ^ 1'b0 ;
  assign n8764 = n8763 ^ n8539 ^ n2381 ;
  assign n8765 = n8764 ^ n3227 ^ n825 ;
  assign n8766 = n5672 ^ n4636 ^ 1'b0 ;
  assign n8767 = n8765 & n8766 ;
  assign n8768 = n5415 ^ n5215 ^ n2569 ;
  assign n8769 = ( ~n1614 & n2512 ) | ( ~n1614 & n8532 ) | ( n2512 & n8532 ) ;
  assign n8770 = ( n1961 & n3521 ) | ( n1961 & ~n5489 ) | ( n3521 & ~n5489 ) ;
  assign n8771 = ( n646 & n8769 ) | ( n646 & n8770 ) | ( n8769 & n8770 ) ;
  assign n8772 = n8768 & n8771 ;
  assign n8773 = ( ~n324 & n5405 ) | ( ~n324 & n6665 ) | ( n5405 & n6665 ) ;
  assign n8774 = x64 & ~n7139 ;
  assign n8775 = n8774 ^ n2610 ^ 1'b0 ;
  assign n8776 = n1521 & n5684 ;
  assign n8777 = n8776 ^ n7127 ^ 1'b0 ;
  assign n8778 = ( ~n6736 & n8775 ) | ( ~n6736 & n8777 ) | ( n8775 & n8777 ) ;
  assign n8781 = n5602 ^ n5412 ^ 1'b0 ;
  assign n8779 = n7952 ^ n3411 ^ 1'b0 ;
  assign n8780 = n8779 ^ n7375 ^ n201 ;
  assign n8782 = n8781 ^ n8780 ^ n6180 ;
  assign n8783 = n3075 ^ n2587 ^ 1'b0 ;
  assign n8784 = ~n3866 & n7527 ;
  assign n8785 = n1334 & n8784 ;
  assign n8786 = n8785 ^ n5862 ^ n313 ;
  assign n8787 = n8786 ^ n6938 ^ n2827 ;
  assign n8788 = n2648 ^ n2417 ^ n726 ;
  assign n8789 = n6010 ^ n337 ^ 1'b0 ;
  assign n8790 = ( ~n7542 & n8788 ) | ( ~n7542 & n8789 ) | ( n8788 & n8789 ) ;
  assign n8791 = ( n2385 & n6896 ) | ( n2385 & n8790 ) | ( n6896 & n8790 ) ;
  assign n8792 = ( n2425 & n4259 ) | ( n2425 & ~n8391 ) | ( n4259 & ~n8391 ) ;
  assign n8793 = n3208 ^ n1959 ^ n340 ;
  assign n8794 = ( n890 & ~n8792 ) | ( n890 & n8793 ) | ( ~n8792 & n8793 ) ;
  assign n8795 = ( x73 & ~n8791 ) | ( x73 & n8794 ) | ( ~n8791 & n8794 ) ;
  assign n8796 = n1815 | n7022 ;
  assign n8797 = n8796 ^ n3158 ^ 1'b0 ;
  assign n8798 = n8797 ^ n8769 ^ n5480 ;
  assign n8799 = x49 & ~n7246 ;
  assign n8800 = ( n1630 & n2941 ) | ( n1630 & n4987 ) | ( n2941 & n4987 ) ;
  assign n8801 = n1127 | n4077 ;
  assign n8802 = n1664 | n8801 ;
  assign n8803 = ( n935 & n1396 ) | ( n935 & n8802 ) | ( n1396 & n8802 ) ;
  assign n8804 = ~n1962 & n8803 ;
  assign n8805 = n7520 & n8804 ;
  assign n8806 = ( n199 & n646 ) | ( n199 & n5004 ) | ( n646 & n5004 ) ;
  assign n8807 = ~n659 & n8806 ;
  assign n8808 = n5339 | n8807 ;
  assign n8809 = ( n5201 & n8453 ) | ( n5201 & n8808 ) | ( n8453 & n8808 ) ;
  assign n8813 = n204 | n4557 ;
  assign n8810 = n3098 & ~n3670 ;
  assign n8811 = ( ~n6495 & n7953 ) | ( ~n6495 & n8810 ) | ( n7953 & n8810 ) ;
  assign n8812 = ( n1483 & n3992 ) | ( n1483 & n8811 ) | ( n3992 & n8811 ) ;
  assign n8814 = n8813 ^ n8812 ^ n3871 ;
  assign n8815 = n7972 ^ n4857 ^ n1557 ;
  assign n8816 = n6167 ^ n4497 ^ n180 ;
  assign n8817 = n8816 ^ n2465 ^ 1'b0 ;
  assign n8818 = n8815 & n8817 ;
  assign n8828 = n3096 ^ n1391 ^ n778 ;
  assign n8826 = ( n1845 & n2311 ) | ( n1845 & n6990 ) | ( n2311 & n6990 ) ;
  assign n8827 = x103 & ~n8826 ;
  assign n8829 = n8828 ^ n8827 ^ n5926 ;
  assign n8819 = n3967 ^ n3302 ^ n428 ;
  assign n8820 = n8819 ^ n2994 ^ n1761 ;
  assign n8821 = n8820 ^ n4350 ^ n1912 ;
  assign n8822 = n8821 ^ n1297 ^ 1'b0 ;
  assign n8823 = n1580 ^ n1027 ^ n725 ;
  assign n8824 = n8823 ^ n335 ^ 1'b0 ;
  assign n8825 = n8822 & ~n8824 ;
  assign n8830 = n8829 ^ n8825 ^ n7858 ;
  assign n8831 = n6544 ^ n4907 ^ 1'b0 ;
  assign n8832 = n8831 ^ n6998 ^ n2854 ;
  assign n8833 = ( ~n2446 & n2720 ) | ( ~n2446 & n6868 ) | ( n2720 & n6868 ) ;
  assign n8834 = ( n1340 & n2686 ) | ( n1340 & ~n5080 ) | ( n2686 & ~n5080 ) ;
  assign n8835 = n8834 ^ n7254 ^ n6810 ;
  assign n8836 = ( n6582 & n8833 ) | ( n6582 & n8835 ) | ( n8833 & n8835 ) ;
  assign n8837 = n989 & ~n5694 ;
  assign n8838 = ~n3413 & n7625 ;
  assign n8839 = n565 & n8838 ;
  assign n8840 = n673 | n8839 ;
  assign n8841 = n8837 & ~n8840 ;
  assign n8842 = n1913 & n3712 ;
  assign n8843 = ~n2242 & n8842 ;
  assign n8844 = ( n2218 & n4667 ) | ( n2218 & n8843 ) | ( n4667 & n8843 ) ;
  assign n8845 = n8844 ^ n1050 ^ 1'b0 ;
  assign n8846 = ~n5848 & n5930 ;
  assign n8847 = ( n6261 & ~n8845 ) | ( n6261 & n8846 ) | ( ~n8845 & n8846 ) ;
  assign n8848 = ( n352 & n3292 ) | ( n352 & ~n3580 ) | ( n3292 & ~n3580 ) ;
  assign n8849 = n4527 ^ n3646 ^ 1'b0 ;
  assign n8850 = ( n565 & n8848 ) | ( n565 & ~n8849 ) | ( n8848 & ~n8849 ) ;
  assign n8851 = ( n2385 & n5291 ) | ( n2385 & ~n5598 ) | ( n5291 & ~n5598 ) ;
  assign n8852 = n8851 ^ n2854 ^ n2124 ;
  assign n8853 = n2031 ^ n1766 ^ n1125 ;
  assign n8854 = ( n2102 & ~n2537 ) | ( n2102 & n4490 ) | ( ~n2537 & n4490 ) ;
  assign n8855 = ( n4384 & n8853 ) | ( n4384 & ~n8854 ) | ( n8853 & ~n8854 ) ;
  assign n8856 = ( n1095 & n5622 ) | ( n1095 & n8855 ) | ( n5622 & n8855 ) ;
  assign n8857 = n8856 ^ n1932 ^ n857 ;
  assign n8858 = ( ~n2145 & n3443 ) | ( ~n2145 & n5537 ) | ( n3443 & n5537 ) ;
  assign n8859 = n8858 ^ n1498 ^ 1'b0 ;
  assign n8860 = n2596 & ~n8744 ;
  assign n8861 = ~n3615 & n8860 ;
  assign n8862 = ( n7098 & ~n7621 ) | ( n7098 & n8393 ) | ( ~n7621 & n8393 ) ;
  assign n8863 = ( n3499 & n8861 ) | ( n3499 & ~n8862 ) | ( n8861 & ~n8862 ) ;
  assign n8868 = x40 & n2842 ;
  assign n8869 = ( ~x12 & n3320 ) | ( ~x12 & n8868 ) | ( n3320 & n8868 ) ;
  assign n8866 = n7323 ^ n2703 ^ n2406 ;
  assign n8864 = n6778 ^ n2862 ^ n571 ;
  assign n8865 = ( n508 & n3175 ) | ( n508 & ~n8864 ) | ( n3175 & ~n8864 ) ;
  assign n8867 = n8866 ^ n8865 ^ x107 ;
  assign n8870 = n8869 ^ n8867 ^ 1'b0 ;
  assign n8871 = ( n3915 & n6720 ) | ( n3915 & n6898 ) | ( n6720 & n6898 ) ;
  assign n8872 = ~n3111 & n5774 ;
  assign n8873 = ~n8871 & n8872 ;
  assign n8874 = n3954 ^ n3922 ^ 1'b0 ;
  assign n8875 = n8874 ^ n6343 ^ n4740 ;
  assign n8876 = n2115 & ~n2780 ;
  assign n8877 = x84 & ~n8876 ;
  assign n8878 = n8877 ^ n5897 ^ 1'b0 ;
  assign n8879 = n4072 & n8878 ;
  assign n8880 = n8879 ^ n6396 ^ 1'b0 ;
  assign n8881 = n1037 & ~n4581 ;
  assign n8882 = n8881 ^ n3657 ^ 1'b0 ;
  assign n8892 = n1930 ^ n972 ^ n479 ;
  assign n8893 = n8892 ^ n820 ^ 1'b0 ;
  assign n8894 = ~n1673 & n8893 ;
  assign n8895 = ~n3773 & n8894 ;
  assign n8896 = ( n1142 & ~n1258 ) | ( n1142 & n8895 ) | ( ~n1258 & n8895 ) ;
  assign n8889 = ( n885 & n2521 ) | ( n885 & ~n3548 ) | ( n2521 & ~n3548 ) ;
  assign n8890 = n8889 ^ n5070 ^ n3169 ;
  assign n8884 = ~n4619 & n5058 ;
  assign n8885 = ( n214 & n1174 ) | ( n214 & n8884 ) | ( n1174 & n8884 ) ;
  assign n8886 = n8885 ^ n1885 ^ 1'b0 ;
  assign n8887 = ( n3375 & n7497 ) | ( n3375 & ~n8886 ) | ( n7497 & ~n8886 ) ;
  assign n8883 = n373 | n7805 ;
  assign n8888 = n8887 ^ n8883 ^ n4593 ;
  assign n8891 = n8890 ^ n8888 ^ n1632 ;
  assign n8897 = n8896 ^ n8891 ^ n4754 ;
  assign n8899 = ( x46 & ~n301 ) | ( x46 & n841 ) | ( ~n301 & n841 ) ;
  assign n8898 = n4428 ^ n3643 ^ n2294 ;
  assign n8900 = n8899 ^ n8898 ^ 1'b0 ;
  assign n8901 = ( n304 & n4868 ) | ( n304 & n8900 ) | ( n4868 & n8900 ) ;
  assign n8902 = n4831 ^ n2554 ^ n2247 ;
  assign n8903 = n6023 ^ n3899 ^ n699 ;
  assign n8904 = n8903 ^ n6825 ^ 1'b0 ;
  assign n8905 = n272 & n4545 ;
  assign n8906 = n6514 & n8905 ;
  assign n8907 = ( n2113 & n7977 ) | ( n2113 & n8906 ) | ( n7977 & n8906 ) ;
  assign n8908 = n1953 | n6508 ;
  assign n8909 = n8908 ^ n8543 ^ 1'b0 ;
  assign n8910 = ( n4858 & ~n5713 ) | ( n4858 & n8909 ) | ( ~n5713 & n8909 ) ;
  assign n8911 = ( x102 & n983 ) | ( x102 & n8072 ) | ( n983 & n8072 ) ;
  assign n8915 = n3688 ^ n998 ^ 1'b0 ;
  assign n8912 = n518 & n2765 ;
  assign n8913 = n8912 ^ n7064 ^ n6363 ;
  assign n8914 = n8913 ^ n6961 ^ n5648 ;
  assign n8916 = n8915 ^ n8914 ^ 1'b0 ;
  assign n8918 = n3726 ^ n2314 ^ n1670 ;
  assign n8917 = n4544 ^ n4505 ^ n3257 ;
  assign n8919 = n8918 ^ n8917 ^ n1779 ;
  assign n8920 = ( n7667 & ~n7937 ) | ( n7667 & n8919 ) | ( ~n7937 & n8919 ) ;
  assign n8921 = n8920 ^ n2196 ^ 1'b0 ;
  assign n8922 = n5205 & n8921 ;
  assign n8923 = ( n1566 & n4477 ) | ( n1566 & n7021 ) | ( n4477 & n7021 ) ;
  assign n8924 = x109 & ~n8923 ;
  assign n8925 = n8924 ^ n2321 ^ 1'b0 ;
  assign n8926 = n4150 ^ n375 ^ 1'b0 ;
  assign n8927 = ~n6928 & n8926 ;
  assign n8928 = ( n3019 & n7459 ) | ( n3019 & ~n8927 ) | ( n7459 & ~n8927 ) ;
  assign n8929 = n8928 ^ n6826 ^ n2350 ;
  assign n8930 = n8207 ^ n4951 ^ n1625 ;
  assign n8931 = n2539 ^ n671 ^ 1'b0 ;
  assign n8932 = n8931 ^ n5821 ^ 1'b0 ;
  assign n8933 = n8930 & ~n8932 ;
  assign n8939 = n1951 | n3463 ;
  assign n8934 = n8270 ^ n3825 ^ n3037 ;
  assign n8935 = n8934 ^ n3940 ^ n1428 ;
  assign n8936 = n4584 | n6103 ;
  assign n8937 = n1535 & ~n8936 ;
  assign n8938 = ( n5476 & ~n8935 ) | ( n5476 & n8937 ) | ( ~n8935 & n8937 ) ;
  assign n8940 = n8939 ^ n8938 ^ n8243 ;
  assign n8941 = n6766 ^ n3450 ^ n721 ;
  assign n8942 = ( n763 & ~n5074 ) | ( n763 & n8941 ) | ( ~n5074 & n8941 ) ;
  assign n8947 = n7488 ^ n2024 ^ n1984 ;
  assign n8943 = n8230 ^ n4383 ^ n1349 ;
  assign n8944 = n8943 ^ n7724 ^ n2894 ;
  assign n8945 = n8944 ^ n5398 ^ 1'b0 ;
  assign n8946 = n935 & ~n8945 ;
  assign n8948 = n8947 ^ n8946 ^ 1'b0 ;
  assign n8951 = n277 | n2211 ;
  assign n8952 = n175 | n8951 ;
  assign n8949 = ( n386 & ~n1284 ) | ( n386 & n3845 ) | ( ~n1284 & n3845 ) ;
  assign n8950 = ( n677 & n2728 ) | ( n677 & ~n8949 ) | ( n2728 & ~n8949 ) ;
  assign n8953 = n8952 ^ n8950 ^ n2779 ;
  assign n8954 = n8953 ^ n7781 ^ n5570 ;
  assign n8955 = n3288 & n3306 ;
  assign n8956 = ~n5945 & n8955 ;
  assign n8957 = n7704 | n8956 ;
  assign n8958 = ( n4239 & n5797 ) | ( n4239 & ~n8957 ) | ( n5797 & ~n8957 ) ;
  assign n8959 = ( n558 & ~n1163 ) | ( n558 & n6983 ) | ( ~n1163 & n6983 ) ;
  assign n8960 = n899 & n6078 ;
  assign n8961 = n8581 ^ n513 ^ 1'b0 ;
  assign n8962 = ~n2439 & n7647 ;
  assign n8963 = ( n1964 & ~n5968 ) | ( n1964 & n8962 ) | ( ~n5968 & n8962 ) ;
  assign n8964 = ~n1912 & n6462 ;
  assign n8965 = n5045 ^ n4992 ^ n1678 ;
  assign n8966 = n4341 ^ n2713 ^ n2660 ;
  assign n8967 = n8966 ^ n3889 ^ n3788 ;
  assign n8968 = n8967 ^ n3093 ^ n2712 ;
  assign n8978 = ( n1381 & n2473 ) | ( n1381 & n3697 ) | ( n2473 & n3697 ) ;
  assign n8969 = n4895 ^ n1013 ^ 1'b0 ;
  assign n8970 = n1496 & n8969 ;
  assign n8971 = n5187 ^ n3871 ^ 1'b0 ;
  assign n8972 = n8390 & n8971 ;
  assign n8973 = ( n589 & ~n8970 ) | ( n589 & n8972 ) | ( ~n8970 & n8972 ) ;
  assign n8974 = n8973 ^ n7106 ^ 1'b0 ;
  assign n8975 = n5731 ^ n4565 ^ 1'b0 ;
  assign n8976 = n8974 | n8975 ;
  assign n8977 = n4028 & ~n8976 ;
  assign n8979 = n8978 ^ n8977 ^ 1'b0 ;
  assign n8980 = n3959 ^ n604 ^ 1'b0 ;
  assign n8981 = ( x116 & ~n1657 ) | ( x116 & n2997 ) | ( ~n1657 & n2997 ) ;
  assign n8983 = x69 & n2014 ;
  assign n8984 = ( n2053 & ~n4284 ) | ( n2053 & n8983 ) | ( ~n4284 & n8983 ) ;
  assign n8982 = n7963 ^ n7441 ^ 1'b0 ;
  assign n8985 = n8984 ^ n8982 ^ n7909 ;
  assign n8986 = n5466 ^ n4466 ^ 1'b0 ;
  assign n8987 = n8986 ^ n4600 ^ n3602 ;
  assign n8988 = n2210 ^ n131 ^ 1'b0 ;
  assign n8989 = ( n4730 & n5248 ) | ( n4730 & ~n8988 ) | ( n5248 & ~n8988 ) ;
  assign n8990 = n8989 ^ n8385 ^ n5079 ;
  assign n8991 = n8990 ^ n3045 ^ n2555 ;
  assign n8992 = n7122 ^ n1614 ^ x83 ;
  assign n8993 = n8992 ^ n7369 ^ 1'b0 ;
  assign n8994 = n6931 ^ n339 ^ 1'b0 ;
  assign n8995 = n2080 & n8994 ;
  assign n8996 = ( n920 & n4600 ) | ( n920 & ~n8995 ) | ( n4600 & ~n8995 ) ;
  assign n8997 = n3250 | n4609 ;
  assign n8998 = n8996 | n8997 ;
  assign n8999 = n984 & n8998 ;
  assign n9000 = n8999 ^ n5582 ^ 1'b0 ;
  assign n9001 = ( n4062 & n4308 ) | ( n4062 & n5041 ) | ( n4308 & n5041 ) ;
  assign n9002 = n9001 ^ n4242 ^ n1381 ;
  assign n9003 = n1893 & ~n4510 ;
  assign n9004 = n9003 ^ x38 ^ 1'b0 ;
  assign n9005 = n926 & ~n8101 ;
  assign n9006 = ~n8970 & n9005 ;
  assign n9007 = n9006 ^ n1657 ^ 1'b0 ;
  assign n9008 = n3428 | n9007 ;
  assign n9009 = n5044 ^ n3150 ^ 1'b0 ;
  assign n9010 = ( n393 & n758 ) | ( n393 & n4918 ) | ( n758 & n4918 ) ;
  assign n9011 = n9010 ^ n7179 ^ n1532 ;
  assign n9012 = ( n2936 & n9009 ) | ( n2936 & n9011 ) | ( n9009 & n9011 ) ;
  assign n9013 = n9012 ^ n356 ^ 1'b0 ;
  assign n9014 = n2339 ^ n1559 ^ n669 ;
  assign n9015 = ( x88 & n304 ) | ( x88 & n2817 ) | ( n304 & n2817 ) ;
  assign n9016 = n9015 ^ n3074 ^ 1'b0 ;
  assign n9017 = ( n7951 & n9014 ) | ( n7951 & n9016 ) | ( n9014 & n9016 ) ;
  assign n9018 = ~n1323 & n5056 ;
  assign n9019 = n680 & n9018 ;
  assign n9020 = n2503 | n3807 ;
  assign n9021 = n4529 | n9020 ;
  assign n9022 = ( n6490 & n9019 ) | ( n6490 & ~n9021 ) | ( n9019 & ~n9021 ) ;
  assign n9023 = ( n1694 & n4876 ) | ( n1694 & n6275 ) | ( n4876 & n6275 ) ;
  assign n9024 = n2513 & ~n9023 ;
  assign n9025 = n1694 & ~n2559 ;
  assign n9026 = n9025 ^ n6792 ^ 1'b0 ;
  assign n9027 = n9026 ^ n2922 ^ n2742 ;
  assign n9032 = ( ~n3130 & n4559 ) | ( ~n3130 & n7014 ) | ( n4559 & n7014 ) ;
  assign n9028 = n586 & n816 ;
  assign n9029 = n3629 ^ n568 ^ n547 ;
  assign n9030 = ( n2421 & n6703 ) | ( n2421 & ~n9029 ) | ( n6703 & ~n9029 ) ;
  assign n9031 = ( x100 & ~n9028 ) | ( x100 & n9030 ) | ( ~n9028 & n9030 ) ;
  assign n9033 = n9032 ^ n9031 ^ n6657 ;
  assign n9037 = ~n865 & n1263 ;
  assign n9034 = n6305 ^ x1 ^ 1'b0 ;
  assign n9035 = n2917 | n9034 ;
  assign n9036 = n306 | n9035 ;
  assign n9038 = n9037 ^ n9036 ^ n7647 ;
  assign n9039 = n5906 & ~n8048 ;
  assign n9040 = ( n5287 & n5922 ) | ( n5287 & ~n9039 ) | ( n5922 & ~n9039 ) ;
  assign n9041 = n9040 ^ n7471 ^ n5234 ;
  assign n9043 = ( n5081 & n5305 ) | ( n5081 & n7613 ) | ( n5305 & n7613 ) ;
  assign n9042 = n158 | n4109 ;
  assign n9044 = n9043 ^ n9042 ^ 1'b0 ;
  assign n9045 = n9044 ^ n2401 ^ 1'b0 ;
  assign n9046 = n7701 & ~n9045 ;
  assign n9047 = ( n467 & ~n1833 ) | ( n467 & n2557 ) | ( ~n1833 & n2557 ) ;
  assign n9048 = n9047 ^ n5121 ^ n3434 ;
  assign n9049 = n2299 ^ n843 ^ 1'b0 ;
  assign n9050 = n9048 & ~n9049 ;
  assign n9051 = n9050 ^ n1997 ^ 1'b0 ;
  assign n9052 = n8813 ^ n5078 ^ n1896 ;
  assign n9053 = n9052 ^ n6921 ^ n6198 ;
  assign n9067 = n8340 ^ n4086 ^ 1'b0 ;
  assign n9066 = ( n3563 & n5398 ) | ( n3563 & ~n6985 ) | ( n5398 & ~n6985 ) ;
  assign n9063 = n1936 ^ n859 ^ 1'b0 ;
  assign n9064 = n4037 | n9063 ;
  assign n9054 = ( n2482 & n3684 ) | ( n2482 & n6225 ) | ( n3684 & n6225 ) ;
  assign n9055 = n9054 ^ n2213 ^ 1'b0 ;
  assign n9056 = ~n2226 & n6052 ;
  assign n9057 = n186 & n9056 ;
  assign n9058 = n9055 | n9057 ;
  assign n9059 = n9058 ^ n6982 ^ 1'b0 ;
  assign n9060 = n7198 ^ n4413 ^ n3738 ;
  assign n9061 = x121 | n9060 ;
  assign n9062 = n9059 | n9061 ;
  assign n9065 = n9064 ^ n9062 ^ n8531 ;
  assign n9068 = n9067 ^ n9066 ^ n9065 ;
  assign n9069 = ( n2937 & n9053 ) | ( n2937 & ~n9068 ) | ( n9053 & ~n9068 ) ;
  assign n9070 = ( n520 & ~n3623 ) | ( n520 & n7677 ) | ( ~n3623 & n7677 ) ;
  assign n9071 = n6094 | n9070 ;
  assign n9072 = n9071 ^ n3977 ^ 1'b0 ;
  assign n9073 = ( n175 & ~n7264 ) | ( n175 & n9072 ) | ( ~n7264 & n9072 ) ;
  assign n9080 = n4553 ^ n2385 ^ 1'b0 ;
  assign n9081 = ~n3630 & n9080 ;
  assign n9076 = ( n471 & n1045 ) | ( n471 & ~n4217 ) | ( n1045 & ~n4217 ) ;
  assign n9074 = n2927 ^ n2134 ^ 1'b0 ;
  assign n9075 = ~n1235 & n9074 ;
  assign n9077 = n9076 ^ n9075 ^ n341 ;
  assign n9078 = n3886 ^ n562 ^ 1'b0 ;
  assign n9079 = n9077 & n9078 ;
  assign n9082 = n9081 ^ n9079 ^ n6024 ;
  assign n9083 = n161 & n7230 ;
  assign n9084 = ~n3029 & n9083 ;
  assign n9085 = n9084 ^ n8493 ^ n5557 ;
  assign n9086 = n4001 ^ n766 ^ 1'b0 ;
  assign n9087 = n9086 ^ n5153 ^ n1118 ;
  assign n9088 = n799 & ~n3155 ;
  assign n9089 = n9088 ^ n6199 ^ 1'b0 ;
  assign n9090 = n1369 | n9089 ;
  assign n9091 = n8383 ^ x68 ^ 1'b0 ;
  assign n9096 = ( n2396 & ~n2506 ) | ( n2396 & n9054 ) | ( ~n2506 & n9054 ) ;
  assign n9095 = n8864 ^ n5303 ^ n2760 ;
  assign n9097 = n9096 ^ n9095 ^ n2701 ;
  assign n9092 = n310 | n1723 ;
  assign n9093 = x109 | n9092 ;
  assign n9094 = ~n1986 & n9093 ;
  assign n9098 = n9097 ^ n9094 ^ 1'b0 ;
  assign n9099 = n9098 ^ n3842 ^ 1'b0 ;
  assign n9100 = ( x75 & ~x90 ) | ( x75 & n4353 ) | ( ~x90 & n4353 ) ;
  assign n9101 = n3705 & ~n9100 ;
  assign n9102 = n9101 ^ n6739 ^ n5594 ;
  assign n9103 = ( n7087 & ~n9068 ) | ( n7087 & n9102 ) | ( ~n9068 & n9102 ) ;
  assign n9104 = n1400 ^ n1236 ^ n783 ;
  assign n9105 = ( n1163 & ~n2534 ) | ( n1163 & n6510 ) | ( ~n2534 & n6510 ) ;
  assign n9106 = n795 & n4228 ;
  assign n9107 = ~n9105 & n9106 ;
  assign n9108 = n9107 ^ n8446 ^ 1'b0 ;
  assign n9109 = ~n9104 & n9108 ;
  assign n9110 = n9109 ^ n645 ^ 1'b0 ;
  assign n9111 = n1394 & n6994 ;
  assign n9112 = n9111 ^ n4285 ^ 1'b0 ;
  assign n9113 = n5553 & n9112 ;
  assign n9114 = n9113 ^ n4743 ^ 1'b0 ;
  assign n9115 = ( ~n811 & n4425 ) | ( ~n811 & n7392 ) | ( n4425 & n7392 ) ;
  assign n9116 = n8082 | n9115 ;
  assign n9117 = n9116 ^ n2826 ^ 1'b0 ;
  assign n9118 = n9117 ^ n7208 ^ n1492 ;
  assign n9120 = n8073 ^ n5783 ^ n2193 ;
  assign n9119 = ( ~n202 & n1306 ) | ( ~n202 & n4547 ) | ( n1306 & n4547 ) ;
  assign n9121 = n9120 ^ n9119 ^ n4532 ;
  assign n9122 = n3283 & ~n9121 ;
  assign n9123 = n925 & ~n1912 ;
  assign n9124 = n9123 ^ n5563 ^ n5050 ;
  assign n9125 = n6972 & n9124 ;
  assign n9126 = ~n4058 & n9125 ;
  assign n9127 = n9126 ^ n4003 ^ 1'b0 ;
  assign n9128 = n5414 ^ n2146 ^ n457 ;
  assign n9129 = n9128 ^ n4626 ^ 1'b0 ;
  assign n9130 = n4392 ^ n2281 ^ 1'b0 ;
  assign n9131 = ~n9129 & n9130 ;
  assign n9132 = ( ~n175 & n3860 ) | ( ~n175 & n9131 ) | ( n3860 & n9131 ) ;
  assign n9133 = ( n1025 & ~n2114 ) | ( n1025 & n4055 ) | ( ~n2114 & n4055 ) ;
  assign n9134 = n9132 | n9133 ;
  assign n9135 = ( n205 & n2946 ) | ( n205 & n3824 ) | ( n2946 & n3824 ) ;
  assign n9136 = n1380 & n9135 ;
  assign n9140 = ( n277 & n1135 ) | ( n277 & n1334 ) | ( n1135 & n1334 ) ;
  assign n9137 = n4223 ^ n925 ^ 1'b0 ;
  assign n9138 = ( ~n1983 & n8233 ) | ( ~n1983 & n9137 ) | ( n8233 & n9137 ) ;
  assign n9139 = n1058 & ~n9138 ;
  assign n9141 = n9140 ^ n9139 ^ 1'b0 ;
  assign n9142 = n7079 ^ n4001 ^ n1568 ;
  assign n9146 = ( n5195 & n5537 ) | ( n5195 & ~n6438 ) | ( n5537 & ~n6438 ) ;
  assign n9147 = n9146 ^ n3351 ^ 1'b0 ;
  assign n9143 = ( n1911 & ~n2608 ) | ( n1911 & n4311 ) | ( ~n2608 & n4311 ) ;
  assign n9144 = ( n2579 & n4078 ) | ( n2579 & ~n9143 ) | ( n4078 & ~n9143 ) ;
  assign n9145 = n9144 ^ n3138 ^ n204 ;
  assign n9148 = n9147 ^ n9145 ^ n2582 ;
  assign n9149 = n7434 ^ n6104 ^ n3205 ;
  assign n9152 = n4640 ^ n4346 ^ 1'b0 ;
  assign n9153 = ~n848 & n9152 ;
  assign n9150 = ( n359 & ~n1075 ) | ( n359 & n3347 ) | ( ~n1075 & n3347 ) ;
  assign n9151 = n2137 & ~n9150 ;
  assign n9154 = n9153 ^ n9151 ^ 1'b0 ;
  assign n9155 = ( n8084 & ~n9149 ) | ( n8084 & n9154 ) | ( ~n9149 & n9154 ) ;
  assign n9156 = ( n1525 & n2817 ) | ( n1525 & n4801 ) | ( n2817 & n4801 ) ;
  assign n9157 = n9156 ^ n1333 ^ 1'b0 ;
  assign n9158 = ~n5545 & n9157 ;
  assign n9159 = ~n5148 & n9158 ;
  assign n9160 = n9159 ^ n8497 ^ 1'b0 ;
  assign n9161 = n2801 ^ n1233 ^ 1'b0 ;
  assign n9162 = n2550 & n9161 ;
  assign n9163 = n9162 ^ n4651 ^ 1'b0 ;
  assign n9164 = ~n902 & n3882 ;
  assign n9165 = n9163 | n9164 ;
  assign n9166 = n705 | n9165 ;
  assign n9167 = n8256 ^ n2218 ^ n1334 ;
  assign n9168 = n7667 & ~n9167 ;
  assign n9169 = n4233 | n9168 ;
  assign n9179 = n8552 ^ n7379 ^ n626 ;
  assign n9176 = ~n2935 & n5201 ;
  assign n9177 = n9176 ^ n5493 ^ n3525 ;
  assign n9172 = n2306 & ~n3202 ;
  assign n9173 = n1957 ^ n1362 ^ 1'b0 ;
  assign n9174 = n9173 ^ n1853 ^ 1'b0 ;
  assign n9175 = ( n6165 & ~n9172 ) | ( n6165 & n9174 ) | ( ~n9172 & n9174 ) ;
  assign n9178 = n9177 ^ n9175 ^ n2915 ;
  assign n9170 = ~n1409 & n4965 ;
  assign n9171 = ~n555 & n9170 ;
  assign n9180 = n9179 ^ n9178 ^ n9171 ;
  assign n9181 = n2377 ^ n1820 ^ 1'b0 ;
  assign n9182 = n3716 | n9181 ;
  assign n9183 = n7845 ^ n2158 ^ x65 ;
  assign n9184 = n7398 ^ x54 ^ 1'b0 ;
  assign n9185 = n9184 ^ n2974 ^ 1'b0 ;
  assign n9186 = ~n8371 & n9185 ;
  assign n9187 = ~n4505 & n5569 ;
  assign n9188 = ~n4398 & n9187 ;
  assign n9189 = ( n5321 & n9186 ) | ( n5321 & n9188 ) | ( n9186 & n9188 ) ;
  assign n9194 = n6013 ^ n4882 ^ 1'b0 ;
  assign n9195 = ( n722 & n1306 ) | ( n722 & ~n9194 ) | ( n1306 & ~n9194 ) ;
  assign n9190 = n8439 ^ n5060 ^ n1642 ;
  assign n9191 = n7952 ^ n4644 ^ n2325 ;
  assign n9192 = n9190 & n9191 ;
  assign n9193 = n5123 & n9192 ;
  assign n9196 = n9195 ^ n9193 ^ n1359 ;
  assign n9197 = n5644 ^ n4944 ^ 1'b0 ;
  assign n9198 = n258 & ~n9197 ;
  assign n9199 = ( n402 & ~n2594 ) | ( n402 & n6251 ) | ( ~n2594 & n6251 ) ;
  assign n9200 = ( ~n1034 & n2887 ) | ( ~n1034 & n3265 ) | ( n2887 & n3265 ) ;
  assign n9201 = n2286 & ~n9200 ;
  assign n9202 = ~n9199 & n9201 ;
  assign n9203 = n9198 & ~n9202 ;
  assign n9204 = n9203 ^ n4770 ^ 1'b0 ;
  assign n9208 = n6546 ^ n1616 ^ 1'b0 ;
  assign n9205 = n2401 & n6213 ;
  assign n9206 = ~n3076 & n9205 ;
  assign n9207 = n9206 ^ n4183 ^ n1315 ;
  assign n9209 = n9208 ^ n9207 ^ 1'b0 ;
  assign n9210 = ( n629 & n2705 ) | ( n629 & n7209 ) | ( n2705 & n7209 ) ;
  assign n9212 = ( n1016 & n4910 ) | ( n1016 & ~n8135 ) | ( n4910 & ~n8135 ) ;
  assign n9211 = ( n3575 & n3737 ) | ( n3575 & ~n6324 ) | ( n3737 & ~n6324 ) ;
  assign n9213 = n9212 ^ n9211 ^ 1'b0 ;
  assign n9216 = n1422 & ~n2206 ;
  assign n9217 = n9216 ^ n2329 ^ x58 ;
  assign n9214 = n3139 ^ n2011 ^ 1'b0 ;
  assign n9215 = n1148 & ~n9214 ;
  assign n9218 = n9217 ^ n9215 ^ n5508 ;
  assign n9219 = n6703 ^ n4953 ^ 1'b0 ;
  assign n9220 = ( n766 & ~n3335 ) | ( n766 & n8390 ) | ( ~n3335 & n8390 ) ;
  assign n9221 = n3520 ^ n2972 ^ 1'b0 ;
  assign n9222 = n2480 & n7316 ;
  assign n9223 = n9222 ^ n1781 ^ n332 ;
  assign n9224 = ( n9220 & n9221 ) | ( n9220 & ~n9223 ) | ( n9221 & ~n9223 ) ;
  assign n9225 = n5372 & n9224 ;
  assign n9226 = ~n9219 & n9225 ;
  assign n9232 = n1123 ^ n462 ^ 1'b0 ;
  assign n9233 = ~n4045 & n9232 ;
  assign n9227 = ~n600 & n3924 ;
  assign n9228 = ~n1512 & n6084 ;
  assign n9229 = n9228 ^ n8478 ^ 1'b0 ;
  assign n9230 = n9227 | n9229 ;
  assign n9231 = n5986 | n9230 ;
  assign n9234 = n9233 ^ n9231 ^ n160 ;
  assign n9235 = n5872 ^ n5214 ^ n3954 ;
  assign n9236 = ~n8229 & n8437 ;
  assign n9251 = n1612 | n2538 ;
  assign n9246 = n2983 ^ n2224 ^ x127 ;
  assign n9243 = n457 & n2346 ;
  assign n9244 = ~n261 & n9243 ;
  assign n9245 = n9244 ^ n1557 ^ n633 ;
  assign n9247 = n9246 ^ n9245 ^ n4692 ;
  assign n9240 = n3431 ^ n880 ^ 1'b0 ;
  assign n9241 = n3937 & ~n9240 ;
  assign n9237 = ( n581 & ~n2369 ) | ( n581 & n2882 ) | ( ~n2369 & n2882 ) ;
  assign n9238 = ( n3688 & ~n6186 ) | ( n3688 & n9237 ) | ( ~n6186 & n9237 ) ;
  assign n9239 = n2506 & ~n9238 ;
  assign n9242 = n9241 ^ n9239 ^ 1'b0 ;
  assign n9248 = n9247 ^ n9242 ^ 1'b0 ;
  assign n9249 = n9248 ^ n582 ^ n544 ;
  assign n9250 = ( ~n5455 & n8092 ) | ( ~n5455 & n9249 ) | ( n8092 & n9249 ) ;
  assign n9252 = n9251 ^ n9250 ^ n6113 ;
  assign n9259 = ( ~n1428 & n1916 ) | ( ~n1428 & n1993 ) | ( n1916 & n1993 ) ;
  assign n9260 = n6027 ^ n3548 ^ 1'b0 ;
  assign n9261 = n9259 & ~n9260 ;
  assign n9256 = ~n3413 & n7155 ;
  assign n9257 = n8608 & n9256 ;
  assign n9258 = ( n3210 & ~n8697 ) | ( n3210 & n9257 ) | ( ~n8697 & n9257 ) ;
  assign n9253 = ~n738 & n795 ;
  assign n9254 = n9253 ^ n3439 ^ 1'b0 ;
  assign n9255 = n9254 ^ n3529 ^ n273 ;
  assign n9262 = n9261 ^ n9258 ^ n9255 ;
  assign n9263 = n9262 ^ n1738 ^ 1'b0 ;
  assign n9264 = n7794 | n9263 ;
  assign n9265 = n825 | n5389 ;
  assign n9266 = n8115 & ~n9265 ;
  assign n9280 = n8949 ^ n2863 ^ n2273 ;
  assign n9267 = n6979 ^ n1999 ^ n1510 ;
  assign n9268 = n137 & n139 ;
  assign n9269 = ~n137 & n9268 ;
  assign n9270 = n1309 & n1395 ;
  assign n9271 = n9269 & n9270 ;
  assign n9272 = n9269 | n9271 ;
  assign n9273 = n9271 & ~n9272 ;
  assign n9274 = n1222 | n9273 ;
  assign n9275 = n1222 & ~n9274 ;
  assign n9276 = n9275 ^ n5969 ^ 1'b0 ;
  assign n9277 = n9267 | n9276 ;
  assign n9278 = n3364 ^ n2992 ^ 1'b0 ;
  assign n9279 = ~n9277 & n9278 ;
  assign n9281 = n9280 ^ n9279 ^ n5518 ;
  assign n9282 = n6845 ^ n1541 ^ 1'b0 ;
  assign n9286 = n5725 ^ n4034 ^ n1184 ;
  assign n9285 = ( n392 & n5278 ) | ( n392 & n6178 ) | ( n5278 & n6178 ) ;
  assign n9287 = n9286 ^ n9285 ^ n5556 ;
  assign n9288 = n9287 ^ n199 ^ 1'b0 ;
  assign n9289 = n4559 & ~n9288 ;
  assign n9290 = ~n8038 & n9289 ;
  assign n9291 = ~n4539 & n9290 ;
  assign n9283 = ( n2214 & ~n3373 ) | ( n2214 & n4087 ) | ( ~n3373 & n4087 ) ;
  assign n9284 = ~n2476 & n9283 ;
  assign n9292 = n9291 ^ n9284 ^ 1'b0 ;
  assign n9294 = x91 ^ x4 ^ 1'b0 ;
  assign n9295 = x83 & n9294 ;
  assign n9293 = n5751 ^ n1867 ^ 1'b0 ;
  assign n9296 = n9295 ^ n9293 ^ n6416 ;
  assign n9297 = ( ~x1 & n6964 ) | ( ~x1 & n9296 ) | ( n6964 & n9296 ) ;
  assign n9298 = n7439 & n8848 ;
  assign n9299 = n1408 & ~n9298 ;
  assign n9301 = ( ~n214 & n2013 ) | ( ~n214 & n5407 ) | ( n2013 & n5407 ) ;
  assign n9302 = n9301 ^ n860 ^ 1'b0 ;
  assign n9303 = ~n5784 & n9302 ;
  assign n9300 = n4966 ^ n4021 ^ n475 ;
  assign n9304 = n9303 ^ n9300 ^ n3126 ;
  assign n9305 = n8498 ^ n3212 ^ 1'b0 ;
  assign n9306 = n6352 ^ n5428 ^ n2775 ;
  assign n9307 = n9306 ^ n6240 ^ n2958 ;
  assign n9309 = ( ~n1947 & n2212 ) | ( ~n1947 & n3579 ) | ( n2212 & n3579 ) ;
  assign n9308 = ( n3139 & ~n3975 ) | ( n3139 & n4080 ) | ( ~n3975 & n4080 ) ;
  assign n9310 = n9309 ^ n9308 ^ 1'b0 ;
  assign n9311 = n2363 | n9310 ;
  assign n9312 = ( ~n1333 & n2734 ) | ( ~n1333 & n8073 ) | ( n2734 & n8073 ) ;
  assign n9313 = n9312 ^ n4088 ^ 1'b0 ;
  assign n9320 = x32 & n2563 ;
  assign n9321 = ~n5032 & n9320 ;
  assign n9319 = n698 & ~n2785 ;
  assign n9322 = n9321 ^ n9319 ^ 1'b0 ;
  assign n9317 = n2803 ^ n2330 ^ n2281 ;
  assign n9318 = n7895 | n9317 ;
  assign n9323 = n9322 ^ n9318 ^ 1'b0 ;
  assign n9314 = ( n3119 & n3456 ) | ( n3119 & ~n6864 ) | ( n3456 & ~n6864 ) ;
  assign n9315 = ( n1643 & n2065 ) | ( n1643 & ~n9314 ) | ( n2065 & ~n9314 ) ;
  assign n9316 = ( ~n270 & n5998 ) | ( ~n270 & n9315 ) | ( n5998 & n9315 ) ;
  assign n9324 = n9323 ^ n9316 ^ n7218 ;
  assign n9325 = n6162 ^ n4427 ^ n1253 ;
  assign n9326 = x117 | n1567 ;
  assign n9327 = n9326 ^ n2087 ^ 1'b0 ;
  assign n9328 = n7588 ^ n1676 ^ 1'b0 ;
  assign n9329 = n2427 | n9328 ;
  assign n9330 = n9329 ^ n6153 ^ 1'b0 ;
  assign n9331 = n9330 ^ n7216 ^ n2338 ;
  assign n9332 = ( n1935 & ~n9327 ) | ( n1935 & n9331 ) | ( ~n9327 & n9331 ) ;
  assign n9333 = n4438 ^ n3295 ^ n548 ;
  assign n9334 = n667 & ~n8736 ;
  assign n9337 = n4764 ^ n4197 ^ 1'b0 ;
  assign n9338 = n9337 ^ n3269 ^ n2029 ;
  assign n9335 = ( n2545 & n5516 ) | ( n2545 & n7625 ) | ( n5516 & n7625 ) ;
  assign n9336 = n5140 & n9335 ;
  assign n9339 = n9338 ^ n9336 ^ 1'b0 ;
  assign n9340 = n8630 ^ n5522 ^ n5507 ;
  assign n9341 = n2219 & ~n5734 ;
  assign n9342 = n9341 ^ n6140 ^ 1'b0 ;
  assign n9343 = ~n4967 & n9342 ;
  assign n9344 = n5685 & n9343 ;
  assign n9345 = n5727 & n8135 ;
  assign n9346 = ~n4116 & n8989 ;
  assign n9347 = ( n1515 & n3117 ) | ( n1515 & ~n9346 ) | ( n3117 & ~n9346 ) ;
  assign n9348 = n7398 ^ n4025 ^ 1'b0 ;
  assign n9349 = ( ~n1874 & n3601 ) | ( ~n1874 & n6352 ) | ( n3601 & n6352 ) ;
  assign n9350 = n9349 ^ n6781 ^ n4325 ;
  assign n9351 = n175 & ~n2470 ;
  assign n9352 = n9351 ^ n569 ^ 1'b0 ;
  assign n9353 = n9352 ^ n5177 ^ 1'b0 ;
  assign n9354 = ( n3227 & n4785 ) | ( n3227 & n6230 ) | ( n4785 & n6230 ) ;
  assign n9355 = n4152 ^ n410 ^ 1'b0 ;
  assign n9356 = n9355 ^ n3529 ^ 1'b0 ;
  assign n9357 = n9354 | n9356 ;
  assign n9358 = ( n2794 & ~n5504 ) | ( n2794 & n5581 ) | ( ~n5504 & n5581 ) ;
  assign n9363 = n4911 ^ n4007 ^ 1'b0 ;
  assign n9361 = ( n1260 & n1877 ) | ( n1260 & n5444 ) | ( n1877 & n5444 ) ;
  assign n9362 = n9361 ^ n4539 ^ n983 ;
  assign n9364 = n9363 ^ n9362 ^ n7260 ;
  assign n9359 = n8174 ^ n7690 ^ 1'b0 ;
  assign n9360 = n9359 ^ n4378 ^ n2622 ;
  assign n9365 = n9364 ^ n9360 ^ 1'b0 ;
  assign n9366 = n2707 & n9365 ;
  assign n9367 = n785 & n4417 ;
  assign n9368 = n9367 ^ n600 ^ 1'b0 ;
  assign n9369 = n6221 & ~n9368 ;
  assign n9370 = n9369 ^ n7688 ^ n3568 ;
  assign n9371 = n4666 & n9370 ;
  assign n9372 = n9371 ^ n1036 ^ 1'b0 ;
  assign n9373 = n8433 ^ x17 ^ 1'b0 ;
  assign n9374 = n2545 | n9373 ;
  assign n9375 = n9374 ^ n3164 ^ n820 ;
  assign n9376 = ~n5864 & n8011 ;
  assign n9377 = n2605 & n9376 ;
  assign n9378 = n5880 ^ n3721 ^ 1'b0 ;
  assign n9379 = ~n1902 & n7765 ;
  assign n9380 = n5054 ^ n3795 ^ n1382 ;
  assign n9381 = n9380 ^ n8086 ^ n1418 ;
  assign n9382 = n1404 ^ n453 ^ 1'b0 ;
  assign n9383 = n4520 & n8970 ;
  assign n9384 = n9382 & n9383 ;
  assign n9385 = n367 & n637 ;
  assign n9388 = n2393 ^ n1062 ^ n357 ;
  assign n9389 = n9388 ^ n2972 ^ x67 ;
  assign n9390 = n6971 & n9389 ;
  assign n9391 = n9390 ^ n3144 ^ 1'b0 ;
  assign n9392 = ( ~n300 & n1663 ) | ( ~n300 & n9391 ) | ( n1663 & n9391 ) ;
  assign n9386 = ( n1045 & n1600 ) | ( n1045 & ~n2443 ) | ( n1600 & ~n2443 ) ;
  assign n9387 = n9280 & ~n9386 ;
  assign n9393 = n9392 ^ n9387 ^ 1'b0 ;
  assign n9394 = n9393 ^ n6838 ^ 1'b0 ;
  assign n9395 = n1518 ^ x100 ^ 1'b0 ;
  assign n9396 = n3397 & ~n6819 ;
  assign n9397 = n9395 & n9396 ;
  assign n9398 = n7149 ^ n2485 ^ n1746 ;
  assign n9399 = ( n5777 & n6959 ) | ( n5777 & ~n9398 ) | ( n6959 & ~n9398 ) ;
  assign n9403 = n6337 ^ n2555 ^ 1'b0 ;
  assign n9404 = n8029 & ~n9403 ;
  assign n9405 = n9404 ^ n3330 ^ n1986 ;
  assign n9406 = n7090 & ~n9405 ;
  assign n9407 = n9406 ^ n2469 ^ 1'b0 ;
  assign n9401 = ~n2317 & n4633 ;
  assign n9402 = n2535 & n9401 ;
  assign n9400 = n2620 | n6368 ;
  assign n9408 = n9407 ^ n9402 ^ n9400 ;
  assign n9409 = ( n1579 & n2921 ) | ( n1579 & ~n3735 ) | ( n2921 & ~n3735 ) ;
  assign n9410 = n9409 ^ n3083 ^ 1'b0 ;
  assign n9411 = n9408 & ~n9410 ;
  assign n9413 = ( n199 & n6898 ) | ( n199 & n8630 ) | ( n6898 & n8630 ) ;
  assign n9412 = n3726 ^ n2700 ^ 1'b0 ;
  assign n9414 = n9413 ^ n9412 ^ n7538 ;
  assign n9415 = n1318 | n6610 ;
  assign n9416 = n9415 ^ n1977 ^ 1'b0 ;
  assign n9417 = n9416 ^ n4081 ^ n308 ;
  assign n9418 = ( n7710 & n8446 ) | ( n7710 & ~n9413 ) | ( n8446 & ~n9413 ) ;
  assign n9419 = ( ~n1569 & n4529 ) | ( ~n1569 & n6181 ) | ( n4529 & n6181 ) ;
  assign n9420 = ( n285 & n1570 ) | ( n285 & n5667 ) | ( n1570 & n5667 ) ;
  assign n9421 = ( ~n2832 & n3242 ) | ( ~n2832 & n9420 ) | ( n3242 & n9420 ) ;
  assign n9422 = n9421 ^ n1298 ^ n1159 ;
  assign n9423 = n4190 & n4903 ;
  assign n9424 = ( n1681 & n5361 ) | ( n1681 & ~n9423 ) | ( n5361 & ~n9423 ) ;
  assign n9425 = n9422 & n9424 ;
  assign n9426 = ( n1165 & n5562 ) | ( n1165 & n9425 ) | ( n5562 & n9425 ) ;
  assign n9427 = ( n4545 & ~n9419 ) | ( n4545 & n9426 ) | ( ~n9419 & n9426 ) ;
  assign n9428 = n9427 ^ n3037 ^ n2839 ;
  assign n9430 = ( n2478 & n4816 ) | ( n2478 & n5296 ) | ( n4816 & n5296 ) ;
  assign n9429 = n5703 & ~n8341 ;
  assign n9431 = n9430 ^ n9429 ^ 1'b0 ;
  assign n9432 = ( n2798 & ~n7320 ) | ( n2798 & n9431 ) | ( ~n7320 & n9431 ) ;
  assign n9433 = n1052 | n1864 ;
  assign n9434 = n9433 ^ x46 ^ 1'b0 ;
  assign n9435 = ~n1416 & n2999 ;
  assign n9436 = ~n5610 & n9435 ;
  assign n9437 = n9434 & ~n9436 ;
  assign n9438 = n3642 & n9437 ;
  assign n9439 = ( n2741 & ~n5284 ) | ( n2741 & n5287 ) | ( ~n5284 & n5287 ) ;
  assign n9440 = n9439 ^ n4177 ^ n2907 ;
  assign n9441 = ( n2140 & n6533 ) | ( n2140 & n9440 ) | ( n6533 & n9440 ) ;
  assign n9442 = ( n131 & ~n1916 ) | ( n131 & n9441 ) | ( ~n1916 & n9441 ) ;
  assign n9449 = ( n234 & ~n3785 ) | ( n234 & n4736 ) | ( ~n3785 & n4736 ) ;
  assign n9450 = n9449 ^ n1810 ^ n1686 ;
  assign n9451 = n9450 ^ n7905 ^ 1'b0 ;
  assign n9446 = ( n979 & n2513 ) | ( n979 & n4081 ) | ( n2513 & n4081 ) ;
  assign n9443 = n3188 ^ n2632 ^ n247 ;
  assign n9444 = ( n3388 & ~n5813 ) | ( n3388 & n9443 ) | ( ~n5813 & n9443 ) ;
  assign n9445 = ( ~n1810 & n2209 ) | ( ~n1810 & n9444 ) | ( n2209 & n9444 ) ;
  assign n9447 = n9446 ^ n9445 ^ 1'b0 ;
  assign n9448 = n9447 ^ n891 ^ x24 ;
  assign n9452 = n9451 ^ n9448 ^ n7805 ;
  assign n9453 = ( n2863 & ~n3357 ) | ( n2863 & n9452 ) | ( ~n3357 & n9452 ) ;
  assign n9454 = n6629 ^ n920 ^ 1'b0 ;
  assign n9455 = n4858 & n9454 ;
  assign n9456 = n5541 ^ n2358 ^ 1'b0 ;
  assign n9457 = n3613 | n9456 ;
  assign n9458 = ( n2495 & n3866 ) | ( n2495 & n4735 ) | ( n3866 & n4735 ) ;
  assign n9459 = ( ~n3240 & n9457 ) | ( ~n3240 & n9458 ) | ( n9457 & n9458 ) ;
  assign n9460 = ( n1500 & ~n5556 ) | ( n1500 & n9459 ) | ( ~n5556 & n9459 ) ;
  assign n9461 = n9460 ^ n5177 ^ n4604 ;
  assign n9462 = n8475 ^ n846 ^ n233 ;
  assign n9463 = n831 & ~n5215 ;
  assign n9464 = ~n9462 & n9463 ;
  assign n9465 = ( n2617 & n9461 ) | ( n2617 & n9464 ) | ( n9461 & n9464 ) ;
  assign n9469 = n3725 ^ n1808 ^ 1'b0 ;
  assign n9470 = n4925 & ~n9469 ;
  assign n9467 = n3508 ^ n3275 ^ 1'b0 ;
  assign n9466 = ( n2557 & n3000 ) | ( n2557 & ~n4782 ) | ( n3000 & ~n4782 ) ;
  assign n9468 = n9467 ^ n9466 ^ n2188 ;
  assign n9471 = n9470 ^ n9468 ^ 1'b0 ;
  assign n9482 = ( n2757 & n3629 ) | ( n2757 & n6185 ) | ( n3629 & n6185 ) ;
  assign n9481 = n8057 ^ n5696 ^ 1'b0 ;
  assign n9472 = ( x66 & n2677 ) | ( x66 & ~n4298 ) | ( n2677 & ~n4298 ) ;
  assign n9473 = ( n7592 & n8810 ) | ( n7592 & ~n9472 ) | ( n8810 & ~n9472 ) ;
  assign n9474 = n600 & ~n3586 ;
  assign n9475 = n9474 ^ n8641 ^ 1'b0 ;
  assign n9476 = n1003 & ~n5849 ;
  assign n9477 = n4687 & n9476 ;
  assign n9478 = n9477 ^ n6477 ^ x13 ;
  assign n9479 = ( n2618 & n9475 ) | ( n2618 & ~n9478 ) | ( n9475 & ~n9478 ) ;
  assign n9480 = ( ~n3499 & n9473 ) | ( ~n3499 & n9479 ) | ( n9473 & n9479 ) ;
  assign n9483 = n9482 ^ n9481 ^ n9480 ;
  assign n9484 = ( n2140 & n7991 ) | ( n2140 & n9483 ) | ( n7991 & n9483 ) ;
  assign n9485 = ( n1809 & ~n9471 ) | ( n1809 & n9484 ) | ( ~n9471 & n9484 ) ;
  assign n9486 = ( n2348 & n2509 ) | ( n2348 & ~n2600 ) | ( n2509 & ~n2600 ) ;
  assign n9488 = ( n753 & n2765 ) | ( n753 & ~n4825 ) | ( n2765 & ~n4825 ) ;
  assign n9487 = ~n4581 & n5044 ;
  assign n9489 = n9488 ^ n9487 ^ 1'b0 ;
  assign n9490 = n9489 ^ n5027 ^ n1511 ;
  assign n9491 = ( n4272 & n9486 ) | ( n4272 & n9490 ) | ( n9486 & n9490 ) ;
  assign n9492 = n9147 ^ n1417 ^ 1'b0 ;
  assign n9493 = n787 & ~n9492 ;
  assign n9494 = n7023 & n9493 ;
  assign n9495 = ~n5648 & n9494 ;
  assign n9498 = n848 | n4359 ;
  assign n9496 = ( n439 & ~n464 ) | ( n439 & n7259 ) | ( ~n464 & n7259 ) ;
  assign n9497 = ( n453 & n6976 ) | ( n453 & n9496 ) | ( n6976 & n9496 ) ;
  assign n9499 = n9498 ^ n9497 ^ 1'b0 ;
  assign n9500 = ~n6635 & n9499 ;
  assign n9507 = n1485 ^ n988 ^ 1'b0 ;
  assign n9508 = n8390 & n9507 ;
  assign n9501 = n537 | n2013 ;
  assign n9502 = ( n1334 & n2955 ) | ( n1334 & ~n5718 ) | ( n2955 & ~n5718 ) ;
  assign n9503 = n7747 | n9502 ;
  assign n9504 = n9501 & ~n9503 ;
  assign n9505 = ( n5056 & n6581 ) | ( n5056 & n9504 ) | ( n6581 & n9504 ) ;
  assign n9506 = n9505 ^ n5411 ^ n1705 ;
  assign n9509 = n9508 ^ n9506 ^ n4349 ;
  assign n9510 = n2373 ^ n2140 ^ n1736 ;
  assign n9511 = n9510 ^ n6408 ^ n3698 ;
  assign n9512 = n1000 & n9511 ;
  assign n9513 = ~n1611 & n9512 ;
  assign n9514 = n708 | n5721 ;
  assign n9515 = n9513 & ~n9514 ;
  assign n9516 = n5199 ^ n1908 ^ 1'b0 ;
  assign n9517 = n8602 & ~n9516 ;
  assign n9518 = n248 & n9517 ;
  assign n9519 = ~n3098 & n3410 ;
  assign n9520 = n9519 ^ n9309 ^ n4591 ;
  assign n9524 = n1975 ^ n1371 ^ n970 ;
  assign n9523 = n2547 | n5523 ;
  assign n9525 = n9524 ^ n9523 ^ 1'b0 ;
  assign n9526 = ( ~n3658 & n8487 ) | ( ~n3658 & n9525 ) | ( n8487 & n9525 ) ;
  assign n9522 = n1306 & n4948 ;
  assign n9521 = n6058 & n8808 ;
  assign n9527 = n9526 ^ n9522 ^ n9521 ;
  assign n9528 = n5071 | n7492 ;
  assign n9529 = ( n3096 & ~n5650 ) | ( n3096 & n9528 ) | ( ~n5650 & n9528 ) ;
  assign n9530 = ( n218 & ~n4278 ) | ( n218 & n7234 ) | ( ~n4278 & n7234 ) ;
  assign n9531 = n2713 | n6713 ;
  assign n9532 = n4831 & ~n9531 ;
  assign n9533 = n4859 | n9532 ;
  assign n9534 = n415 & n2621 ;
  assign n9535 = n217 & n9534 ;
  assign n9536 = ~n5400 & n9535 ;
  assign n9537 = ( n2340 & n5523 ) | ( n2340 & ~n9536 ) | ( n5523 & ~n9536 ) ;
  assign n9538 = n9537 ^ n2236 ^ n1953 ;
  assign n9539 = n9538 ^ n3738 ^ n3460 ;
  assign n9540 = ( n9530 & ~n9533 ) | ( n9530 & n9539 ) | ( ~n9533 & n9539 ) ;
  assign n9541 = n9540 ^ n4687 ^ n2959 ;
  assign n9542 = ( n955 & ~n2706 ) | ( n955 & n4684 ) | ( ~n2706 & n4684 ) ;
  assign n9543 = n1171 & n3029 ;
  assign n9544 = ~n3541 & n9543 ;
  assign n9545 = ~n1228 & n1570 ;
  assign n9546 = n9544 & n9545 ;
  assign n9547 = ( n1092 & n9542 ) | ( n1092 & ~n9546 ) | ( n9542 & ~n9546 ) ;
  assign n9548 = n4227 ^ n3746 ^ 1'b0 ;
  assign n9549 = ~n3081 & n9548 ;
  assign n9550 = n8615 ^ n8298 ^ n2047 ;
  assign n9551 = ( n540 & ~n9179 ) | ( n540 & n9550 ) | ( ~n9179 & n9550 ) ;
  assign n9552 = ( n7056 & n9549 ) | ( n7056 & ~n9551 ) | ( n9549 & ~n9551 ) ;
  assign n9553 = ( ~n328 & n2425 ) | ( ~n328 & n4437 ) | ( n2425 & n4437 ) ;
  assign n9554 = n5558 & ~n9553 ;
  assign n9555 = n5632 ^ n472 ^ 1'b0 ;
  assign n9556 = n2681 & ~n9555 ;
  assign n9557 = n2140 & ~n9556 ;
  assign n9558 = ( n373 & n2243 ) | ( n373 & ~n4702 ) | ( n2243 & ~n4702 ) ;
  assign n9559 = n1110 & ~n3800 ;
  assign n9560 = ( n8715 & ~n9558 ) | ( n8715 & n9559 ) | ( ~n9558 & n9559 ) ;
  assign n9561 = ( n4896 & ~n5980 ) | ( n4896 & n9560 ) | ( ~n5980 & n9560 ) ;
  assign n9562 = n4804 ^ n3931 ^ n1416 ;
  assign n9563 = ~n3503 & n9562 ;
  assign n9564 = n9561 & n9563 ;
  assign n9568 = ~n282 & n2621 ;
  assign n9569 = ~n2091 & n9568 ;
  assign n9565 = n580 & n4739 ;
  assign n9566 = n3017 | n9565 ;
  assign n9567 = n8387 & ~n9566 ;
  assign n9570 = n9569 ^ n9567 ^ n5318 ;
  assign n9571 = n6499 & ~n7211 ;
  assign n9572 = n9571 ^ n7582 ^ 1'b0 ;
  assign n9573 = n2816 ^ n2373 ^ 1'b0 ;
  assign n9574 = n9573 ^ n8521 ^ n429 ;
  assign n9575 = ~n9572 & n9574 ;
  assign n9576 = ( n1207 & ~n3251 ) | ( n1207 & n4010 ) | ( ~n3251 & n4010 ) ;
  assign n9579 = n2242 ^ n2144 ^ n950 ;
  assign n9577 = n6186 ^ n6038 ^ 1'b0 ;
  assign n9578 = n489 & n9577 ;
  assign n9580 = n9579 ^ n9578 ^ n3651 ;
  assign n9581 = n4843 & n9409 ;
  assign n9585 = ~n335 & n2402 ;
  assign n9586 = ~n2467 & n9585 ;
  assign n9587 = ( n3364 & ~n6037 ) | ( n3364 & n9586 ) | ( ~n6037 & n9586 ) ;
  assign n9583 = n4168 & n7337 ;
  assign n9584 = n9583 ^ n3898 ^ 1'b0 ;
  assign n9582 = n4371 ^ n3815 ^ n2351 ;
  assign n9588 = n9587 ^ n9584 ^ n9582 ;
  assign n9589 = n9581 | n9588 ;
  assign n9594 = n2785 ^ n1428 ^ 1'b0 ;
  assign n9595 = n2065 & n9594 ;
  assign n9593 = n5333 ^ n3888 ^ n661 ;
  assign n9591 = ( ~n2145 & n4795 ) | ( ~n2145 & n4846 ) | ( n4795 & n4846 ) ;
  assign n9590 = ( n3677 & n4159 ) | ( n3677 & n9140 ) | ( n4159 & n9140 ) ;
  assign n9592 = n9591 ^ n9590 ^ n608 ;
  assign n9596 = n9595 ^ n9593 ^ n9592 ;
  assign n9597 = n2195 ^ n2139 ^ n869 ;
  assign n9598 = n9597 ^ n2358 ^ 1'b0 ;
  assign n9599 = ( n1119 & n9037 ) | ( n1119 & n9598 ) | ( n9037 & n9598 ) ;
  assign n9600 = n9423 ^ n4464 ^ n3557 ;
  assign n9601 = ~n3666 & n7141 ;
  assign n9602 = ~n9600 & n9601 ;
  assign n9603 = ( ~n1998 & n9599 ) | ( ~n1998 & n9602 ) | ( n9599 & n9602 ) ;
  assign n9604 = ( n2637 & n3887 ) | ( n2637 & ~n6113 ) | ( n3887 & ~n6113 ) ;
  assign n9605 = ~n9372 & n9604 ;
  assign n9606 = n9605 ^ n8182 ^ 1'b0 ;
  assign n9607 = ( n541 & ~n2066 ) | ( n541 & n3586 ) | ( ~n2066 & n3586 ) ;
  assign n9608 = n4855 ^ n3814 ^ n2713 ;
  assign n9609 = n9608 ^ n378 ^ 1'b0 ;
  assign n9610 = n9607 & ~n9609 ;
  assign n9615 = n6054 ^ n4046 ^ n2467 ;
  assign n9611 = n3568 ^ n2618 ^ n2383 ;
  assign n9612 = ( ~n4130 & n8028 ) | ( ~n4130 & n9611 ) | ( n8028 & n9611 ) ;
  assign n9613 = n9612 ^ n4607 ^ 1'b0 ;
  assign n9614 = ( ~n4870 & n9544 ) | ( ~n4870 & n9613 ) | ( n9544 & n9613 ) ;
  assign n9616 = n9615 ^ n9614 ^ 1'b0 ;
  assign n9617 = ( n357 & n389 ) | ( n357 & n1300 ) | ( n389 & n1300 ) ;
  assign n9618 = n9617 ^ n4366 ^ n841 ;
  assign n9619 = ( n2509 & ~n2791 ) | ( n2509 & n3513 ) | ( ~n2791 & n3513 ) ;
  assign n9620 = n9619 ^ n4796 ^ n2356 ;
  assign n9621 = n9620 ^ n3188 ^ 1'b0 ;
  assign n9622 = n9618 & n9621 ;
  assign n9623 = n1082 | n1400 ;
  assign n9624 = n1611 | n9623 ;
  assign n9625 = ~n6072 & n9624 ;
  assign n9626 = n9625 ^ n6653 ^ n5612 ;
  assign n9627 = n9622 & ~n9626 ;
  assign n9628 = n8460 & n9627 ;
  assign n9629 = n3056 & n3391 ;
  assign n9630 = n9629 ^ n5381 ^ 1'b0 ;
  assign n9632 = ( ~n3433 & n3582 ) | ( ~n3433 & n7588 ) | ( n3582 & n7588 ) ;
  assign n9631 = n1966 & ~n5073 ;
  assign n9633 = n9632 ^ n9631 ^ 1'b0 ;
  assign n9636 = n2963 ^ n2113 ^ 1'b0 ;
  assign n9634 = n1967 & n6045 ;
  assign n9635 = n2749 & n9634 ;
  assign n9637 = n9636 ^ n9635 ^ n7485 ;
  assign n9638 = n9637 ^ n8541 ^ 1'b0 ;
  assign n9639 = ( n9630 & n9633 ) | ( n9630 & ~n9638 ) | ( n9633 & ~n9638 ) ;
  assign n9640 = n3698 | n4375 ;
  assign n9641 = ( n1211 & n2703 ) | ( n1211 & ~n4184 ) | ( n2703 & ~n4184 ) ;
  assign n9642 = ( ~n1315 & n9640 ) | ( ~n1315 & n9641 ) | ( n9640 & n9641 ) ;
  assign n9643 = n9642 ^ n1218 ^ 1'b0 ;
  assign n9644 = n8996 & ~n9643 ;
  assign n9645 = n9295 ^ n540 ^ x122 ;
  assign n9647 = ~n1919 & n4510 ;
  assign n9646 = ~n4956 & n8624 ;
  assign n9648 = n9647 ^ n9646 ^ 1'b0 ;
  assign n9649 = n8787 & n9648 ;
  assign n9650 = n9649 ^ n2902 ^ 1'b0 ;
  assign n9651 = ( ~n2139 & n2293 ) | ( ~n2139 & n4425 ) | ( n2293 & n4425 ) ;
  assign n9652 = ( n7703 & n8487 ) | ( n7703 & ~n9651 ) | ( n8487 & ~n9651 ) ;
  assign n9653 = n1434 & ~n9652 ;
  assign n9654 = n9653 ^ n2846 ^ 1'b0 ;
  assign n9655 = n1705 | n9654 ;
  assign n9656 = n9510 ^ n4581 ^ n724 ;
  assign n9657 = n4973 ^ n214 ^ 1'b0 ;
  assign n9658 = ( n1119 & n6002 ) | ( n1119 & n9657 ) | ( n6002 & n9657 ) ;
  assign n9659 = n9658 ^ n5545 ^ n2335 ;
  assign n9660 = n1809 & n3474 ;
  assign n9661 = n9660 ^ n2708 ^ 1'b0 ;
  assign n9662 = ( n1771 & n3880 ) | ( n1771 & ~n9661 ) | ( n3880 & ~n9661 ) ;
  assign n9663 = ( n901 & n9659 ) | ( n901 & ~n9662 ) | ( n9659 & ~n9662 ) ;
  assign n9665 = ( n184 & ~n2827 ) | ( n184 & n6781 ) | ( ~n2827 & n6781 ) ;
  assign n9664 = n8829 ^ n4022 ^ n962 ;
  assign n9666 = n9665 ^ n9664 ^ n7896 ;
  assign n9667 = ( n6749 & n6883 ) | ( n6749 & n9666 ) | ( n6883 & n9666 ) ;
  assign n9668 = ( n2308 & n3424 ) | ( n2308 & ~n8627 ) | ( n3424 & ~n8627 ) ;
  assign n9669 = n8058 ^ n3225 ^ n2554 ;
  assign n9670 = ( n408 & n6013 ) | ( n408 & n7259 ) | ( n6013 & n7259 ) ;
  assign n9672 = n1487 ^ n1430 ^ 1'b0 ;
  assign n9671 = n3768 ^ n2817 ^ n379 ;
  assign n9673 = n9672 ^ n9671 ^ 1'b0 ;
  assign n9674 = n9670 | n9673 ;
  assign n9675 = n2636 & ~n9674 ;
  assign n9676 = ( n638 & n1490 ) | ( n638 & ~n2876 ) | ( n1490 & ~n2876 ) ;
  assign n9677 = ( n2642 & n3821 ) | ( n2642 & n8295 ) | ( n3821 & n8295 ) ;
  assign n9678 = n9677 ^ n5525 ^ n1967 ;
  assign n9679 = ( n1478 & n9676 ) | ( n1478 & n9678 ) | ( n9676 & n9678 ) ;
  assign n9680 = ( n2053 & n4746 ) | ( n2053 & n8917 ) | ( n4746 & n8917 ) ;
  assign n9681 = n8843 & n9680 ;
  assign n9689 = n353 & n8813 ;
  assign n9690 = n9689 ^ n3740 ^ n129 ;
  assign n9691 = n9690 ^ n8478 ^ n3223 ;
  assign n9684 = n2381 | n3443 ;
  assign n9685 = n1176 & ~n9684 ;
  assign n9686 = n9685 ^ n1403 ^ 1'b0 ;
  assign n9687 = n2235 & n9686 ;
  assign n9682 = n3626 ^ n1393 ^ n1194 ;
  assign n9683 = n8620 & ~n9682 ;
  assign n9688 = n9687 ^ n9683 ^ 1'b0 ;
  assign n9692 = n9691 ^ n9688 ^ n6246 ;
  assign n9693 = ~n826 & n1704 ;
  assign n9694 = ( n4124 & ~n7090 ) | ( n4124 & n7577 ) | ( ~n7090 & n7577 ) ;
  assign n9695 = ( n3926 & ~n9693 ) | ( n3926 & n9694 ) | ( ~n9693 & n9694 ) ;
  assign n9696 = n3610 ^ x22 ^ 1'b0 ;
  assign n9697 = n9696 ^ n1559 ^ 1'b0 ;
  assign n9698 = ~n3580 & n9697 ;
  assign n9699 = ( n598 & n2865 ) | ( n598 & n3093 ) | ( n2865 & n3093 ) ;
  assign n9700 = ( n3914 & n9361 ) | ( n3914 & ~n9699 ) | ( n9361 & ~n9699 ) ;
  assign n9701 = ( n924 & ~n933 ) | ( n924 & n1335 ) | ( ~n933 & n1335 ) ;
  assign n9702 = n9701 ^ n2882 ^ n976 ;
  assign n9703 = n9702 ^ n4967 ^ n766 ;
  assign n9704 = ~n4910 & n9703 ;
  assign n9705 = n9704 ^ n7412 ^ 1'b0 ;
  assign n9707 = n7735 | n8444 ;
  assign n9708 = n2949 & ~n9707 ;
  assign n9706 = n3900 | n5068 ;
  assign n9709 = n9708 ^ n9706 ^ 1'b0 ;
  assign n9710 = n1984 & ~n9709 ;
  assign n9711 = n9710 ^ n3267 ^ 1'b0 ;
  assign n9712 = ~n9705 & n9711 ;
  assign n9717 = n9223 ^ n8623 ^ n6261 ;
  assign n9713 = n1457 & n1891 ;
  assign n9714 = n3836 & ~n9713 ;
  assign n9715 = n3807 & n9714 ;
  assign n9716 = ( n6933 & n7704 ) | ( n6933 & n9715 ) | ( n7704 & n9715 ) ;
  assign n9718 = n9717 ^ n9716 ^ n2147 ;
  assign n9719 = n7231 ^ n5523 ^ n2625 ;
  assign n9720 = n9719 ^ n7335 ^ 1'b0 ;
  assign n9721 = n3008 & ~n9720 ;
  assign n9726 = ( n901 & ~n3467 ) | ( n901 & n4090 ) | ( ~n3467 & n4090 ) ;
  assign n9723 = ( ~n1644 & n2169 ) | ( ~n1644 & n7900 ) | ( n2169 & n7900 ) ;
  assign n9722 = ( n1045 & n2473 ) | ( n1045 & ~n3145 ) | ( n2473 & ~n3145 ) ;
  assign n9724 = n9723 ^ n9722 ^ 1'b0 ;
  assign n9725 = n9149 | n9724 ;
  assign n9727 = n9726 ^ n9725 ^ n8624 ;
  assign n9729 = ( n861 & n4247 ) | ( n861 & ~n4650 ) | ( n4247 & ~n4650 ) ;
  assign n9728 = n8738 ^ n4886 ^ n583 ;
  assign n9730 = n9729 ^ n9728 ^ n2426 ;
  assign n9731 = ~n7634 & n9730 ;
  assign n9732 = n9731 ^ n4055 ^ 1'b0 ;
  assign n9733 = ( ~n6892 & n9727 ) | ( ~n6892 & n9732 ) | ( n9727 & n9732 ) ;
  assign n9734 = n1977 & ~n6489 ;
  assign n9735 = ( ~x0 & n3525 ) | ( ~x0 & n9734 ) | ( n3525 & n9734 ) ;
  assign n9736 = n7407 ^ n1084 ^ n453 ;
  assign n9737 = n2213 | n9736 ;
  assign n9738 = n7701 | n9737 ;
  assign n9739 = ( n1912 & n2311 ) | ( n1912 & n9738 ) | ( n2311 & n9738 ) ;
  assign n9740 = n9739 ^ n4345 ^ 1'b0 ;
  assign n9741 = ( ~n4188 & n4264 ) | ( ~n4188 & n6316 ) | ( n4264 & n6316 ) ;
  assign n9742 = ( n3522 & n5790 ) | ( n3522 & ~n9741 ) | ( n5790 & ~n9741 ) ;
  assign n9743 = ( n5613 & ~n8292 ) | ( n5613 & n9742 ) | ( ~n8292 & n9742 ) ;
  assign n9746 = ( n2105 & n2126 ) | ( n2105 & n2542 ) | ( n2126 & n2542 ) ;
  assign n9744 = ~n2145 & n4836 ;
  assign n9745 = n7974 & ~n9744 ;
  assign n9747 = n9746 ^ n9745 ^ 1'b0 ;
  assign n9751 = n5078 ^ n3893 ^ 1'b0 ;
  assign n9752 = n9751 ^ n4234 ^ n1112 ;
  assign n9753 = n9752 ^ n3929 ^ 1'b0 ;
  assign n9748 = ( n830 & ~n1443 ) | ( n830 & n3251 ) | ( ~n1443 & n3251 ) ;
  assign n9749 = n7546 ^ n1460 ^ n937 ;
  assign n9750 = n9748 | n9749 ;
  assign n9754 = n9753 ^ n9750 ^ 1'b0 ;
  assign n9755 = n7575 ^ n6123 ^ 1'b0 ;
  assign n9756 = ~n1183 & n9755 ;
  assign n9757 = n9756 ^ n2243 ^ n1032 ;
  assign n9758 = n9757 ^ n3174 ^ n643 ;
  assign n9759 = n9758 ^ n4292 ^ x99 ;
  assign n9760 = ( ~n758 & n1088 ) | ( ~n758 & n8565 ) | ( n1088 & n8565 ) ;
  assign n9761 = n1172 & n9760 ;
  assign n9762 = n6494 ^ n2606 ^ n916 ;
  assign n9763 = n9762 ^ n9060 ^ 1'b0 ;
  assign n9769 = ( n1388 & n1581 ) | ( n1388 & ~n1625 ) | ( n1581 & ~n1625 ) ;
  assign n9770 = ~n8543 & n9769 ;
  assign n9771 = n2928 & n9770 ;
  assign n9768 = n8235 ^ n3619 ^ n2039 ;
  assign n9764 = n5611 ^ n4164 ^ 1'b0 ;
  assign n9765 = n2954 | n9764 ;
  assign n9766 = ( n1487 & n3675 ) | ( n1487 & ~n9708 ) | ( n3675 & ~n9708 ) ;
  assign n9767 = ( n3267 & n9765 ) | ( n3267 & n9766 ) | ( n9765 & n9766 ) ;
  assign n9772 = n9771 ^ n9768 ^ n9767 ;
  assign n9773 = n9741 ^ n6353 ^ n767 ;
  assign n9774 = n9773 ^ n8343 ^ 1'b0 ;
  assign n9775 = n3473 ^ n2279 ^ 1'b0 ;
  assign n9776 = n4031 & n9775 ;
  assign n9777 = n9776 ^ n6105 ^ n335 ;
  assign n9780 = ( n1054 & n1086 ) | ( n1054 & ~n1652 ) | ( n1086 & ~n1652 ) ;
  assign n9781 = n3209 ^ n1534 ^ 1'b0 ;
  assign n9782 = ~n9780 & n9781 ;
  assign n9778 = n4692 ^ n655 ^ 1'b0 ;
  assign n9779 = x103 & ~n9778 ;
  assign n9783 = n9782 ^ n9779 ^ 1'b0 ;
  assign n9784 = ~n5049 & n9783 ;
  assign n9787 = n4170 ^ n921 ^ n604 ;
  assign n9788 = ( n1299 & n1557 ) | ( n1299 & n9787 ) | ( n1557 & n9787 ) ;
  assign n9785 = x92 & ~n7476 ;
  assign n9786 = ~n4072 & n9785 ;
  assign n9789 = n9788 ^ n9786 ^ n2570 ;
  assign n9790 = n1233 ^ n271 ^ 1'b0 ;
  assign n9791 = n9790 ^ n5599 ^ 1'b0 ;
  assign n9792 = n7963 & n9791 ;
  assign n9793 = ( n3304 & ~n9207 ) | ( n3304 & n9792 ) | ( ~n9207 & n9792 ) ;
  assign n9794 = n6956 ^ n4155 ^ n605 ;
  assign n9795 = n9793 & n9794 ;
  assign n9796 = n9702 ^ n7815 ^ n1085 ;
  assign n9797 = ( n4282 & n5552 ) | ( n4282 & n5578 ) | ( n5552 & n5578 ) ;
  assign n9798 = ( n131 & n4145 ) | ( n131 & n9797 ) | ( n4145 & n9797 ) ;
  assign n9799 = ( n1532 & n2933 ) | ( n1532 & ~n6662 ) | ( n2933 & ~n6662 ) ;
  assign n9800 = n3910 ^ n1359 ^ n1294 ;
  assign n9801 = n9585 & n9800 ;
  assign n9802 = n2729 & n3490 ;
  assign n9803 = n9802 ^ n2483 ^ n766 ;
  assign n9804 = n9803 ^ n4416 ^ n330 ;
  assign n9805 = n5522 ^ n2419 ^ n2116 ;
  assign n9806 = n9805 ^ n4278 ^ n822 ;
  assign n9807 = n471 & ~n2712 ;
  assign n9808 = n9807 ^ n5736 ^ 1'b0 ;
  assign n9809 = n9808 ^ n9109 ^ n5025 ;
  assign n9810 = ( n561 & ~n9806 ) | ( n561 & n9809 ) | ( ~n9806 & n9809 ) ;
  assign n9811 = n5616 ^ n1271 ^ n632 ;
  assign n9812 = n2184 & n5150 ;
  assign n9813 = n9812 ^ n6938 ^ n2912 ;
  assign n9814 = n9813 ^ n9137 ^ 1'b0 ;
  assign n9815 = n9811 | n9814 ;
  assign n9816 = n4813 | n9815 ;
  assign n9817 = n8295 ^ n4965 ^ 1'b0 ;
  assign n9818 = ( n2118 & ~n7954 ) | ( n2118 & n9817 ) | ( ~n7954 & n9817 ) ;
  assign n9819 = n7706 ^ n5331 ^ 1'b0 ;
  assign n9820 = n7407 & ~n9819 ;
  assign n9821 = n4581 | n9133 ;
  assign n9822 = ( ~n3113 & n5451 ) | ( ~n3113 & n9821 ) | ( n5451 & n9821 ) ;
  assign n9823 = ( ~n2406 & n5153 ) | ( ~n2406 & n5715 ) | ( n5153 & n5715 ) ;
  assign n9824 = ( ~n5148 & n6189 ) | ( ~n5148 & n8086 ) | ( n6189 & n8086 ) ;
  assign n9825 = n973 & ~n9824 ;
  assign n9826 = ~n3110 & n9050 ;
  assign n9827 = n9826 ^ n3183 ^ 1'b0 ;
  assign n9828 = n9096 | n9827 ;
  assign n9829 = n6226 ^ n2366 ^ n1276 ;
  assign n9830 = n9829 ^ n865 ^ 1'b0 ;
  assign n9831 = n7231 | n9830 ;
  assign n9832 = n6347 ^ n1377 ^ n1012 ;
  assign n9833 = ( ~n1994 & n2405 ) | ( ~n1994 & n2581 ) | ( n2405 & n2581 ) ;
  assign n9834 = n2002 | n3852 ;
  assign n9835 = ~n9833 & n9834 ;
  assign n9836 = n9832 | n9835 ;
  assign n9837 = n9831 & ~n9836 ;
  assign n9838 = ( n900 & n1484 ) | ( n900 & n5635 ) | ( n1484 & n5635 ) ;
  assign n9839 = ( ~n6357 & n7996 ) | ( ~n6357 & n9838 ) | ( n7996 & n9838 ) ;
  assign n9840 = n5305 ^ n3038 ^ n1910 ;
  assign n9841 = n8662 ^ n4735 ^ n456 ;
  assign n9842 = ( ~n7515 & n9840 ) | ( ~n7515 & n9841 ) | ( n9840 & n9841 ) ;
  assign n9843 = ( n7094 & n9839 ) | ( n7094 & n9842 ) | ( n9839 & n9842 ) ;
  assign n9844 = n8890 ^ n3316 ^ n2554 ;
  assign n9845 = n9844 ^ n3323 ^ 1'b0 ;
  assign n9846 = ( n7155 & ~n8215 ) | ( n7155 & n9845 ) | ( ~n8215 & n9845 ) ;
  assign n9847 = ( n2372 & ~n2599 ) | ( n2372 & n4447 ) | ( ~n2599 & n4447 ) ;
  assign n9848 = n2066 ^ n850 ^ 1'b0 ;
  assign n9849 = n1308 ^ n890 ^ 1'b0 ;
  assign n9850 = n6414 | n9849 ;
  assign n9851 = ( ~n4147 & n9848 ) | ( ~n4147 & n9850 ) | ( n9848 & n9850 ) ;
  assign n9852 = ( n1994 & n6480 ) | ( n1994 & ~n9851 ) | ( n6480 & ~n9851 ) ;
  assign n9853 = n6043 ^ n4878 ^ 1'b0 ;
  assign n9854 = ~n670 & n4520 ;
  assign n9855 = ( n3885 & ~n5095 ) | ( n3885 & n9854 ) | ( ~n5095 & n9854 ) ;
  assign n9856 = ( n1532 & n6164 ) | ( n1532 & n9855 ) | ( n6164 & n9855 ) ;
  assign n9857 = n9853 & n9856 ;
  assign n9858 = ~n4155 & n9857 ;
  assign n9859 = n5122 & ~n6033 ;
  assign n9860 = n9859 ^ n1605 ^ 1'b0 ;
  assign n9861 = n9860 ^ n9073 ^ n2712 ;
  assign n9863 = n3208 ^ n1677 ^ 1'b0 ;
  assign n9862 = n6068 & ~n6133 ;
  assign n9864 = n9863 ^ n9862 ^ 1'b0 ;
  assign n9870 = n805 | n1790 ;
  assign n9871 = n1055 | n9870 ;
  assign n9872 = ( n649 & n4078 ) | ( n649 & n9840 ) | ( n4078 & n9840 ) ;
  assign n9873 = ( ~n9449 & n9871 ) | ( ~n9449 & n9872 ) | ( n9871 & n9872 ) ;
  assign n9869 = n3496 ^ n2539 ^ 1'b0 ;
  assign n9874 = n9873 ^ n9869 ^ n1856 ;
  assign n9865 = n6288 ^ n1672 ^ n518 ;
  assign n9866 = ~n701 & n9865 ;
  assign n9867 = n9866 ^ n4742 ^ 1'b0 ;
  assign n9868 = n3812 | n9867 ;
  assign n9875 = n9874 ^ n9868 ^ 1'b0 ;
  assign n9876 = n8240 ^ n6200 ^ n2474 ;
  assign n9877 = n7052 ^ n6528 ^ 1'b0 ;
  assign n9878 = ~n9876 & n9877 ;
  assign n9879 = n5054 & ~n9626 ;
  assign n9880 = ~n9075 & n9879 ;
  assign n9881 = ( ~n1877 & n8162 ) | ( ~n1877 & n9880 ) | ( n8162 & n9880 ) ;
  assign n9882 = n9131 ^ n8136 ^ x38 ;
  assign n9887 = n7430 ^ n3825 ^ n1511 ;
  assign n9883 = n2828 ^ n2393 ^ n1122 ;
  assign n9884 = n9883 ^ n3764 ^ 1'b0 ;
  assign n9885 = n2270 & n9884 ;
  assign n9886 = n9885 ^ n4966 ^ n1436 ;
  assign n9888 = n9887 ^ n9886 ^ n1594 ;
  assign n9891 = n2239 ^ n663 ^ 1'b0 ;
  assign n9892 = n593 & ~n9891 ;
  assign n9889 = n231 | n1445 ;
  assign n9890 = n9889 ^ n3422 ^ 1'b0 ;
  assign n9893 = n9892 ^ n9890 ^ n2794 ;
  assign n9894 = ~n2437 & n3824 ;
  assign n9895 = ( ~n870 & n2450 ) | ( ~n870 & n9894 ) | ( n2450 & n9894 ) ;
  assign n9896 = n4633 ^ n3009 ^ n1605 ;
  assign n9897 = n9896 ^ n4636 ^ n1043 ;
  assign n9898 = n332 & n8241 ;
  assign n9899 = ~n9897 & n9898 ;
  assign n9900 = ~n7545 & n9899 ;
  assign n9901 = n1485 & ~n9900 ;
  assign n9902 = n9901 ^ n424 ^ 1'b0 ;
  assign n9903 = n9902 ^ n3187 ^ 1'b0 ;
  assign n9904 = n4318 | n9903 ;
  assign n9909 = ( x55 & n1479 ) | ( x55 & n3523 ) | ( n1479 & n3523 ) ;
  assign n9906 = ( n1741 & n2953 ) | ( n1741 & n5711 ) | ( n2953 & n5711 ) ;
  assign n9907 = n2302 | n2345 ;
  assign n9908 = ( ~n4619 & n9906 ) | ( ~n4619 & n9907 ) | ( n9906 & n9907 ) ;
  assign n9905 = n4817 ^ n4021 ^ n2493 ;
  assign n9910 = n9909 ^ n9908 ^ n9905 ;
  assign n9911 = ( n944 & ~n3955 ) | ( n944 & n8749 ) | ( ~n3955 & n8749 ) ;
  assign n9912 = n3275 & n7413 ;
  assign n9913 = ~n9911 & n9912 ;
  assign n9914 = ( n5622 & ~n7952 ) | ( n5622 & n9913 ) | ( ~n7952 & n9913 ) ;
  assign n9915 = n1311 | n4948 ;
  assign n9916 = n9915 ^ n2774 ^ 1'b0 ;
  assign n9917 = n4352 ^ n2168 ^ n2063 ;
  assign n9918 = n662 | n1550 ;
  assign n9919 = n5397 & ~n9918 ;
  assign n9920 = n9919 ^ n9120 ^ 1'b0 ;
  assign n9921 = ~n9917 & n9920 ;
  assign n9922 = n9921 ^ n1021 ^ 1'b0 ;
  assign n9923 = x1 & n9922 ;
  assign n9924 = n1554 ^ n647 ^ 1'b0 ;
  assign n9925 = ( ~n1444 & n1799 ) | ( ~n1444 & n8711 ) | ( n1799 & n8711 ) ;
  assign n9926 = n1762 & n9925 ;
  assign n9927 = n7905 & n9926 ;
  assign n9934 = ( n820 & n1051 ) | ( n820 & n4147 ) | ( n1051 & n4147 ) ;
  assign n9931 = ( n995 & ~n2869 ) | ( n995 & n2916 ) | ( ~n2869 & n2916 ) ;
  assign n9932 = n9395 | n9931 ;
  assign n9933 = n9932 ^ n3885 ^ 1'b0 ;
  assign n9928 = n5434 | n9863 ;
  assign n9929 = ( n2113 & n4954 ) | ( n2113 & ~n9928 ) | ( n4954 & ~n9928 ) ;
  assign n9930 = n9929 ^ n1015 ^ 1'b0 ;
  assign n9935 = n9934 ^ n9933 ^ n9930 ;
  assign n9936 = ( n677 & ~n1956 ) | ( n677 & n8471 ) | ( ~n1956 & n8471 ) ;
  assign n9937 = n9936 ^ n4120 ^ n2090 ;
  assign n9938 = ( n397 & n3281 ) | ( n397 & ~n8487 ) | ( n3281 & ~n8487 ) ;
  assign n9939 = ( n5390 & ~n9937 ) | ( n5390 & n9938 ) | ( ~n9937 & n9938 ) ;
  assign n9940 = n2794 & ~n9939 ;
  assign n9941 = ( n2581 & n3283 ) | ( n2581 & ~n8058 ) | ( n3283 & ~n8058 ) ;
  assign n9942 = n7040 ^ n3659 ^ x99 ;
  assign n9943 = n9941 & ~n9942 ;
  assign n9944 = n6548 | n9943 ;
  assign n9945 = ~n913 & n2038 ;
  assign n9946 = ( ~n925 & n1698 ) | ( ~n925 & n2759 ) | ( n1698 & n2759 ) ;
  assign n9950 = n379 | n508 ;
  assign n9951 = n8727 & ~n9950 ;
  assign n9952 = n9951 ^ n3620 ^ n457 ;
  assign n9953 = n2590 ^ n634 ^ 1'b0 ;
  assign n9954 = ( n2939 & n5629 ) | ( n2939 & n9953 ) | ( n5629 & n9953 ) ;
  assign n9955 = ( n2716 & ~n3950 ) | ( n2716 & n9954 ) | ( ~n3950 & n9954 ) ;
  assign n9956 = ~n9952 & n9955 ;
  assign n9957 = n9956 ^ n8033 ^ 1'b0 ;
  assign n9947 = n4234 ^ n2052 ^ n1367 ;
  assign n9948 = n9947 ^ n4384 ^ n2003 ;
  assign n9949 = ~n4736 & n9948 ;
  assign n9958 = n9957 ^ n9949 ^ n1188 ;
  assign n9959 = ( n9945 & ~n9946 ) | ( n9945 & n9958 ) | ( ~n9946 & n9958 ) ;
  assign n9960 = n7215 ^ n3193 ^ 1'b0 ;
  assign n9961 = n700 & n9960 ;
  assign n9962 = ~n280 & n9961 ;
  assign n9963 = n9962 ^ n6490 ^ 1'b0 ;
  assign n9964 = n6333 ^ n5303 ^ 1'b0 ;
  assign n9965 = ~n2830 & n9964 ;
  assign n9966 = n9965 ^ n2995 ^ 1'b0 ;
  assign n9967 = ( ~n514 & n2024 ) | ( ~n514 & n6080 ) | ( n2024 & n6080 ) ;
  assign n9968 = ( n3708 & n9355 ) | ( n3708 & n9967 ) | ( n9355 & n9967 ) ;
  assign n9969 = n5383 ^ n2695 ^ 1'b0 ;
  assign n9970 = ~n353 & n9969 ;
  assign n9973 = ( n754 & n1193 ) | ( n754 & n5364 ) | ( n1193 & n5364 ) ;
  assign n9974 = ~n4930 & n9973 ;
  assign n9975 = n9974 ^ n889 ^ 1'b0 ;
  assign n9971 = n5110 ^ n728 ^ 1'b0 ;
  assign n9972 = n398 & ~n9971 ;
  assign n9976 = n9975 ^ n9972 ^ n199 ;
  assign n9977 = ( x34 & ~n9687 ) | ( x34 & n9976 ) | ( ~n9687 & n9976 ) ;
  assign n9978 = n1088 ^ n245 ^ 1'b0 ;
  assign n9979 = n4877 & ~n9978 ;
  assign n9980 = n9979 ^ n6539 ^ n1609 ;
  assign n9981 = n2998 & ~n7249 ;
  assign n9982 = ~n6602 & n6861 ;
  assign n9983 = ~n9981 & n9982 ;
  assign n9984 = ( n139 & n6418 ) | ( n139 & n7555 ) | ( n6418 & n7555 ) ;
  assign n9985 = ( n7739 & ~n7901 ) | ( n7739 & n9984 ) | ( ~n7901 & n9984 ) ;
  assign n9986 = n9985 ^ n816 ^ 1'b0 ;
  assign n9987 = ~n1349 & n7272 ;
  assign n9988 = ( n393 & n4330 ) | ( n393 & ~n9987 ) | ( n4330 & ~n9987 ) ;
  assign n9989 = n9988 ^ n6598 ^ 1'b0 ;
  assign n9990 = ( x49 & n6279 ) | ( x49 & n9206 ) | ( n6279 & n9206 ) ;
  assign n9991 = ( n2773 & n5206 ) | ( n2773 & n6437 ) | ( n5206 & n6437 ) ;
  assign n9992 = n762 & n1554 ;
  assign n9993 = n919 & n1210 ;
  assign n9994 = ( n1822 & n4926 ) | ( n1822 & ~n5644 ) | ( n4926 & ~n5644 ) ;
  assign n9995 = ( n9992 & n9993 ) | ( n9992 & ~n9994 ) | ( n9993 & ~n9994 ) ;
  assign n9996 = n9995 ^ n4032 ^ n2776 ;
  assign n9997 = n650 ^ n341 ^ 1'b0 ;
  assign n9998 = n9997 ^ n8740 ^ n5332 ;
  assign n10002 = ( x39 & n2727 ) | ( x39 & ~n3056 ) | ( n2727 & ~n3056 ) ;
  assign n9999 = ( n2842 & n5559 ) | ( n2842 & n6607 ) | ( n5559 & n6607 ) ;
  assign n10000 = n9999 ^ n6572 ^ 1'b0 ;
  assign n10001 = n2224 & ~n10000 ;
  assign n10003 = n10002 ^ n10001 ^ n8144 ;
  assign n10004 = n10003 ^ n7905 ^ 1'b0 ;
  assign n10005 = n9998 & ~n10004 ;
  assign n10006 = n6601 ^ n5817 ^ n2461 ;
  assign n10007 = n7752 ^ n6023 ^ n5976 ;
  assign n10008 = n10006 & n10007 ;
  assign n10009 = ~n9958 & n10008 ;
  assign n10010 = ( n2482 & n5178 ) | ( n2482 & n5641 ) | ( n5178 & n5641 ) ;
  assign n10011 = ( n3370 & n7264 ) | ( n3370 & n10010 ) | ( n7264 & n10010 ) ;
  assign n10016 = n5813 ^ n3049 ^ n2043 ;
  assign n10012 = n8988 ^ n7002 ^ n6961 ;
  assign n10013 = n169 | n3666 ;
  assign n10014 = n10013 ^ n2669 ^ 1'b0 ;
  assign n10015 = n10012 | n10014 ;
  assign n10017 = n10016 ^ n10015 ^ 1'b0 ;
  assign n10018 = ~n5704 & n10017 ;
  assign n10021 = n3617 ^ n2545 ^ n844 ;
  assign n10020 = ( n2788 & n5065 ) | ( n2788 & n7370 ) | ( n5065 & n7370 ) ;
  assign n10019 = ( n924 & n9101 ) | ( n924 & n9954 ) | ( n9101 & n9954 ) ;
  assign n10022 = n10021 ^ n10020 ^ n10019 ;
  assign n10023 = ( n2092 & ~n7259 ) | ( n2092 & n7347 ) | ( ~n7259 & n7347 ) ;
  assign n10024 = n9361 ^ n8177 ^ n511 ;
  assign n10025 = ( n7082 & n10023 ) | ( n7082 & ~n10024 ) | ( n10023 & ~n10024 ) ;
  assign n10026 = n3557 & n8487 ;
  assign n10027 = ~n2280 & n10026 ;
  assign n10028 = n4622 ^ n4228 ^ n3822 ;
  assign n10029 = ( n3789 & n9636 ) | ( n3789 & n10028 ) | ( n9636 & n10028 ) ;
  assign n10030 = ( ~x124 & n582 ) | ( ~x124 & n2995 ) | ( n582 & n2995 ) ;
  assign n10031 = n10030 ^ n3704 ^ n3375 ;
  assign n10032 = ( n9539 & n10029 ) | ( n9539 & ~n10031 ) | ( n10029 & ~n10031 ) ;
  assign n10033 = ( ~n768 & n1466 ) | ( ~n768 & n1840 ) | ( n1466 & n1840 ) ;
  assign n10034 = ( n4225 & ~n6684 ) | ( n4225 & n10033 ) | ( ~n6684 & n10033 ) ;
  assign n10035 = n8470 ^ n5351 ^ 1'b0 ;
  assign n10036 = n7056 & n10035 ;
  assign n10042 = ~n1748 & n5100 ;
  assign n10040 = n6907 ^ n1266 ^ 1'b0 ;
  assign n10041 = n4350 & ~n10040 ;
  assign n10037 = ( n5892 & n6288 ) | ( n5892 & n7479 ) | ( n6288 & n7479 ) ;
  assign n10038 = n10037 ^ n5260 ^ n2767 ;
  assign n10039 = n7916 & ~n10038 ;
  assign n10043 = n10042 ^ n10041 ^ n10039 ;
  assign n10044 = n10043 ^ n5011 ^ 1'b0 ;
  assign n10045 = n2504 & n10044 ;
  assign n10046 = ( ~n1839 & n1868 ) | ( ~n1839 & n4976 ) | ( n1868 & n4976 ) ;
  assign n10047 = n3661 ^ n859 ^ 1'b0 ;
  assign n10048 = ~n2105 & n10047 ;
  assign n10049 = n10025 & n10048 ;
  assign n10050 = n8226 & ~n10049 ;
  assign n10051 = ( n1676 & n4284 ) | ( n1676 & ~n10050 ) | ( n4284 & ~n10050 ) ;
  assign n10052 = n7067 ^ n3895 ^ 1'b0 ;
  assign n10053 = n2117 | n10052 ;
  assign n10055 = ( n245 & ~n1573 ) | ( n245 & n6280 ) | ( ~n1573 & n6280 ) ;
  assign n10054 = n5430 & n9738 ;
  assign n10056 = n10055 ^ n10054 ^ 1'b0 ;
  assign n10057 = n5458 ^ n1466 ^ 1'b0 ;
  assign n10058 = n1849 & n2250 ;
  assign n10059 = n10058 ^ n826 ^ n797 ;
  assign n10060 = ( n1362 & ~n10057 ) | ( n1362 & n10059 ) | ( ~n10057 & n10059 ) ;
  assign n10061 = ~n9572 & n10060 ;
  assign n10063 = n1785 ^ n1609 ^ 1'b0 ;
  assign n10064 = n9199 & ~n10063 ;
  assign n10062 = n5244 ^ n5027 ^ 1'b0 ;
  assign n10065 = n10064 ^ n10062 ^ n6508 ;
  assign n10066 = ( ~n6200 & n7738 ) | ( ~n6200 & n10065 ) | ( n7738 & n10065 ) ;
  assign n10067 = n8470 ^ n3890 ^ x9 ;
  assign n10068 = n10066 | n10067 ;
  assign n10071 = n8123 ^ n7370 ^ 1'b0 ;
  assign n10072 = ~n3100 & n10071 ;
  assign n10073 = ~n3472 & n10072 ;
  assign n10069 = ( n1122 & n1618 ) | ( n1122 & ~n3201 ) | ( n1618 & ~n3201 ) ;
  assign n10070 = ( n1109 & n9261 ) | ( n1109 & ~n10069 ) | ( n9261 & ~n10069 ) ;
  assign n10074 = n10073 ^ n10070 ^ 1'b0 ;
  assign n10075 = n2362 & ~n10074 ;
  assign n10076 = n5099 & ~n10075 ;
  assign n10079 = n1629 ^ n751 ^ x106 ;
  assign n10077 = n2518 ^ n1993 ^ n329 ;
  assign n10078 = ( n423 & ~n9833 ) | ( n423 & n10077 ) | ( ~n9833 & n10077 ) ;
  assign n10080 = n10079 ^ n10078 ^ n6706 ;
  assign n10081 = n10080 ^ n5152 ^ 1'b0 ;
  assign n10082 = n3103 & n10081 ;
  assign n10083 = ( ~x105 & n1125 ) | ( ~x105 & n2038 ) | ( n1125 & n2038 ) ;
  assign n10084 = ( n3122 & n6592 ) | ( n3122 & ~n10083 ) | ( n6592 & ~n10083 ) ;
  assign n10085 = n2449 ^ n1996 ^ x83 ;
  assign n10086 = n10085 ^ n3278 ^ 1'b0 ;
  assign n10087 = n2791 & ~n10086 ;
  assign n10088 = n10087 ^ n2170 ^ 1'b0 ;
  assign n10089 = ~n8615 & n10088 ;
  assign n10090 = n1211 & n4966 ;
  assign n10091 = n7509 ^ n6384 ^ n655 ;
  assign n10092 = ~n1595 & n6218 ;
  assign n10093 = x112 & n10092 ;
  assign n10094 = ~n2561 & n10093 ;
  assign n10095 = n2264 | n10094 ;
  assign n10096 = n10095 ^ n342 ^ 1'b0 ;
  assign n10097 = ( n10090 & n10091 ) | ( n10090 & n10096 ) | ( n10091 & n10096 ) ;
  assign n10098 = ( n359 & n3017 ) | ( n359 & ~n8623 ) | ( n3017 & ~n8623 ) ;
  assign n10099 = ( n5805 & ~n8121 ) | ( n5805 & n10098 ) | ( ~n8121 & n10098 ) ;
  assign n10104 = n4405 ^ n2249 ^ 1'b0 ;
  assign n10100 = ( ~n2570 & n3586 ) | ( ~n2570 & n6128 ) | ( n3586 & n6128 ) ;
  assign n10101 = ( n2615 & n4275 ) | ( n2615 & ~n10100 ) | ( n4275 & ~n10100 ) ;
  assign n10102 = n10101 ^ n2221 ^ n1901 ;
  assign n10103 = n10102 ^ n7820 ^ n7575 ;
  assign n10105 = n10104 ^ n10103 ^ 1'b0 ;
  assign n10106 = n8894 ^ n4134 ^ n1023 ;
  assign n10107 = ( n1932 & ~n10104 ) | ( n1932 & n10106 ) | ( ~n10104 & n10106 ) ;
  assign n10108 = ( ~n924 & n5225 ) | ( ~n924 & n9007 ) | ( n5225 & n9007 ) ;
  assign n10109 = n1868 & ~n4878 ;
  assign n10110 = n1575 & n10109 ;
  assign n10111 = ( ~n2759 & n10039 ) | ( ~n2759 & n10110 ) | ( n10039 & n10110 ) ;
  assign n10112 = n10111 ^ n3932 ^ 1'b0 ;
  assign n10113 = n10108 | n10112 ;
  assign n10119 = n1578 | n5560 ;
  assign n10120 = n10119 ^ n1135 ^ 1'b0 ;
  assign n10121 = ~n7357 & n10120 ;
  assign n10122 = n6816 & n10121 ;
  assign n10123 = n3752 ^ n1005 ^ 1'b0 ;
  assign n10124 = ( n201 & n4142 ) | ( n201 & n10123 ) | ( n4142 & n10123 ) ;
  assign n10125 = ( n9618 & n10122 ) | ( n9618 & n10124 ) | ( n10122 & n10124 ) ;
  assign n10114 = n6494 ^ n2960 ^ n1597 ;
  assign n10115 = n3619 ^ n1149 ^ n328 ;
  assign n10116 = ( ~n858 & n7956 ) | ( ~n858 & n10115 ) | ( n7956 & n10115 ) ;
  assign n10117 = ~n10114 & n10116 ;
  assign n10118 = n6138 & n10117 ;
  assign n10126 = n10125 ^ n10118 ^ n2944 ;
  assign n10127 = ( n704 & n2450 ) | ( n704 & ~n6184 ) | ( n2450 & ~n6184 ) ;
  assign n10128 = n8644 ^ n2101 ^ n2075 ;
  assign n10129 = n10128 ^ n6266 ^ x75 ;
  assign n10130 = ( n9955 & n10127 ) | ( n9955 & ~n10129 ) | ( n10127 & ~n10129 ) ;
  assign n10135 = n1416 | n3430 ;
  assign n10136 = n10135 ^ n6961 ^ 1'b0 ;
  assign n10131 = n8167 ^ n7365 ^ n1155 ;
  assign n10132 = ~n1579 & n5710 ;
  assign n10133 = n10131 & ~n10132 ;
  assign n10134 = n5298 & n10133 ;
  assign n10137 = n10136 ^ n10134 ^ 1'b0 ;
  assign n10138 = n1998 ^ n410 ^ 1'b0 ;
  assign n10139 = n5476 & n10138 ;
  assign n10140 = n7336 ^ n2697 ^ n2503 ;
  assign n10141 = n8490 ^ n1472 ^ 1'b0 ;
  assign n10142 = n1698 & ~n10141 ;
  assign n10143 = ~n10140 & n10142 ;
  assign n10144 = n10073 ^ n870 ^ 1'b0 ;
  assign n10146 = ( n3265 & n5562 ) | ( n3265 & n8821 ) | ( n5562 & n8821 ) ;
  assign n10145 = n8865 ^ x59 ^ 1'b0 ;
  assign n10147 = n10146 ^ n10145 ^ 1'b0 ;
  assign n10148 = n4890 & ~n10147 ;
  assign n10149 = n141 | n2892 ;
  assign n10150 = n6495 | n8289 ;
  assign n10151 = n2311 & ~n10150 ;
  assign n10152 = ( n5808 & n10149 ) | ( n5808 & n10151 ) | ( n10149 & n10151 ) ;
  assign n10153 = x80 ^ x66 ^ 1'b0 ;
  assign n10154 = n5324 & n10153 ;
  assign n10155 = n5880 & n10154 ;
  assign n10156 = n10152 & n10155 ;
  assign n10157 = ~n3072 & n5445 ;
  assign n10158 = ( n5474 & n8312 ) | ( n5474 & ~n10157 ) | ( n8312 & ~n10157 ) ;
  assign n10159 = ( n1146 & n2025 ) | ( n1146 & ~n10158 ) | ( n2025 & ~n10158 ) ;
  assign n10163 = n8808 ^ n1566 ^ 1'b0 ;
  assign n10160 = n6116 ^ n4540 ^ 1'b0 ;
  assign n10161 = ~n9722 & n10160 ;
  assign n10162 = n10161 ^ n5848 ^ n3062 ;
  assign n10164 = n10163 ^ n10162 ^ n795 ;
  assign n10165 = n9177 ^ n2663 ^ n843 ;
  assign n10166 = n8777 ^ n7110 ^ 1'b0 ;
  assign n10167 = n10165 & ~n10166 ;
  assign n10168 = n1944 | n3197 ;
  assign n10169 = n5531 & ~n10168 ;
  assign n10170 = n2280 & ~n2767 ;
  assign n10171 = n3910 & n9147 ;
  assign n10172 = n386 & n10171 ;
  assign n10176 = n1735 | n3001 ;
  assign n10177 = ( x45 & n1042 ) | ( x45 & n10176 ) | ( n1042 & n10176 ) ;
  assign n10175 = n1231 & n1340 ;
  assign n10178 = n10177 ^ n10175 ^ 1'b0 ;
  assign n10173 = ~n2478 & n6049 ;
  assign n10174 = n6564 & n10173 ;
  assign n10179 = n10178 ^ n10174 ^ n2336 ;
  assign n10180 = n10179 ^ n9697 ^ 1'b0 ;
  assign n10183 = n1543 | n2714 ;
  assign n10184 = ( n2736 & ~n2875 ) | ( n2736 & n10183 ) | ( ~n2875 & n10183 ) ;
  assign n10182 = n2412 & ~n9032 ;
  assign n10185 = n10184 ^ n10182 ^ 1'b0 ;
  assign n10181 = n6302 ^ n4962 ^ n4627 ;
  assign n10186 = n10185 ^ n10181 ^ n9602 ;
  assign n10187 = n7858 & ~n8553 ;
  assign n10188 = ( n934 & n3076 ) | ( n934 & n7497 ) | ( n3076 & n7497 ) ;
  assign n10189 = n4667 & n10188 ;
  assign n10190 = n10189 ^ n8480 ^ 1'b0 ;
  assign n10202 = n1390 & ~n1613 ;
  assign n10200 = ( ~n289 & n2555 ) | ( ~n289 & n8864 ) | ( n2555 & n8864 ) ;
  assign n10198 = n5507 & ~n9128 ;
  assign n10199 = n4727 & n10198 ;
  assign n10201 = n10200 ^ n10199 ^ n3641 ;
  assign n10196 = n6401 ^ n5243 ^ x60 ;
  assign n10191 = n4279 ^ n3855 ^ n2299 ;
  assign n10192 = n2030 | n2939 ;
  assign n10193 = x24 | n10192 ;
  assign n10194 = ( n3693 & n10191 ) | ( n3693 & n10193 ) | ( n10191 & n10193 ) ;
  assign n10195 = ( n3176 & ~n6165 ) | ( n3176 & n10194 ) | ( ~n6165 & n10194 ) ;
  assign n10197 = n10196 ^ n10195 ^ n6648 ;
  assign n10203 = n10202 ^ n10201 ^ n10197 ;
  assign n10204 = ~n10190 & n10203 ;
  assign n10205 = n10204 ^ n7076 ^ 1'b0 ;
  assign n10206 = ~n2719 & n10205 ;
  assign n10207 = n1529 & ~n3242 ;
  assign n10208 = n10207 ^ n1096 ^ 1'b0 ;
  assign n10209 = n10206 & ~n10208 ;
  assign n10214 = n4779 ^ n3072 ^ 1'b0 ;
  assign n10210 = ( x71 & n510 ) | ( x71 & ~n6591 ) | ( n510 & ~n6591 ) ;
  assign n10211 = n1984 & n5023 ;
  assign n10212 = ~n8949 & n10211 ;
  assign n10213 = n10210 & ~n10212 ;
  assign n10215 = n10214 ^ n10213 ^ 1'b0 ;
  assign n10216 = n10215 ^ n7350 ^ n3935 ;
  assign n10217 = n3311 & ~n7777 ;
  assign n10218 = n5710 & n10217 ;
  assign n10219 = n233 & ~n1114 ;
  assign n10220 = n10219 ^ n5598 ^ 1'b0 ;
  assign n10221 = n9636 ^ n1643 ^ 1'b0 ;
  assign n10222 = n517 & n2758 ;
  assign n10223 = n10222 ^ n4072 ^ n3472 ;
  assign n10224 = n234 & ~n4272 ;
  assign n10225 = ~n7824 & n10224 ;
  assign n10226 = ( n6019 & n10223 ) | ( n6019 & ~n10225 ) | ( n10223 & ~n10225 ) ;
  assign n10227 = ( n1257 & ~n10221 ) | ( n1257 & n10226 ) | ( ~n10221 & n10226 ) ;
  assign n10229 = ( ~n206 & n4627 ) | ( ~n206 & n9402 ) | ( n4627 & n9402 ) ;
  assign n10228 = n1857 | n3966 ;
  assign n10230 = n10229 ^ n10228 ^ 1'b0 ;
  assign n10231 = ( n626 & n4011 ) | ( n626 & ~n4291 ) | ( n4011 & ~n4291 ) ;
  assign n10232 = n9619 ^ n3677 ^ n458 ;
  assign n10233 = n10073 | n10232 ;
  assign n10234 = ~n3075 & n4565 ;
  assign n10235 = n7330 ^ n293 ^ 1'b0 ;
  assign n10236 = n9689 | n10235 ;
  assign n10237 = n3827 ^ n334 ^ x121 ;
  assign n10238 = ( n1785 & n5276 ) | ( n1785 & n10237 ) | ( n5276 & n10237 ) ;
  assign n10242 = n4645 ^ n917 ^ n596 ;
  assign n10239 = n1967 | n6680 ;
  assign n10240 = n1321 & ~n10239 ;
  assign n10241 = ( n5472 & n8679 ) | ( n5472 & n10240 ) | ( n8679 & n10240 ) ;
  assign n10243 = n10242 ^ n10241 ^ n3773 ;
  assign n10244 = n1335 ^ n837 ^ x42 ;
  assign n10245 = n2135 & n9162 ;
  assign n10246 = n10245 ^ n2827 ^ 1'b0 ;
  assign n10247 = n10246 ^ n7515 ^ n4097 ;
  assign n10248 = ( ~n5060 & n10244 ) | ( ~n5060 & n10247 ) | ( n10244 & n10247 ) ;
  assign n10249 = ( n10238 & n10243 ) | ( n10238 & ~n10248 ) | ( n10243 & ~n10248 ) ;
  assign n10250 = n4317 ^ n1289 ^ 1'b0 ;
  assign n10251 = n5651 ^ n5434 ^ n2253 ;
  assign n10252 = x7 & ~n8983 ;
  assign n10253 = ~n10251 & n10252 ;
  assign n10254 = n4290 ^ n1025 ^ 1'b0 ;
  assign n10255 = ~n2614 & n10254 ;
  assign n10256 = n10253 & n10255 ;
  assign n10257 = n10256 ^ n4701 ^ 1'b0 ;
  assign n10258 = n10257 ^ n5012 ^ 1'b0 ;
  assign n10259 = n5330 & ~n10258 ;
  assign n10260 = n3023 & n9089 ;
  assign n10261 = n10260 ^ n7215 ^ 1'b0 ;
  assign n10262 = ( n7813 & n8233 ) | ( n7813 & n10261 ) | ( n8233 & n10261 ) ;
  assign n10263 = n5578 | n10262 ;
  assign n10264 = n10259 | n10263 ;
  assign n10267 = ( ~n2792 & n9065 ) | ( ~n2792 & n9308 ) | ( n9065 & n9308 ) ;
  assign n10265 = n1379 ^ n430 ^ 1'b0 ;
  assign n10266 = n5906 & ~n10265 ;
  assign n10268 = n10267 ^ n10266 ^ n5133 ;
  assign n10269 = n894 ^ n520 ^ 1'b0 ;
  assign n10270 = ( n1560 & n3738 ) | ( n1560 & ~n5080 ) | ( n3738 & ~n5080 ) ;
  assign n10271 = n10270 ^ n2357 ^ n2230 ;
  assign n10272 = ( ~n851 & n10269 ) | ( ~n851 & n10271 ) | ( n10269 & n10271 ) ;
  assign n10276 = n6760 ^ n6209 ^ 1'b0 ;
  assign n10277 = n10276 ^ n3515 ^ n2925 ;
  assign n10273 = n1381 | n4612 ;
  assign n10274 = n4442 ^ n192 ^ 1'b0 ;
  assign n10275 = ( n4556 & n10273 ) | ( n4556 & ~n10274 ) | ( n10273 & ~n10274 ) ;
  assign n10278 = n10277 ^ n10275 ^ n1959 ;
  assign n10279 = n10278 ^ n1131 ^ 1'b0 ;
  assign n10283 = n8181 ^ n7063 ^ n1418 ;
  assign n10280 = n4464 ^ n3757 ^ n1193 ;
  assign n10281 = n3776 & n4590 ;
  assign n10282 = n10280 & n10281 ;
  assign n10284 = n10283 ^ n10282 ^ n5509 ;
  assign n10285 = n1442 & n1893 ;
  assign n10286 = ~n10284 & n10285 ;
  assign n10287 = ( n298 & n1374 ) | ( n298 & ~n2098 ) | ( n1374 & ~n2098 ) ;
  assign n10288 = ( n2216 & ~n2457 ) | ( n2216 & n6603 ) | ( ~n2457 & n6603 ) ;
  assign n10289 = n10288 ^ n5665 ^ n5001 ;
  assign n10290 = n8715 ^ n6574 ^ n1682 ;
  assign n10291 = n10290 ^ n9952 ^ n5531 ;
  assign n10292 = n5913 & ~n10291 ;
  assign n10293 = n9501 ^ n1651 ^ 1'b0 ;
  assign n10294 = ( ~n8395 & n8839 ) | ( ~n8395 & n10293 ) | ( n8839 & n10293 ) ;
  assign n10295 = ( n2693 & n6414 ) | ( n2693 & ~n10294 ) | ( n6414 & ~n10294 ) ;
  assign n10296 = n8982 ^ n8116 ^ n3043 ;
  assign n10297 = n10296 ^ n2058 ^ 1'b0 ;
  assign n10298 = n2844 & n3711 ;
  assign n10299 = n10298 ^ n3916 ^ n2493 ;
  assign n10300 = ( n2922 & n4934 ) | ( n2922 & n10299 ) | ( n4934 & n10299 ) ;
  assign n10301 = ~n3703 & n10089 ;
  assign n10302 = ~n2360 & n10301 ;
  assign n10303 = ( n1039 & ~n2470 ) | ( n1039 & n2798 ) | ( ~n2470 & n2798 ) ;
  assign n10304 = ( x41 & n4968 ) | ( x41 & ~n10303 ) | ( n4968 & ~n10303 ) ;
  assign n10305 = n10304 ^ n3063 ^ n494 ;
  assign n10306 = ( n1239 & n1966 ) | ( n1239 & ~n7585 ) | ( n1966 & ~n7585 ) ;
  assign n10307 = n5295 & ~n10306 ;
  assign n10308 = ( n1996 & n7359 ) | ( n1996 & n10307 ) | ( n7359 & n10307 ) ;
  assign n10309 = n9736 ^ n2124 ^ n1868 ;
  assign n10310 = n10309 ^ n5112 ^ n3603 ;
  assign n10317 = n4502 ^ n1710 ^ x121 ;
  assign n10318 = n6324 & ~n10317 ;
  assign n10319 = ( n148 & n1719 ) | ( n148 & ~n10318 ) | ( n1719 & ~n10318 ) ;
  assign n10311 = n1802 ^ n201 ^ 1'b0 ;
  assign n10312 = n10311 ^ n7439 ^ n620 ;
  assign n10313 = n2369 ^ n2018 ^ 1'b0 ;
  assign n10314 = n10313 ^ n6484 ^ 1'b0 ;
  assign n10315 = n10312 & n10314 ;
  assign n10316 = n10315 ^ n9439 ^ n3271 ;
  assign n10320 = n10319 ^ n10316 ^ 1'b0 ;
  assign n10321 = n8280 & n10320 ;
  assign n10322 = ( n1690 & n6476 ) | ( n1690 & n7290 ) | ( n6476 & n7290 ) ;
  assign n10323 = ( n2611 & ~n8861 ) | ( n2611 & n10322 ) | ( ~n8861 & n10322 ) ;
  assign n10326 = n636 ^ x91 ^ 1'b0 ;
  assign n10324 = n1467 | n7579 ;
  assign n10325 = n10324 ^ n6658 ^ n818 ;
  assign n10327 = n10326 ^ n10325 ^ n2077 ;
  assign n10328 = n10149 ^ n197 ^ 1'b0 ;
  assign n10329 = ( n4794 & ~n5172 ) | ( n4794 & n10328 ) | ( ~n5172 & n10328 ) ;
  assign n10330 = n10329 ^ n8470 ^ n7108 ;
  assign n10333 = n8715 ^ n3778 ^ n1346 ;
  assign n10331 = n7059 ^ n1413 ^ n1217 ;
  assign n10332 = n10331 ^ n5270 ^ n3748 ;
  assign n10334 = n10333 ^ n10332 ^ n451 ;
  assign n10335 = n6128 ^ n3809 ^ 1'b0 ;
  assign n10336 = n1400 | n10335 ;
  assign n10337 = n10336 ^ n320 ^ 1'b0 ;
  assign n10338 = n7584 & n10337 ;
  assign n10339 = n6896 ^ n4569 ^ n1550 ;
  assign n10340 = n10339 ^ n2313 ^ n518 ;
  assign n10341 = n5736 ^ n4110 ^ n2301 ;
  assign n10342 = n10341 ^ n4567 ^ 1'b0 ;
  assign n10343 = ~n1515 & n10342 ;
  assign n10344 = n6034 & ~n6064 ;
  assign n10348 = n5411 ^ n5333 ^ 1'b0 ;
  assign n10349 = n5644 | n10348 ;
  assign n10350 = n10349 ^ n1989 ^ 1'b0 ;
  assign n10345 = ~n164 & n1650 ;
  assign n10346 = n10345 ^ n8669 ^ 1'b0 ;
  assign n10347 = n6054 & ~n10346 ;
  assign n10351 = n10350 ^ n10347 ^ 1'b0 ;
  assign n10352 = ~n1474 & n10351 ;
  assign n10353 = n10352 ^ x72 ^ 1'b0 ;
  assign n10354 = n2390 | n10353 ;
  assign n10355 = n10344 & ~n10354 ;
  assign n10356 = ( n7841 & n10343 ) | ( n7841 & ~n10355 ) | ( n10343 & ~n10355 ) ;
  assign n10357 = n9769 ^ n1444 ^ n1290 ;
  assign n10358 = ( ~n130 & n1228 ) | ( ~n130 & n3068 ) | ( n1228 & n3068 ) ;
  assign n10359 = n10358 ^ n4953 ^ n4342 ;
  assign n10360 = ( n2934 & ~n10357 ) | ( n2934 & n10359 ) | ( ~n10357 & n10359 ) ;
  assign n10361 = n362 | n6282 ;
  assign n10362 = n10361 ^ n9447 ^ 1'b0 ;
  assign n10363 = ~n830 & n3145 ;
  assign n10364 = n9237 & n10363 ;
  assign n10365 = n7509 ^ n6626 ^ n6569 ;
  assign n10366 = ( n10214 & ~n10364 ) | ( n10214 & n10365 ) | ( ~n10364 & n10365 ) ;
  assign n10367 = n7913 ^ n6740 ^ 1'b0 ;
  assign n10368 = n269 & ~n10367 ;
  assign n10369 = n8162 ^ n6409 ^ n2919 ;
  assign n10370 = n10368 & n10369 ;
  assign n10371 = ~x70 & n10370 ;
  assign n10373 = n5679 ^ n216 ^ 1'b0 ;
  assign n10374 = n7394 & ~n10373 ;
  assign n10372 = ~n5169 & n5718 ;
  assign n10375 = n10374 ^ n10372 ^ 1'b0 ;
  assign n10376 = n2696 | n2794 ;
  assign n10377 = n5644 & ~n10376 ;
  assign n10378 = n10377 ^ n6792 ^ n3242 ;
  assign n10379 = ( n927 & ~n2281 ) | ( n927 & n5360 ) | ( ~n2281 & n5360 ) ;
  assign n10382 = x10 & n8400 ;
  assign n10383 = ~n6314 & n10382 ;
  assign n10380 = ( n835 & n2022 ) | ( n835 & n3523 ) | ( n2022 & n3523 ) ;
  assign n10381 = ( n1005 & n2578 ) | ( n1005 & ~n10380 ) | ( n2578 & ~n10380 ) ;
  assign n10384 = n10383 ^ n10381 ^ n2772 ;
  assign n10385 = ( ~n10378 & n10379 ) | ( ~n10378 & n10384 ) | ( n10379 & n10384 ) ;
  assign n10386 = n6596 ^ n3314 ^ n1528 ;
  assign n10387 = n5572 | n10386 ;
  assign n10388 = n10387 ^ n4192 ^ 1'b0 ;
  assign n10392 = n10309 ^ n5206 ^ n1116 ;
  assign n10390 = ( n177 & ~n7381 ) | ( n177 & n10201 ) | ( ~n7381 & n10201 ) ;
  assign n10391 = ( n5621 & n10033 ) | ( n5621 & n10390 ) | ( n10033 & n10390 ) ;
  assign n10389 = n9534 ^ n9367 ^ 1'b0 ;
  assign n10393 = n10392 ^ n10391 ^ n10389 ;
  assign n10394 = n4577 ^ n4015 ^ 1'b0 ;
  assign n10395 = ( n2276 & n2916 ) | ( n2276 & ~n10394 ) | ( n2916 & ~n10394 ) ;
  assign n10396 = n2904 ^ n2736 ^ n2568 ;
  assign n10398 = ~n1079 & n1946 ;
  assign n10397 = n4186 ^ n2866 ^ n1395 ;
  assign n10399 = n10398 ^ n10397 ^ n5659 ;
  assign n10400 = n833 | n10399 ;
  assign n10401 = n9894 ^ n795 ^ 1'b0 ;
  assign n10402 = n2934 | n10401 ;
  assign n10403 = n10402 ^ n5494 ^ x87 ;
  assign n10404 = n5582 ^ n2331 ^ n1313 ;
  assign n10405 = n10404 ^ n2740 ^ n604 ;
  assign n10406 = n10405 ^ n920 ^ 1'b0 ;
  assign n10407 = ( n5594 & n10403 ) | ( n5594 & n10406 ) | ( n10403 & n10406 ) ;
  assign n10408 = ( ~n8597 & n9526 ) | ( ~n8597 & n9925 ) | ( n9526 & n9925 ) ;
  assign n10409 = ~n3689 & n5295 ;
  assign n10411 = n3901 & ~n5306 ;
  assign n10412 = n3198 & n10411 ;
  assign n10413 = ( ~x64 & n3538 ) | ( ~x64 & n10412 ) | ( n3538 & n10412 ) ;
  assign n10410 = ( n1758 & n2427 ) | ( n1758 & ~n3221 ) | ( n2427 & ~n3221 ) ;
  assign n10414 = n10413 ^ n10410 ^ x40 ;
  assign n10415 = n4100 & n4366 ;
  assign n10416 = n6785 ^ n6164 ^ 1'b0 ;
  assign n10417 = ( n335 & ~n4169 ) | ( n335 & n10416 ) | ( ~n4169 & n10416 ) ;
  assign n10418 = ~n1694 & n2825 ;
  assign n10419 = ~n2774 & n6230 ;
  assign n10420 = n9993 ^ n2190 ^ 1'b0 ;
  assign n10421 = ~n10419 & n10420 ;
  assign n10422 = n10418 & ~n10421 ;
  assign n10423 = n10422 ^ n7435 ^ n326 ;
  assign n10424 = n10423 ^ n2386 ^ x5 ;
  assign n10425 = n4383 ^ n2631 ^ n1018 ;
  assign n10426 = n10425 ^ n3570 ^ 1'b0 ;
  assign n10427 = n10165 ^ n352 ^ n211 ;
  assign n10429 = n4654 ^ n3812 ^ n2376 ;
  assign n10430 = n10429 ^ n4117 ^ n1371 ;
  assign n10428 = x3 & ~n5624 ;
  assign n10431 = n10430 ^ n10428 ^ 1'b0 ;
  assign n10432 = n571 & ~n947 ;
  assign n10433 = n10432 ^ n10357 ^ 1'b0 ;
  assign n10434 = n4952 & ~n6215 ;
  assign n10435 = n10434 ^ n1312 ^ 1'b0 ;
  assign n10437 = n1873 ^ n845 ^ 1'b0 ;
  assign n10436 = ( n693 & n3127 ) | ( n693 & n5170 ) | ( n3127 & n5170 ) ;
  assign n10438 = n10437 ^ n10436 ^ 1'b0 ;
  assign n10439 = n8074 ^ n5392 ^ 1'b0 ;
  assign n10441 = n1461 & n3762 ;
  assign n10440 = n4628 ^ n3850 ^ 1'b0 ;
  assign n10442 = n10441 ^ n10440 ^ n7959 ;
  assign n10443 = n9450 ^ n8281 ^ n1250 ;
  assign n10444 = n2473 & ~n10443 ;
  assign n10445 = n10444 ^ n371 ^ 1'b0 ;
  assign n10448 = ~n445 & n728 ;
  assign n10446 = n7943 ^ n1307 ^ n878 ;
  assign n10447 = n10446 ^ n3166 ^ n410 ;
  assign n10449 = n10448 ^ n10447 ^ n3821 ;
  assign n10450 = ( n746 & n10445 ) | ( n746 & n10449 ) | ( n10445 & n10449 ) ;
  assign n10452 = n5962 ^ n2785 ^ 1'b0 ;
  assign n10451 = ( n3214 & ~n4907 ) | ( n3214 & n6250 ) | ( ~n4907 & n6250 ) ;
  assign n10453 = n10452 ^ n10451 ^ n9124 ;
  assign n10454 = n4663 ^ n1251 ^ 1'b0 ;
  assign n10455 = n3153 & ~n10454 ;
  assign n10456 = n10455 ^ n4930 ^ 1'b0 ;
  assign n10457 = n10456 ^ n7917 ^ 1'b0 ;
  assign n10458 = n10237 ^ n7747 ^ 1'b0 ;
  assign n10460 = n1680 ^ n1313 ^ 1'b0 ;
  assign n10459 = n7891 ^ n5604 ^ n1633 ;
  assign n10461 = n10460 ^ n10459 ^ n2460 ;
  assign n10462 = ( n9574 & ~n9666 ) | ( n9574 & n10461 ) | ( ~n9666 & n10461 ) ;
  assign n10463 = n7088 ^ n2026 ^ n1718 ;
  assign n10464 = ~n8214 & n9317 ;
  assign n10465 = n195 & ~n7059 ;
  assign n10466 = n7517 & ~n10465 ;
  assign n10467 = n2968 & n10466 ;
  assign n10468 = n4014 ^ n2099 ^ 1'b0 ;
  assign n10469 = n10468 ^ n4507 ^ n3409 ;
  assign n10470 = n10469 ^ x74 ^ 1'b0 ;
  assign n10471 = ( ~n2225 & n2733 ) | ( ~n2225 & n10470 ) | ( n2733 & n10470 ) ;
  assign n10472 = ( n235 & ~n5574 ) | ( n235 & n10471 ) | ( ~n5574 & n10471 ) ;
  assign n10473 = n9670 ^ n5147 ^ 1'b0 ;
  assign n10474 = n3736 | n5490 ;
  assign n10475 = n2403 | n10474 ;
  assign n10476 = n2205 & n10475 ;
  assign n10479 = n10021 ^ n2990 ^ 1'b0 ;
  assign n10480 = n3005 & n10479 ;
  assign n10477 = ~n3069 & n4608 ;
  assign n10478 = n10477 ^ x33 ^ 1'b0 ;
  assign n10481 = n10480 ^ n10478 ^ n3941 ;
  assign n10482 = n3033 ^ n725 ^ 1'b0 ;
  assign n10483 = n10282 | n10482 ;
  assign n10484 = n2560 ^ n1232 ^ n296 ;
  assign n10488 = ( n2403 & n3748 ) | ( n2403 & n9286 ) | ( n3748 & n9286 ) ;
  assign n10485 = n2849 & n5726 ;
  assign n10486 = n10485 ^ n572 ^ 1'b0 ;
  assign n10487 = ( ~n2278 & n6242 ) | ( ~n2278 & n10486 ) | ( n6242 & n10486 ) ;
  assign n10489 = n10488 ^ n10487 ^ 1'b0 ;
  assign n10490 = ( ~n9031 & n10484 ) | ( ~n9031 & n10489 ) | ( n10484 & n10489 ) ;
  assign n10491 = ( x12 & ~n5242 ) | ( x12 & n6145 ) | ( ~n5242 & n6145 ) ;
  assign n10494 = n7928 ^ n5894 ^ 1'b0 ;
  assign n10492 = ( ~n2204 & n4502 ) | ( ~n2204 & n6548 ) | ( n4502 & n6548 ) ;
  assign n10493 = ( ~n3033 & n8909 ) | ( ~n3033 & n10492 ) | ( n8909 & n10492 ) ;
  assign n10495 = n10494 ^ n10493 ^ n9489 ;
  assign n10496 = ~n4427 & n9031 ;
  assign n10497 = n2810 ^ n1617 ^ n203 ;
  assign n10498 = ~n3495 & n10497 ;
  assign n10499 = n10498 ^ n10432 ^ n2820 ;
  assign n10501 = n666 & n2373 ;
  assign n10502 = n10501 ^ n2941 ^ 1'b0 ;
  assign n10500 = n4989 ^ n4525 ^ n3173 ;
  assign n10503 = n10502 ^ n10500 ^ n189 ;
  assign n10504 = ( n869 & n3217 ) | ( n869 & n5053 ) | ( n3217 & n5053 ) ;
  assign n10505 = ( n600 & n3283 ) | ( n600 & ~n7811 ) | ( n3283 & ~n7811 ) ;
  assign n10506 = n10505 ^ n10162 ^ n7407 ;
  assign n10507 = ( n6225 & ~n10504 ) | ( n6225 & n10506 ) | ( ~n10504 & n10506 ) ;
  assign n10508 = n1082 & ~n6402 ;
  assign n10514 = n10037 ^ n3574 ^ n1932 ;
  assign n10509 = ~n3804 & n6366 ;
  assign n10510 = n10509 ^ n9097 ^ 1'b0 ;
  assign n10511 = n2083 & n10510 ;
  assign n10512 = ( ~n6403 & n8198 ) | ( ~n6403 & n10511 ) | ( n8198 & n10511 ) ;
  assign n10513 = n10512 ^ n6527 ^ n449 ;
  assign n10515 = n10514 ^ n10513 ^ 1'b0 ;
  assign n10516 = n10508 | n10515 ;
  assign n10517 = ~n3259 & n6222 ;
  assign n10518 = n10517 ^ n5717 ^ n5136 ;
  assign n10519 = n7277 ^ n7138 ^ 1'b0 ;
  assign n10522 = n2754 ^ n2570 ^ n418 ;
  assign n10521 = n5945 ^ n2536 ^ 1'b0 ;
  assign n10520 = n3851 ^ n3505 ^ 1'b0 ;
  assign n10523 = n10522 ^ n10521 ^ n10520 ;
  assign n10524 = ~n2375 & n3207 ;
  assign n10525 = n10524 ^ n1783 ^ n683 ;
  assign n10526 = n2479 | n10525 ;
  assign n10527 = ( n7703 & n10523 ) | ( n7703 & ~n10526 ) | ( n10523 & ~n10526 ) ;
  assign n10528 = n5024 ^ n201 ^ 1'b0 ;
  assign n10529 = ( n4145 & n7631 ) | ( n4145 & ~n10528 ) | ( n7631 & ~n10528 ) ;
  assign n10530 = n7262 ^ n2658 ^ n2356 ;
  assign n10531 = n592 & ~n4362 ;
  assign n10532 = n10531 ^ n1173 ^ 1'b0 ;
  assign n10533 = n2020 & ~n4481 ;
  assign n10534 = ( n3718 & n10532 ) | ( n3718 & n10533 ) | ( n10532 & n10533 ) ;
  assign n10535 = n7513 ^ n131 ^ 1'b0 ;
  assign n10536 = n10535 ^ n5780 ^ n1877 ;
  assign n10537 = n3954 ^ n2169 ^ 1'b0 ;
  assign n10538 = n6362 & n10537 ;
  assign n10539 = n10538 ^ n4913 ^ 1'b0 ;
  assign n10540 = ( ~n7106 & n7673 ) | ( ~n7106 & n8584 ) | ( n7673 & n8584 ) ;
  assign n10541 = ( n485 & n1072 ) | ( n485 & ~n3156 ) | ( n1072 & ~n3156 ) ;
  assign n10542 = n10541 ^ n7060 ^ n1994 ;
  assign n10543 = ~n3361 & n9447 ;
  assign n10544 = ( ~n8273 & n10542 ) | ( ~n8273 & n10543 ) | ( n10542 & n10543 ) ;
  assign n10545 = ~n1828 & n7427 ;
  assign n10546 = n5998 & ~n10545 ;
  assign n10547 = n10546 ^ n7683 ^ 1'b0 ;
  assign n10548 = ( n5464 & n5490 ) | ( n5464 & n10547 ) | ( n5490 & n10547 ) ;
  assign n10549 = n1151 & ~n10548 ;
  assign n10550 = n10549 ^ n7585 ^ n334 ;
  assign n10551 = n2912 ^ n2895 ^ 1'b0 ;
  assign n10552 = n2807 | n10551 ;
  assign n10555 = n1186 | n2306 ;
  assign n10553 = n3202 & ~n5053 ;
  assign n10554 = ~n1297 & n10553 ;
  assign n10556 = n10555 ^ n10554 ^ n165 ;
  assign n10557 = n8314 ^ n587 ^ 1'b0 ;
  assign n10558 = n3328 & n10557 ;
  assign n10561 = ( x37 & n854 ) | ( x37 & n1201 ) | ( n854 & n1201 ) ;
  assign n10562 = n10561 ^ n1848 ^ n1025 ;
  assign n10563 = ( n582 & n1795 ) | ( n582 & ~n10562 ) | ( n1795 & ~n10562 ) ;
  assign n10559 = n4412 & ~n4456 ;
  assign n10560 = n10559 ^ n5713 ^ n3264 ;
  assign n10564 = n10563 ^ n10560 ^ n5937 ;
  assign n10565 = n6974 ^ n4891 ^ 1'b0 ;
  assign n10566 = n2689 | n2965 ;
  assign n10567 = ( n5084 & n5735 ) | ( n5084 & n10566 ) | ( n5735 & n10566 ) ;
  assign n10568 = n4704 ^ n942 ^ 1'b0 ;
  assign n10569 = n10567 & n10568 ;
  assign n10570 = n9016 ^ n3982 ^ n2092 ;
  assign n10571 = n8918 ^ n7778 ^ n5415 ;
  assign n10572 = n10571 ^ n7141 ^ n304 ;
  assign n10573 = n4951 ^ n2939 ^ n596 ;
  assign n10574 = n10573 ^ n7304 ^ 1'b0 ;
  assign n10575 = n10522 | n10574 ;
  assign n10576 = n10575 ^ n9968 ^ n4883 ;
  assign n10577 = n3320 ^ n2528 ^ 1'b0 ;
  assign n10578 = ( n710 & n1694 ) | ( n710 & ~n10577 ) | ( n1694 & ~n10577 ) ;
  assign n10579 = n10578 ^ n1226 ^ 1'b0 ;
  assign n10580 = n10579 ^ n8789 ^ n5521 ;
  assign n10581 = n6198 ^ n4079 ^ 1'b0 ;
  assign n10582 = ( n2594 & n4555 ) | ( n2594 & n8912 ) | ( n4555 & n8912 ) ;
  assign n10583 = n9728 ^ n4008 ^ 1'b0 ;
  assign n10584 = ( n1971 & ~n9537 ) | ( n1971 & n10583 ) | ( ~n9537 & n10583 ) ;
  assign n10585 = n10582 | n10584 ;
  assign n10586 = ( n7638 & n10581 ) | ( n7638 & ~n10585 ) | ( n10581 & ~n10585 ) ;
  assign n10587 = ~n751 & n7098 ;
  assign n10588 = n10586 & ~n10587 ;
  assign n10605 = n9447 ^ n8312 ^ n4939 ;
  assign n10589 = n8305 ^ n5815 ^ 1'b0 ;
  assign n10590 = n2921 & ~n10589 ;
  assign n10591 = n4474 & n10590 ;
  assign n10592 = n10591 ^ n7891 ^ 1'b0 ;
  assign n10593 = n8011 & n10592 ;
  assign n10594 = n6953 & n10593 ;
  assign n10595 = ( n818 & n2811 ) | ( n818 & ~n5954 ) | ( n2811 & ~n5954 ) ;
  assign n10596 = x113 & n10595 ;
  assign n10597 = ~n397 & n10596 ;
  assign n10598 = n1863 ^ n1828 ^ 1'b0 ;
  assign n10599 = n2660 ^ n1470 ^ n1141 ;
  assign n10600 = ( n4098 & n10598 ) | ( n4098 & n10599 ) | ( n10598 & n10599 ) ;
  assign n10601 = ~n10597 & n10600 ;
  assign n10602 = n3738 ^ n1713 ^ 1'b0 ;
  assign n10603 = n10601 | n10602 ;
  assign n10604 = n10594 | n10603 ;
  assign n10606 = n10605 ^ n10604 ^ 1'b0 ;
  assign n10607 = ( n2231 & n4623 ) | ( n2231 & n8421 ) | ( n4623 & n8421 ) ;
  assign n10608 = n3506 | n6087 ;
  assign n10609 = n1569 & ~n10608 ;
  assign n10610 = n10607 & ~n10609 ;
  assign n10611 = ~n5726 & n10610 ;
  assign n10612 = n5802 ^ n3498 ^ n801 ;
  assign n10613 = n10612 ^ n301 ^ 1'b0 ;
  assign n10614 = n3467 & n10613 ;
  assign n10617 = n1263 & ~n10524 ;
  assign n10618 = n10617 ^ n7200 ^ 1'b0 ;
  assign n10619 = n10618 ^ n7082 ^ n4358 ;
  assign n10620 = ( n5259 & n8166 ) | ( n5259 & ~n10619 ) | ( n8166 & ~n10619 ) ;
  assign n10615 = n6375 ^ n3807 ^ 1'b0 ;
  assign n10616 = n2515 | n10615 ;
  assign n10621 = n10620 ^ n10616 ^ n1220 ;
  assign n10625 = n1125 & n8156 ;
  assign n10626 = n10625 ^ n2003 ^ 1'b0 ;
  assign n10627 = ( n7632 & ~n9132 ) | ( n7632 & n10626 ) | ( ~n9132 & n10626 ) ;
  assign n10623 = n10448 ^ n3554 ^ n485 ;
  assign n10622 = ( n371 & ~n1134 ) | ( n371 & n7290 ) | ( ~n1134 & n7290 ) ;
  assign n10624 = n10623 ^ n10622 ^ n3948 ;
  assign n10628 = n10627 ^ n10624 ^ n5000 ;
  assign n10629 = ( n1386 & n3422 ) | ( n1386 & ~n9600 ) | ( n3422 & ~n9600 ) ;
  assign n10630 = n622 | n7803 ;
  assign n10631 = n10629 & ~n10630 ;
  assign n10632 = n10559 ^ n7002 ^ 1'b0 ;
  assign n10633 = n10632 ^ n791 ^ n475 ;
  assign n10635 = n3461 & ~n6574 ;
  assign n10636 = ( n4804 & n7481 ) | ( n4804 & ~n10635 ) | ( n7481 & ~n10635 ) ;
  assign n10634 = n9496 ^ n9031 ^ 1'b0 ;
  assign n10637 = n10636 ^ n10634 ^ n8116 ;
  assign n10638 = n5005 & ~n5133 ;
  assign n10640 = ( n1551 & ~n2070 ) | ( n1551 & n2900 ) | ( ~n2070 & n2900 ) ;
  assign n10641 = ( n2164 & ~n7274 ) | ( n2164 & n10640 ) | ( ~n7274 & n10640 ) ;
  assign n10639 = n5738 ^ n4773 ^ n1370 ;
  assign n10642 = n10641 ^ n10639 ^ n8813 ;
  assign n10643 = ( n593 & n3460 ) | ( n593 & ~n10642 ) | ( n3460 & ~n10642 ) ;
  assign n10644 = ( ~n1095 & n3600 ) | ( ~n1095 & n5723 ) | ( n3600 & n5723 ) ;
  assign n10645 = n3701 & n3959 ;
  assign n10646 = ~x22 & n10645 ;
  assign n10647 = n10646 ^ n7601 ^ n5195 ;
  assign n10648 = n10647 ^ n9359 ^ n964 ;
  assign n10649 = n6375 ^ n5840 ^ 1'b0 ;
  assign n10650 = n7819 & ~n10649 ;
  assign n10651 = n2299 ^ n336 ^ n151 ;
  assign n10652 = ( n324 & n1886 ) | ( n324 & n6544 ) | ( n1886 & n6544 ) ;
  assign n10653 = n3141 & n9946 ;
  assign n10654 = n10652 & n10653 ;
  assign n10655 = ~n10452 & n10654 ;
  assign n10656 = ( n10085 & ~n10651 ) | ( n10085 & n10655 ) | ( ~n10651 & n10655 ) ;
  assign n10657 = n10656 ^ n418 ^ 1'b0 ;
  assign n10658 = n8981 & n10657 ;
  assign n10659 = n8142 ^ n4790 ^ 1'b0 ;
  assign n10660 = n10659 ^ n9851 ^ n5521 ;
  assign n10661 = ( n180 & n6925 ) | ( n180 & n9748 ) | ( n6925 & n9748 ) ;
  assign n10662 = ( ~n1135 & n1829 ) | ( ~n1135 & n3288 ) | ( n1829 & n3288 ) ;
  assign n10663 = n10662 ^ n10023 ^ 1'b0 ;
  assign n10666 = n277 & ~n1213 ;
  assign n10665 = n8737 ^ n5416 ^ n1810 ;
  assign n10664 = n5048 ^ n2032 ^ n1619 ;
  assign n10667 = n10666 ^ n10665 ^ n10664 ;
  assign n10668 = ( n2185 & n8837 ) | ( n2185 & ~n10667 ) | ( n8837 & ~n10667 ) ;
  assign n10669 = ( n2602 & n7811 ) | ( n2602 & ~n10651 ) | ( n7811 & ~n10651 ) ;
  assign n10670 = n2692 ^ n187 ^ 1'b0 ;
  assign n10671 = ~n5097 & n10670 ;
  assign n10672 = n10671 ^ n2340 ^ 1'b0 ;
  assign n10673 = ( n802 & n3337 ) | ( n802 & n7757 ) | ( n3337 & n7757 ) ;
  assign n10674 = ( n1510 & n4080 ) | ( n1510 & ~n5213 ) | ( n4080 & ~n5213 ) ;
  assign n10675 = n10674 ^ n2541 ^ n2242 ;
  assign n10676 = ( n2151 & n10673 ) | ( n2151 & n10675 ) | ( n10673 & n10675 ) ;
  assign n10677 = ( n10669 & n10672 ) | ( n10669 & n10676 ) | ( n10672 & n10676 ) ;
  assign n10678 = ~n763 & n9573 ;
  assign n10679 = ~n2384 & n10678 ;
  assign n10682 = n5097 ^ n194 ^ 1'b0 ;
  assign n10681 = ( ~n3208 & n4467 ) | ( ~n3208 & n8042 ) | ( n4467 & n8042 ) ;
  assign n10680 = ( n1547 & n6560 ) | ( n1547 & n10524 ) | ( n6560 & n10524 ) ;
  assign n10683 = n10682 ^ n10681 ^ n10680 ;
  assign n10684 = ( n1728 & n5967 ) | ( n1728 & n9006 ) | ( n5967 & n9006 ) ;
  assign n10685 = ( n1447 & n8589 ) | ( n1447 & n10684 ) | ( n8589 & n10684 ) ;
  assign n10686 = n5037 & ~n9553 ;
  assign n10687 = n5034 ^ n1451 ^ n1141 ;
  assign n10688 = n8402 ^ n2931 ^ 1'b0 ;
  assign n10689 = ( n9854 & n10687 ) | ( n9854 & n10688 ) | ( n10687 & n10688 ) ;
  assign n10690 = ( n1666 & n1797 ) | ( n1666 & ~n6739 ) | ( n1797 & ~n6739 ) ;
  assign n10691 = n10690 ^ n8380 ^ n2482 ;
  assign n10692 = n10689 | n10691 ;
  assign n10693 = ( n780 & n3446 ) | ( n780 & n6871 ) | ( n3446 & n6871 ) ;
  assign n10694 = ( n306 & n6018 ) | ( n306 & n10693 ) | ( n6018 & n10693 ) ;
  assign n10695 = n524 & ~n1413 ;
  assign n10696 = ~n584 & n10695 ;
  assign n10697 = n10696 ^ n6189 ^ n1409 ;
  assign n10698 = n4076 & n10697 ;
  assign n10699 = n3485 ^ n3046 ^ 1'b0 ;
  assign n10700 = n2059 & ~n4064 ;
  assign n10701 = ~n10699 & n10700 ;
  assign n10702 = ~n4992 & n10149 ;
  assign n10703 = ( n259 & ~n4740 ) | ( n259 & n10702 ) | ( ~n4740 & n10702 ) ;
  assign n10704 = ( ~n10698 & n10701 ) | ( ~n10698 & n10703 ) | ( n10701 & n10703 ) ;
  assign n10705 = n3190 | n3320 ;
  assign n10706 = n10705 ^ n3638 ^ 1'b0 ;
  assign n10707 = ( n334 & ~n1639 ) | ( n334 & n4107 ) | ( ~n1639 & n4107 ) ;
  assign n10708 = ( n3823 & n10377 ) | ( n3823 & n10707 ) | ( n10377 & n10707 ) ;
  assign n10709 = ( n2542 & n10706 ) | ( n2542 & ~n10708 ) | ( n10706 & ~n10708 ) ;
  assign n10710 = n2230 & ~n5426 ;
  assign n10711 = ~n3032 & n10710 ;
  assign n10712 = n2430 | n4425 ;
  assign n10713 = n10711 & ~n10712 ;
  assign n10714 = n6483 ^ n4967 ^ n1885 ;
  assign n10715 = ~n458 & n4086 ;
  assign n10716 = ( n2608 & n10714 ) | ( n2608 & n10715 ) | ( n10714 & n10715 ) ;
  assign n10720 = n2428 ^ n2023 ^ 1'b0 ;
  assign n10721 = n10720 ^ n3998 ^ n2606 ;
  assign n10717 = n4116 ^ n3804 ^ 1'b0 ;
  assign n10718 = ~n194 & n10717 ;
  assign n10719 = n10718 ^ n8727 ^ n5031 ;
  assign n10722 = n10721 ^ n10719 ^ n7947 ;
  assign n10731 = n4819 ^ n552 ^ 1'b0 ;
  assign n10732 = n4028 & n10731 ;
  assign n10733 = n9277 & n10732 ;
  assign n10729 = n3319 ^ n963 ^ 1'b0 ;
  assign n10723 = x32 & ~n2351 ;
  assign n10724 = n10723 ^ n1390 ^ 1'b0 ;
  assign n10725 = ~n4834 & n10724 ;
  assign n10726 = n5455 & n7065 ;
  assign n10727 = ~n10725 & n10726 ;
  assign n10728 = n7613 & ~n10727 ;
  assign n10730 = n10729 ^ n10728 ^ 1'b0 ;
  assign n10734 = n10733 ^ n10730 ^ n3588 ;
  assign n10735 = n7256 & n8892 ;
  assign n10736 = ~n10734 & n10735 ;
  assign n10737 = ( ~n889 & n6740 ) | ( ~n889 & n10736 ) | ( n6740 & n10736 ) ;
  assign n10738 = ( n563 & n8946 ) | ( n563 & n9894 ) | ( n8946 & n9894 ) ;
  assign n10739 = ( n866 & n2116 ) | ( n866 & n7576 ) | ( n2116 & n7576 ) ;
  assign n10740 = n10739 ^ n10514 ^ n7779 ;
  assign n10741 = ~n1896 & n4292 ;
  assign n10742 = ~n1966 & n10741 ;
  assign n10743 = ~n1858 & n5172 ;
  assign n10748 = n3001 ^ x89 ^ 1'b0 ;
  assign n10744 = n7641 ^ n6008 ^ 1'b0 ;
  assign n10745 = n4480 ^ n347 ^ 1'b0 ;
  assign n10746 = ( n538 & n1442 ) | ( n538 & ~n10745 ) | ( n1442 & ~n10745 ) ;
  assign n10747 = ( n10196 & n10744 ) | ( n10196 & n10746 ) | ( n10744 & n10746 ) ;
  assign n10749 = n10748 ^ n10747 ^ n4137 ;
  assign n10750 = n4442 & ~n5609 ;
  assign n10751 = n10750 ^ n6251 ^ 1'b0 ;
  assign n10752 = ( ~n775 & n7705 ) | ( ~n775 & n10627 ) | ( n7705 & n10627 ) ;
  assign n10753 = ( n8947 & ~n9811 ) | ( n8947 & n10752 ) | ( ~n9811 & n10752 ) ;
  assign n10754 = n8833 ^ n5644 ^ n2474 ;
  assign n10755 = ( n649 & ~n6077 ) | ( n649 & n7494 ) | ( ~n6077 & n7494 ) ;
  assign n10756 = ( n2813 & n4121 ) | ( n2813 & n10755 ) | ( n4121 & n10755 ) ;
  assign n10757 = n10754 & n10756 ;
  assign n10758 = ( ~n680 & n2760 ) | ( ~n680 & n5651 ) | ( n2760 & n5651 ) ;
  assign n10759 = n5644 | n10758 ;
  assign n10760 = n10739 ^ n4114 ^ x18 ;
  assign n10761 = n10760 ^ n10418 ^ n4308 ;
  assign n10762 = n10761 ^ n6168 ^ n3083 ;
  assign n10763 = ( n2086 & n2465 ) | ( n2086 & ~n10206 ) | ( n2465 & ~n10206 ) ;
  assign n10764 = n4964 ^ n4386 ^ n141 ;
  assign n10765 = n2152 & ~n4850 ;
  assign n10766 = ( ~n8371 & n10764 ) | ( ~n8371 & n10765 ) | ( n10764 & n10765 ) ;
  assign n10767 = n10766 ^ n7927 ^ n3646 ;
  assign n10768 = ( n154 & ~n1775 ) | ( n154 & n4101 ) | ( ~n1775 & n4101 ) ;
  assign n10769 = n10768 ^ n10012 ^ n280 ;
  assign n10770 = ( n635 & n10767 ) | ( n635 & ~n10769 ) | ( n10767 & ~n10769 ) ;
  assign n10771 = ~n158 & n963 ;
  assign n10772 = n5259 & n10771 ;
  assign n10773 = n9510 ^ n7702 ^ n6628 ;
  assign n10774 = n10773 ^ n9898 ^ n3366 ;
  assign n10775 = ( n3166 & n10772 ) | ( n3166 & ~n10774 ) | ( n10772 & ~n10774 ) ;
  assign n10776 = n7968 & n10607 ;
  assign n10777 = n4209 & n10776 ;
  assign n10778 = ( n352 & n2340 ) | ( n352 & ~n10777 ) | ( n2340 & ~n10777 ) ;
  assign n10779 = n8663 & n10778 ;
  assign n10780 = ~n10071 & n10779 ;
  assign n10781 = n9115 ^ n4566 ^ n2401 ;
  assign n10782 = n5469 ^ n3924 ^ 1'b0 ;
  assign n10783 = ( n2801 & ~n10781 ) | ( n2801 & n10782 ) | ( ~n10781 & n10782 ) ;
  assign n10786 = n779 | n1964 ;
  assign n10784 = ( n773 & n2632 ) | ( n773 & ~n2946 ) | ( n2632 & ~n2946 ) ;
  assign n10785 = ( ~n1679 & n8202 ) | ( ~n1679 & n10784 ) | ( n8202 & n10784 ) ;
  assign n10787 = n10786 ^ n10785 ^ n10020 ;
  assign n10788 = ( x21 & n768 ) | ( x21 & ~n7680 ) | ( n768 & ~n7680 ) ;
  assign n10789 = ~n9941 & n10788 ;
  assign n10790 = n10789 ^ n5226 ^ 1'b0 ;
  assign n10791 = n10319 ^ n5659 ^ 1'b0 ;
  assign n10792 = n10791 ^ n5694 ^ n1462 ;
  assign n10793 = ~n5048 & n7398 ;
  assign n10794 = n10793 ^ n8345 ^ n5659 ;
  assign n10796 = n6938 ^ n4459 ^ n2498 ;
  assign n10795 = ( n4921 & n6352 ) | ( n4921 & ~n10559 ) | ( n6352 & ~n10559 ) ;
  assign n10797 = n10796 ^ n10795 ^ n6158 ;
  assign n10798 = n5300 | n9867 ;
  assign n10799 = n9558 ^ n5128 ^ 1'b0 ;
  assign n10800 = ( n3696 & n7415 ) | ( n3696 & n7501 ) | ( n7415 & n7501 ) ;
  assign n10801 = n3448 ^ n917 ^ 1'b0 ;
  assign n10802 = n10801 ^ n7132 ^ n3947 ;
  assign n10803 = ( n1956 & n2019 ) | ( n1956 & ~n6141 ) | ( n2019 & ~n6141 ) ;
  assign n10804 = ( n1351 & ~n7083 ) | ( n1351 & n10803 ) | ( ~n7083 & n10803 ) ;
  assign n10805 = n9326 ^ n1301 ^ 1'b0 ;
  assign n10806 = n1565 & ~n7429 ;
  assign n10807 = ( n1363 & n2315 ) | ( n1363 & n10806 ) | ( n2315 & n10806 ) ;
  assign n10808 = ( n7988 & n10805 ) | ( n7988 & n10807 ) | ( n10805 & n10807 ) ;
  assign n10809 = n10808 ^ n3794 ^ n2408 ;
  assign n10810 = n223 | n2309 ;
  assign n10811 = n10809 & ~n10810 ;
  assign n10812 = ~n684 & n9521 ;
  assign n10813 = n10812 ^ n1298 ^ 1'b0 ;
  assign n10820 = x103 & ~n4041 ;
  assign n10821 = ( ~n2156 & n8703 ) | ( ~n2156 & n10820 ) | ( n8703 & n10820 ) ;
  assign n10815 = n5546 ^ n5390 ^ 1'b0 ;
  assign n10816 = ~n6178 & n10815 ;
  assign n10817 = n10816 ^ n2542 ^ 1'b0 ;
  assign n10818 = ~n3807 & n10817 ;
  assign n10819 = ~n2386 & n10818 ;
  assign n10814 = n1838 & ~n2299 ;
  assign n10822 = n10821 ^ n10819 ^ n10814 ;
  assign n10824 = n3612 | n6561 ;
  assign n10825 = n10824 ^ n6939 ^ n3247 ;
  assign n10826 = n10825 ^ n7556 ^ n5788 ;
  assign n10823 = ( ~n5658 & n6304 ) | ( ~n5658 & n6850 ) | ( n6304 & n6850 ) ;
  assign n10827 = n10826 ^ n10823 ^ 1'b0 ;
  assign n10830 = n8588 ^ n3704 ^ n2646 ;
  assign n10829 = ( n467 & n2074 ) | ( n467 & n4357 ) | ( n2074 & n4357 ) ;
  assign n10828 = n1734 & ~n7689 ;
  assign n10831 = n10830 ^ n10829 ^ n10828 ;
  assign n10832 = n10831 ^ n541 ^ 1'b0 ;
  assign n10833 = n5286 & n10832 ;
  assign n10834 = n10101 ^ n176 ^ 1'b0 ;
  assign n10835 = n9237 ^ n7135 ^ n5680 ;
  assign n10836 = n10835 ^ n7868 ^ n5558 ;
  assign n10837 = n10836 ^ n8087 ^ n2803 ;
  assign n10838 = n8533 ^ n8025 ^ n6493 ;
  assign n10839 = n2821 | n10838 ;
  assign n10840 = n6785 & ~n10839 ;
  assign n10841 = n10312 ^ n7342 ^ 1'b0 ;
  assign n10846 = ( ~n301 & n1931 ) | ( ~n301 & n2045 ) | ( n1931 & n2045 ) ;
  assign n10842 = ~n4059 & n5245 ;
  assign n10843 = ~n1107 & n1972 ;
  assign n10844 = n10843 ^ n7607 ^ n7002 ;
  assign n10845 = ( n10535 & ~n10842 ) | ( n10535 & n10844 ) | ( ~n10842 & n10844 ) ;
  assign n10847 = n10846 ^ n10845 ^ n9736 ;
  assign n10848 = n4770 ^ n3482 ^ 1'b0 ;
  assign n10849 = n6829 ^ n679 ^ 1'b0 ;
  assign n10850 = n10848 & n10849 ;
  assign n10851 = n6778 & n7351 ;
  assign n10852 = n5833 & n10851 ;
  assign n10853 = ( n5848 & n6476 ) | ( n5848 & ~n10852 ) | ( n6476 & ~n10852 ) ;
  assign n10854 = ~n3990 & n9790 ;
  assign n10855 = ~n200 & n10854 ;
  assign n10856 = n10855 ^ n7088 ^ n5927 ;
  assign n10858 = n7620 ^ n7406 ^ 1'b0 ;
  assign n10859 = n624 | n6251 ;
  assign n10860 = n10858 | n10859 ;
  assign n10857 = ( n1932 & n6287 ) | ( n1932 & ~n10609 ) | ( n6287 & ~n10609 ) ;
  assign n10861 = n10860 ^ n10857 ^ n4670 ;
  assign n10862 = ( n4128 & ~n10856 ) | ( n4128 & n10861 ) | ( ~n10856 & n10861 ) ;
  assign n10865 = n784 | n4611 ;
  assign n10866 = n2314 & ~n10865 ;
  assign n10867 = n10866 ^ n5996 ^ 1'b0 ;
  assign n10868 = ~n10560 & n10867 ;
  assign n10863 = n4732 & n7809 ;
  assign n10864 = ~n4271 & n10863 ;
  assign n10869 = n10868 ^ n10864 ^ x59 ;
  assign n10870 = n633 & n6562 ;
  assign n10871 = n4515 & n10870 ;
  assign n10872 = ~n925 & n954 ;
  assign n10873 = n10872 ^ n8263 ^ 1'b0 ;
  assign n10874 = n10297 ^ n9407 ^ 1'b0 ;
  assign n10875 = n5525 ^ n4039 ^ 1'b0 ;
  assign n10876 = n10875 ^ n4134 ^ n3970 ;
  assign n10877 = n1239 & ~n10876 ;
  assign n10878 = ~n9420 & n10877 ;
  assign n10879 = n1148 & ~n10878 ;
  assign n10880 = n10879 ^ n6996 ^ 1'b0 ;
  assign n10881 = ( n864 & ~n3301 ) | ( n864 & n10880 ) | ( ~n3301 & n10880 ) ;
  assign n10882 = n465 & n8692 ;
  assign n10883 = n10882 ^ n146 ^ 1'b0 ;
  assign n10884 = ( n2818 & n8956 ) | ( n2818 & n10883 ) | ( n8956 & n10883 ) ;
  assign n10885 = ( n2090 & n7990 ) | ( n2090 & ~n10884 ) | ( n7990 & ~n10884 ) ;
  assign n10886 = n3489 ^ n2625 ^ 1'b0 ;
  assign n10887 = ( ~n270 & n8016 ) | ( ~n270 & n10886 ) | ( n8016 & n10886 ) ;
  assign n10888 = n10887 ^ x10 ^ 1'b0 ;
  assign n10892 = n4077 ^ n2464 ^ n1739 ;
  assign n10891 = ( ~n1519 & n1965 ) | ( ~n1519 & n1977 ) | ( n1965 & n1977 ) ;
  assign n10889 = n4307 ^ n1698 ^ 1'b0 ;
  assign n10890 = x32 & n10889 ;
  assign n10893 = n10892 ^ n10891 ^ n10890 ;
  assign n10894 = x80 & n10893 ;
  assign n10895 = n10888 & n10894 ;
  assign n10896 = n5637 ^ n337 ^ 1'b0 ;
  assign n10897 = n2679 | n3307 ;
  assign n10898 = n3311 | n10897 ;
  assign n10902 = ~n2679 & n6298 ;
  assign n10903 = n2817 & n10902 ;
  assign n10899 = ( n666 & n1226 ) | ( n666 & n3544 ) | ( n1226 & n3544 ) ;
  assign n10900 = ( n4421 & ~n7583 ) | ( n4421 & n10899 ) | ( ~n7583 & n10899 ) ;
  assign n10901 = n4377 | n10900 ;
  assign n10904 = n10903 ^ n10901 ^ n6916 ;
  assign n10905 = n10904 ^ n10845 ^ n4230 ;
  assign n10906 = n5565 & n9179 ;
  assign n10907 = ( n347 & n7615 ) | ( n347 & ~n10906 ) | ( n7615 & ~n10906 ) ;
  assign n10908 = ( n2555 & n8229 ) | ( n2555 & ~n10907 ) | ( n8229 & ~n10907 ) ;
  assign n10910 = n5702 ^ n5169 ^ 1'b0 ;
  assign n10909 = n702 & ~n1806 ;
  assign n10911 = n10910 ^ n10909 ^ n1747 ;
  assign n10912 = n5095 & ~n8449 ;
  assign n10913 = ~n4322 & n10912 ;
  assign n10914 = n10913 ^ n2619 ^ 1'b0 ;
  assign n10919 = n1794 | n7944 ;
  assign n10920 = n10919 ^ n3676 ^ n3405 ;
  assign n10921 = n1012 & ~n10920 ;
  assign n10915 = n8393 ^ n3066 ^ 1'b0 ;
  assign n10916 = n2523 | n10915 ;
  assign n10917 = n499 & ~n10916 ;
  assign n10918 = n6392 & n10917 ;
  assign n10922 = n10921 ^ n10918 ^ 1'b0 ;
  assign n10924 = n486 & ~n3686 ;
  assign n10925 = n10924 ^ x5 ^ 1'b0 ;
  assign n10926 = n10925 ^ n6657 ^ n1638 ;
  assign n10923 = n1982 & n4148 ;
  assign n10927 = n10926 ^ n10923 ^ 1'b0 ;
  assign n10930 = n8052 ^ n3929 ^ n320 ;
  assign n10928 = n369 | n8340 ;
  assign n10929 = n10928 ^ n5510 ^ 1'b0 ;
  assign n10931 = n10930 ^ n10929 ^ n3049 ;
  assign n10932 = n5813 & ~n7341 ;
  assign n10933 = n4770 & n10932 ;
  assign n10934 = n10933 ^ n7543 ^ n4012 ;
  assign n10935 = n10934 ^ n10412 ^ n4132 ;
  assign n10936 = n1428 ^ n355 ^ 1'b0 ;
  assign n10937 = n9771 | n10936 ;
  assign n10938 = n10937 ^ n1184 ^ n333 ;
  assign n10939 = n8073 & n10938 ;
  assign n10940 = ~n5324 & n10939 ;
  assign n10941 = n10940 ^ n6167 ^ n4229 ;
  assign n10942 = n2799 | n5186 ;
  assign n10943 = n10942 ^ n9938 ^ n3268 ;
  assign n10944 = ( n6927 & n10941 ) | ( n6927 & ~n10943 ) | ( n10941 & ~n10943 ) ;
  assign n10945 = n4027 ^ x3 ^ 1'b0 ;
  assign n10946 = n10945 ^ n5942 ^ 1'b0 ;
  assign n10947 = n10946 ^ n5935 ^ 1'b0 ;
  assign n10948 = n2942 & n6677 ;
  assign n10949 = n10948 ^ n2391 ^ 1'b0 ;
  assign n10950 = n2550 & ~n10949 ;
  assign n10951 = n10950 ^ n4072 ^ 1'b0 ;
  assign n10952 = ( n3955 & ~n6213 ) | ( n3955 & n6540 ) | ( ~n6213 & n6540 ) ;
  assign n10953 = ~n1719 & n9848 ;
  assign n10954 = n10953 ^ n6565 ^ 1'b0 ;
  assign n10955 = ( n2951 & ~n3989 ) | ( n2951 & n10954 ) | ( ~n3989 & n10954 ) ;
  assign n10956 = n10952 & n10955 ;
  assign n10957 = ~n10411 & n10956 ;
  assign n10958 = n10957 ^ n6013 ^ 1'b0 ;
  assign n10961 = ( n200 & n1052 ) | ( n200 & n5462 ) | ( n1052 & n5462 ) ;
  assign n10959 = n3984 ^ n3355 ^ n3139 ;
  assign n10960 = n2710 | n10959 ;
  assign n10962 = n10961 ^ n10960 ^ 1'b0 ;
  assign n10963 = n5144 ^ n4839 ^ n4446 ;
  assign n10964 = n10962 | n10963 ;
  assign n10965 = ~n916 & n9719 ;
  assign n10966 = n10965 ^ n904 ^ 1'b0 ;
  assign n10967 = n10966 ^ n6428 ^ 1'b0 ;
  assign n10968 = n6733 ^ n6103 ^ n5071 ;
  assign n10969 = n3854 ^ n3161 ^ 1'b0 ;
  assign n10970 = n6601 | n10969 ;
  assign n10971 = ( n2309 & ~n7680 ) | ( n2309 & n9662 ) | ( ~n7680 & n9662 ) ;
  assign n10973 = ~n236 & n2900 ;
  assign n10972 = n2707 & ~n6639 ;
  assign n10974 = n10973 ^ n10972 ^ 1'b0 ;
  assign n10975 = n5416 ^ n4236 ^ n706 ;
  assign n10976 = ( ~n3145 & n6389 ) | ( ~n3145 & n10975 ) | ( n6389 & n10975 ) ;
  assign n10977 = n6399 ^ n1688 ^ 1'b0 ;
  assign n10978 = n4971 | n10977 ;
  assign n10979 = ~n10976 & n10978 ;
  assign n10980 = n9850 | n10979 ;
  assign n10981 = n10974 | n10980 ;
  assign n10982 = ( n4659 & ~n4802 ) | ( n4659 & n10981 ) | ( ~n4802 & n10981 ) ;
  assign n10991 = ( n779 & ~n1359 ) | ( n779 & n7812 ) | ( ~n1359 & n7812 ) ;
  assign n10985 = ~n1079 & n1117 ;
  assign n10986 = n10985 ^ n5549 ^ n4053 ;
  assign n10987 = ~n3480 & n10986 ;
  assign n10988 = n10987 ^ n2013 ^ 1'b0 ;
  assign n10989 = n10988 ^ n1969 ^ 1'b0 ;
  assign n10990 = n2446 | n10989 ;
  assign n10983 = n6765 ^ n1428 ^ 1'b0 ;
  assign n10984 = n3104 & n10983 ;
  assign n10992 = n10991 ^ n10990 ^ n10984 ;
  assign n10993 = n7553 ^ n1566 ^ 1'b0 ;
  assign n10994 = n10993 ^ n5272 ^ n4628 ;
  assign n10995 = ( n6868 & n9173 ) | ( n6868 & ~n9257 ) | ( n9173 & ~n9257 ) ;
  assign n10996 = ( x9 & n1739 ) | ( x9 & ~n3772 ) | ( n1739 & ~n3772 ) ;
  assign n10997 = n10996 ^ n8507 ^ n1579 ;
  assign n10998 = ( ~n1092 & n10995 ) | ( ~n1092 & n10997 ) | ( n10995 & n10997 ) ;
  assign n10999 = n10998 ^ n2534 ^ n1377 ;
  assign n11000 = n10760 ^ n10636 ^ n5919 ;
  assign n11001 = n190 | n4003 ;
  assign n11002 = n5132 | n11001 ;
  assign n11003 = n1382 & n11002 ;
  assign n11004 = n157 & n11003 ;
  assign n11005 = n3130 ^ n1682 ^ 1'b0 ;
  assign n11006 = n1781 ^ n733 ^ 1'b0 ;
  assign n11007 = n523 & n11006 ;
  assign n11008 = n11007 ^ n10026 ^ 1'b0 ;
  assign n11009 = n5100 ^ x27 ^ 1'b0 ;
  assign n11010 = ( x18 & n10253 ) | ( x18 & ~n11009 ) | ( n10253 & ~n11009 ) ;
  assign n11011 = n11010 ^ n8954 ^ 1'b0 ;
  assign n11012 = x96 & n3018 ;
  assign n11013 = ( n6825 & ~n7135 ) | ( n6825 & n11012 ) | ( ~n7135 & n11012 ) ;
  assign n11014 = n11013 ^ n7913 ^ n2517 ;
  assign n11015 = ( n1248 & n2934 ) | ( n1248 & ~n6280 ) | ( n2934 & ~n6280 ) ;
  assign n11016 = n11015 ^ n8734 ^ n4781 ;
  assign n11017 = n5383 & n11016 ;
  assign n11018 = n11017 ^ n5740 ^ 1'b0 ;
  assign n11019 = ( n549 & ~n8495 ) | ( n549 & n10597 ) | ( ~n8495 & n10597 ) ;
  assign n11020 = ~n3602 & n8666 ;
  assign n11021 = n11019 & n11020 ;
  assign n11022 = n913 | n5659 ;
  assign n11023 = n11022 ^ n6120 ^ 1'b0 ;
  assign n11024 = n11023 ^ n5160 ^ n2650 ;
  assign n11025 = ( ~n2617 & n4918 ) | ( ~n2617 & n11024 ) | ( n4918 & n11024 ) ;
  assign n11026 = ( ~n10701 & n10702 ) | ( ~n10701 & n11025 ) | ( n10702 & n11025 ) ;
  assign n11027 = n11026 ^ n9687 ^ n8617 ;
  assign n11028 = n8520 ^ n6495 ^ 1'b0 ;
  assign n11029 = n11028 ^ n5948 ^ 1'b0 ;
  assign n11030 = n6840 & n11029 ;
  assign n11031 = ( x63 & n3671 ) | ( x63 & ~n11030 ) | ( n3671 & ~n11030 ) ;
  assign n11032 = n8729 ^ n6407 ^ n1692 ;
  assign n11033 = n1212 ^ n910 ^ 1'b0 ;
  assign n11034 = n11033 ^ n1304 ^ 1'b0 ;
  assign n11035 = ~n11032 & n11034 ;
  assign n11036 = n11035 ^ n5220 ^ 1'b0 ;
  assign n11037 = n2695 & ~n7280 ;
  assign n11038 = ~n7233 & n11037 ;
  assign n11039 = n4592 ^ n2418 ^ 1'b0 ;
  assign n11040 = ~n11038 & n11039 ;
  assign n11041 = ~n6298 & n9143 ;
  assign n11042 = ( n3319 & n6388 ) | ( n3319 & n11041 ) | ( n6388 & n11041 ) ;
  assign n11043 = ( n5782 & n11040 ) | ( n5782 & n11042 ) | ( n11040 & n11042 ) ;
  assign n11044 = ~n8746 & n8748 ;
  assign n11045 = ( n1875 & n2176 ) | ( n1875 & ~n2721 ) | ( n2176 & ~n2721 ) ;
  assign n11046 = ~n8200 & n9701 ;
  assign n11047 = n4933 & n11046 ;
  assign n11048 = ( n8394 & n11045 ) | ( n8394 & ~n11047 ) | ( n11045 & ~n11047 ) ;
  assign n11049 = n10920 ^ n7601 ^ n2140 ;
  assign n11052 = ( n2206 & n7511 ) | ( n2206 & ~n9534 ) | ( n7511 & ~n9534 ) ;
  assign n11050 = n1442 & n9738 ;
  assign n11051 = n11050 ^ n9787 ^ 1'b0 ;
  assign n11053 = n11052 ^ n11051 ^ n2511 ;
  assign n11054 = n3036 ^ n387 ^ 1'b0 ;
  assign n11055 = ~n6508 & n11054 ;
  assign n11056 = n11055 ^ n4789 ^ n3697 ;
  assign n11057 = ( n1551 & n5589 ) | ( n1551 & ~n10962 ) | ( n5589 & ~n10962 ) ;
  assign n11058 = ( ~n3126 & n8696 ) | ( ~n3126 & n9277 ) | ( n8696 & n9277 ) ;
  assign n11059 = ~n1556 & n11058 ;
  assign n11060 = n11059 ^ n10445 ^ n1815 ;
  assign n11061 = ( n1573 & ~n3766 ) | ( n1573 & n4190 ) | ( ~n3766 & n4190 ) ;
  assign n11062 = ( n955 & n1706 ) | ( n955 & n11061 ) | ( n1706 & n11061 ) ;
  assign n11063 = ( n4340 & n8393 ) | ( n4340 & ~n11062 ) | ( n8393 & ~n11062 ) ;
  assign n11067 = n365 & n2124 ;
  assign n11064 = ( n1220 & ~n3259 ) | ( n1220 & n3587 ) | ( ~n3259 & n3587 ) ;
  assign n11065 = x0 & n690 ;
  assign n11066 = n11064 & ~n11065 ;
  assign n11068 = n11067 ^ n11066 ^ 1'b0 ;
  assign n11069 = n2250 & ~n11068 ;
  assign n11070 = ( n617 & ~n11063 ) | ( n617 & n11069 ) | ( ~n11063 & n11069 ) ;
  assign n11071 = n7100 ^ n293 ^ 1'b0 ;
  assign n11072 = n5578 ^ n4921 ^ n1679 ;
  assign n11073 = n11072 ^ n3738 ^ n1136 ;
  assign n11080 = n5124 ^ n3601 ^ n1158 ;
  assign n11075 = ( ~n2557 & n2816 ) | ( ~n2557 & n4590 ) | ( n2816 & n4590 ) ;
  assign n11076 = n2961 | n3941 ;
  assign n11077 = n1334 & ~n11076 ;
  assign n11078 = ( n4577 & n5655 ) | ( n4577 & n11077 ) | ( n5655 & n11077 ) ;
  assign n11079 = ( n9238 & n11075 ) | ( n9238 & n11078 ) | ( n11075 & n11078 ) ;
  assign n11074 = n7678 ^ n2135 ^ 1'b0 ;
  assign n11081 = n11080 ^ n11079 ^ n11074 ;
  assign n11082 = n809 | n8769 ;
  assign n11083 = n10151 & ~n11082 ;
  assign n11084 = n11083 ^ n6504 ^ 1'b0 ;
  assign n11085 = ~n1254 & n8813 ;
  assign n11086 = ~x99 & n11085 ;
  assign n11087 = n11086 ^ n3624 ^ n1125 ;
  assign n11088 = ~n1929 & n11087 ;
  assign n11089 = ( n1673 & n9618 ) | ( n1673 & n9841 ) | ( n9618 & n9841 ) ;
  assign n11090 = n11089 ^ n2097 ^ n1839 ;
  assign n11092 = n482 ^ x3 ^ 1'b0 ;
  assign n11093 = n326 & n11092 ;
  assign n11091 = ~n2041 & n5677 ;
  assign n11094 = n11093 ^ n11091 ^ n3768 ;
  assign n11095 = n9036 & n11094 ;
  assign n11096 = n11095 ^ n7288 ^ 1'b0 ;
  assign n11097 = n11090 & n11096 ;
  assign n11098 = ( ~n3600 & n4039 ) | ( ~n3600 & n7120 ) | ( n4039 & n7120 ) ;
  assign n11099 = ~n2348 & n4713 ;
  assign n11100 = ( n1607 & n2452 ) | ( n1607 & ~n6222 ) | ( n2452 & ~n6222 ) ;
  assign n11101 = n11100 ^ n5449 ^ n1802 ;
  assign n11102 = n3117 ^ n670 ^ 1'b0 ;
  assign n11103 = x2 & n11102 ;
  assign n11104 = n10520 & n11103 ;
  assign n11105 = n6740 ^ n5334 ^ n324 ;
  assign n11106 = n7088 ^ n7082 ^ n976 ;
  assign n11111 = n1828 | n2701 ;
  assign n11107 = n10582 ^ n986 ^ 1'b0 ;
  assign n11108 = n935 & ~n11107 ;
  assign n11109 = n6943 ^ n2720 ^ 1'b0 ;
  assign n11110 = n11108 & ~n11109 ;
  assign n11112 = n11111 ^ n11110 ^ n6649 ;
  assign n11113 = n11112 ^ n267 ^ 1'b0 ;
  assign n11114 = ( n11105 & ~n11106 ) | ( n11105 & n11113 ) | ( ~n11106 & n11113 ) ;
  assign n11115 = ( ~n425 & n741 ) | ( ~n425 & n4625 ) | ( n741 & n4625 ) ;
  assign n11116 = n1645 | n9838 ;
  assign n11117 = n11115 & ~n11116 ;
  assign n11118 = n146 & n10196 ;
  assign n11119 = n1378 & n8981 ;
  assign n11120 = n11119 ^ n4702 ^ 1'b0 ;
  assign n11121 = n11120 ^ n8312 ^ n2214 ;
  assign n11122 = n1007 & n11121 ;
  assign n11123 = ~n11118 & n11122 ;
  assign n11124 = n1092 | n9933 ;
  assign n11127 = n1262 ^ n321 ^ 1'b0 ;
  assign n11128 = n10299 & ~n11127 ;
  assign n11125 = n1833 & n2401 ;
  assign n11126 = n11125 ^ n5385 ^ 1'b0 ;
  assign n11129 = n11128 ^ n11126 ^ n2227 ;
  assign n11130 = ( n2561 & n5442 ) | ( n2561 & n11129 ) | ( n5442 & n11129 ) ;
  assign n11131 = n4830 ^ n3495 ^ n853 ;
  assign n11134 = ( n463 & n807 ) | ( n463 & n4873 ) | ( n807 & n4873 ) ;
  assign n11132 = n1751 & ~n4269 ;
  assign n11133 = n11132 ^ n7383 ^ 1'b0 ;
  assign n11135 = n11134 ^ n11133 ^ 1'b0 ;
  assign n11136 = n11131 & n11135 ;
  assign n11137 = n10934 & n11136 ;
  assign n11139 = n10690 ^ n3300 ^ n735 ;
  assign n11140 = n11139 ^ n4067 ^ n2777 ;
  assign n11138 = ~n466 & n8571 ;
  assign n11141 = n11140 ^ n11138 ^ 1'b0 ;
  assign n11143 = n3410 & n5741 ;
  assign n11144 = ~x27 & n11143 ;
  assign n11142 = ( n2550 & n3328 ) | ( n2550 & n3667 ) | ( n3328 & n3667 ) ;
  assign n11145 = n11144 ^ n11142 ^ 1'b0 ;
  assign n11148 = n462 & n8881 ;
  assign n11146 = n2877 ^ n2066 ^ n1321 ;
  assign n11147 = n11146 ^ n8811 ^ n3461 ;
  assign n11149 = n11148 ^ n11147 ^ n1181 ;
  assign n11150 = ( n357 & n4095 ) | ( n357 & ~n7791 ) | ( n4095 & ~n7791 ) ;
  assign n11151 = n11150 ^ n1259 ^ 1'b0 ;
  assign n11152 = ~n6251 & n11151 ;
  assign n11153 = n11152 ^ n3533 ^ 1'b0 ;
  assign n11154 = n11153 ^ n10406 ^ n831 ;
  assign n11168 = x109 & ~n2517 ;
  assign n11169 = n2863 & n11168 ;
  assign n11170 = ( n2692 & n5848 ) | ( n2692 & ~n6088 ) | ( n5848 & ~n6088 ) ;
  assign n11171 = n4381 | n11170 ;
  assign n11172 = n189 | n11171 ;
  assign n11173 = n11172 ^ n547 ^ 1'b0 ;
  assign n11174 = n11169 & n11173 ;
  assign n11155 = ( ~n1614 & n1865 ) | ( ~n1614 & n3778 ) | ( n1865 & n3778 ) ;
  assign n11156 = n377 & n6667 ;
  assign n11157 = ~n11155 & n11156 ;
  assign n11158 = n11157 ^ n1560 ^ 1'b0 ;
  assign n11159 = n6578 | n11158 ;
  assign n11160 = ( n1369 & ~n2677 ) | ( n1369 & n3425 ) | ( ~n2677 & n3425 ) ;
  assign n11161 = ( n1643 & n4015 ) | ( n1643 & n5469 ) | ( n4015 & n5469 ) ;
  assign n11163 = ( ~n4971 & n5315 ) | ( ~n4971 & n7268 ) | ( n5315 & n7268 ) ;
  assign n11162 = n719 & ~n4410 ;
  assign n11164 = n11163 ^ n11162 ^ 1'b0 ;
  assign n11165 = n11161 & n11164 ;
  assign n11166 = ~n11160 & n11165 ;
  assign n11167 = n11159 | n11166 ;
  assign n11175 = n11174 ^ n11167 ^ 1'b0 ;
  assign n11176 = ( n3652 & n10575 ) | ( n3652 & n11095 ) | ( n10575 & n11095 ) ;
  assign n11177 = n3291 ^ n840 ^ 1'b0 ;
  assign n11178 = n6914 & n10525 ;
  assign n11179 = ( n1977 & n4591 ) | ( n1977 & ~n7560 ) | ( n4591 & ~n7560 ) ;
  assign n11180 = n11179 ^ n9123 ^ n8970 ;
  assign n11181 = n8837 | n11180 ;
  assign n11182 = ( n5885 & n11178 ) | ( n5885 & n11181 ) | ( n11178 & n11181 ) ;
  assign n11183 = n11177 & n11182 ;
  assign n11184 = n9452 ^ n545 ^ n315 ;
  assign n11185 = n917 & n7443 ;
  assign n11186 = ( ~n1042 & n2225 ) | ( ~n1042 & n11185 ) | ( n2225 & n11185 ) ;
  assign n11187 = n5256 ^ n508 ^ 1'b0 ;
  assign n11188 = n10638 | n11187 ;
  assign n11189 = n5075 ^ n3728 ^ 1'b0 ;
  assign n11190 = n8454 & n11108 ;
  assign n11191 = ~n11189 & n11190 ;
  assign n11192 = n11191 ^ n9526 ^ n3178 ;
  assign n11193 = n9479 ^ n5003 ^ n1221 ;
  assign n11194 = n545 ^ n172 ^ 1'b0 ;
  assign n11195 = n11194 ^ n8394 ^ n2838 ;
  assign n11196 = n393 | n7844 ;
  assign n11197 = n3485 ^ x63 ^ 1'b0 ;
  assign n11198 = n11197 ^ n3469 ^ n1528 ;
  assign n11199 = ( n3140 & ~n4812 ) | ( n3140 & n11198 ) | ( ~n4812 & n11198 ) ;
  assign n11200 = ~n5525 & n11199 ;
  assign n11201 = ~n9112 & n11200 ;
  assign n11208 = n7265 ^ n1341 ^ 1'b0 ;
  assign n11205 = ( n3202 & n3830 ) | ( n3202 & ~n6120 ) | ( n3830 & ~n6120 ) ;
  assign n11203 = n8556 & ~n9140 ;
  assign n11204 = n11203 ^ n6622 ^ 1'b0 ;
  assign n11206 = n11205 ^ n11204 ^ n8556 ;
  assign n11202 = n5817 ^ n3339 ^ 1'b0 ;
  assign n11207 = n11206 ^ n11202 ^ n8435 ;
  assign n11209 = n11208 ^ n11207 ^ n9945 ;
  assign n11210 = ( n2125 & n5842 ) | ( n2125 & ~n8316 ) | ( n5842 & ~n8316 ) ;
  assign n11211 = ( n252 & ~n697 ) | ( n252 & n1951 ) | ( ~n697 & n1951 ) ;
  assign n11212 = ( ~n3494 & n8519 ) | ( ~n3494 & n11211 ) | ( n8519 & n11211 ) ;
  assign n11213 = ( n4279 & n11210 ) | ( n4279 & ~n11212 ) | ( n11210 & ~n11212 ) ;
  assign n11214 = ~n10349 & n11213 ;
  assign n11215 = n1946 & n7549 ;
  assign n11216 = n11215 ^ n2065 ^ 1'b0 ;
  assign n11217 = ( n4100 & n4538 ) | ( n4100 & ~n11216 ) | ( n4538 & ~n11216 ) ;
  assign n11218 = n8317 ^ n3130 ^ 1'b0 ;
  assign n11219 = n7724 ^ n2191 ^ n2149 ;
  assign n11220 = ( n510 & ~n3009 ) | ( n510 & n11219 ) | ( ~n3009 & n11219 ) ;
  assign n11221 = ( ~n7706 & n11218 ) | ( ~n7706 & n11220 ) | ( n11218 & n11220 ) ;
  assign n11222 = n5945 ^ n1291 ^ 1'b0 ;
  assign n11223 = n11222 ^ n6551 ^ 1'b0 ;
  assign n11224 = n6424 & ~n11223 ;
  assign n11225 = n9029 ^ n7427 ^ n2337 ;
  assign n11230 = n2139 ^ n1034 ^ 1'b0 ;
  assign n11231 = n7497 & ~n11230 ;
  assign n11226 = n2116 & n5149 ;
  assign n11227 = n11226 ^ n4365 ^ 1'b0 ;
  assign n11228 = ~n6364 & n11227 ;
  assign n11229 = n11228 ^ n1343 ^ 1'b0 ;
  assign n11232 = n11231 ^ n11229 ^ n5083 ;
  assign n11233 = ( n4292 & n11225 ) | ( n4292 & n11232 ) | ( n11225 & n11232 ) ;
  assign n11234 = ( n354 & ~n2799 ) | ( n354 & n4588 ) | ( ~n2799 & n4588 ) ;
  assign n11235 = n9510 ^ n1537 ^ n1386 ;
  assign n11236 = n2247 | n11235 ;
  assign n11237 = ( ~n1867 & n11234 ) | ( ~n1867 & n11236 ) | ( n11234 & n11236 ) ;
  assign n11238 = n4178 & ~n4475 ;
  assign n11239 = n11140 ^ n6013 ^ n259 ;
  assign n11240 = ~n9488 & n11239 ;
  assign n11241 = n2763 ^ n2179 ^ n1133 ;
  assign n11242 = ( n902 & ~n6354 ) | ( n902 & n11241 ) | ( ~n6354 & n11241 ) ;
  assign n11243 = ( n4484 & n5514 ) | ( n4484 & n6622 ) | ( n5514 & n6622 ) ;
  assign n11244 = ( ~n1710 & n8906 ) | ( ~n1710 & n11243 ) | ( n8906 & n11243 ) ;
  assign n11245 = n7882 ^ n217 ^ 1'b0 ;
  assign n11246 = n2126 | n11245 ;
  assign n11247 = n11246 ^ n7230 ^ n831 ;
  assign n11248 = n7260 & ~n11247 ;
  assign n11254 = ~n2800 & n3600 ;
  assign n11255 = n11254 ^ n2163 ^ 1'b0 ;
  assign n11249 = n7431 ^ n1740 ^ n1647 ;
  assign n11250 = n11249 ^ n6456 ^ x119 ;
  assign n11251 = n6933 ^ n6887 ^ 1'b0 ;
  assign n11252 = n11250 & n11251 ;
  assign n11253 = ~n2770 & n11252 ;
  assign n11256 = n11255 ^ n11253 ^ 1'b0 ;
  assign n11257 = ~n791 & n3955 ;
  assign n11258 = n11257 ^ n1400 ^ 1'b0 ;
  assign n11259 = n6918 ^ n1780 ^ 1'b0 ;
  assign n11260 = n6181 | n11259 ;
  assign n11261 = ( ~n649 & n11258 ) | ( ~n649 & n11260 ) | ( n11258 & n11260 ) ;
  assign n11262 = n8692 ^ n8319 ^ n3234 ;
  assign n11263 = n1441 & n11262 ;
  assign n11264 = n805 & n11263 ;
  assign n11265 = ( ~n8652 & n10246 ) | ( ~n8652 & n11264 ) | ( n10246 & n11264 ) ;
  assign n11266 = ~n690 & n7857 ;
  assign n11267 = n11266 ^ n2679 ^ 1'b0 ;
  assign n11268 = n1490 & n1963 ;
  assign n11269 = ~n11267 & n11268 ;
  assign n11274 = n8402 ^ n7495 ^ 1'b0 ;
  assign n11275 = ~n5586 & n11274 ;
  assign n11276 = n11275 ^ n4879 ^ n4008 ;
  assign n11277 = n6833 | n11276 ;
  assign n11270 = ( n870 & ~n1162 ) | ( n870 & n2335 ) | ( ~n1162 & n2335 ) ;
  assign n11271 = n11270 ^ n7683 ^ n3953 ;
  assign n11272 = n8676 ^ n6707 ^ n3665 ;
  assign n11273 = ~n11271 & n11272 ;
  assign n11278 = n11277 ^ n11273 ^ n8983 ;
  assign n11279 = n11278 ^ n9817 ^ n2790 ;
  assign n11280 = n7334 ^ n2524 ^ 1'b0 ;
  assign n11281 = ( n234 & ~n7775 ) | ( n234 & n11280 ) | ( ~n7775 & n11280 ) ;
  assign n11282 = n7243 ^ n1929 ^ 1'b0 ;
  assign n11283 = n2665 & n11282 ;
  assign n11284 = n11283 ^ n10867 ^ 1'b0 ;
  assign n11285 = n201 | n11284 ;
  assign n11286 = ( n1959 & ~n6860 ) | ( n1959 & n10559 ) | ( ~n6860 & n10559 ) ;
  assign n11287 = ~n8314 & n11286 ;
  assign n11288 = n11285 & n11287 ;
  assign n11289 = n7605 ^ n7314 ^ 1'b0 ;
  assign n11290 = n2842 & ~n11289 ;
  assign n11291 = n10690 ^ n5241 ^ 1'b0 ;
  assign n11292 = ( n1561 & n6760 ) | ( n1561 & ~n11291 ) | ( n6760 & ~n11291 ) ;
  assign n11293 = n11292 ^ n7683 ^ 1'b0 ;
  assign n11294 = ( ~n1972 & n10179 ) | ( ~n1972 & n10607 ) | ( n10179 & n10607 ) ;
  assign n11295 = n7350 ^ n4634 ^ 1'b0 ;
  assign n11296 = n3024 & ~n11295 ;
  assign n11297 = ( n1911 & n4851 ) | ( n1911 & n11296 ) | ( n4851 & n11296 ) ;
  assign n11298 = ( n6260 & ~n9935 ) | ( n6260 & n11297 ) | ( ~n9935 & n11297 ) ;
  assign n11299 = n5053 ^ n3888 ^ n2371 ;
  assign n11300 = ( n4022 & n6396 ) | ( n4022 & n11009 ) | ( n6396 & n11009 ) ;
  assign n11301 = n4349 & n11300 ;
  assign n11302 = n7564 ^ n4583 ^ 1'b0 ;
  assign n11303 = ~n482 & n4855 ;
  assign n11304 = ( n1751 & n8207 ) | ( n1751 & n11303 ) | ( n8207 & n11303 ) ;
  assign n11305 = n9014 ^ n7337 ^ n5761 ;
  assign n11306 = n3265 ^ n1795 ^ n267 ;
  assign n11307 = ( n11304 & n11305 ) | ( n11304 & n11306 ) | ( n11305 & n11306 ) ;
  assign n11308 = n2220 & n8085 ;
  assign n11309 = ~n9712 & n11308 ;
  assign n11310 = n5364 ^ n3704 ^ 1'b0 ;
  assign n11311 = n1494 & ~n11310 ;
  assign n11312 = n11311 ^ n4401 ^ n952 ;
  assign n11313 = ( n352 & ~n5117 ) | ( n352 & n5616 ) | ( ~n5117 & n5616 ) ;
  assign n11314 = ( ~n6407 & n11312 ) | ( ~n6407 & n11313 ) | ( n11312 & n11313 ) ;
  assign n11315 = n11314 ^ n2948 ^ n156 ;
  assign n11316 = n6754 ^ n4107 ^ n282 ;
  assign n11317 = ( ~n5759 & n6077 ) | ( ~n5759 & n11316 ) | ( n6077 & n11316 ) ;
  assign n11318 = ( ~n902 & n1181 ) | ( ~n902 & n11317 ) | ( n1181 & n11317 ) ;
  assign n11319 = n7601 ^ n3082 ^ n2801 ;
  assign n11320 = n11319 ^ n7407 ^ x117 ;
  assign n11321 = n5858 ^ n2445 ^ n1448 ;
  assign n11322 = ( n5826 & n9496 ) | ( n5826 & n11321 ) | ( n9496 & n11321 ) ;
  assign n11323 = ( ~n11318 & n11320 ) | ( ~n11318 & n11322 ) | ( n11320 & n11322 ) ;
  assign n11324 = ( n7542 & ~n8791 ) | ( n7542 & n11323 ) | ( ~n8791 & n11323 ) ;
  assign n11326 = ( n791 & n2807 ) | ( n791 & n5136 ) | ( n2807 & n5136 ) ;
  assign n11327 = n3126 & ~n11326 ;
  assign n11328 = n11327 ^ n848 ^ 1'b0 ;
  assign n11329 = n11328 ^ n6431 ^ n1522 ;
  assign n11325 = n9100 ^ n7895 ^ n3609 ;
  assign n11330 = n11329 ^ n11325 ^ n3641 ;
  assign n11331 = n10931 | n11330 ;
  assign n11332 = n1880 | n11331 ;
  assign n11333 = ( n2775 & n5176 ) | ( n2775 & ~n9637 ) | ( n5176 & ~n9637 ) ;
  assign n11334 = n6297 ^ n3601 ^ 1'b0 ;
  assign n11335 = n11334 ^ n10985 ^ n10803 ;
  assign n11336 = n2103 & n11093 ;
  assign n11337 = n3899 & n11336 ;
  assign n11338 = n11337 ^ n8490 ^ n2213 ;
  assign n11339 = n1651 ^ n799 ^ 1'b0 ;
  assign n11340 = n11338 & ~n11339 ;
  assign n11341 = ~n1410 & n11340 ;
  assign n11342 = ( n170 & n1286 ) | ( n170 & ~n11341 ) | ( n1286 & ~n11341 ) ;
  assign n11343 = ~n277 & n11342 ;
  assign n11344 = n11343 ^ n3131 ^ 1'b0 ;
  assign n11345 = n3156 ^ n1522 ^ 1'b0 ;
  assign n11346 = n10405 ^ n6773 ^ n2728 ;
  assign n11347 = ( n4319 & ~n11345 ) | ( n4319 & n11346 ) | ( ~n11345 & n11346 ) ;
  assign n11351 = ( n1372 & n3178 ) | ( n1372 & ~n8028 ) | ( n3178 & ~n8028 ) ;
  assign n11348 = n6128 ^ n5021 ^ n2980 ;
  assign n11349 = n11348 ^ n5887 ^ n4083 ;
  assign n11350 = n11349 ^ n5661 ^ n3251 ;
  assign n11352 = n11351 ^ n11350 ^ n5760 ;
  assign n11353 = n9855 ^ n2646 ^ 1'b0 ;
  assign n11354 = ~n11352 & n11353 ;
  assign n11355 = n3464 ^ n1005 ^ n998 ;
  assign n11356 = n11355 ^ n11318 ^ 1'b0 ;
  assign n11357 = n11354 & ~n11356 ;
  assign n11358 = ( n2149 & n5232 ) | ( n2149 & n11357 ) | ( n5232 & n11357 ) ;
  assign n11359 = n406 ^ n265 ^ 1'b0 ;
  assign n11361 = x117 & ~n1261 ;
  assign n11362 = n990 & n11361 ;
  assign n11363 = n11362 ^ n9917 ^ n810 ;
  assign n11360 = n2154 & n5100 ;
  assign n11364 = n11363 ^ n11360 ^ 1'b0 ;
  assign n11365 = n8996 ^ n6672 ^ 1'b0 ;
  assign n11366 = ( n11359 & n11364 ) | ( n11359 & ~n11365 ) | ( n11364 & ~n11365 ) ;
  assign n11367 = ( ~n8728 & n10398 ) | ( ~n8728 & n11366 ) | ( n10398 & n11366 ) ;
  assign n11368 = ~n466 & n4093 ;
  assign n11369 = ~n6063 & n11368 ;
  assign n11370 = n4600 ^ n680 ^ 1'b0 ;
  assign n11371 = n11369 & ~n11370 ;
  assign n11376 = n8315 ^ n6077 ^ n1363 ;
  assign n11377 = ~n4886 & n11376 ;
  assign n11378 = n9100 & n11377 ;
  assign n11372 = n6039 ^ n3339 ^ 1'b0 ;
  assign n11373 = n4111 & n11372 ;
  assign n11374 = n10732 & n11373 ;
  assign n11375 = n7710 & n11374 ;
  assign n11379 = n11378 ^ n11375 ^ n6743 ;
  assign n11383 = ( n593 & ~n2611 ) | ( n593 & n9241 ) | ( ~n2611 & n9241 ) ;
  assign n11381 = n1342 ^ n1305 ^ 1'b0 ;
  assign n11380 = ( n1000 & n2904 ) | ( n1000 & ~n5353 ) | ( n2904 & ~n5353 ) ;
  assign n11382 = n11381 ^ n11380 ^ n1258 ;
  assign n11384 = n11383 ^ n11382 ^ n7800 ;
  assign n11385 = n8295 ^ n4259 ^ 1'b0 ;
  assign n11386 = n3792 & ~n11385 ;
  assign n11391 = n4765 ^ n1595 ^ 1'b0 ;
  assign n11392 = x83 & ~n11391 ;
  assign n11387 = ( n3656 & n6322 ) | ( n3656 & ~n9120 ) | ( n6322 & ~n9120 ) ;
  assign n11388 = ~n5630 & n11387 ;
  assign n11389 = n11388 ^ n4907 ^ 1'b0 ;
  assign n11390 = n7940 & ~n11389 ;
  assign n11393 = n11392 ^ n11390 ^ 1'b0 ;
  assign n11394 = n3391 ^ x4 ^ 1'b0 ;
  assign n11395 = n11394 ^ n1603 ^ n394 ;
  assign n11396 = n11395 ^ n3491 ^ n2260 ;
  assign n11397 = n2302 ^ n2185 ^ 1'b0 ;
  assign n11398 = ( n197 & n1939 ) | ( n197 & ~n11397 ) | ( n1939 & ~n11397 ) ;
  assign n11399 = n11398 ^ n7111 ^ n3948 ;
  assign n11400 = n7582 & n7744 ;
  assign n11401 = n9995 ^ n8275 ^ 1'b0 ;
  assign n11402 = ( n7068 & n8041 ) | ( n7068 & ~n8080 ) | ( n8041 & ~n8080 ) ;
  assign n11403 = n4531 & ~n5124 ;
  assign n11404 = n5671 ^ n1095 ^ 1'b0 ;
  assign n11405 = n11404 ^ n5264 ^ n753 ;
  assign n11406 = n3716 ^ n1490 ^ 1'b0 ;
  assign n11407 = n5285 & ~n11406 ;
  assign n11408 = n11405 & n11407 ;
  assign n11409 = ( ~n1120 & n2825 ) | ( ~n1120 & n6520 ) | ( n2825 & n6520 ) ;
  assign n11410 = n5328 ^ n1293 ^ 1'b0 ;
  assign n11411 = ~n11409 & n11410 ;
  assign n11412 = n2551 | n11411 ;
  assign n11413 = ( n1376 & ~n8615 ) | ( n1376 & n8696 ) | ( ~n8615 & n8696 ) ;
  assign n11414 = n11413 ^ n11398 ^ n475 ;
  assign n11415 = n11414 ^ n6973 ^ 1'b0 ;
  assign n11416 = n2689 & ~n11415 ;
  assign n11417 = n607 & n2467 ;
  assign n11418 = n8327 ^ n857 ^ 1'b0 ;
  assign n11419 = ~n7211 & n11418 ;
  assign n11420 = n11419 ^ n3396 ^ 1'b0 ;
  assign n11421 = ( n1258 & n7984 ) | ( n1258 & ~n11420 ) | ( n7984 & ~n11420 ) ;
  assign n11422 = ( ~n3102 & n3946 ) | ( ~n3102 & n4027 ) | ( n3946 & n4027 ) ;
  assign n11423 = n4189 & n11422 ;
  assign n11424 = ~n1765 & n4453 ;
  assign n11425 = n7483 & n11424 ;
  assign n11426 = ( ~x54 & n1117 ) | ( ~x54 & n4107 ) | ( n1117 & n4107 ) ;
  assign n11427 = ( ~n2727 & n3905 ) | ( ~n2727 & n11426 ) | ( n3905 & n11426 ) ;
  assign n11429 = n8692 ^ n4900 ^ 1'b0 ;
  assign n11430 = n724 & ~n11429 ;
  assign n11428 = n5406 & ~n10684 ;
  assign n11431 = n11430 ^ n11428 ^ 1'b0 ;
  assign n11432 = n3215 & n8763 ;
  assign n11433 = ( n11427 & n11431 ) | ( n11427 & ~n11432 ) | ( n11431 & ~n11432 ) ;
  assign n11434 = n11433 ^ n9593 ^ 1'b0 ;
  assign n11435 = ( ~n669 & n8257 ) | ( ~n669 & n11225 ) | ( n8257 & n11225 ) ;
  assign n11436 = n11435 ^ n4494 ^ n2097 ;
  assign n11437 = n2609 | n8082 ;
  assign n11438 = n11437 ^ n4396 ^ 1'b0 ;
  assign n11439 = n11438 ^ n5655 ^ n697 ;
  assign n11440 = n1304 & ~n10280 ;
  assign n11441 = ~n1167 & n11440 ;
  assign n11442 = n11441 ^ n643 ^ 1'b0 ;
  assign n11443 = n11442 ^ n10950 ^ n10643 ;
  assign n11444 = ~n1563 & n2624 ;
  assign n11445 = ( n2396 & n11055 ) | ( n2396 & ~n11444 ) | ( n11055 & ~n11444 ) ;
  assign n11446 = ( n908 & ~n5079 ) | ( n908 & n11445 ) | ( ~n5079 & n11445 ) ;
  assign n11450 = n3381 ^ n1729 ^ n1513 ;
  assign n11447 = n4588 ^ n2014 ^ n1708 ;
  assign n11448 = ( n5032 & n8197 ) | ( n5032 & n11447 ) | ( n8197 & n11447 ) ;
  assign n11449 = n7180 | n11448 ;
  assign n11451 = n11450 ^ n11449 ^ 1'b0 ;
  assign n11452 = n7337 ^ n3368 ^ 1'b0 ;
  assign n11453 = n822 & ~n11452 ;
  assign n11454 = n11453 ^ n6873 ^ n2957 ;
  assign n11455 = n11454 ^ n8322 ^ n3768 ;
  assign n11456 = n180 & ~n1765 ;
  assign n11457 = x25 & ~n5601 ;
  assign n11458 = n11457 ^ n2058 ^ 1'b0 ;
  assign n11459 = n10974 & n11458 ;
  assign n11460 = n7900 & n11459 ;
  assign n11461 = n1121 & ~n11460 ;
  assign n11462 = n335 | n1093 ;
  assign n11463 = n11462 ^ n7661 ^ 1'b0 ;
  assign n11464 = ~n1234 & n6454 ;
  assign n11465 = n11464 ^ n1727 ^ 1'b0 ;
  assign n11466 = ( n2576 & n11463 ) | ( n2576 & n11465 ) | ( n11463 & n11465 ) ;
  assign n11467 = n4806 ^ n4495 ^ n2724 ;
  assign n11468 = ( n466 & n1506 ) | ( n466 & ~n2253 ) | ( n1506 & ~n2253 ) ;
  assign n11469 = n11468 ^ n9367 ^ n5125 ;
  assign n11470 = n11469 ^ n9620 ^ n2976 ;
  assign n11471 = ( ~n11055 & n11467 ) | ( ~n11055 & n11470 ) | ( n11467 & n11470 ) ;
  assign n11472 = ( ~n2026 & n2838 ) | ( ~n2026 & n4553 ) | ( n2838 & n4553 ) ;
  assign n11473 = ( n3613 & ~n3642 ) | ( n3613 & n11472 ) | ( ~n3642 & n11472 ) ;
  assign n11474 = n6572 ^ n1308 ^ 1'b0 ;
  assign n11475 = ( n6722 & ~n11473 ) | ( n6722 & n11474 ) | ( ~n11473 & n11474 ) ;
  assign n11476 = n2200 & ~n8729 ;
  assign n11477 = n11476 ^ n1396 ^ 1'b0 ;
  assign n11478 = n10024 & ~n11477 ;
  assign n11479 = ( n367 & ~n3440 ) | ( n367 & n11478 ) | ( ~n3440 & n11478 ) ;
  assign n11480 = n7771 ^ n6813 ^ n4735 ;
  assign n11481 = n4760 & n11164 ;
  assign n11482 = ~n11480 & n11481 ;
  assign n11489 = n5552 ^ n5215 ^ n1104 ;
  assign n11490 = n2269 | n11489 ;
  assign n11486 = ( n613 & ~n2654 ) | ( n613 & n7990 ) | ( ~n2654 & n7990 ) ;
  assign n11487 = n11486 ^ n6389 ^ n4879 ;
  assign n11483 = n1254 & ~n2007 ;
  assign n11484 = n11483 ^ n8127 ^ 1'b0 ;
  assign n11485 = ~n2916 & n11484 ;
  assign n11488 = n11487 ^ n11485 ^ 1'b0 ;
  assign n11491 = n11490 ^ n11488 ^ n3606 ;
  assign n11492 = n5184 ^ n4431 ^ n2141 ;
  assign n11493 = ( n4706 & n8692 ) | ( n4706 & n11492 ) | ( n8692 & n11492 ) ;
  assign n11495 = n8433 ^ n4352 ^ 1'b0 ;
  assign n11496 = n9420 & ~n11495 ;
  assign n11494 = n8618 ^ n3167 ^ n1587 ;
  assign n11497 = n11496 ^ n11494 ^ n10605 ;
  assign n11499 = n3058 ^ n1554 ^ 1'b0 ;
  assign n11498 = ( n3942 & n4486 ) | ( n3942 & ~n11318 ) | ( n4486 & ~n11318 ) ;
  assign n11500 = n11499 ^ n11498 ^ n11179 ;
  assign n11501 = n11500 ^ n4191 ^ n2036 ;
  assign n11502 = ( n288 & ~n5748 ) | ( n288 & n11501 ) | ( ~n5748 & n11501 ) ;
  assign n11503 = n5428 ^ n3589 ^ n2765 ;
  assign n11504 = n11503 ^ n1168 ^ 1'b0 ;
  assign n11505 = n8532 ^ n1407 ^ 1'b0 ;
  assign n11506 = n2554 & ~n11505 ;
  assign n11507 = ~n11504 & n11506 ;
  assign n11508 = n3191 & n11507 ;
  assign n11509 = n10296 ^ n3026 ^ 1'b0 ;
  assign n11510 = ( n6028 & ~n11508 ) | ( n6028 & n11509 ) | ( ~n11508 & n11509 ) ;
  assign n11512 = ( ~n845 & n3282 ) | ( ~n845 & n9947 ) | ( n3282 & n9947 ) ;
  assign n11511 = ( n252 & n814 ) | ( n252 & ~n6273 ) | ( n814 & ~n6273 ) ;
  assign n11513 = n11512 ^ n11511 ^ n319 ;
  assign n11514 = n801 | n883 ;
  assign n11515 = n4141 | n11514 ;
  assign n11516 = n10106 | n11515 ;
  assign n11517 = ~n8514 & n11516 ;
  assign n11518 = ( n252 & ~n4303 ) | ( n252 & n6580 ) | ( ~n4303 & n6580 ) ;
  assign n11519 = n839 | n11518 ;
  assign n11520 = n11517 | n11519 ;
  assign n11521 = n4592 & n10448 ;
  assign n11522 = n11521 ^ n9829 ^ n6874 ;
  assign n11523 = n1793 ^ n553 ^ 1'b0 ;
  assign n11524 = n9149 ^ n6603 ^ 1'b0 ;
  assign n11525 = n758 & ~n11524 ;
  assign n11526 = n11525 ^ n9147 ^ 1'b0 ;
  assign n11527 = n4965 & n11526 ;
  assign n11528 = n1359 ^ n653 ^ x112 ;
  assign n11529 = n11528 ^ n3870 ^ n2534 ;
  assign n11530 = n7003 ^ n6247 ^ n6024 ;
  assign n11531 = n11530 ^ n7081 ^ n2251 ;
  assign n11532 = ( n11527 & n11529 ) | ( n11527 & ~n11531 ) | ( n11529 & ~n11531 ) ;
  assign n11533 = n425 & n4392 ;
  assign n11534 = n11533 ^ n1029 ^ 1'b0 ;
  assign n11535 = n8931 ^ n3595 ^ n966 ;
  assign n11536 = ( n3147 & n11413 ) | ( n3147 & ~n11535 ) | ( n11413 & ~n11535 ) ;
  assign n11537 = ( n567 & n9190 ) | ( n567 & n11536 ) | ( n9190 & n11536 ) ;
  assign n11538 = n7264 | n8953 ;
  assign n11539 = ( n889 & n11537 ) | ( n889 & n11538 ) | ( n11537 & n11538 ) ;
  assign n11544 = ( n3135 & n3314 ) | ( n3135 & n7254 ) | ( n3314 & n7254 ) ;
  assign n11545 = n11544 ^ n8883 ^ n4821 ;
  assign n11546 = ( ~n3621 & n9598 ) | ( ~n3621 & n11545 ) | ( n9598 & n11545 ) ;
  assign n11540 = n7596 ^ n6184 ^ n4712 ;
  assign n11541 = ( n1283 & n5131 ) | ( n1283 & ~n11540 ) | ( n5131 & ~n11540 ) ;
  assign n11542 = n1893 & n11541 ;
  assign n11543 = ~n8929 & n11542 ;
  assign n11547 = n11546 ^ n11543 ^ n4181 ;
  assign n11548 = n9591 ^ n8839 ^ n5291 ;
  assign n11549 = n11548 ^ n9742 ^ n6039 ;
  assign n11550 = n10557 ^ n7134 ^ x10 ;
  assign n11551 = ~n495 & n11550 ;
  assign n11552 = n11551 ^ n10232 ^ 1'b0 ;
  assign n11553 = n6656 & ~n10191 ;
  assign n11554 = ( ~n4943 & n6667 ) | ( ~n4943 & n11553 ) | ( n6667 & n11553 ) ;
  assign n11555 = ( ~n2458 & n3888 ) | ( ~n2458 & n3928 ) | ( n3888 & n3928 ) ;
  assign n11556 = n11555 ^ n910 ^ n371 ;
  assign n11557 = n608 | n5778 ;
  assign n11558 = n11557 ^ n6474 ^ 1'b0 ;
  assign n11559 = ( ~n4034 & n9722 ) | ( ~n4034 & n11558 ) | ( n9722 & n11558 ) ;
  assign n11560 = n1274 & n9409 ;
  assign n11561 = n1931 & n11560 ;
  assign n11562 = ( n3469 & n4786 ) | ( n3469 & n11561 ) | ( n4786 & n11561 ) ;
  assign n11563 = ( ~x37 & n1925 ) | ( ~x37 & n3296 ) | ( n1925 & n3296 ) ;
  assign n11564 = n11563 ^ n7210 ^ x111 ;
  assign n11565 = n5722 | n11564 ;
  assign n11566 = n11565 ^ n5269 ^ 1'b0 ;
  assign n11567 = n8828 ^ n7021 ^ n3513 ;
  assign n11568 = n2616 ^ n953 ^ x16 ;
  assign n11569 = n11568 ^ n1637 ^ n389 ;
  assign n11570 = n11569 ^ n9534 ^ 1'b0 ;
  assign n11571 = n1845 | n11570 ;
  assign n11572 = ( n11207 & n11567 ) | ( n11207 & ~n11571 ) | ( n11567 & ~n11571 ) ;
  assign n11573 = n9059 ^ n6473 ^ 1'b0 ;
  assign n11574 = n8057 ^ n6883 ^ 1'b0 ;
  assign n11575 = ( n2060 & n3881 ) | ( n2060 & ~n4020 ) | ( n3881 & ~n4020 ) ;
  assign n11576 = n7996 & ~n11575 ;
  assign n11577 = n11576 ^ n4983 ^ 1'b0 ;
  assign n11578 = ( n8794 & n11574 ) | ( n8794 & n11577 ) | ( n11574 & n11577 ) ;
  assign n11579 = ~n3861 & n10718 ;
  assign n11580 = n11579 ^ n11025 ^ n2280 ;
  assign n11581 = n3330 ^ n1357 ^ 1'b0 ;
  assign n11582 = ~n11580 & n11581 ;
  assign n11583 = n8854 ^ n5205 ^ n2029 ;
  assign n11584 = ~n3851 & n5802 ;
  assign n11585 = n11584 ^ n9779 ^ n2980 ;
  assign n11586 = n11585 ^ n5954 ^ n5813 ;
  assign n11587 = ( n3679 & n11583 ) | ( n3679 & n11586 ) | ( n11583 & n11586 ) ;
  assign n11588 = ( n3565 & ~n4275 ) | ( n3565 & n4900 ) | ( ~n4275 & n4900 ) ;
  assign n11589 = n10639 ^ n4021 ^ n1399 ;
  assign n11590 = n11589 ^ n3561 ^ 1'b0 ;
  assign n11591 = n11588 | n11590 ;
  assign n11592 = n6990 ^ n3565 ^ n3515 ;
  assign n11593 = n3222 ^ n1983 ^ n529 ;
  assign n11594 = ( n1758 & n11592 ) | ( n1758 & n11593 ) | ( n11592 & n11593 ) ;
  assign n11595 = ( n10176 & n11591 ) | ( n10176 & ~n11594 ) | ( n11591 & ~n11594 ) ;
  assign n11596 = ( n429 & n726 ) | ( n429 & ~n758 ) | ( n726 & ~n758 ) ;
  assign n11597 = ( n1274 & n2221 ) | ( n1274 & ~n11596 ) | ( n2221 & ~n11596 ) ;
  assign n11598 = ( n901 & n1451 ) | ( n901 & ~n11597 ) | ( n1451 & ~n11597 ) ;
  assign n11599 = n3731 | n3860 ;
  assign n11600 = n11599 ^ n1592 ^ 1'b0 ;
  assign n11601 = n11600 ^ n7392 ^ 1'b0 ;
  assign n11602 = ~n11598 & n11601 ;
  assign n11603 = ( n6782 & ~n8442 ) | ( n6782 & n11602 ) | ( ~n8442 & n11602 ) ;
  assign n11604 = n3249 & n11413 ;
  assign n11605 = n11604 ^ n10240 ^ 1'b0 ;
  assign n11606 = ( n7275 & n9987 ) | ( n7275 & ~n11605 ) | ( n9987 & ~n11605 ) ;
  assign n11607 = ( n7148 & n7467 ) | ( n7148 & n8319 ) | ( n7467 & n8319 ) ;
  assign n11608 = n3070 & n11607 ;
  assign n11609 = n11608 ^ n5504 ^ 1'b0 ;
  assign n11610 = n1541 & ~n11609 ;
  assign n11611 = ( x112 & n604 ) | ( x112 & n4049 ) | ( n604 & n4049 ) ;
  assign n11612 = ~n5472 & n11611 ;
  assign n11613 = ~n940 & n11612 ;
  assign n11614 = n11613 ^ n6290 ^ n2615 ;
  assign n11615 = n7405 ^ n3754 ^ n565 ;
  assign n11616 = n6514 ^ n2957 ^ n2535 ;
  assign n11617 = n131 & ~n3384 ;
  assign n11618 = n6611 & n11617 ;
  assign n11619 = n11616 | n11618 ;
  assign n11620 = ( n1847 & n5402 ) | ( n1847 & n5808 ) | ( n5402 & n5808 ) ;
  assign n11621 = n11620 ^ n5436 ^ 1'b0 ;
  assign n11622 = n5916 & n11621 ;
  assign n11623 = n5312 ^ n3279 ^ 1'b0 ;
  assign n11624 = ( n2142 & n8388 ) | ( n2142 & n11623 ) | ( n8388 & n11623 ) ;
  assign n11626 = n8641 ^ n7441 ^ 1'b0 ;
  assign n11627 = n7416 | n11626 ;
  assign n11625 = n3983 & ~n8990 ;
  assign n11628 = n11627 ^ n11625 ^ n8018 ;
  assign n11629 = n7673 ^ n5882 ^ n3144 ;
  assign n11636 = n3538 ^ n845 ^ 1'b0 ;
  assign n11637 = ~n8829 & n11636 ;
  assign n11630 = n2174 ^ n826 ^ 1'b0 ;
  assign n11631 = n1282 | n11630 ;
  assign n11632 = n11631 ^ n5539 ^ n1686 ;
  assign n11633 = n11632 ^ n900 ^ n387 ;
  assign n11634 = n2980 & ~n11633 ;
  assign n11635 = n7895 & n11634 ;
  assign n11638 = n11637 ^ n11635 ^ n11320 ;
  assign n11639 = ~n11629 & n11638 ;
  assign n11640 = n11639 ^ n8569 ^ 1'b0 ;
  assign n11641 = ( n1993 & n6508 ) | ( n1993 & ~n6964 ) | ( n6508 & ~n6964 ) ;
  assign n11642 = n3919 ^ n3387 ^ n3155 ;
  assign n11643 = n11641 & n11642 ;
  assign n11644 = ~n184 & n415 ;
  assign n11645 = n5052 ^ n2138 ^ n1701 ;
  assign n11646 = ( n449 & n3695 ) | ( n449 & n11645 ) | ( n3695 & n11645 ) ;
  assign n11647 = ( n6809 & ~n7060 ) | ( n6809 & n11646 ) | ( ~n7060 & n11646 ) ;
  assign n11648 = n11647 ^ n3807 ^ 1'b0 ;
  assign n11650 = n453 & n1677 ;
  assign n11651 = ~n5945 & n11650 ;
  assign n11649 = n1371 & n1889 ;
  assign n11652 = n11651 ^ n11649 ^ 1'b0 ;
  assign n11653 = n2813 ^ x119 ^ 1'b0 ;
  assign n11654 = ( ~n1764 & n4159 ) | ( ~n1764 & n11653 ) | ( n4159 & n11653 ) ;
  assign n11657 = n3460 ^ n2671 ^ n1500 ;
  assign n11658 = n11657 ^ n4109 ^ n3356 ;
  assign n11655 = n9580 ^ n7448 ^ n6377 ;
  assign n11656 = ( n1481 & n6886 ) | ( n1481 & ~n11655 ) | ( n6886 & ~n11655 ) ;
  assign n11659 = n11658 ^ n11656 ^ 1'b0 ;
  assign n11660 = n11654 & ~n11659 ;
  assign n11661 = n11660 ^ n3965 ^ n2252 ;
  assign n11662 = n9100 ^ n8676 ^ n4284 ;
  assign n11663 = ( n1373 & n2130 ) | ( n1373 & ~n11662 ) | ( n2130 & ~n11662 ) ;
  assign n11664 = ( n748 & n840 ) | ( n748 & ~n3883 ) | ( n840 & ~n3883 ) ;
  assign n11665 = n6607 | n11664 ;
  assign n11666 = n11665 ^ n9338 ^ 1'b0 ;
  assign n11667 = ( ~n971 & n3069 ) | ( ~n971 & n8867 ) | ( n3069 & n8867 ) ;
  assign n11668 = n11667 ^ n6700 ^ n549 ;
  assign n11669 = ( ~n1493 & n1581 ) | ( ~n1493 & n10402 ) | ( n1581 & n10402 ) ;
  assign n11670 = ~n5459 & n11669 ;
  assign n11671 = n8866 ^ n6111 ^ 1'b0 ;
  assign n11672 = ( n6055 & n7814 ) | ( n6055 & ~n11671 ) | ( n7814 & ~n11671 ) ;
  assign n11673 = n6982 ^ n6330 ^ n6202 ;
  assign n11677 = n4739 | n6350 ;
  assign n11674 = n3747 ^ n689 ^ 1'b0 ;
  assign n11675 = n7686 | n11674 ;
  assign n11676 = n3264 | n11675 ;
  assign n11678 = n11677 ^ n11676 ^ 1'b0 ;
  assign n11679 = n8615 ^ n3304 ^ 1'b0 ;
  assign n11680 = n6795 ^ n1172 ^ 1'b0 ;
  assign n11681 = n11679 & ~n11680 ;
  assign n11682 = ( n3892 & n6776 ) | ( n3892 & n11681 ) | ( n6776 & n11681 ) ;
  assign n11683 = n7811 ^ n6700 ^ n1712 ;
  assign n11684 = n11683 ^ n9802 ^ n365 ;
  assign n11685 = n7502 & n11609 ;
  assign n11686 = n11685 ^ n3884 ^ 1'b0 ;
  assign n11687 = n10225 ^ n3684 ^ n889 ;
  assign n11688 = n2117 ^ n478 ^ 1'b0 ;
  assign n11689 = ~n11687 & n11688 ;
  assign n11690 = ~n9207 & n11689 ;
  assign n11691 = n10463 ^ n2136 ^ 1'b0 ;
  assign n11692 = ( ~n1082 & n7359 ) | ( ~n1082 & n11691 ) | ( n7359 & n11691 ) ;
  assign n11701 = n1848 & n5279 ;
  assign n11702 = n5073 & ~n11701 ;
  assign n11693 = n9555 ^ n5093 ^ n4485 ;
  assign n11694 = ~n1194 & n5801 ;
  assign n11695 = n11694 ^ n6816 ^ 1'b0 ;
  assign n11697 = ( n1210 & ~n3050 ) | ( n1210 & n3268 ) | ( ~n3050 & n3268 ) ;
  assign n11696 = n3515 & ~n7752 ;
  assign n11698 = n11697 ^ n11696 ^ 1'b0 ;
  assign n11699 = ( n5871 & ~n11695 ) | ( n5871 & n11698 ) | ( ~n11695 & n11698 ) ;
  assign n11700 = ( n10176 & ~n11693 ) | ( n10176 & n11699 ) | ( ~n11693 & n11699 ) ;
  assign n11703 = n11702 ^ n11700 ^ x89 ;
  assign n11704 = n6661 & ~n10919 ;
  assign n11705 = ~n2276 & n11704 ;
  assign n11706 = n1954 | n2551 ;
  assign n11707 = n11706 ^ n8307 ^ n2450 ;
  assign n11708 = ( n7079 & n11705 ) | ( n7079 & ~n11707 ) | ( n11705 & ~n11707 ) ;
  assign n11709 = n11708 ^ n3396 ^ n2868 ;
  assign n11710 = n2517 & n3470 ;
  assign n11711 = n5232 ^ n1309 ^ 1'b0 ;
  assign n11712 = n5546 & ~n11711 ;
  assign n11717 = n5285 ^ n2327 ^ 1'b0 ;
  assign n11718 = n1692 | n11717 ;
  assign n11716 = x74 & ~n9869 ;
  assign n11713 = n1179 & n10860 ;
  assign n11714 = n11713 ^ n10429 ^ n966 ;
  assign n11715 = ( n770 & ~n5609 ) | ( n770 & n11714 ) | ( ~n5609 & n11714 ) ;
  assign n11719 = n11718 ^ n11716 ^ n11715 ;
  assign n11720 = ( n648 & ~n1225 ) | ( n648 & n6635 ) | ( ~n1225 & n6635 ) ;
  assign n11721 = n11720 ^ n2859 ^ 1'b0 ;
  assign n11722 = ( n4076 & n6917 ) | ( n4076 & n11721 ) | ( n6917 & n11721 ) ;
  assign n11723 = n11722 ^ n11516 ^ 1'b0 ;
  assign n11724 = ( n1340 & n5871 ) | ( n1340 & ~n11723 ) | ( n5871 & ~n11723 ) ;
  assign n11725 = ( n3526 & n4415 ) | ( n3526 & ~n6257 ) | ( n4415 & ~n6257 ) ;
  assign n11726 = n11725 ^ n8005 ^ n6433 ;
  assign n11727 = n3783 ^ n2457 ^ n315 ;
  assign n11728 = n296 & n7155 ;
  assign n11729 = ~n11727 & n11728 ;
  assign n11730 = ( ~n1208 & n6975 ) | ( ~n1208 & n11729 ) | ( n6975 & n11729 ) ;
  assign n11731 = n9504 ^ n8939 ^ n6553 ;
  assign n11732 = ( n10389 & n11345 ) | ( n10389 & ~n11731 ) | ( n11345 & ~n11731 ) ;
  assign n11734 = n9809 ^ n8344 ^ n775 ;
  assign n11735 = ( n322 & ~n8723 ) | ( n322 & n11734 ) | ( ~n8723 & n11734 ) ;
  assign n11733 = n4310 & ~n9669 ;
  assign n11736 = n11735 ^ n11733 ^ 1'b0 ;
  assign n11737 = n386 | n4577 ;
  assign n11738 = ( n1020 & ~n8139 ) | ( n1020 & n8996 ) | ( ~n8139 & n8996 ) ;
  assign n11739 = n11738 ^ n5535 ^ n1466 ;
  assign n11740 = n11739 ^ n7882 ^ n2702 ;
  assign n11741 = ( n1345 & n4404 ) | ( n1345 & ~n5698 ) | ( n4404 & ~n5698 ) ;
  assign n11742 = n7954 & ~n11741 ;
  assign n11743 = ( ~n1542 & n1716 ) | ( ~n1542 & n11742 ) | ( n1716 & n11742 ) ;
  assign n11744 = ( n2894 & n8426 ) | ( n2894 & n11743 ) | ( n8426 & n11743 ) ;
  assign n11745 = ( n669 & n780 ) | ( n669 & n5955 ) | ( n780 & n5955 ) ;
  assign n11746 = n9508 & ~n11745 ;
  assign n11747 = n11746 ^ n10687 ^ 1'b0 ;
  assign n11748 = n11747 ^ n8569 ^ n809 ;
  assign n11749 = ( ~n5848 & n8156 ) | ( ~n5848 & n10754 ) | ( n8156 & n10754 ) ;
  assign n11750 = ~n9729 & n11749 ;
  assign n11753 = n10331 ^ n464 ^ 1'b0 ;
  assign n11754 = x26 & ~n11753 ;
  assign n11751 = ( ~n1619 & n4396 ) | ( ~n1619 & n6816 ) | ( n4396 & n6816 ) ;
  assign n11752 = n1109 | n11751 ;
  assign n11755 = n11754 ^ n11752 ^ 1'b0 ;
  assign n11756 = n1431 ^ n721 ^ n502 ;
  assign n11757 = ( n225 & n308 ) | ( n225 & ~n11756 ) | ( n308 & ~n11756 ) ;
  assign n11758 = n11757 ^ n1652 ^ n237 ;
  assign n11759 = n11758 ^ n11059 ^ n7147 ;
  assign n11760 = n6024 ^ n4138 ^ n1935 ;
  assign n11761 = ( n1437 & ~n2016 ) | ( n1437 & n11760 ) | ( ~n2016 & n11760 ) ;
  assign n11762 = n7474 ^ n4855 ^ 1'b0 ;
  assign n11763 = n6057 ^ n2654 ^ n1620 ;
  assign n11764 = ( n2581 & n5601 ) | ( n2581 & ~n11763 ) | ( n5601 & ~n11763 ) ;
  assign n11765 = n11764 ^ n10399 ^ 1'b0 ;
  assign n11766 = n11762 | n11765 ;
  assign n11767 = n8154 ^ n992 ^ 1'b0 ;
  assign n11768 = n1050 | n11767 ;
  assign n11777 = n5987 ^ n3167 ^ 1'b0 ;
  assign n11775 = n7842 ^ n3790 ^ 1'b0 ;
  assign n11776 = n11775 ^ n11381 ^ n1738 ;
  assign n11771 = n5061 ^ n2470 ^ 1'b0 ;
  assign n11772 = n1779 & n11771 ;
  assign n11769 = n6979 ^ n3241 ^ n1912 ;
  assign n11770 = ( n771 & n9301 ) | ( n771 & n11769 ) | ( n9301 & n11769 ) ;
  assign n11773 = n11772 ^ n11770 ^ n11671 ;
  assign n11774 = ( n2608 & n8895 ) | ( n2608 & n11773 ) | ( n8895 & n11773 ) ;
  assign n11778 = n11777 ^ n11776 ^ n11774 ;
  assign n11779 = n6357 ^ n900 ^ x77 ;
  assign n11780 = n2560 ^ n1110 ^ n713 ;
  assign n11781 = ( n1655 & ~n3646 ) | ( n1655 & n11780 ) | ( ~n3646 & n11780 ) ;
  assign n11782 = ~n2923 & n11781 ;
  assign n11783 = ~n3789 & n11782 ;
  assign n11784 = ( n6213 & n11779 ) | ( n6213 & n11783 ) | ( n11779 & n11783 ) ;
  assign n11785 = n4639 ^ n3893 ^ n1945 ;
  assign n11786 = ( n2873 & ~n9959 ) | ( n2873 & n11785 ) | ( ~n9959 & n11785 ) ;
  assign n11787 = n10577 & n11786 ;
  assign n11789 = n3598 ^ n2188 ^ n463 ;
  assign n11788 = ( n1474 & n4970 ) | ( n1474 & ~n5296 ) | ( n4970 & ~n5296 ) ;
  assign n11790 = n11789 ^ n11788 ^ n5292 ;
  assign n11791 = n2730 & n3973 ;
  assign n11792 = n5515 & n11791 ;
  assign n11793 = ~n7520 & n11792 ;
  assign n11794 = n1207 & n1276 ;
  assign n11795 = ( n4833 & n5037 ) | ( n4833 & n11794 ) | ( n5037 & n11794 ) ;
  assign n11796 = n11795 ^ n5564 ^ n2865 ;
  assign n11797 = n1570 & ~n7505 ;
  assign n11798 = n7734 ^ n2142 ^ 1'b0 ;
  assign n11799 = ~n11797 & n11798 ;
  assign n11800 = ~n8477 & n11799 ;
  assign n11801 = ~n11796 & n11800 ;
  assign n11802 = n4564 ^ n4080 ^ 1'b0 ;
  assign n11803 = n10037 & n11802 ;
  assign n11804 = n11803 ^ n2319 ^ 1'b0 ;
  assign n11805 = n8599 ^ n5658 ^ n1380 ;
  assign n11806 = n2980 ^ x125 ^ 1'b0 ;
  assign n11807 = n11806 ^ n1541 ^ n904 ;
  assign n11808 = ( n4836 & ~n11805 ) | ( n4836 & n11807 ) | ( ~n11805 & n11807 ) ;
  assign n11809 = n3317 | n10346 ;
  assign n11810 = n11809 ^ n9470 ^ 1'b0 ;
  assign n11811 = n11810 ^ n3101 ^ n2250 ;
  assign n11812 = n11811 ^ n7716 ^ n6786 ;
  assign n11813 = n902 | n1555 ;
  assign n11814 = n11813 ^ n680 ^ 1'b0 ;
  assign n11815 = n2720 & ~n11814 ;
  assign n11816 = n10509 | n11815 ;
  assign n11817 = n1511 | n5960 ;
  assign n11818 = n11817 ^ n5963 ^ 1'b0 ;
  assign n11819 = ~n4689 & n6666 ;
  assign n11820 = n380 | n10039 ;
  assign n11821 = n11819 & ~n11820 ;
  assign n11822 = ( n4228 & n11818 ) | ( n4228 & n11821 ) | ( n11818 & n11821 ) ;
  assign n11824 = ( ~x59 & n511 ) | ( ~x59 & n4135 ) | ( n511 & n4135 ) ;
  assign n11825 = n11824 ^ n11504 ^ n259 ;
  assign n11823 = ~n1179 & n6513 ;
  assign n11826 = n11825 ^ n11823 ^ n9544 ;
  assign n11827 = n3424 ^ x116 ^ 1'b0 ;
  assign n11828 = ~n8111 & n11827 ;
  assign n11829 = ( x76 & n10903 ) | ( x76 & ~n11828 ) | ( n10903 & ~n11828 ) ;
  assign n11830 = ( n7826 & n9173 ) | ( n7826 & ~n11829 ) | ( n9173 & ~n11829 ) ;
  assign n11831 = n2922 | n11830 ;
  assign n11832 = n11831 ^ n6724 ^ 1'b0 ;
  assign n11833 = n11832 ^ n9410 ^ 1'b0 ;
  assign n11834 = n11833 ^ n11620 ^ n9067 ;
  assign n11835 = n8164 & n11834 ;
  assign n11836 = n458 & ~n3714 ;
  assign n11837 = n211 & n11836 ;
  assign n11838 = ( ~n2050 & n2982 ) | ( ~n2050 & n11837 ) | ( n2982 & n11837 ) ;
  assign n11839 = n8380 ^ n5164 ^ 1'b0 ;
  assign n11840 = n11839 ^ n8023 ^ n3799 ;
  assign n11841 = ~n11838 & n11840 ;
  assign n11842 = n11841 ^ n11146 ^ 1'b0 ;
  assign n11843 = n10322 ^ n6856 ^ 1'b0 ;
  assign n11844 = n10820 ^ n2273 ^ n1047 ;
  assign n11845 = n8730 ^ n7724 ^ 1'b0 ;
  assign n11846 = n11844 | n11845 ;
  assign n11847 = n11846 ^ n9032 ^ 1'b0 ;
  assign n11848 = ~n4319 & n4424 ;
  assign n11849 = ~n3034 & n11848 ;
  assign n11850 = n11849 ^ n5777 ^ 1'b0 ;
  assign n11851 = ( n10662 & n11847 ) | ( n10662 & n11850 ) | ( n11847 & n11850 ) ;
  assign n11852 = n2680 ^ n1986 ^ 1'b0 ;
  assign n11853 = ~n1433 & n2295 ;
  assign n11854 = ( n5150 & n11852 ) | ( n5150 & n11853 ) | ( n11852 & n11853 ) ;
  assign n11859 = n2663 ^ n510 ^ 1'b0 ;
  assign n11857 = ~n6754 & n9508 ;
  assign n11858 = ~n2360 & n11857 ;
  assign n11855 = n3623 ^ n3301 ^ 1'b0 ;
  assign n11856 = n11855 ^ n10165 ^ n447 ;
  assign n11860 = n11859 ^ n11858 ^ n11856 ;
  assign n11861 = ( n619 & ~n10403 ) | ( n619 & n11447 ) | ( ~n10403 & n11447 ) ;
  assign n11862 = n7382 ^ n6218 ^ n4273 ;
  assign n11863 = ( n3358 & n11861 ) | ( n3358 & ~n11862 ) | ( n11861 & ~n11862 ) ;
  assign n11864 = n11863 ^ n11009 ^ n8612 ;
  assign n11865 = n6216 | n11864 ;
  assign n11866 = ~n4362 & n5767 ;
  assign n11867 = n11866 ^ x41 ^ 1'b0 ;
  assign n11868 = ~n3750 & n11867 ;
  assign n11869 = n853 & ~n11868 ;
  assign n11873 = n8825 ^ n6852 ^ n6092 ;
  assign n11870 = ~n2459 & n6476 ;
  assign n11871 = ( ~n924 & n7466 ) | ( ~n924 & n11870 ) | ( n7466 & n11870 ) ;
  assign n11872 = ( n4979 & n7547 ) | ( n4979 & n11871 ) | ( n7547 & n11871 ) ;
  assign n11874 = n11873 ^ n11872 ^ 1'b0 ;
  assign n11875 = n6722 ^ n321 ^ 1'b0 ;
  assign n11876 = n2590 & ~n11875 ;
  assign n11877 = n11876 ^ n11575 ^ n10784 ;
  assign n11878 = n1963 | n6192 ;
  assign n11879 = n11878 ^ n9559 ^ n7903 ;
  assign n11885 = ( n149 & ~n1849 ) | ( n149 & n4167 ) | ( ~n1849 & n4167 ) ;
  assign n11880 = ( ~n3960 & n6677 ) | ( ~n3960 & n7734 ) | ( n6677 & n7734 ) ;
  assign n11881 = n11880 ^ n3824 ^ n3139 ;
  assign n11882 = ( n928 & n1633 ) | ( n928 & ~n2497 ) | ( n1633 & ~n2497 ) ;
  assign n11883 = ~n1207 & n11882 ;
  assign n11884 = n11881 & ~n11883 ;
  assign n11886 = n11885 ^ n11884 ^ 1'b0 ;
  assign n11887 = ( n4513 & n9555 ) | ( n4513 & ~n11886 ) | ( n9555 & ~n11886 ) ;
  assign n11888 = n8883 ^ n3620 ^ 1'b0 ;
  assign n11889 = ( n3532 & n7320 ) | ( n3532 & n11888 ) | ( n7320 & n11888 ) ;
  assign n11890 = n10753 & ~n11889 ;
  assign n11891 = ( n5506 & ~n5629 ) | ( n5506 & n7991 ) | ( ~n5629 & n7991 ) ;
  assign n11892 = n1034 & n1166 ;
  assign n11893 = ( n6065 & n7120 ) | ( n6065 & ~n11892 ) | ( n7120 & ~n11892 ) ;
  assign n11898 = x26 & ~n9115 ;
  assign n11899 = n1340 & n11898 ;
  assign n11894 = n2900 | n6182 ;
  assign n11895 = n9386 ^ n6900 ^ n970 ;
  assign n11896 = ( n2187 & n11894 ) | ( n2187 & ~n11895 ) | ( n11894 & ~n11895 ) ;
  assign n11897 = ( n7811 & n10151 ) | ( n7811 & ~n11896 ) | ( n10151 & ~n11896 ) ;
  assign n11900 = n11899 ^ n11897 ^ n9089 ;
  assign n11902 = n9067 ^ n4434 ^ n3485 ;
  assign n11903 = n11902 ^ n10641 ^ n6369 ;
  assign n11901 = n3391 & n7398 ;
  assign n11904 = n11903 ^ n11901 ^ 1'b0 ;
  assign n11905 = n11900 | n11904 ;
  assign n11906 = n11504 ^ n4711 ^ n2558 ;
  assign n11907 = ( n4307 & n4544 ) | ( n4307 & n11906 ) | ( n4544 & n11906 ) ;
  assign n11908 = n11907 ^ n6000 ^ n1854 ;
  assign n11909 = n11908 ^ n6728 ^ n4575 ;
  assign n11910 = n582 ^ n581 ^ 1'b0 ;
  assign n11911 = n11909 & ~n11910 ;
  assign n11912 = n11041 ^ n5819 ^ n3746 ;
  assign n11913 = n5746 ^ n4388 ^ 1'b0 ;
  assign n11921 = n2931 & ~n7717 ;
  assign n11922 = n11921 ^ n6713 ^ 1'b0 ;
  assign n11918 = n1251 | n3377 ;
  assign n11919 = n5935 | n11918 ;
  assign n11916 = ( n620 & n1678 ) | ( n620 & ~n3275 ) | ( n1678 & ~n3275 ) ;
  assign n11917 = ( n1017 & n1916 ) | ( n1017 & n11916 ) | ( n1916 & n11916 ) ;
  assign n11920 = n11919 ^ n11917 ^ n5279 ;
  assign n11914 = ( n2891 & n7638 ) | ( n2891 & n8159 ) | ( n7638 & n8159 ) ;
  assign n11915 = n11914 ^ n1990 ^ 1'b0 ;
  assign n11923 = n11922 ^ n11920 ^ n11915 ;
  assign n11924 = ~n1176 & n4943 ;
  assign n11925 = n11924 ^ n1259 ^ 1'b0 ;
  assign n11926 = n8384 ^ n2287 ^ 1'b0 ;
  assign n11927 = n11925 & ~n11926 ;
  assign n11928 = ( n779 & ~n4105 ) | ( n779 & n11927 ) | ( ~n4105 & n11927 ) ;
  assign n11931 = n5097 ^ n4006 ^ n2515 ;
  assign n11929 = n6734 ^ n4490 ^ n3031 ;
  assign n11930 = n945 & ~n11929 ;
  assign n11932 = n11931 ^ n11930 ^ 1'b0 ;
  assign n11938 = ( n5321 & ~n5421 ) | ( n5321 & n7033 ) | ( ~n5421 & n7033 ) ;
  assign n11939 = ( n1088 & n4493 ) | ( n1088 & n11938 ) | ( n4493 & n11938 ) ;
  assign n11940 = n6596 ^ n3022 ^ 1'b0 ;
  assign n11941 = n11939 & n11940 ;
  assign n11942 = n11941 ^ n11045 ^ 1'b0 ;
  assign n11933 = n11359 ^ n8164 ^ x36 ;
  assign n11934 = n11933 ^ n8387 ^ n5503 ;
  assign n11935 = n11934 ^ n5602 ^ n2118 ;
  assign n11936 = ~n1056 & n3935 ;
  assign n11937 = n11935 & n11936 ;
  assign n11943 = n11942 ^ n11937 ^ n2964 ;
  assign n11944 = n4964 ^ n4130 ^ 1'b0 ;
  assign n11945 = ( n441 & ~n827 ) | ( n441 & n1461 ) | ( ~n827 & n1461 ) ;
  assign n11946 = n1444 | n11945 ;
  assign n11947 = ( n4590 & n4903 ) | ( n4590 & n11946 ) | ( n4903 & n11946 ) ;
  assign n11948 = ( n3815 & n6658 ) | ( n3815 & ~n11947 ) | ( n6658 & ~n11947 ) ;
  assign n11949 = n11948 ^ n11204 ^ n7398 ;
  assign n11950 = ( n2928 & ~n5093 ) | ( n2928 & n11949 ) | ( ~n5093 & n11949 ) ;
  assign n11951 = n9615 ^ n3046 ^ 1'b0 ;
  assign n11952 = ( n624 & ~n4756 ) | ( n624 & n11951 ) | ( ~n4756 & n11951 ) ;
  assign n11953 = n8249 ^ n4490 ^ 1'b0 ;
  assign n11954 = n11337 ^ n8052 ^ 1'b0 ;
  assign n11955 = ~n4878 & n11954 ;
  assign n11956 = n3911 & ~n6815 ;
  assign n11957 = ~n1538 & n11956 ;
  assign n11958 = ( n3685 & ~n5471 ) | ( n3685 & n11957 ) | ( ~n5471 & n11957 ) ;
  assign n11959 = n1108 & n3193 ;
  assign n11960 = ~n1978 & n11959 ;
  assign n11961 = n11960 ^ n7951 ^ 1'b0 ;
  assign n11962 = ( ~n8052 & n11958 ) | ( ~n8052 & n11961 ) | ( n11958 & n11961 ) ;
  assign n11966 = n10443 ^ n1714 ^ 1'b0 ;
  assign n11963 = n2244 ^ n975 ^ 1'b0 ;
  assign n11964 = n11218 & n11963 ;
  assign n11965 = ~n8788 & n11964 ;
  assign n11967 = n11966 ^ n11965 ^ n498 ;
  assign n11968 = n7082 | n10880 ;
  assign n11970 = n2722 | n4253 ;
  assign n11969 = ( n2052 & ~n6351 ) | ( n2052 & n7704 ) | ( ~n6351 & n7704 ) ;
  assign n11971 = n11970 ^ n11969 ^ 1'b0 ;
  assign n11972 = ( n4392 & ~n6991 ) | ( n4392 & n7717 ) | ( ~n6991 & n7717 ) ;
  assign n11973 = ( n1326 & n6460 ) | ( n1326 & n11258 ) | ( n6460 & n11258 ) ;
  assign n11974 = n4113 ^ n4058 ^ 1'b0 ;
  assign n11975 = ( n1037 & n4623 ) | ( n1037 & n11974 ) | ( n4623 & n11974 ) ;
  assign n11976 = n3888 | n6852 ;
  assign n11977 = n9378 | n11976 ;
  assign n11978 = n3619 ^ n1568 ^ n332 ;
  assign n11979 = ( n2692 & ~n4607 ) | ( n2692 & n11978 ) | ( ~n4607 & n11978 ) ;
  assign n11980 = ( n1029 & n8124 ) | ( n1029 & n11979 ) | ( n8124 & n11979 ) ;
  assign n11981 = n9211 ^ n555 ^ 1'b0 ;
  assign n11982 = n2151 | n11981 ;
  assign n11983 = ( n3582 & ~n8167 ) | ( n3582 & n11982 ) | ( ~n8167 & n11982 ) ;
  assign n11984 = ( n321 & ~n4115 ) | ( n321 & n4446 ) | ( ~n4115 & n4446 ) ;
  assign n11985 = n11984 ^ n179 ^ 1'b0 ;
  assign n11986 = n11985 ^ n10868 ^ 1'b0 ;
  assign n11987 = ( n4223 & n6065 ) | ( n4223 & ~n11986 ) | ( n6065 & ~n11986 ) ;
  assign n11988 = n10699 ^ n4925 ^ n2428 ;
  assign n11989 = n3790 ^ n3700 ^ 1'b0 ;
  assign n11990 = ~n11988 & n11989 ;
  assign n11994 = n148 & ~n11326 ;
  assign n11995 = ~n5916 & n11994 ;
  assign n11991 = n10398 ^ n4307 ^ n2440 ;
  assign n11992 = ~n10629 & n11991 ;
  assign n11993 = n11992 ^ n8462 ^ 1'b0 ;
  assign n11996 = n11995 ^ n11993 ^ n2049 ;
  assign n11997 = ( n5813 & ~n11990 ) | ( n5813 & n11996 ) | ( ~n11990 & n11996 ) ;
  assign n11998 = n7734 ^ n2280 ^ n671 ;
  assign n11999 = n11998 ^ n10318 ^ n8460 ;
  assign n12000 = ( n6098 & n6956 ) | ( n6098 & n11430 ) | ( n6956 & n11430 ) ;
  assign n12001 = n11074 | n12000 ;
  assign n12002 = ( n4896 & ~n7749 ) | ( n4896 & n11838 ) | ( ~n7749 & n11838 ) ;
  assign n12003 = ~n3446 & n5690 ;
  assign n12004 = ( ~x25 & n9335 ) | ( ~x25 & n12003 ) | ( n9335 & n12003 ) ;
  assign n12005 = n12004 ^ n5736 ^ n4570 ;
  assign n12006 = n12005 ^ n4674 ^ 1'b0 ;
  assign n12007 = ~n12002 & n12006 ;
  assign n12008 = n2547 ^ n1266 ^ x73 ;
  assign n12009 = n10456 | n12008 ;
  assign n12012 = n2889 ^ n2049 ^ 1'b0 ;
  assign n12013 = n441 & n12012 ;
  assign n12014 = n12013 ^ n8509 ^ 1'b0 ;
  assign n12015 = n7862 & ~n12014 ;
  assign n12016 = n12015 ^ n11463 ^ n7867 ;
  assign n12010 = n7565 ^ n7160 ^ x20 ;
  assign n12011 = ( ~n1694 & n9451 ) | ( ~n1694 & n12010 ) | ( n9451 & n12010 ) ;
  assign n12017 = n12016 ^ n12011 ^ n7757 ;
  assign n12018 = n975 | n3985 ;
  assign n12019 = n11083 & ~n12018 ;
  assign n12020 = n3656 ^ n2469 ^ 1'b0 ;
  assign n12021 = n8322 | n12020 ;
  assign n12022 = n5717 ^ x13 ^ 1'b0 ;
  assign n12023 = ~n8615 & n12022 ;
  assign n12024 = n12023 ^ n5058 ^ n4651 ;
  assign n12025 = ( ~n3631 & n5123 ) | ( ~n3631 & n12024 ) | ( n5123 & n12024 ) ;
  assign n12026 = ( ~n3186 & n10050 ) | ( ~n3186 & n12025 ) | ( n10050 & n12025 ) ;
  assign n12028 = n7972 ^ n3781 ^ 1'b0 ;
  assign n12029 = n1161 & ~n12028 ;
  assign n12030 = n12029 ^ n2865 ^ n2402 ;
  assign n12027 = n2995 | n11586 ;
  assign n12031 = n12030 ^ n12027 ^ n10597 ;
  assign n12032 = n8344 ^ n5818 ^ 1'b0 ;
  assign n12033 = n345 & ~n6175 ;
  assign n12034 = ~n12032 & n12033 ;
  assign n12035 = ( ~n1461 & n11108 ) | ( ~n1461 & n12034 ) | ( n11108 & n12034 ) ;
  assign n12036 = n1303 | n12035 ;
  assign n12037 = n8803 & ~n9844 ;
  assign n12038 = n1880 & n2167 ;
  assign n12039 = ~n1958 & n12038 ;
  assign n12040 = ( n1301 & ~n3881 ) | ( n1301 & n7259 ) | ( ~n3881 & n7259 ) ;
  assign n12041 = n4541 ^ n2018 ^ n698 ;
  assign n12042 = n4986 | n12041 ;
  assign n12043 = ( n12039 & n12040 ) | ( n12039 & n12042 ) | ( n12040 & n12042 ) ;
  assign n12044 = n12043 ^ n10096 ^ 1'b0 ;
  assign n12045 = ( ~n9835 & n10548 ) | ( ~n9835 & n12044 ) | ( n10548 & n12044 ) ;
  assign n12046 = ~n1875 & n3413 ;
  assign n12047 = n4427 | n12046 ;
  assign n12048 = n4765 | n12047 ;
  assign n12049 = ( n4361 & n5699 ) | ( n4361 & n12048 ) | ( n5699 & n12048 ) ;
  assign n12050 = ( n5490 & ~n5601 ) | ( n5490 & n12049 ) | ( ~n5601 & n12049 ) ;
  assign n12051 = n7627 ^ n7596 ^ 1'b0 ;
  assign n12052 = ( n2847 & n12050 ) | ( n2847 & n12051 ) | ( n12050 & n12051 ) ;
  assign n12057 = ( ~n423 & n926 ) | ( ~n423 & n2643 ) | ( n926 & n2643 ) ;
  assign n12058 = ( n5061 & n9014 ) | ( n5061 & n12057 ) | ( n9014 & n12057 ) ;
  assign n12053 = n5046 ^ n3079 ^ n719 ;
  assign n12054 = ~n1645 & n12053 ;
  assign n12055 = n12054 ^ n8109 ^ n566 ;
  assign n12056 = n12055 ^ n4867 ^ n3963 ;
  assign n12059 = n12058 ^ n12056 ^ n8055 ;
  assign n12060 = ( ~n2029 & n3008 ) | ( ~n2029 & n4079 ) | ( n3008 & n4079 ) ;
  assign n12061 = n12060 ^ n4452 ^ x43 ;
  assign n12062 = n1003 & n5149 ;
  assign n12063 = n8547 & n12062 ;
  assign n12064 = n2388 & ~n12063 ;
  assign n12065 = n9032 ^ n5721 ^ 1'b0 ;
  assign n12066 = ~n8537 & n12065 ;
  assign n12067 = n5052 | n5263 ;
  assign n12068 = n6123 ^ n1343 ^ n1322 ;
  assign n12069 = ( n664 & ~n8312 ) | ( n664 & n10201 ) | ( ~n8312 & n10201 ) ;
  assign n12070 = n7867 & ~n12069 ;
  assign n12071 = n12070 ^ x18 ^ 1'b0 ;
  assign n12072 = n6029 ^ n2995 ^ n2857 ;
  assign n12073 = n12071 | n12072 ;
  assign n12074 = n12073 ^ n5016 ^ 1'b0 ;
  assign n12075 = ( n2664 & n3308 ) | ( n2664 & ~n4866 ) | ( n3308 & ~n4866 ) ;
  assign n12076 = n12075 ^ n8976 ^ n3666 ;
  assign n12077 = ( n12068 & n12074 ) | ( n12068 & n12076 ) | ( n12074 & n12076 ) ;
  assign n12078 = ~n9938 & n12077 ;
  assign n12079 = n12078 ^ n7949 ^ 1'b0 ;
  assign n12080 = n2034 | n12079 ;
  assign n12081 = ( n1541 & n2954 ) | ( n1541 & ~n6233 ) | ( n2954 & ~n6233 ) ;
  assign n12082 = ( n8054 & n11184 ) | ( n8054 & n12081 ) | ( n11184 & n12081 ) ;
  assign n12083 = n12082 ^ n8152 ^ n2236 ;
  assign n12085 = n4074 ^ n2322 ^ 1'b0 ;
  assign n12084 = n6582 ^ n5778 ^ n3904 ;
  assign n12086 = n12085 ^ n12084 ^ 1'b0 ;
  assign n12087 = n10146 ^ n8342 ^ 1'b0 ;
  assign n12088 = n6551 ^ n710 ^ 1'b0 ;
  assign n12090 = n3988 ^ n866 ^ n562 ;
  assign n12089 = ( n617 & n3351 ) | ( n617 & ~n3411 ) | ( n3351 & ~n3411 ) ;
  assign n12091 = n12090 ^ n12089 ^ 1'b0 ;
  assign n12092 = n12091 ^ n5819 ^ n4755 ;
  assign n12093 = n243 | n1556 ;
  assign n12094 = n507 & ~n12093 ;
  assign n12095 = ( n1518 & n2439 ) | ( n1518 & n12094 ) | ( n2439 & n12094 ) ;
  assign n12096 = ( ~n1527 & n3090 ) | ( ~n1527 & n6010 ) | ( n3090 & n6010 ) ;
  assign n12097 = n12096 ^ n4878 ^ n4843 ;
  assign n12098 = ( ~n4687 & n5604 ) | ( ~n4687 & n12097 ) | ( n5604 & n12097 ) ;
  assign n12099 = n5525 | n12098 ;
  assign n12100 = n12099 ^ n5624 ^ 1'b0 ;
  assign n12101 = ( n1242 & n12095 ) | ( n1242 & ~n12100 ) | ( n12095 & ~n12100 ) ;
  assign n12102 = n12101 ^ n4308 ^ 1'b0 ;
  assign n12103 = n9067 | n11794 ;
  assign n12104 = n12103 ^ n6533 ^ 1'b0 ;
  assign n12105 = ~n4610 & n5013 ;
  assign n12106 = n12105 ^ n11258 ^ n8612 ;
  assign n12107 = ( n2138 & n12104 ) | ( n2138 & ~n12106 ) | ( n12104 & ~n12106 ) ;
  assign n12111 = n330 & ~n1655 ;
  assign n12108 = ( n1891 & n5091 ) | ( n1891 & ~n9782 ) | ( n5091 & ~n9782 ) ;
  assign n12109 = n8019 ^ n3607 ^ 1'b0 ;
  assign n12110 = ~n12108 & n12109 ;
  assign n12112 = n12111 ^ n12110 ^ n2978 ;
  assign n12113 = n1126 & ~n9072 ;
  assign n12114 = n12113 ^ n8496 ^ 1'b0 ;
  assign n12115 = ~n11773 & n12114 ;
  assign n12116 = ( n1669 & ~n4874 ) | ( n1669 & n8621 ) | ( ~n4874 & n8621 ) ;
  assign n12117 = ( n1239 & n6186 ) | ( n1239 & n8099 ) | ( n6186 & n8099 ) ;
  assign n12118 = n7795 ^ n326 ^ 1'b0 ;
  assign n12119 = n1422 ^ n129 ^ 1'b0 ;
  assign n12120 = ( ~n7824 & n12118 ) | ( ~n7824 & n12119 ) | ( n12118 & n12119 ) ;
  assign n12121 = ( x105 & n8127 ) | ( x105 & n9865 ) | ( n8127 & n9865 ) ;
  assign n12122 = ( n2996 & ~n6395 ) | ( n2996 & n9295 ) | ( ~n6395 & n9295 ) ;
  assign n12123 = n12122 ^ n5302 ^ 1'b0 ;
  assign n12129 = n1778 ^ n1460 ^ n137 ;
  assign n12130 = n4805 | n12129 ;
  assign n12131 = n12130 ^ n3173 ^ 1'b0 ;
  assign n12132 = n12131 ^ n12085 ^ n1925 ;
  assign n12133 = n12132 ^ n1460 ^ 1'b0 ;
  assign n12134 = n2624 & n12133 ;
  assign n12124 = ( n2313 & n2671 ) | ( n2313 & ~n2810 ) | ( n2671 & ~n2810 ) ;
  assign n12125 = x3 & ~n10806 ;
  assign n12126 = n12125 ^ n4402 ^ 1'b0 ;
  assign n12127 = ( n2802 & n4176 ) | ( n2802 & n12126 ) | ( n4176 & n12126 ) ;
  assign n12128 = ~n12124 & n12127 ;
  assign n12135 = n12134 ^ n12128 ^ 1'b0 ;
  assign n12136 = n5259 | n9800 ;
  assign n12137 = ( ~n7810 & n9245 ) | ( ~n7810 & n10634 ) | ( n9245 & n10634 ) ;
  assign n12138 = n11488 ^ n3617 ^ n2038 ;
  assign n12143 = ( x85 & ~n2403 ) | ( x85 & n4175 ) | ( ~n2403 & n4175 ) ;
  assign n12144 = ( n7441 & n7626 ) | ( n7441 & n12143 ) | ( n7626 & n12143 ) ;
  assign n12139 = n8649 ^ n2175 ^ x127 ;
  assign n12140 = n7030 ^ n3147 ^ n370 ;
  assign n12141 = ( n1414 & n12139 ) | ( n1414 & n12140 ) | ( n12139 & n12140 ) ;
  assign n12142 = ( n3702 & n6460 ) | ( n3702 & n12141 ) | ( n6460 & n12141 ) ;
  assign n12145 = n12144 ^ n12142 ^ 1'b0 ;
  assign n12146 = n10842 ^ n587 ^ 1'b0 ;
  assign n12147 = ~n1501 & n12146 ;
  assign n12150 = n8886 ^ n8808 ^ n3001 ;
  assign n12148 = n5897 | n8444 ;
  assign n12149 = ( n2785 & n11219 ) | ( n2785 & ~n12148 ) | ( n11219 & ~n12148 ) ;
  assign n12151 = n12150 ^ n12149 ^ n1276 ;
  assign n12152 = n3351 | n12151 ;
  assign n12153 = n7888 | n12152 ;
  assign n12154 = ( n1694 & n2449 ) | ( n1694 & n4606 ) | ( n2449 & n4606 ) ;
  assign n12155 = n12154 ^ n4751 ^ 1'b0 ;
  assign n12157 = n2851 | n4242 ;
  assign n12158 = n4915 & ~n12157 ;
  assign n12156 = n10843 ^ n10358 ^ n8591 ;
  assign n12159 = n12158 ^ n12156 ^ n4365 ;
  assign n12160 = n8738 ^ n4972 ^ 1'b0 ;
  assign n12161 = x126 & n12160 ;
  assign n12162 = ~n3718 & n12161 ;
  assign n12163 = n12162 ^ n5917 ^ 1'b0 ;
  assign n12164 = n12163 ^ n1916 ^ n1239 ;
  assign n12166 = n3178 ^ n1794 ^ n605 ;
  assign n12165 = ( x95 & n582 ) | ( x95 & ~n1982 ) | ( n582 & ~n1982 ) ;
  assign n12167 = n12166 ^ n12165 ^ n2357 ;
  assign n12168 = ( n2859 & ~n6990 ) | ( n2859 & n12108 ) | ( ~n6990 & n12108 ) ;
  assign n12169 = n12168 ^ n5260 ^ n1975 ;
  assign n12170 = n1262 & ~n6094 ;
  assign n12171 = n2918 ^ n1563 ^ n1533 ;
  assign n12172 = n3592 ^ n2058 ^ n1470 ;
  assign n12173 = ( n1234 & n1932 ) | ( n1234 & ~n12172 ) | ( n1932 & ~n12172 ) ;
  assign n12174 = ( n4779 & ~n7553 ) | ( n4779 & n12173 ) | ( ~n7553 & n12173 ) ;
  assign n12175 = ( n8399 & n12171 ) | ( n8399 & n12174 ) | ( n12171 & n12174 ) ;
  assign n12176 = n8744 ^ n8007 ^ n7809 ;
  assign n12177 = n12176 ^ n10136 ^ n7292 ;
  assign n12178 = n12177 ^ n3850 ^ n3788 ;
  assign n12179 = n6091 & n11895 ;
  assign n12180 = n1628 & n12179 ;
  assign n12183 = n7788 ^ n6240 ^ n740 ;
  assign n12181 = n3416 ^ n282 ^ 1'b0 ;
  assign n12182 = ( ~n551 & n12132 ) | ( ~n551 & n12181 ) | ( n12132 & n12181 ) ;
  assign n12184 = n12183 ^ n12182 ^ n2208 ;
  assign n12186 = n1047 | n7845 ;
  assign n12187 = n12186 ^ n3364 ^ 1'b0 ;
  assign n12188 = ( n889 & n1056 ) | ( n889 & n12187 ) | ( n1056 & n12187 ) ;
  assign n12189 = n1975 ^ n1838 ^ n403 ;
  assign n12190 = n12189 ^ n7514 ^ n6228 ;
  assign n12191 = n12190 ^ n4083 ^ n2471 ;
  assign n12192 = n12188 | n12191 ;
  assign n12193 = n12192 ^ n2834 ^ 1'b0 ;
  assign n12185 = n4750 & ~n9468 ;
  assign n12194 = n12193 ^ n12185 ^ n1126 ;
  assign n12195 = n4378 ^ n3473 ^ n1199 ;
  assign n12196 = ~n6477 & n12195 ;
  assign n12197 = n870 & n10023 ;
  assign n12198 = n12196 & n12197 ;
  assign n12199 = n12198 ^ n6494 ^ n1291 ;
  assign n12200 = n9992 ^ n4486 ^ n493 ;
  assign n12201 = n524 & n2923 ;
  assign n12202 = n3211 ^ n1238 ^ 1'b0 ;
  assign n12203 = ~n7192 & n12202 ;
  assign n12204 = ~n12201 & n12203 ;
  assign n12205 = n12204 ^ n4943 ^ 1'b0 ;
  assign n12206 = n12205 ^ n6063 ^ n2316 ;
  assign n12207 = n12206 ^ n8566 ^ 1'b0 ;
  assign n12208 = n12207 ^ n7905 ^ n2153 ;
  assign n12209 = ( ~n151 & n12200 ) | ( ~n151 & n12208 ) | ( n12200 & n12208 ) ;
  assign n12210 = ( ~n9539 & n12199 ) | ( ~n9539 & n12209 ) | ( n12199 & n12209 ) ;
  assign n12211 = n8359 ^ n2853 ^ n1874 ;
  assign n12212 = ( ~n10887 & n11698 ) | ( ~n10887 & n12211 ) | ( n11698 & n12211 ) ;
  assign n12213 = n997 & n7908 ;
  assign n12214 = ( n258 & n8180 ) | ( n258 & ~n12213 ) | ( n8180 & ~n12213 ) ;
  assign n12215 = n840 & n10901 ;
  assign n12216 = n12215 ^ n4342 ^ n2381 ;
  assign n12220 = n1704 & n3569 ;
  assign n12217 = n5794 ^ n3032 ^ 1'b0 ;
  assign n12218 = n6870 | n12217 ;
  assign n12219 = n12218 ^ n8403 ^ n4862 ;
  assign n12221 = n12220 ^ n12219 ^ 1'b0 ;
  assign n12231 = n4492 ^ n3208 ^ 1'b0 ;
  assign n12224 = ( n2978 & n4352 ) | ( n2978 & ~n6606 ) | ( n4352 & ~n6606 ) ;
  assign n12222 = n5381 ^ n5375 ^ n4749 ;
  assign n12223 = n11042 | n12222 ;
  assign n12225 = n12224 ^ n12223 ^ 1'b0 ;
  assign n12226 = ( ~n1963 & n4348 ) | ( ~n1963 & n9805 ) | ( n4348 & n9805 ) ;
  assign n12227 = ~n1210 & n5429 ;
  assign n12228 = ( ~n1799 & n8025 ) | ( ~n1799 & n12227 ) | ( n8025 & n12227 ) ;
  assign n12229 = n12226 & n12228 ;
  assign n12230 = ~n12225 & n12229 ;
  assign n12232 = n12231 ^ n12230 ^ n9505 ;
  assign n12233 = n9727 ^ n6835 ^ n5578 ;
  assign n12234 = n10079 ^ n2111 ^ 1'b0 ;
  assign n12235 = n12234 ^ n5890 ^ 1'b0 ;
  assign n12236 = n12233 & n12235 ;
  assign n12237 = n2101 ^ n1627 ^ x45 ;
  assign n12238 = ( n2289 & n4876 ) | ( n2289 & n8437 ) | ( n4876 & n8437 ) ;
  assign n12239 = n12237 & n12238 ;
  assign n12240 = ~n2256 & n12239 ;
  assign n12241 = ( ~n4322 & n10488 ) | ( ~n4322 & n12240 ) | ( n10488 & n12240 ) ;
  assign n12242 = n8976 ^ n7792 ^ n7059 ;
  assign n12243 = ( ~n3408 & n7465 ) | ( ~n3408 & n9769 ) | ( n7465 & n9769 ) ;
  assign n12244 = n8641 ^ n7674 ^ 1'b0 ;
  assign n12245 = n12243 & n12244 ;
  assign n12246 = ( n9335 & n12242 ) | ( n9335 & n12245 ) | ( n12242 & n12245 ) ;
  assign n12251 = n1527 | n7344 ;
  assign n12249 = ( n2295 & ~n4252 ) | ( n2295 & n10041 ) | ( ~n4252 & n10041 ) ;
  assign n12247 = n3565 & ~n10283 ;
  assign n12248 = n4285 & n12247 ;
  assign n12250 = n12249 ^ n12248 ^ n1086 ;
  assign n12252 = n12251 ^ n12250 ^ 1'b0 ;
  assign n12253 = ~n4497 & n12252 ;
  assign n12254 = ( n1575 & n5106 ) | ( n1575 & ~n11744 ) | ( n5106 & ~n11744 ) ;
  assign n12255 = ( n2763 & ~n6494 ) | ( n2763 & n8043 ) | ( ~n6494 & n8043 ) ;
  assign n12265 = ~n3922 & n5376 ;
  assign n12266 = n12265 ^ n1131 ^ 1'b0 ;
  assign n12263 = n10221 ^ n10020 ^ n3046 ;
  assign n12264 = ~n8309 & n12263 ;
  assign n12267 = n12266 ^ n12264 ^ 1'b0 ;
  assign n12256 = ~n1986 & n4925 ;
  assign n12257 = n3655 & n6344 ;
  assign n12258 = n12257 ^ n2375 ^ 1'b0 ;
  assign n12259 = n12256 & n12258 ;
  assign n12260 = n10598 & n12259 ;
  assign n12261 = n12260 ^ n11525 ^ n5948 ;
  assign n12262 = ( n1265 & ~n11041 ) | ( n1265 & n12261 ) | ( ~n11041 & n12261 ) ;
  assign n12268 = n12267 ^ n12262 ^ 1'b0 ;
  assign n12269 = n10379 ^ n6828 ^ n2965 ;
  assign n12271 = n7601 ^ n1549 ^ n1265 ;
  assign n12272 = ( ~n2602 & n4739 ) | ( ~n2602 & n12271 ) | ( n4739 & n12271 ) ;
  assign n12270 = ~n352 & n5432 ;
  assign n12273 = n12272 ^ n12270 ^ 1'b0 ;
  assign n12274 = n12273 ^ n1789 ^ 1'b0 ;
  assign n12275 = n10241 ^ n6100 ^ 1'b0 ;
  assign n12276 = n12275 ^ n5526 ^ n392 ;
  assign n12277 = n5150 ^ n4659 ^ 1'b0 ;
  assign n12278 = n7065 & ~n12277 ;
  assign n12279 = n8553 ^ n2483 ^ 1'b0 ;
  assign n12280 = n12278 & ~n12279 ;
  assign n12281 = n9202 ^ n3438 ^ 1'b0 ;
  assign n12282 = n6183 & ~n12281 ;
  assign n12283 = n10875 ^ n3464 ^ 1'b0 ;
  assign n12284 = ~n2654 & n12283 ;
  assign n12285 = n5740 ^ n4072 ^ n528 ;
  assign n12286 = n4517 & n5269 ;
  assign n12287 = n12286 ^ n2255 ^ 1'b0 ;
  assign n12288 = ( n5494 & n6951 ) | ( n5494 & ~n12287 ) | ( n6951 & ~n12287 ) ;
  assign n12289 = ( ~n4234 & n4948 ) | ( ~n4234 & n6029 ) | ( n4948 & n6029 ) ;
  assign n12290 = n12289 ^ n3530 ^ 1'b0 ;
  assign n12291 = ~n1617 & n12290 ;
  assign n12292 = ( n4326 & n12288 ) | ( n4326 & ~n12291 ) | ( n12288 & ~n12291 ) ;
  assign n12293 = n5738 & n11120 ;
  assign n12294 = ~n439 & n12293 ;
  assign n12295 = n1998 | n11683 ;
  assign n12296 = n11799 | n12295 ;
  assign n12297 = n12296 ^ n8620 ^ n1212 ;
  assign n12298 = ( n4299 & ~n7936 ) | ( n4299 & n12297 ) | ( ~n7936 & n12297 ) ;
  assign n12299 = ( n4915 & n6471 ) | ( n4915 & n12298 ) | ( n6471 & n12298 ) ;
  assign n12300 = n8903 ^ n4855 ^ 1'b0 ;
  assign n12301 = n12300 ^ n8358 ^ n1290 ;
  assign n12302 = n10350 ^ n9607 ^ n8282 ;
  assign n12303 = n7620 ^ n6114 ^ 1'b0 ;
  assign n12304 = n9184 & n12303 ;
  assign n12305 = n3966 | n9120 ;
  assign n12306 = n12305 ^ n10860 ^ 1'b0 ;
  assign n12307 = ( n3454 & ~n7350 ) | ( n3454 & n10963 ) | ( ~n7350 & n10963 ) ;
  assign n12308 = n12306 & ~n12307 ;
  assign n12309 = n12308 ^ n11682 ^ 1'b0 ;
  assign n12314 = n4292 ^ n2512 ^ 1'b0 ;
  assign n12315 = ~n4935 & n12314 ;
  assign n12310 = n170 | n2965 ;
  assign n12311 = n12310 ^ n8316 ^ 1'b0 ;
  assign n12312 = n12311 ^ n7435 ^ n4662 ;
  assign n12313 = n9361 & n12312 ;
  assign n12316 = n12315 ^ n12313 ^ 1'b0 ;
  assign n12317 = n2279 & n12316 ;
  assign n12318 = n789 & n12317 ;
  assign n12319 = n12318 ^ n9124 ^ n3247 ;
  assign n12320 = ( n1882 & n7017 ) | ( n1882 & n11505 ) | ( n7017 & n11505 ) ;
  assign n12321 = ( n774 & n10468 ) | ( n774 & n12320 ) | ( n10468 & n12320 ) ;
  assign n12322 = n4455 ^ n603 ^ 1'b0 ;
  assign n12323 = n3940 & n12322 ;
  assign n12324 = n4088 ^ n3276 ^ n2600 ;
  assign n12325 = ( n2101 & ~n4655 ) | ( n2101 & n12324 ) | ( ~n4655 & n12324 ) ;
  assign n12326 = n12325 ^ n10488 ^ n459 ;
  assign n12327 = n12326 ^ n6140 ^ 1'b0 ;
  assign n12328 = n12327 ^ n8652 ^ n6516 ;
  assign n12329 = n12328 ^ n2066 ^ 1'b0 ;
  assign n12330 = n8421 | n12329 ;
  assign n12331 = ( n2596 & n4832 ) | ( n2596 & ~n5493 ) | ( n4832 & ~n5493 ) ;
  assign n12332 = n7194 ^ n907 ^ x109 ;
  assign n12333 = n4628 | n12332 ;
  assign n12334 = n12333 ^ n11579 ^ n2202 ;
  assign n12335 = n5644 ^ n5638 ^ n4579 ;
  assign n12336 = n12334 & n12335 ;
  assign n12337 = ~n12331 & n12336 ;
  assign n12338 = n3925 | n12337 ;
  assign n12339 = n866 & ~n12338 ;
  assign n12340 = n12339 ^ n8710 ^ n3905 ;
  assign n12341 = n6299 ^ n4937 ^ 1'b0 ;
  assign n12342 = n2377 | n12341 ;
  assign n12343 = n12342 ^ n8170 ^ n5956 ;
  assign n12344 = n12343 ^ n4300 ^ 1'b0 ;
  assign n12345 = ~n4646 & n12344 ;
  assign n12351 = ( n1136 & n3653 ) | ( n1136 & n6136 ) | ( n3653 & n6136 ) ;
  assign n12352 = n6136 | n7234 ;
  assign n12353 = ( n6754 & ~n12351 ) | ( n6754 & n12352 ) | ( ~n12351 & n12352 ) ;
  assign n12354 = ( n6792 & n7788 ) | ( n6792 & n12353 ) | ( n7788 & n12353 ) ;
  assign n12346 = ( n415 & ~n838 ) | ( n415 & n3081 ) | ( ~n838 & n3081 ) ;
  assign n12347 = n12346 ^ n3096 ^ 1'b0 ;
  assign n12348 = n12347 ^ n4588 ^ n1998 ;
  assign n12349 = n12348 ^ n9999 ^ 1'b0 ;
  assign n12350 = n6923 & n12349 ;
  assign n12355 = n12354 ^ n12350 ^ 1'b0 ;
  assign n12364 = n5547 ^ n1024 ^ 1'b0 ;
  assign n12365 = n3788 & n12364 ;
  assign n12361 = ( ~n223 & n1228 ) | ( ~n223 & n3117 ) | ( n1228 & n3117 ) ;
  assign n12356 = n994 ^ n693 ^ n264 ;
  assign n12357 = n12356 ^ n7146 ^ n2179 ;
  assign n12358 = n5616 & n12357 ;
  assign n12359 = n12358 ^ n6714 ^ 1'b0 ;
  assign n12360 = ( n1391 & ~n4369 ) | ( n1391 & n12359 ) | ( ~n4369 & n12359 ) ;
  assign n12362 = n12361 ^ n12360 ^ n4567 ;
  assign n12363 = n12362 ^ n9826 ^ n7214 ;
  assign n12366 = n12365 ^ n12363 ^ 1'b0 ;
  assign n12367 = ~n8128 & n12102 ;
  assign n12368 = n12367 ^ n1574 ^ 1'b0 ;
  assign n12369 = n10623 ^ n10090 ^ 1'b0 ;
  assign n12370 = ~n2383 & n2419 ;
  assign n12371 = n2576 & n12370 ;
  assign n12372 = ( x81 & n151 ) | ( x81 & n3821 ) | ( n151 & n3821 ) ;
  assign n12373 = n12372 ^ n1031 ^ 1'b0 ;
  assign n12374 = n540 | n12373 ;
  assign n12375 = ( n632 & n5232 ) | ( n632 & ~n10210 ) | ( n5232 & ~n10210 ) ;
  assign n12376 = n12375 ^ n9736 ^ n6386 ;
  assign n12377 = n12376 ^ n7134 ^ n5376 ;
  assign n12378 = n12374 & n12377 ;
  assign n12380 = n435 & n3654 ;
  assign n12381 = n3385 & ~n12380 ;
  assign n12382 = n12381 ^ n3536 ^ 1'b0 ;
  assign n12379 = n5892 | n7481 ;
  assign n12383 = n12382 ^ n12379 ^ 1'b0 ;
  assign n12384 = n6165 ^ n5074 ^ 1'b0 ;
  assign n12385 = n7613 ^ n4352 ^ n1655 ;
  assign n12386 = n1984 & n3045 ;
  assign n12387 = ( n12384 & n12385 ) | ( n12384 & ~n12386 ) | ( n12385 & ~n12386 ) ;
  assign n12388 = n12387 ^ n9941 ^ n6746 ;
  assign n12389 = ( n421 & n7701 ) | ( n421 & n8961 ) | ( n7701 & n8961 ) ;
  assign n12390 = ( n5788 & n6126 ) | ( n5788 & n9101 ) | ( n6126 & n9101 ) ;
  assign n12391 = ( n217 & ~n486 ) | ( n217 & n2230 ) | ( ~n486 & n2230 ) ;
  assign n12392 = n4711 ^ n3532 ^ 1'b0 ;
  assign n12393 = n8105 ^ n613 ^ 1'b0 ;
  assign n12394 = ( n6746 & n12392 ) | ( n6746 & n12393 ) | ( n12392 & n12393 ) ;
  assign n12395 = n12394 ^ n11799 ^ n723 ;
  assign n12396 = n11579 ^ n11317 ^ n9140 ;
  assign n12397 = n6514 ^ n1878 ^ 1'b0 ;
  assign n12398 = n745 | n12397 ;
  assign n12399 = ( n711 & n1096 ) | ( n711 & n12398 ) | ( n1096 & n12398 ) ;
  assign n12400 = ( n2798 & ~n4424 ) | ( n2798 & n12399 ) | ( ~n4424 & n12399 ) ;
  assign n12401 = ~n1482 & n12400 ;
  assign n12402 = n12396 & n12401 ;
  assign n12403 = ( ~n7170 & n9582 ) | ( ~n7170 & n10748 ) | ( n9582 & n10748 ) ;
  assign n12404 = n8282 ^ n5854 ^ 1'b0 ;
  assign n12405 = ~n2045 & n12404 ;
  assign n12406 = ( n6481 & ~n12403 ) | ( n6481 & n12405 ) | ( ~n12403 & n12405 ) ;
  assign n12407 = ( n2972 & n4159 ) | ( n2972 & ~n10222 ) | ( n4159 & ~n10222 ) ;
  assign n12408 = n205 & ~n12407 ;
  assign n12409 = ~x38 & n12408 ;
  assign n12410 = ( n4034 & n4674 ) | ( n4034 & n12409 ) | ( n4674 & n12409 ) ;
  assign n12411 = n5564 ^ n2660 ^ 1'b0 ;
  assign n12412 = n5439 ^ n1634 ^ n1262 ;
  assign n12413 = n12412 ^ n10566 ^ n4216 ;
  assign n12414 = n12413 ^ n11561 ^ 1'b0 ;
  assign n12415 = n12414 ^ n12085 ^ n2644 ;
  assign n12416 = n237 & ~n6037 ;
  assign n12417 = ( n549 & ~n1181 ) | ( n549 & n12416 ) | ( ~n1181 & n12416 ) ;
  assign n12418 = ( ~n3194 & n9672 ) | ( ~n3194 & n11553 ) | ( n9672 & n11553 ) ;
  assign n12419 = ( n4114 & n9409 ) | ( n4114 & n12418 ) | ( n9409 & n12418 ) ;
  assign n12429 = n12124 ^ n3331 ^ n2423 ;
  assign n12420 = ( n3997 & ~n4547 ) | ( n3997 & n12003 ) | ( ~n4547 & n12003 ) ;
  assign n12421 = ( n845 & n896 ) | ( n845 & ~n6073 ) | ( n896 & ~n6073 ) ;
  assign n12422 = n12421 ^ n8468 ^ n2140 ;
  assign n12423 = n8660 | n12422 ;
  assign n12424 = n12423 ^ n6642 ^ 1'b0 ;
  assign n12425 = x114 & n11961 ;
  assign n12426 = n12425 ^ n8475 ^ 1'b0 ;
  assign n12427 = n12424 | n12426 ;
  assign n12428 = ( n1633 & ~n12420 ) | ( n1633 & n12427 ) | ( ~n12420 & n12427 ) ;
  assign n12430 = n12429 ^ n12428 ^ n6864 ;
  assign n12431 = n12419 & n12430 ;
  assign n12432 = ( ~n4848 & n11568 ) | ( ~n4848 & n11947 ) | ( n11568 & n11947 ) ;
  assign n12433 = ( n4641 & ~n5702 ) | ( n4641 & n9931 ) | ( ~n5702 & n9931 ) ;
  assign n12434 = n12433 ^ n6314 ^ n5462 ;
  assign n12435 = n10403 | n12434 ;
  assign n12436 = n12432 | n12435 ;
  assign n12437 = ~n3408 & n10898 ;
  assign n12438 = n12437 ^ n4988 ^ 1'b0 ;
  assign n12439 = n1551 | n1644 ;
  assign n12440 = n12172 | n12439 ;
  assign n12441 = n2306 & n12440 ;
  assign n12442 = x72 & n8786 ;
  assign n12443 = n12442 ^ n981 ^ 1'b0 ;
  assign n12444 = n1623 & n4802 ;
  assign n12445 = n12444 ^ n379 ^ 1'b0 ;
  assign n12446 = n5866 ^ n3898 ^ 1'b0 ;
  assign n12447 = ( n3766 & ~n4943 ) | ( n3766 & n9102 ) | ( ~n4943 & n9102 ) ;
  assign n12448 = ( ~n3620 & n4761 ) | ( ~n3620 & n5070 ) | ( n4761 & n5070 ) ;
  assign n12449 = n12448 ^ n9475 ^ n2898 ;
  assign n12450 = ( n8658 & n12447 ) | ( n8658 & ~n12449 ) | ( n12447 & ~n12449 ) ;
  assign n12451 = ( ~n811 & n1055 ) | ( ~n811 & n1862 ) | ( n1055 & n1862 ) ;
  assign n12452 = n12451 ^ x1 ^ 1'b0 ;
  assign n12453 = n12450 & ~n12452 ;
  assign n12454 = ( ~x121 & n2025 ) | ( ~x121 & n7031 ) | ( n2025 & n7031 ) ;
  assign n12455 = n410 & n573 ;
  assign n12456 = ~n1784 & n12455 ;
  assign n12457 = n12456 ^ n12230 ^ n4848 ;
  assign n12458 = ~n1739 & n5075 ;
  assign n12459 = ( n2417 & n6543 ) | ( n2417 & n12458 ) | ( n6543 & n12458 ) ;
  assign n12460 = ( n6524 & n12457 ) | ( n6524 & ~n12459 ) | ( n12457 & ~n12459 ) ;
  assign n12461 = n3852 ^ n1900 ^ n258 ;
  assign n12463 = n2097 & ~n7003 ;
  assign n12464 = n12463 ^ n5892 ^ 1'b0 ;
  assign n12465 = n12464 ^ n10073 ^ n5433 ;
  assign n12462 = ~n7855 & n12001 ;
  assign n12466 = n12465 ^ n12462 ^ 1'b0 ;
  assign n12467 = n3021 & ~n3557 ;
  assign n12468 = ( ~n1941 & n8043 ) | ( ~n1941 & n12467 ) | ( n8043 & n12467 ) ;
  assign n12469 = ( n844 & n1261 ) | ( n844 & n6471 ) | ( n1261 & n6471 ) ;
  assign n12470 = ( n5718 & n11845 ) | ( n5718 & n12469 ) | ( n11845 & n12469 ) ;
  assign n12471 = n1932 & n2480 ;
  assign n12472 = n12471 ^ n8315 ^ n5139 ;
  assign n12473 = ( n2258 & n9656 ) | ( n2258 & n12472 ) | ( n9656 & n12472 ) ;
  assign n12478 = n7280 ^ n2389 ^ n201 ;
  assign n12479 = n12478 ^ n5969 ^ n2081 ;
  assign n12474 = ~n1784 & n9449 ;
  assign n12475 = n5910 & n12474 ;
  assign n12476 = n8166 ^ n5937 ^ 1'b0 ;
  assign n12477 = ~n12475 & n12476 ;
  assign n12480 = n12479 ^ n12477 ^ 1'b0 ;
  assign n12482 = n12260 ^ n8223 ^ 1'b0 ;
  assign n12483 = n1459 & n12482 ;
  assign n12481 = ( n349 & ~n4777 ) | ( n349 & n6238 ) | ( ~n4777 & n6238 ) ;
  assign n12484 = n12483 ^ n12481 ^ 1'b0 ;
  assign n12485 = n12480 & n12484 ;
  assign n12486 = n10251 ^ n9678 ^ n2712 ;
  assign n12487 = n12486 ^ n8032 ^ n2607 ;
  assign n12488 = n12487 ^ n1750 ^ n1025 ;
  assign n12489 = ( n250 & n1367 ) | ( n250 & ~n9619 ) | ( n1367 & ~n9619 ) ;
  assign n12490 = n1809 | n9735 ;
  assign n12491 = ( n1013 & n12489 ) | ( n1013 & ~n12490 ) | ( n12489 & ~n12490 ) ;
  assign n12493 = n10620 ^ n7912 ^ n2058 ;
  assign n12492 = n8701 & ~n12393 ;
  assign n12494 = n12493 ^ n12492 ^ 1'b0 ;
  assign n12495 = n11312 ^ n4446 ^ 1'b0 ;
  assign n12501 = ( n2896 & ~n6967 ) | ( n2896 & n8147 ) | ( ~n6967 & n8147 ) ;
  assign n12498 = ~n545 & n3017 ;
  assign n12499 = ( n1050 & n1512 ) | ( n1050 & n12498 ) | ( n1512 & n12498 ) ;
  assign n12500 = n12499 ^ n8797 ^ n1056 ;
  assign n12502 = n12501 ^ n12500 ^ n3391 ;
  assign n12496 = n2751 ^ n1036 ^ 1'b0 ;
  assign n12497 = n8751 | n12496 ;
  assign n12503 = n12502 ^ n12497 ^ n1330 ;
  assign n12504 = ( n1420 & n2541 ) | ( n1420 & n6065 ) | ( n2541 & n6065 ) ;
  assign n12505 = n3433 | n7608 ;
  assign n12506 = ~n2216 & n12505 ;
  assign n12507 = ( n1195 & n12504 ) | ( n1195 & ~n12506 ) | ( n12504 & ~n12506 ) ;
  assign n12508 = n1889 & ~n11774 ;
  assign n12509 = ( n4046 & n7896 ) | ( n4046 & n8806 ) | ( n7896 & n8806 ) ;
  assign n12510 = ~n3952 & n12509 ;
  assign n12511 = n12510 ^ n5807 ^ 1'b0 ;
  assign n12512 = n223 | n1563 ;
  assign n12513 = ( n553 & n6669 ) | ( n553 & ~n8639 ) | ( n6669 & ~n8639 ) ;
  assign n12514 = ( n528 & n12512 ) | ( n528 & n12513 ) | ( n12512 & n12513 ) ;
  assign n12515 = n5980 ^ n1734 ^ 1'b0 ;
  assign n12516 = n8633 | n12515 ;
  assign n12517 = n12514 | n12516 ;
  assign n12518 = n12517 ^ n8859 ^ 1'b0 ;
  assign n12519 = ~n2951 & n12518 ;
  assign n12520 = n6503 ^ n4093 ^ n2919 ;
  assign n12521 = n12520 ^ n10339 ^ n2078 ;
  assign n12522 = n2418 ^ n1805 ^ n641 ;
  assign n12523 = n12522 ^ n4176 ^ n500 ;
  assign n12524 = n12523 ^ n9730 ^ n2428 ;
  assign n12525 = n3737 & ~n7891 ;
  assign n12526 = n12525 ^ n11701 ^ n3266 ;
  assign n12527 = n12526 ^ n8920 ^ n6478 ;
  assign n12528 = n3927 ^ x74 ^ 1'b0 ;
  assign n12529 = n12528 ^ n5595 ^ n3744 ;
  assign n12534 = ( n1177 & n2834 ) | ( n1177 & ~n6951 ) | ( n2834 & ~n6951 ) ;
  assign n12533 = n10226 ^ n1981 ^ n1911 ;
  assign n12530 = n8198 ^ n1360 ^ 1'b0 ;
  assign n12531 = x75 & ~n12530 ;
  assign n12532 = ( ~x112 & n4496 ) | ( ~x112 & n12531 ) | ( n4496 & n12531 ) ;
  assign n12535 = n12534 ^ n12533 ^ n12532 ;
  assign n12536 = n12398 ^ n1966 ^ 1'b0 ;
  assign n12537 = n7174 | n12536 ;
  assign n12538 = n2331 ^ n919 ^ 1'b0 ;
  assign n12539 = ~n1002 & n12538 ;
  assign n12540 = n12539 ^ n2506 ^ 1'b0 ;
  assign n12541 = n4478 & ~n12540 ;
  assign n12542 = n12541 ^ n9644 ^ 1'b0 ;
  assign n12543 = ~n3439 & n12542 ;
  assign n12546 = n10916 ^ n4359 ^ n646 ;
  assign n12547 = n6900 & n12546 ;
  assign n12548 = n12547 ^ n2780 ^ 1'b0 ;
  assign n12544 = n5984 ^ n3381 ^ 1'b0 ;
  assign n12545 = n12544 ^ n4430 ^ n4070 ;
  assign n12549 = n12548 ^ n12545 ^ 1'b0 ;
  assign n12550 = n2060 | n5699 ;
  assign n12554 = n2421 & ~n10058 ;
  assign n12555 = n12554 ^ n5753 ^ 1'b0 ;
  assign n12553 = n9544 ^ n3340 ^ n2261 ;
  assign n12551 = ( n3689 & ~n6348 ) | ( n3689 & n10521 ) | ( ~n6348 & n10521 ) ;
  assign n12552 = n12551 ^ n3935 ^ n653 ;
  assign n12556 = n12555 ^ n12553 ^ n12552 ;
  assign n12557 = n12556 ^ n4304 ^ 1'b0 ;
  assign n12558 = n559 & ~n5053 ;
  assign n12559 = n1845 & n12558 ;
  assign n12560 = n12559 ^ n3270 ^ 1'b0 ;
  assign n12561 = ( n4098 & ~n8088 ) | ( n4098 & n12560 ) | ( ~n8088 & n12560 ) ;
  assign n12562 = n923 & n10946 ;
  assign n12563 = n12562 ^ n6304 ^ 1'b0 ;
  assign n12564 = n7306 | n12108 ;
  assign n12565 = n12564 ^ n3693 ^ 1'b0 ;
  assign n12566 = ( ~n2372 & n6675 ) | ( ~n2372 & n12565 ) | ( n6675 & n12565 ) ;
  assign n12567 = n12566 ^ n4270 ^ 1'b0 ;
  assign n12568 = ~n8420 & n12567 ;
  assign n12569 = n5391 ^ n3817 ^ n3243 ;
  assign n12570 = n11363 ^ n9973 ^ 1'b0 ;
  assign n12571 = n12570 ^ n9990 ^ 1'b0 ;
  assign n12572 = n12569 | n12571 ;
  assign n12576 = ( ~n793 & n2969 ) | ( ~n793 & n3710 ) | ( n2969 & n3710 ) ;
  assign n12577 = ( ~n4305 & n8503 ) | ( ~n4305 & n12576 ) | ( n8503 & n12576 ) ;
  assign n12578 = ( ~n1890 & n4128 ) | ( ~n1890 & n12577 ) | ( n4128 & n12577 ) ;
  assign n12573 = n153 | n8652 ;
  assign n12574 = n9331 & ~n12573 ;
  assign n12575 = n1878 & n12574 ;
  assign n12579 = n12578 ^ n12575 ^ 1'b0 ;
  assign n12580 = x33 & n12579 ;
  assign n12581 = n1340 & n5753 ;
  assign n12582 = ( n4569 & ~n8469 ) | ( n4569 & n8931 ) | ( ~n8469 & n8931 ) ;
  assign n12585 = n9805 ^ n2928 ^ 1'b0 ;
  assign n12586 = n9037 ^ n2727 ^ 1'b0 ;
  assign n12587 = n12586 ^ n1709 ^ 1'b0 ;
  assign n12588 = n12585 | n12587 ;
  assign n12583 = ( n2074 & n5032 ) | ( n2074 & n5199 ) | ( n5032 & n5199 ) ;
  assign n12584 = n11985 & n12583 ;
  assign n12589 = n12588 ^ n12584 ^ 1'b0 ;
  assign n12590 = n12332 ^ n2136 ^ 1'b0 ;
  assign n12591 = n12590 ^ n5822 ^ n3115 ;
  assign n12592 = ( n5738 & n9098 ) | ( n5738 & ~n10764 ) | ( n9098 & ~n10764 ) ;
  assign n12593 = n8892 ^ n7359 ^ n6713 ;
  assign n12594 = ( n461 & ~n7546 ) | ( n461 & n12593 ) | ( ~n7546 & n12593 ) ;
  assign n12595 = n9793 | n12594 ;
  assign n12596 = n5601 | n12595 ;
  assign n12597 = n6397 & ~n12596 ;
  assign n12598 = ( n1951 & n4467 ) | ( n1951 & n8383 ) | ( n4467 & n8383 ) ;
  assign n12599 = ( n4846 & ~n7780 ) | ( n4846 & n12598 ) | ( ~n7780 & n12598 ) ;
  assign n12600 = ( n5968 & n6365 ) | ( n5968 & n8146 ) | ( n6365 & n8146 ) ;
  assign n12601 = n9701 ^ n3878 ^ 1'b0 ;
  assign n12602 = n651 & ~n12601 ;
  assign n12603 = ( n3592 & n11024 ) | ( n3592 & n12602 ) | ( n11024 & n12602 ) ;
  assign n12604 = ( n525 & n668 ) | ( n525 & n5152 ) | ( n668 & n5152 ) ;
  assign n12605 = n12604 ^ n12555 ^ n3065 ;
  assign n12606 = ( n11853 & n12323 ) | ( n11853 & ~n12605 ) | ( n12323 & ~n12605 ) ;
  assign n12607 = n12606 ^ n12343 ^ n8201 ;
  assign n12608 = n12275 ^ n9749 ^ n255 ;
  assign n12609 = ( n2663 & ~n7094 ) | ( n2663 & n12608 ) | ( ~n7094 & n12608 ) ;
  assign n12610 = n9447 ^ n4346 ^ n275 ;
  assign n12611 = n11698 ^ n1878 ^ n337 ;
  assign n12622 = n9247 & ~n10809 ;
  assign n12612 = n9677 ^ n847 ^ 1'b0 ;
  assign n12613 = n4637 & ~n12612 ;
  assign n12615 = n7400 & n7977 ;
  assign n12614 = n1677 & ~n6956 ;
  assign n12616 = n12615 ^ n12614 ^ 1'b0 ;
  assign n12617 = ( ~n5744 & n11108 ) | ( ~n5744 & n12616 ) | ( n11108 & n12616 ) ;
  assign n12618 = n12617 ^ n9156 ^ n3123 ;
  assign n12619 = ( n9602 & n12613 ) | ( n9602 & n12618 ) | ( n12613 & n12618 ) ;
  assign n12620 = n4779 ^ n1975 ^ 1'b0 ;
  assign n12621 = ~n12619 & n12620 ;
  assign n12623 = n12622 ^ n12621 ^ 1'b0 ;
  assign n12624 = n12611 & n12623 ;
  assign n12625 = n10207 ^ n6102 ^ n2467 ;
  assign n12630 = n1162 & ~n12544 ;
  assign n12626 = n10973 ^ n5152 ^ n3851 ;
  assign n12627 = n12626 ^ n6598 ^ n5732 ;
  assign n12628 = n1267 & n12627 ;
  assign n12629 = n12628 ^ n2482 ^ 1'b0 ;
  assign n12631 = n12630 ^ n12629 ^ n2821 ;
  assign n12633 = n1399 & n2224 ;
  assign n12634 = ~n4728 & n12633 ;
  assign n12635 = ( n1362 & n4819 ) | ( n1362 & n12634 ) | ( n4819 & n12634 ) ;
  assign n12636 = n12635 ^ n5270 ^ 1'b0 ;
  assign n12632 = n10739 ^ n9611 ^ n5488 ;
  assign n12637 = n12636 ^ n12632 ^ n4813 ;
  assign n12638 = ( ~n3339 & n6240 ) | ( ~n3339 & n11907 ) | ( n6240 & n11907 ) ;
  assign n12639 = ( n1573 & n6445 ) | ( n1573 & ~n11388 ) | ( n6445 & ~n11388 ) ;
  assign n12640 = n6581 | n11885 ;
  assign n12641 = n12639 & ~n12640 ;
  assign n12642 = ~n4003 & n4242 ;
  assign n12643 = n4034 ^ n645 ^ 1'b0 ;
  assign n12644 = ( n569 & n1366 ) | ( n569 & n12643 ) | ( n1366 & n12643 ) ;
  assign n12645 = n12642 & ~n12644 ;
  assign n12650 = n5851 ^ n4241 ^ n1936 ;
  assign n12646 = ( ~n328 & n2898 ) | ( ~n328 & n7988 ) | ( n2898 & n7988 ) ;
  assign n12647 = n11317 | n12646 ;
  assign n12648 = n12647 ^ n8140 ^ 1'b0 ;
  assign n12649 = ~n7294 & n12648 ;
  assign n12651 = n12650 ^ n12649 ^ n3053 ;
  assign n12652 = n4129 & ~n8307 ;
  assign n12653 = n6946 | n8081 ;
  assign n12654 = n12653 ^ n5308 ^ 1'b0 ;
  assign n12655 = n3271 & n8641 ;
  assign n12656 = ~n4719 & n12655 ;
  assign n12657 = n12656 ^ n9254 ^ 1'b0 ;
  assign n12658 = n1359 | n12657 ;
  assign n12659 = ( ~n6243 & n12654 ) | ( ~n6243 & n12658 ) | ( n12654 & n12658 ) ;
  assign n12660 = n12652 & ~n12659 ;
  assign n12661 = n12660 ^ n9194 ^ n6818 ;
  assign n12662 = n9193 ^ n8697 ^ n2999 ;
  assign n12663 = n12662 ^ n6481 ^ n847 ;
  assign n12664 = n6324 ^ n6165 ^ 1'b0 ;
  assign n12665 = ~n12663 & n12664 ;
  assign n12666 = n9001 ^ n4470 ^ n3654 ;
  assign n12667 = n7746 ^ n439 ^ 1'b0 ;
  assign n12668 = n12666 & n12667 ;
  assign n12669 = ( ~n1749 & n3750 ) | ( ~n1749 & n12438 ) | ( n3750 & n12438 ) ;
  assign n12670 = n4622 & ~n11115 ;
  assign n12671 = n12670 ^ n12411 ^ n9066 ;
  assign n12672 = n9865 ^ n2479 ^ n2313 ;
  assign n12673 = ( n4562 & n6881 ) | ( n4562 & n9502 ) | ( n6881 & n9502 ) ;
  assign n12679 = ( n2809 & ~n3748 ) | ( n2809 & n5954 ) | ( ~n3748 & n5954 ) ;
  assign n12674 = n9728 ^ n4477 ^ n2819 ;
  assign n12675 = n10087 & n12674 ;
  assign n12676 = ( n2863 & n4651 ) | ( n2863 & ~n12675 ) | ( n4651 & ~n12675 ) ;
  assign n12677 = ~n6442 & n12676 ;
  assign n12678 = n12677 ^ n3006 ^ 1'b0 ;
  assign n12680 = n12679 ^ n12678 ^ 1'b0 ;
  assign n12681 = n5767 ^ n3761 ^ n1798 ;
  assign n12682 = n2311 ^ n1104 ^ 1'b0 ;
  assign n12683 = n5697 & ~n12682 ;
  assign n12684 = n12683 ^ x72 ^ 1'b0 ;
  assign n12685 = n8648 ^ n2292 ^ n1007 ;
  assign n12686 = n11611 ^ n6971 ^ n1152 ;
  assign n12687 = n12686 ^ n4729 ^ 1'b0 ;
  assign n12688 = n8256 | n12687 ;
  assign n12689 = n8104 ^ n1000 ^ 1'b0 ;
  assign n12691 = n10793 ^ n8853 ^ 1'b0 ;
  assign n12692 = n9534 & ~n12691 ;
  assign n12693 = n12692 ^ n715 ^ 1'b0 ;
  assign n12694 = n12693 ^ n1915 ^ 1'b0 ;
  assign n12690 = ( n928 & n3828 ) | ( n928 & ~n3986 ) | ( n3828 & ~n3986 ) ;
  assign n12695 = n12694 ^ n12690 ^ 1'b0 ;
  assign n12696 = n12307 ^ n11640 ^ x39 ;
  assign n12697 = n8286 ^ n6414 ^ x64 ;
  assign n12698 = n12697 ^ n4833 ^ 1'b0 ;
  assign n12699 = n2645 & n12698 ;
  assign n12700 = n2215 ^ n480 ^ x62 ;
  assign n12701 = n2389 ^ n141 ^ 1'b0 ;
  assign n12702 = ~n8047 & n12701 ;
  assign n12703 = n12702 ^ n9723 ^ n188 ;
  assign n12704 = n12703 ^ n4162 ^ 1'b0 ;
  assign n12705 = ~n3132 & n12704 ;
  assign n12706 = n8881 ^ n2212 ^ 1'b0 ;
  assign n12707 = n2200 & ~n12706 ;
  assign n12709 = ~n3641 & n8207 ;
  assign n12710 = n12709 ^ n5451 ^ 1'b0 ;
  assign n12711 = n12710 ^ n1501 ^ 1'b0 ;
  assign n12708 = n5697 ^ n3250 ^ 1'b0 ;
  assign n12712 = n12711 ^ n12708 ^ 1'b0 ;
  assign n12713 = ( ~n12705 & n12707 ) | ( ~n12705 & n12712 ) | ( n12707 & n12712 ) ;
  assign n12714 = n12700 & ~n12713 ;
  assign n12715 = ~n12699 & n12714 ;
  assign n12716 = ( n3989 & ~n8181 ) | ( n3989 & n8885 ) | ( ~n8181 & n8885 ) ;
  assign n12731 = n5327 & ~n11499 ;
  assign n12732 = n12731 ^ n3300 ^ 1'b0 ;
  assign n12733 = n12732 ^ n8480 ^ n3935 ;
  assign n12728 = n325 & ~n3336 ;
  assign n12729 = n12728 ^ n6651 ^ 1'b0 ;
  assign n12727 = n10244 ^ n5367 ^ 1'b0 ;
  assign n12730 = n12729 ^ n12727 ^ n2574 ;
  assign n12734 = n12733 ^ n12730 ^ n6042 ;
  assign n12735 = n12734 ^ n5316 ^ n1665 ;
  assign n12723 = n6860 ^ n1775 ^ n1376 ;
  assign n12724 = n7792 ^ n5371 ^ 1'b0 ;
  assign n12725 = n12724 ^ n5213 ^ n4400 ;
  assign n12726 = ( n500 & ~n12723 ) | ( n500 & n12725 ) | ( ~n12723 & n12725 ) ;
  assign n12717 = n7841 ^ n3635 ^ n284 ;
  assign n12718 = n12717 ^ n400 ^ 1'b0 ;
  assign n12719 = n1692 | n12718 ;
  assign n12720 = n2725 & ~n8534 ;
  assign n12721 = n12719 & n12720 ;
  assign n12722 = n12721 ^ n11868 ^ n11564 ;
  assign n12736 = n12735 ^ n12726 ^ n12722 ;
  assign n12737 = ( x8 & x111 ) | ( x8 & ~n200 ) | ( x111 & ~n200 ) ;
  assign n12743 = n4532 ^ n3831 ^ n759 ;
  assign n12744 = n8365 & n12743 ;
  assign n12739 = x112 & ~n1114 ;
  assign n12740 = ~n2065 & n12739 ;
  assign n12741 = ( ~n424 & n5337 ) | ( ~n424 & n7105 ) | ( n5337 & n7105 ) ;
  assign n12742 = ( n10127 & ~n12740 ) | ( n10127 & n12741 ) | ( ~n12740 & n12741 ) ;
  assign n12738 = ( n5052 & n8475 ) | ( n5052 & ~n12215 ) | ( n8475 & ~n12215 ) ;
  assign n12745 = n12744 ^ n12742 ^ n12738 ;
  assign n12746 = ~n6444 & n12745 ;
  assign n12747 = ~n12737 & n12746 ;
  assign n12748 = n3188 ^ n2943 ^ n2450 ;
  assign n12749 = n12748 ^ n10006 ^ n1384 ;
  assign n12750 = ( n3899 & n8077 ) | ( n3899 & ~n8534 ) | ( n8077 & ~n8534 ) ;
  assign n12751 = ( n369 & n5426 ) | ( n369 & ~n12750 ) | ( n5426 & ~n12750 ) ;
  assign n12752 = ( ~n3256 & n4868 ) | ( ~n3256 & n5266 ) | ( n4868 & n5266 ) ;
  assign n12753 = ~n870 & n12752 ;
  assign n12754 = n3279 ^ n1229 ^ n647 ;
  assign n12755 = n11139 ^ n10524 ^ n7338 ;
  assign n12756 = ( n8819 & ~n12754 ) | ( n8819 & n12755 ) | ( ~n12754 & n12755 ) ;
  assign n12757 = ~n12753 & n12756 ;
  assign n12758 = n12757 ^ n3831 ^ n2257 ;
  assign n12759 = ( n5684 & n8048 ) | ( n5684 & ~n10123 ) | ( n8048 & ~n10123 ) ;
  assign n12760 = n11074 ^ n6539 ^ n863 ;
  assign n12761 = ( n4634 & n12759 ) | ( n4634 & n12760 ) | ( n12759 & n12760 ) ;
  assign n12762 = ( n2486 & n3316 ) | ( n2486 & n5038 ) | ( n3316 & n5038 ) ;
  assign n12763 = n12181 ^ n8335 ^ n3606 ;
  assign n12764 = n12763 ^ n2812 ^ n218 ;
  assign n12765 = ( n1403 & ~n12762 ) | ( n1403 & n12764 ) | ( ~n12762 & n12764 ) ;
  assign n12766 = n9886 ^ x24 ^ 1'b0 ;
  assign n12767 = n3219 & n12766 ;
  assign n12768 = n6520 ^ n1971 ^ 1'b0 ;
  assign n12769 = n8623 | n8769 ;
  assign n12770 = n3736 & ~n12769 ;
  assign n12771 = n12770 ^ n5416 ^ 1'b0 ;
  assign n12772 = n12768 & n12771 ;
  assign n12773 = ~n11219 & n12772 ;
  assign n12774 = n9556 ^ n2581 ^ 1'b0 ;
  assign n12775 = ~n5424 & n12774 ;
  assign n12776 = n10161 ^ n9231 ^ n4421 ;
  assign n12777 = n1253 & ~n1350 ;
  assign n12778 = n1776 & n12777 ;
  assign n12779 = n12778 ^ n2101 ^ 1'b0 ;
  assign n12780 = n2191 | n11752 ;
  assign n12781 = n12780 ^ n3151 ^ 1'b0 ;
  assign n12782 = n9688 & ~n12781 ;
  assign n12787 = n1411 & n2788 ;
  assign n12785 = n7077 ^ n6953 ^ 1'b0 ;
  assign n12786 = n1913 & n12785 ;
  assign n12788 = n12787 ^ n12786 ^ n2218 ;
  assign n12783 = n11961 ^ n9220 ^ n6707 ;
  assign n12784 = ( ~n940 & n5993 ) | ( ~n940 & n12783 ) | ( n5993 & n12783 ) ;
  assign n12789 = n12788 ^ n12784 ^ n4011 ;
  assign n12790 = ( x6 & n5784 ) | ( x6 & n10714 ) | ( n5784 & n10714 ) ;
  assign n12791 = n3698 & n8696 ;
  assign n12792 = ~n4404 & n12791 ;
  assign n12793 = ( n1996 & n5947 ) | ( n1996 & ~n12792 ) | ( n5947 & ~n12792 ) ;
  assign n12796 = ( n408 & n4541 ) | ( n408 & n5919 ) | ( n4541 & n5919 ) ;
  assign n12797 = n12796 ^ n11852 ^ n5125 ;
  assign n12798 = n12797 ^ n4380 ^ n3979 ;
  assign n12799 = n6318 | n12798 ;
  assign n12800 = n3243 | n12799 ;
  assign n12794 = n10275 ^ n7435 ^ 1'b0 ;
  assign n12795 = n3159 | n12794 ;
  assign n12801 = n12800 ^ n12795 ^ n2401 ;
  assign n12802 = ( n7084 & ~n12793 ) | ( n7084 & n12801 ) | ( ~n12793 & n12801 ) ;
  assign n12803 = n10773 & n12802 ;
  assign n12804 = n1583 & n12803 ;
  assign n12805 = n3831 ^ n2860 ^ 1'b0 ;
  assign n12806 = n6802 & ~n12805 ;
  assign n12807 = n12806 ^ n243 ^ 1'b0 ;
  assign n12808 = ~n8490 & n12692 ;
  assign n12809 = n12808 ^ n5701 ^ 1'b0 ;
  assign n12810 = n1117 & n12809 ;
  assign n12811 = n12810 ^ n7392 ^ 1'b0 ;
  assign n12812 = n9451 ^ n9175 ^ n6203 ;
  assign n12813 = ( n3309 & n12811 ) | ( n3309 & ~n12812 ) | ( n12811 & ~n12812 ) ;
  assign n12814 = ( n4289 & ~n7125 ) | ( n4289 & n8632 ) | ( ~n7125 & n8632 ) ;
  assign n12818 = ( ~n2305 & n3131 ) | ( ~n2305 & n4062 ) | ( n3131 & n4062 ) ;
  assign n12819 = n11040 & ~n12818 ;
  assign n12820 = n12819 ^ n6951 ^ 1'b0 ;
  assign n12821 = ( n1630 & ~n4475 ) | ( n1630 & n12820 ) | ( ~n4475 & n12820 ) ;
  assign n12815 = n1483 & ~n4455 ;
  assign n12816 = ~n3244 & n12815 ;
  assign n12817 = n12816 ^ n6751 ^ n5248 ;
  assign n12822 = n12821 ^ n12817 ^ n676 ;
  assign n12823 = n6034 ^ n568 ^ 1'b0 ;
  assign n12824 = n7572 ^ n920 ^ n798 ;
  assign n12827 = n7369 ^ n1206 ^ 1'b0 ;
  assign n12828 = n11210 & n12827 ;
  assign n12829 = n4976 & n12828 ;
  assign n12826 = ~n295 & n4307 ;
  assign n12830 = n12829 ^ n12826 ^ 1'b0 ;
  assign n12825 = n11916 ^ n5078 ^ n256 ;
  assign n12831 = n12830 ^ n12825 ^ 1'b0 ;
  assign n12832 = ( n3276 & n5050 ) | ( n3276 & n6660 ) | ( n5050 & n6660 ) ;
  assign n12833 = n5545 & n12722 ;
  assign n12834 = n6077 & ~n7148 ;
  assign n12835 = n10056 ^ n6013 ^ n3997 ;
  assign n12836 = ( n1551 & ~n12834 ) | ( n1551 & n12835 ) | ( ~n12834 & n12835 ) ;
  assign n12837 = n7527 ^ n1971 ^ 1'b0 ;
  assign n12838 = ~n7982 & n12837 ;
  assign n12842 = n9863 ^ n8828 ^ 1'b0 ;
  assign n12843 = ( n1442 & n11916 ) | ( n1442 & ~n12842 ) | ( n11916 & ~n12842 ) ;
  assign n12844 = ( ~n7511 & n10196 ) | ( ~n7511 & n12843 ) | ( n10196 & n12843 ) ;
  assign n12839 = n2483 & ~n4114 ;
  assign n12840 = n12839 ^ n3892 ^ 1'b0 ;
  assign n12841 = n12840 ^ n9565 ^ n5053 ;
  assign n12845 = n12844 ^ n12841 ^ n1861 ;
  assign n12846 = n12845 ^ n9048 ^ n2043 ;
  assign n12847 = ( ~n3885 & n7515 ) | ( ~n3885 & n8947 ) | ( n7515 & n8947 ) ;
  assign n12848 = n7759 ^ n4557 ^ 1'b0 ;
  assign n12849 = n3234 ^ n941 ^ 1'b0 ;
  assign n12850 = n205 & ~n12849 ;
  assign n12851 = n11369 ^ n2388 ^ n2022 ;
  assign n12852 = n8869 ^ n7339 ^ n1778 ;
  assign n12853 = n1619 | n5084 ;
  assign n12854 = ( ~n586 & n12852 ) | ( ~n586 & n12853 ) | ( n12852 & n12853 ) ;
  assign n12855 = ( n3093 & n7343 ) | ( n3093 & ~n12174 ) | ( n7343 & ~n12174 ) ;
  assign n12856 = ( n12851 & n12854 ) | ( n12851 & n12855 ) | ( n12854 & n12855 ) ;
  assign n12857 = n12856 ^ n9473 ^ 1'b0 ;
  assign n12858 = n1463 & n12857 ;
  assign n12859 = n5800 | n6107 ;
  assign n12860 = n2948 & ~n12859 ;
  assign n12861 = x48 & n2417 ;
  assign n12862 = n12860 & n12861 ;
  assign n12863 = n12862 ^ n10116 ^ n1409 ;
  assign n12864 = ~n2081 & n3321 ;
  assign n12865 = ( ~n1078 & n7696 ) | ( ~n1078 & n12864 ) | ( n7696 & n12864 ) ;
  assign n12866 = n12565 ^ n4044 ^ x100 ;
  assign n12868 = n2880 & n10115 ;
  assign n12869 = n12868 ^ n2617 ^ 1'b0 ;
  assign n12867 = n4646 ^ n3854 ^ n3044 ;
  assign n12870 = n12869 ^ n12867 ^ x8 ;
  assign n12871 = n12870 ^ n3935 ^ 1'b0 ;
  assign n12872 = n11258 ^ n8289 ^ n7862 ;
  assign n12873 = n12872 ^ n12332 ^ n4442 ;
  assign n12874 = n12873 ^ n7705 ^ n5433 ;
  assign n12875 = n1917 ^ n1114 ^ 1'b0 ;
  assign n12877 = ( n2825 & ~n3164 ) | ( n2825 & n11669 ) | ( ~n3164 & n11669 ) ;
  assign n12878 = ~n6590 & n12877 ;
  assign n12876 = ~n1996 & n4856 ;
  assign n12879 = n12878 ^ n12876 ^ n1617 ;
  assign n12885 = n9400 ^ n2550 ^ n2409 ;
  assign n12880 = n2480 ^ n1953 ^ n418 ;
  assign n12881 = n1062 ^ n456 ^ x98 ;
  assign n12882 = n12881 ^ n2145 ^ 1'b0 ;
  assign n12883 = n8541 & n12882 ;
  assign n12884 = ( ~n2736 & n12880 ) | ( ~n2736 & n12883 ) | ( n12880 & n12883 ) ;
  assign n12886 = n12885 ^ n12884 ^ n10071 ;
  assign n12887 = ~n1436 & n11780 ;
  assign n12888 = n12887 ^ n7322 ^ 1'b0 ;
  assign n12889 = n6407 ^ n5135 ^ 1'b0 ;
  assign n12890 = n12889 ^ n7853 ^ n697 ;
  assign n12891 = n3024 & ~n11212 ;
  assign n12896 = ( n924 & ~n1637 ) | ( n924 & n3438 ) | ( ~n1637 & n3438 ) ;
  assign n12892 = n4862 ^ n1784 ^ x94 ;
  assign n12893 = ~n3764 & n10651 ;
  assign n12894 = n4356 & n12893 ;
  assign n12895 = ( n11498 & n12892 ) | ( n11498 & ~n12894 ) | ( n12892 & ~n12894 ) ;
  assign n12897 = n12896 ^ n12895 ^ n1110 ;
  assign n12900 = n10312 ^ n9156 ^ n4144 ;
  assign n12901 = n12900 ^ n10926 ^ 1'b0 ;
  assign n12898 = ( ~n3857 & n3929 ) | ( ~n3857 & n5259 ) | ( n3929 & n5259 ) ;
  assign n12899 = n12898 ^ n8974 ^ n8043 ;
  assign n12902 = n12901 ^ n12899 ^ n2850 ;
  assign n12903 = n4381 ^ n3516 ^ n1500 ;
  assign n12904 = n7669 ^ n3239 ^ n1106 ;
  assign n12905 = ( n3474 & n12903 ) | ( n3474 & ~n12904 ) | ( n12903 & ~n12904 ) ;
  assign n12906 = n12905 ^ n12419 ^ n4015 ;
  assign n12907 = n12906 ^ n7962 ^ n5817 ;
  assign n12908 = n2315 & n12256 ;
  assign n12909 = n12908 ^ n6826 ^ 1'b0 ;
  assign n12910 = n12829 ^ n11311 ^ n1409 ;
  assign n12911 = n8602 ^ n2073 ^ n1813 ;
  assign n12912 = ( n6275 & n12910 ) | ( n6275 & ~n12911 ) | ( n12910 & ~n12911 ) ;
  assign n12913 = ( n2573 & n6995 ) | ( n2573 & ~n8454 ) | ( n6995 & ~n8454 ) ;
  assign n12914 = ( n5957 & n10384 ) | ( n5957 & n12913 ) | ( n10384 & n12913 ) ;
  assign n12915 = ( ~n12909 & n12912 ) | ( ~n12909 & n12914 ) | ( n12912 & n12914 ) ;
  assign n12916 = n10947 & ~n10968 ;
  assign n12917 = n12916 ^ n10157 ^ 1'b0 ;
  assign n12918 = ( ~n4344 & n5400 ) | ( ~n4344 & n9622 ) | ( n5400 & n9622 ) ;
  assign n12919 = ( ~n2465 & n4263 ) | ( ~n2465 & n12918 ) | ( n4263 & n12918 ) ;
  assign n12922 = n3588 ^ n1652 ^ n1475 ;
  assign n12920 = n7545 ^ n5999 ^ 1'b0 ;
  assign n12921 = n3651 & ~n12920 ;
  assign n12923 = n12922 ^ n12921 ^ n3292 ;
  assign n12924 = n8494 & n9508 ;
  assign n12925 = n12923 & n12924 ;
  assign n12926 = n6873 ^ n2441 ^ n642 ;
  assign n12927 = n2921 ^ n2644 ^ n568 ;
  assign n12928 = ( n1460 & ~n1763 ) | ( n1460 & n12927 ) | ( ~n1763 & n12927 ) ;
  assign n12929 = n12926 | n12928 ;
  assign n12930 = n12929 ^ n1220 ^ 1'b0 ;
  assign n12931 = ( n898 & ~n5031 ) | ( n898 & n11978 ) | ( ~n5031 & n11978 ) ;
  assign n12932 = ( n182 & n251 ) | ( n182 & ~n867 ) | ( n251 & ~n867 ) ;
  assign n12933 = ~n7141 & n12932 ;
  assign n12934 = ~n12931 & n12933 ;
  assign n12935 = ( n1694 & n4058 ) | ( n1694 & ~n4359 ) | ( n4058 & ~n4359 ) ;
  assign n12936 = n9729 | n11179 ;
  assign n12937 = n7275 & ~n12936 ;
  assign n12938 = ( n1347 & n12935 ) | ( n1347 & n12937 ) | ( n12935 & n12937 ) ;
  assign n12939 = ( n6808 & ~n8277 ) | ( n6808 & n12938 ) | ( ~n8277 & n12938 ) ;
  assign n12940 = n3271 & ~n7268 ;
  assign n12941 = n12940 ^ n9070 ^ 1'b0 ;
  assign n12942 = ~n8752 & n9542 ;
  assign n12943 = n12942 ^ n8450 ^ 1'b0 ;
  assign n12944 = ( n1880 & n4159 ) | ( n1880 & ~n5333 ) | ( n4159 & ~n5333 ) ;
  assign n12945 = n4072 & ~n12944 ;
  assign n12946 = ( n6449 & ~n9104 ) | ( n6449 & n12945 ) | ( ~n9104 & n12945 ) ;
  assign n12947 = ( ~n1620 & n4332 ) | ( ~n1620 & n11651 ) | ( n4332 & n11651 ) ;
  assign n12948 = n11960 ^ n4412 ^ n1888 ;
  assign n12949 = n12948 ^ n7058 ^ n1312 ;
  assign n12950 = ( n2058 & n6425 ) | ( n2058 & n12949 ) | ( n6425 & n12949 ) ;
  assign n12951 = ( n7520 & n11780 ) | ( n7520 & ~n12950 ) | ( n11780 & ~n12950 ) ;
  assign n12952 = n8298 ^ n8254 ^ n7049 ;
  assign n12953 = n11701 ^ n1785 ^ n973 ;
  assign n12954 = n8530 ^ n5406 ^ n2526 ;
  assign n12955 = n9734 ^ n8103 ^ 1'b0 ;
  assign n12956 = n12954 & ~n12955 ;
  assign n12960 = n7426 ^ n6361 ^ n5525 ;
  assign n12961 = ( ~n2355 & n2656 ) | ( ~n2355 & n12960 ) | ( n2656 & n12960 ) ;
  assign n12957 = ( n4318 & n4574 ) | ( n4318 & ~n7457 ) | ( n4574 & ~n7457 ) ;
  assign n12958 = n6692 ^ n4422 ^ n2705 ;
  assign n12959 = ( n11134 & n12957 ) | ( n11134 & ~n12958 ) | ( n12957 & ~n12958 ) ;
  assign n12962 = n12961 ^ n12959 ^ n7575 ;
  assign n12963 = ( n485 & n3087 ) | ( n485 & ~n9029 ) | ( n3087 & ~n9029 ) ;
  assign n12964 = ( n3074 & ~n11490 ) | ( n3074 & n12963 ) | ( ~n11490 & n12963 ) ;
  assign n12965 = n7063 ^ n4264 ^ 1'b0 ;
  assign n12970 = n3185 | n5892 ;
  assign n12971 = n12970 ^ n7791 ^ 1'b0 ;
  assign n12966 = n10244 ^ n9138 ^ x86 ;
  assign n12967 = n12966 ^ n4970 ^ n2009 ;
  assign n12968 = n12967 ^ n6322 ^ n146 ;
  assign n12969 = ( ~n379 & n1552 ) | ( ~n379 & n12968 ) | ( n1552 & n12968 ) ;
  assign n12972 = n12971 ^ n12969 ^ 1'b0 ;
  assign n12973 = n10938 ^ n6970 ^ n2459 ;
  assign n12975 = ( n347 & n8136 ) | ( n347 & n8218 ) | ( n8136 & n8218 ) ;
  assign n12974 = n2250 | n3757 ;
  assign n12976 = n12975 ^ n12974 ^ 1'b0 ;
  assign n12977 = ( n10636 & n12973 ) | ( n10636 & n12976 ) | ( n12973 & n12976 ) ;
  assign n12978 = n6565 ^ n4480 ^ 1'b0 ;
  assign n12979 = ( n7040 & n7419 ) | ( n7040 & n12978 ) | ( n7419 & n12978 ) ;
  assign n12980 = n4227 ^ n1361 ^ x51 ;
  assign n12981 = n6671 | n12980 ;
  assign n12982 = ( n8048 & n12979 ) | ( n8048 & ~n12981 ) | ( n12979 & ~n12981 ) ;
  assign n12983 = ( n5956 & ~n8704 ) | ( n5956 & n9206 ) | ( ~n8704 & n9206 ) ;
  assign n12984 = n11383 ^ n708 ^ 1'b0 ;
  assign n12985 = ~n4086 & n8080 ;
  assign n12986 = n6143 & ~n10253 ;
  assign n12987 = n359 & ~n11041 ;
  assign n12988 = n12760 ^ n12457 ^ n4374 ;
  assign n12989 = n3127 & n6023 ;
  assign n12990 = n4396 & n12989 ;
  assign n12991 = n12990 ^ n5873 ^ 1'b0 ;
  assign n12992 = n8202 & n12991 ;
  assign n12999 = ( n547 & ~n11185 ) | ( n547 & n11246 ) | ( ~n11185 & n11246 ) ;
  assign n13000 = n7148 ^ n353 ^ 1'b0 ;
  assign n13001 = n12999 & ~n13000 ;
  assign n12996 = ( x33 & x50 ) | ( x33 & n366 ) | ( x50 & n366 ) ;
  assign n12994 = n509 & n10325 ;
  assign n12995 = n12994 ^ n2364 ^ n409 ;
  assign n12993 = n3288 & ~n5474 ;
  assign n12997 = n12996 ^ n12995 ^ n12993 ;
  assign n12998 = n12997 ^ n1746 ^ 1'b0 ;
  assign n13002 = n13001 ^ n12998 ^ n1176 ;
  assign n13003 = ( n2677 & n7350 ) | ( n2677 & ~n11991 ) | ( n7350 & ~n11991 ) ;
  assign n13004 = n4575 | n11580 ;
  assign n13005 = n7908 ^ n1475 ^ 1'b0 ;
  assign n13006 = n5886 | n13005 ;
  assign n13007 = n9129 | n13006 ;
  assign n13008 = n13007 ^ n5254 ^ 1'b0 ;
  assign n13009 = n589 | n13008 ;
  assign n13010 = n7340 | n13009 ;
  assign n13011 = n3442 ^ n1748 ^ 1'b0 ;
  assign n13012 = ( n2205 & n8650 ) | ( n2205 & n13011 ) | ( n8650 & n13011 ) ;
  assign n13013 = n3950 | n6745 ;
  assign n13014 = n1309 | n13013 ;
  assign n13015 = n9421 ^ n4973 ^ 1'b0 ;
  assign n13016 = n13014 & ~n13015 ;
  assign n13017 = n13012 | n13016 ;
  assign n13018 = n5659 ^ n2935 ^ 1'b0 ;
  assign n13019 = n1712 | n13018 ;
  assign n13020 = ( n3438 & n7375 ) | ( n3438 & ~n13019 ) | ( n7375 & ~n13019 ) ;
  assign n13021 = ~n1605 & n11463 ;
  assign n13022 = ( n4025 & n10590 ) | ( n4025 & n13021 ) | ( n10590 & n13021 ) ;
  assign n13023 = n1781 & ~n10973 ;
  assign n13024 = n9771 & n13023 ;
  assign n13025 = ~n13022 & n13024 ;
  assign n13026 = n9175 ^ n4013 ^ 1'b0 ;
  assign n13027 = n5384 & ~n13026 ;
  assign n13028 = ( n718 & n2328 ) | ( n718 & n7844 ) | ( n2328 & n7844 ) ;
  assign n13029 = ( n8990 & n13027 ) | ( n8990 & ~n13028 ) | ( n13027 & ~n13028 ) ;
  assign n13030 = n2303 | n6150 ;
  assign n13031 = n6905 & ~n13030 ;
  assign n13032 = n3657 ^ n1696 ^ 1'b0 ;
  assign n13033 = n13031 | n13032 ;
  assign n13034 = n1255 & n10732 ;
  assign n13041 = n315 | n4897 ;
  assign n13042 = n13041 ^ n4190 ^ 1'b0 ;
  assign n13043 = n3728 & ~n7950 ;
  assign n13044 = ~n2363 & n13043 ;
  assign n13045 = ~n13042 & n13044 ;
  assign n13035 = n8478 ^ n8282 ^ n5448 ;
  assign n13036 = ( n2844 & n3950 ) | ( n2844 & n8340 ) | ( n3950 & n8340 ) ;
  assign n13037 = n13036 ^ n3516 ^ n1218 ;
  assign n13038 = n13037 ^ n4944 ^ n3795 ;
  assign n13039 = ~n13035 & n13038 ;
  assign n13040 = n13039 ^ n2612 ^ 1'b0 ;
  assign n13046 = n13045 ^ n13040 ^ n1535 ;
  assign n13047 = ~n13034 & n13046 ;
  assign n13048 = n13047 ^ n4888 ^ 1'b0 ;
  assign n13050 = n2360 | n3131 ;
  assign n13051 = n13050 ^ n1623 ^ 1'b0 ;
  assign n13052 = ( n4589 & n5813 ) | ( n4589 & ~n13051 ) | ( n5813 & ~n13051 ) ;
  assign n13049 = n5696 | n11405 ;
  assign n13053 = n13052 ^ n13049 ^ n4353 ;
  assign n13054 = n13053 ^ n2931 ^ n2292 ;
  assign n13060 = n4819 ^ n4153 ^ n1482 ;
  assign n13059 = n681 | n2032 ;
  assign n13061 = n13060 ^ n13059 ^ 1'b0 ;
  assign n13062 = n3330 | n6146 ;
  assign n13063 = n13061 & ~n13062 ;
  assign n13056 = n3603 ^ n2393 ^ n1366 ;
  assign n13055 = n813 & n4752 ;
  assign n13057 = n13056 ^ n13055 ^ 1'b0 ;
  assign n13058 = n13057 ^ n9246 ^ n6917 ;
  assign n13064 = n13063 ^ n13058 ^ 1'b0 ;
  assign n13065 = n13054 & n13064 ;
  assign n13066 = n12944 ^ n9641 ^ n2801 ;
  assign n13067 = n4223 ^ n1867 ^ 1'b0 ;
  assign n13068 = n13066 | n13067 ;
  assign n13069 = n4785 | n11701 ;
  assign n13070 = n13068 & ~n13069 ;
  assign n13071 = n4302 ^ n4101 ^ n1297 ;
  assign n13072 = n4650 ^ n2480 ^ 1'b0 ;
  assign n13073 = ( n508 & n9050 ) | ( n508 & ~n13072 ) | ( n9050 & ~n13072 ) ;
  assign n13074 = ( n7914 & n11334 ) | ( n7914 & ~n13073 ) | ( n11334 & ~n13073 ) ;
  assign n13075 = n6343 ^ n5578 ^ n1533 ;
  assign n13076 = n10207 ^ n6591 ^ n1148 ;
  assign n13077 = n5783 ^ n1574 ^ 1'b0 ;
  assign n13078 = n13077 ^ n6732 ^ 1'b0 ;
  assign n13079 = ( n12690 & n13076 ) | ( n12690 & n13078 ) | ( n13076 & n13078 ) ;
  assign n13080 = ( n2219 & n4732 ) | ( n2219 & n13079 ) | ( n4732 & n13079 ) ;
  assign n13081 = n594 & n3702 ;
  assign n13082 = ~n13080 & n13081 ;
  assign n13083 = n7869 ^ n6240 ^ n572 ;
  assign n13084 = ~n1715 & n8429 ;
  assign n13085 = n13084 ^ x121 ^ 1'b0 ;
  assign n13086 = n11487 ^ n11118 ^ 1'b0 ;
  assign n13087 = x23 & ~n1962 ;
  assign n13088 = n5172 & n13087 ;
  assign n13089 = ( ~n2888 & n10471 ) | ( ~n2888 & n13088 ) | ( n10471 & n13088 ) ;
  assign n13090 = n13089 ^ n9207 ^ 1'b0 ;
  assign n13091 = n6071 ^ n3421 ^ n3129 ;
  assign n13092 = n9727 | n13091 ;
  assign n13093 = n4494 | n13092 ;
  assign n13094 = ( n3254 & n13090 ) | ( n3254 & n13093 ) | ( n13090 & n13093 ) ;
  assign n13095 = n5773 & ~n13094 ;
  assign n13096 = n5730 ^ n3229 ^ n490 ;
  assign n13097 = n11540 ^ n8540 ^ 1'b0 ;
  assign n13098 = n12384 | n13097 ;
  assign n13099 = n7744 | n13098 ;
  assign n13100 = n13099 ^ n8306 ^ 1'b0 ;
  assign n13101 = n13100 ^ n11182 ^ n11044 ;
  assign n13103 = n6347 ^ n1038 ^ 1'b0 ;
  assign n13102 = ( n2232 & ~n3324 ) | ( n2232 & n4375 ) | ( ~n3324 & n4375 ) ;
  assign n13104 = n13103 ^ n13102 ^ n9706 ;
  assign n13105 = ( n1062 & n1163 ) | ( n1062 & ~n12001 ) | ( n1163 & ~n12001 ) ;
  assign n13106 = n4175 ^ n2326 ^ n822 ;
  assign n13107 = ~n6867 & n13106 ;
  assign n13111 = n4941 ^ n3311 ^ 1'b0 ;
  assign n13112 = n13111 ^ n5292 ^ n3343 ;
  assign n13108 = n794 & n2565 ;
  assign n13109 = n13108 ^ n5066 ^ 1'b0 ;
  assign n13110 = ~n12416 & n13109 ;
  assign n13113 = n13112 ^ n13110 ^ 1'b0 ;
  assign n13114 = n12035 ^ n6910 ^ n3563 ;
  assign n13115 = n13114 ^ n4470 ^ 1'b0 ;
  assign n13116 = n10228 ^ n2411 ^ 1'b0 ;
  assign n13117 = ( x118 & n212 ) | ( x118 & ~n13116 ) | ( n212 & ~n13116 ) ;
  assign n13118 = ~n5405 & n8949 ;
  assign n13119 = n13118 ^ n3550 ^ 1'b0 ;
  assign n13120 = ( n12132 & ~n12222 ) | ( n12132 & n13119 ) | ( ~n12222 & n13119 ) ;
  assign n13133 = n2238 & ~n6466 ;
  assign n13134 = n13133 ^ n8748 ^ n3035 ;
  assign n13129 = n1849 & n1861 ;
  assign n13130 = n12372 ^ n7601 ^ n3375 ;
  assign n13131 = ~n13129 & n13130 ;
  assign n13132 = ~n1834 & n13131 ;
  assign n13135 = n13134 ^ n13132 ^ n10161 ;
  assign n13136 = n13135 ^ n1862 ^ 1'b0 ;
  assign n13121 = ~n3641 & n5149 ;
  assign n13122 = ~n9701 & n13121 ;
  assign n13123 = ( n2904 & ~n7743 ) | ( n2904 & n13122 ) | ( ~n7743 & n13122 ) ;
  assign n13124 = ~n7607 & n13123 ;
  assign n13126 = ( ~n3577 & n6364 ) | ( ~n3577 & n6861 ) | ( n6364 & n6861 ) ;
  assign n13125 = n7783 ^ n3509 ^ 1'b0 ;
  assign n13127 = n13126 ^ n13125 ^ n9525 ;
  assign n13128 = n13124 & ~n13127 ;
  assign n13137 = n13136 ^ n13128 ^ 1'b0 ;
  assign n13138 = ~n10862 & n12275 ;
  assign n13139 = n13138 ^ n9911 ^ 1'b0 ;
  assign n13140 = ~n5629 & n11774 ;
  assign n13142 = n11153 ^ n3366 ^ 1'b0 ;
  assign n13143 = n1787 & ~n13142 ;
  assign n13141 = ( ~n4375 & n6471 ) | ( ~n4375 & n9633 ) | ( n6471 & n9633 ) ;
  assign n13144 = n13143 ^ n13141 ^ n11708 ;
  assign n13146 = n1143 & ~n8869 ;
  assign n13147 = n13146 ^ n10079 ^ 1'b0 ;
  assign n13145 = n3392 & n4704 ;
  assign n13148 = n13147 ^ n13145 ^ 1'b0 ;
  assign n13149 = n13148 ^ n9178 ^ n4891 ;
  assign n13153 = n6228 ^ n4944 ^ 1'b0 ;
  assign n13154 = n7246 & ~n13153 ;
  assign n13150 = n12296 ^ n11435 ^ n3467 ;
  assign n13151 = n3233 | n13150 ;
  assign n13152 = n13151 ^ n9207 ^ 1'b0 ;
  assign n13155 = n13154 ^ n13152 ^ 1'b0 ;
  assign n13156 = n9906 ^ n4697 ^ 1'b0 ;
  assign n13157 = n1758 ^ n1032 ^ 1'b0 ;
  assign n13158 = n10720 ^ n2955 ^ 1'b0 ;
  assign n13159 = n10115 & ~n13158 ;
  assign n13160 = ( n7179 & ~n13157 ) | ( n7179 & n13159 ) | ( ~n13157 & n13159 ) ;
  assign n13161 = ( ~n2580 & n8082 ) | ( ~n2580 & n13160 ) | ( n8082 & n13160 ) ;
  assign n13162 = n4061 ^ n334 ^ x2 ;
  assign n13163 = n13162 ^ n8018 ^ n1614 ;
  assign n13164 = n10542 ^ n8697 ^ 1'b0 ;
  assign n13165 = ( n7992 & n13163 ) | ( n7992 & n13164 ) | ( n13163 & n13164 ) ;
  assign n13166 = ( n7651 & n8286 ) | ( n7651 & ~n9611 ) | ( n8286 & ~n9611 ) ;
  assign n13167 = n7040 & n8854 ;
  assign n13168 = ~n5024 & n13167 ;
  assign n13169 = n13166 & ~n13168 ;
  assign n13170 = n13169 ^ n2952 ^ 1'b0 ;
  assign n13171 = n4365 | n6116 ;
  assign n13173 = n4787 ^ n4656 ^ n2294 ;
  assign n13172 = ( n459 & n4930 ) | ( n459 & ~n8231 ) | ( n4930 & ~n8231 ) ;
  assign n13174 = n13173 ^ n13172 ^ n5480 ;
  assign n13175 = n12465 ^ n3275 ^ 1'b0 ;
  assign n13176 = n7414 & ~n13175 ;
  assign n13177 = ( n13171 & n13174 ) | ( n13171 & ~n13176 ) | ( n13174 & ~n13176 ) ;
  assign n13181 = n2605 ^ n378 ^ n141 ;
  assign n13182 = ( n1976 & n6480 ) | ( n1976 & ~n13181 ) | ( n6480 & ~n13181 ) ;
  assign n13178 = n11319 ^ n8886 ^ n3196 ;
  assign n13179 = ( n367 & n2252 ) | ( n367 & n9938 ) | ( n2252 & n9938 ) ;
  assign n13180 = n13178 & ~n13179 ;
  assign n13183 = n13182 ^ n13180 ^ 1'b0 ;
  assign n13184 = n13183 ^ n9115 ^ n3360 ;
  assign n13185 = ( n1236 & n13177 ) | ( n1236 & n13184 ) | ( n13177 & n13184 ) ;
  assign n13186 = n4374 ^ n1583 ^ 1'b0 ;
  assign n13187 = n13186 ^ n10199 ^ 1'b0 ;
  assign n13188 = n178 & n13187 ;
  assign n13189 = n10890 ^ n10257 ^ 1'b0 ;
  assign n13190 = ~n9277 & n13189 ;
  assign n13191 = ( ~n355 & n6838 ) | ( ~n355 & n13190 ) | ( n6838 & n13190 ) ;
  assign n13192 = ( ~n597 & n2164 ) | ( ~n597 & n3214 ) | ( n2164 & n3214 ) ;
  assign n13193 = n6770 & ~n13192 ;
  assign n13194 = n9725 & n13193 ;
  assign n13195 = n13194 ^ n6997 ^ 1'b0 ;
  assign n13196 = n6380 ^ n4435 ^ n1583 ;
  assign n13197 = n8632 ^ n4878 ^ 1'b0 ;
  assign n13198 = n13196 | n13197 ;
  assign n13199 = n13198 ^ n8028 ^ 1'b0 ;
  assign n13200 = n1865 | n13199 ;
  assign n13201 = n6711 ^ n449 ^ 1'b0 ;
  assign n13202 = ~n2851 & n13201 ;
  assign n13204 = n12968 ^ n5632 ^ 1'b0 ;
  assign n13205 = n4384 | n13204 ;
  assign n13203 = ~n5520 & n7858 ;
  assign n13206 = n13205 ^ n13203 ^ 1'b0 ;
  assign n13207 = ( ~n231 & n10334 ) | ( ~n231 & n13206 ) | ( n10334 & n13206 ) ;
  assign n13208 = n3551 ^ n686 ^ 1'b0 ;
  assign n13209 = ~n6594 & n13208 ;
  assign n13210 = n13209 ^ n9869 ^ 1'b0 ;
  assign n13211 = ~n5551 & n5594 ;
  assign n13212 = n13211 ^ n9309 ^ 1'b0 ;
  assign n13214 = n7280 ^ n613 ^ 1'b0 ;
  assign n13213 = n2222 & ~n4128 ;
  assign n13215 = n13214 ^ n13213 ^ 1'b0 ;
  assign n13216 = n13215 ^ n10324 ^ n4813 ;
  assign n13217 = n2274 ^ n1079 ^ 1'b0 ;
  assign n13218 = ( n418 & n3401 ) | ( n418 & ~n5687 ) | ( n3401 & ~n5687 ) ;
  assign n13219 = n13218 ^ n6201 ^ n2191 ;
  assign n13220 = n624 & ~n13219 ;
  assign n13221 = ( n6148 & n13217 ) | ( n6148 & n13220 ) | ( n13217 & n13220 ) ;
  assign n13222 = n9871 ^ n8552 ^ 1'b0 ;
  assign n13223 = n2801 & n13222 ;
  assign n13224 = n8934 ^ n7174 ^ n4931 ;
  assign n13225 = n13224 ^ n11929 ^ n7319 ;
  assign n13226 = n9678 & n13225 ;
  assign n13227 = n13226 ^ n11642 ^ 1'b0 ;
  assign n13228 = ( n5285 & ~n5771 ) | ( n5285 & n10030 ) | ( ~n5771 & n10030 ) ;
  assign n13229 = n13228 ^ n725 ^ 1'b0 ;
  assign n13230 = n9792 ^ n8527 ^ n6927 ;
  assign n13231 = ~n809 & n4218 ;
  assign n13232 = ~n11624 & n13231 ;
  assign n13233 = n13232 ^ n9019 ^ n8729 ;
  assign n13234 = ~n693 & n4058 ;
  assign n13235 = n13234 ^ n3011 ^ 1'b0 ;
  assign n13236 = n2252 | n13235 ;
  assign n13237 = ( n6509 & n10136 ) | ( n6509 & ~n13236 ) | ( n10136 & ~n13236 ) ;
  assign n13238 = n3087 ^ n1989 ^ n1734 ;
  assign n13239 = ( n5075 & n12944 ) | ( n5075 & ~n13238 ) | ( n12944 & ~n13238 ) ;
  assign n13240 = n13239 ^ n1630 ^ n158 ;
  assign n13241 = n13240 ^ n5782 ^ 1'b0 ;
  assign n13242 = ( n1492 & ~n3210 ) | ( n1492 & n6402 ) | ( ~n3210 & n6402 ) ;
  assign n13243 = ( n4169 & n9410 ) | ( n4169 & n11102 ) | ( n9410 & n11102 ) ;
  assign n13244 = n13243 ^ n9657 ^ n3959 ;
  assign n13245 = ( n409 & n13242 ) | ( n409 & ~n13244 ) | ( n13242 & ~n13244 ) ;
  assign n13246 = n9758 ^ n5385 ^ n4681 ;
  assign n13247 = n2181 | n5918 ;
  assign n13248 = n13247 ^ n13006 ^ 1'b0 ;
  assign n13249 = n13248 ^ n12499 ^ n9292 ;
  assign n13250 = ( n3681 & n13246 ) | ( n3681 & ~n13249 ) | ( n13246 & ~n13249 ) ;
  assign n13251 = ( n1567 & ~n4428 ) | ( n1567 & n10665 ) | ( ~n4428 & n10665 ) ;
  assign n13252 = n13251 ^ n861 ^ n828 ;
  assign n13253 = ( n4044 & ~n7415 ) | ( n4044 & n9943 ) | ( ~n7415 & n9943 ) ;
  assign n13262 = n5487 ^ n5114 ^ 1'b0 ;
  assign n13263 = x118 & ~n13262 ;
  assign n13264 = n13263 ^ n12111 ^ n1950 ;
  assign n13258 = n4053 | n4117 ;
  assign n13259 = n7339 | n13258 ;
  assign n13260 = n13259 ^ n2570 ^ 1'b0 ;
  assign n13257 = n6598 ^ n5223 ^ 1'b0 ;
  assign n13261 = n13260 ^ n13257 ^ 1'b0 ;
  assign n13254 = n11394 ^ n4548 ^ 1'b0 ;
  assign n13255 = n13254 ^ n1459 ^ n1264 ;
  assign n13256 = n13255 ^ n9488 ^ n6580 ;
  assign n13265 = n13264 ^ n13261 ^ n13256 ;
  assign n13266 = n10719 ^ n4489 ^ 1'b0 ;
  assign n13267 = n4314 & ~n13266 ;
  assign n13268 = n3707 & n9077 ;
  assign n13269 = n6159 & n6963 ;
  assign n13270 = n6628 & n11296 ;
  assign n13271 = n5400 & ~n7880 ;
  assign n13272 = n6013 | n13271 ;
  assign n13273 = ( n3092 & ~n13270 ) | ( n3092 & n13272 ) | ( ~n13270 & n13272 ) ;
  assign n13274 = n13269 | n13273 ;
  assign n13276 = ( n11206 & n11945 ) | ( n11206 & ~n12885 ) | ( n11945 & ~n12885 ) ;
  assign n13275 = n8989 ^ n4252 ^ n3994 ;
  assign n13277 = n13276 ^ n13275 ^ n6829 ;
  assign n13279 = n6915 ^ n3237 ^ n885 ;
  assign n13278 = n1901 ^ n1479 ^ 1'b0 ;
  assign n13280 = n13279 ^ n13278 ^ n2834 ;
  assign n13281 = n4883 ^ n1141 ^ 1'b0 ;
  assign n13282 = n13273 ^ n10660 ^ 1'b0 ;
  assign n13283 = n4895 | n13282 ;
  assign n13284 = ( n1189 & ~n2683 ) | ( n1189 & n5351 ) | ( ~n2683 & n5351 ) ;
  assign n13285 = n13284 ^ n3444 ^ 1'b0 ;
  assign n13286 = n2650 & n13285 ;
  assign n13287 = ~n8553 & n13286 ;
  assign n13288 = n13287 ^ n5168 ^ 1'b0 ;
  assign n13301 = ~n838 & n3533 ;
  assign n13299 = n9526 ^ n5909 ^ n1545 ;
  assign n13297 = n6720 ^ n2805 ^ n1723 ;
  assign n13298 = n9178 | n13297 ;
  assign n13300 = n13299 ^ n13298 ^ n10206 ;
  assign n13290 = n5193 ^ n4221 ^ n3291 ;
  assign n13291 = n2682 & n13290 ;
  assign n13292 = n13291 ^ n12257 ^ 1'b0 ;
  assign n13289 = ~n3951 & n11653 ;
  assign n13293 = n13292 ^ n13289 ^ 1'b0 ;
  assign n13294 = n2739 ^ n2236 ^ n2070 ;
  assign n13295 = n13294 ^ n10201 ^ n10188 ;
  assign n13296 = n13293 & ~n13295 ;
  assign n13302 = n13301 ^ n13300 ^ n13296 ;
  assign n13303 = n192 & n1312 ;
  assign n13304 = n13303 ^ n11953 ^ 1'b0 ;
  assign n13308 = n4461 ^ n271 ^ 1'b0 ;
  assign n13309 = n6714 | n13308 ;
  assign n13305 = n10324 ^ n7519 ^ n5293 ;
  assign n13306 = ( n9015 & ~n12627 ) | ( n9015 & n13305 ) | ( ~n12627 & n13305 ) ;
  assign n13307 = n13306 ^ n9095 ^ n1948 ;
  assign n13310 = n13309 ^ n13307 ^ n8848 ;
  assign n13313 = n6289 ^ n5973 ^ n648 ;
  assign n13311 = n5873 ^ n994 ^ 1'b0 ;
  assign n13312 = ~n2007 & n13311 ;
  assign n13314 = n13313 ^ n13312 ^ n1442 ;
  assign n13315 = ( n1490 & n1969 ) | ( n1490 & n4581 ) | ( n1969 & n4581 ) ;
  assign n13316 = n10358 | n13315 ;
  assign n13317 = n13316 ^ n1483 ^ 1'b0 ;
  assign n13318 = x83 & ~n2858 ;
  assign n13319 = ~n4970 & n13318 ;
  assign n13320 = ( n3288 & n13317 ) | ( n3288 & n13319 ) | ( n13317 & n13319 ) ;
  assign n13321 = n7890 ^ n4081 ^ 1'b0 ;
  assign n13323 = n9722 ^ n6908 ^ n260 ;
  assign n13322 = x34 & n1743 ;
  assign n13324 = n13323 ^ n13322 ^ 1'b0 ;
  assign n13325 = ~n8577 & n12876 ;
  assign n13326 = ( n2065 & n13324 ) | ( n2065 & ~n13325 ) | ( n13324 & ~n13325 ) ;
  assign n13327 = ( n6661 & n13321 ) | ( n6661 & n13326 ) | ( n13321 & n13326 ) ;
  assign n13328 = ( ~n3279 & n8514 ) | ( ~n3279 & n9011 ) | ( n8514 & n9011 ) ;
  assign n13329 = n3221 & ~n7471 ;
  assign n13330 = ~n2394 & n4762 ;
  assign n13331 = n484 & n13330 ;
  assign n13332 = n13331 ^ n9328 ^ 1'b0 ;
  assign n13335 = n11086 ^ n5897 ^ n394 ;
  assign n13333 = n11061 ^ n3397 ^ n1972 ;
  assign n13334 = ( n1971 & ~n2178 ) | ( n1971 & n13333 ) | ( ~n2178 & n13333 ) ;
  assign n13336 = n13335 ^ n13334 ^ n4534 ;
  assign n13338 = n1314 ^ n976 ^ 1'b0 ;
  assign n13337 = n5222 ^ n2961 ^ n1257 ;
  assign n13339 = n13338 ^ n13337 ^ n1848 ;
  assign n13340 = n10339 ^ n6215 ^ n3792 ;
  assign n13341 = ( n920 & ~n1907 ) | ( n920 & n13340 ) | ( ~n1907 & n13340 ) ;
  assign n13342 = n8984 ^ n8431 ^ n7572 ;
  assign n13343 = n13342 ^ n4272 ^ n545 ;
  assign n13344 = n644 & ~n2912 ;
  assign n13345 = n467 & ~n13344 ;
  assign n13346 = n13345 ^ n7336 ^ n6778 ;
  assign n13347 = n1793 ^ n651 ^ 1'b0 ;
  assign n13348 = n3751 & ~n13347 ;
  assign n13349 = n13348 ^ n1017 ^ x19 ;
  assign n13350 = n3999 ^ n1977 ^ 1'b0 ;
  assign n13351 = n13350 ^ n6818 ^ n2419 ;
  assign n13354 = n5686 ^ n1283 ^ n1149 ;
  assign n13355 = ( n703 & n1767 ) | ( n703 & n13354 ) | ( n1767 & n13354 ) ;
  assign n13352 = ( n288 & n1559 ) | ( n288 & ~n5868 ) | ( n1559 & ~n5868 ) ;
  assign n13353 = n3401 & n13352 ;
  assign n13356 = n13355 ^ n13353 ^ 1'b0 ;
  assign n13360 = n8128 | n10122 ;
  assign n13357 = n9129 ^ n8159 ^ n1785 ;
  assign n13358 = n13357 ^ n3078 ^ n1556 ;
  assign n13359 = ( n6304 & ~n8180 ) | ( n6304 & n13358 ) | ( ~n8180 & n13358 ) ;
  assign n13361 = n13360 ^ n13359 ^ n13276 ;
  assign n13362 = n12134 ^ n6711 ^ n1930 ;
  assign n13363 = ( ~n6344 & n13361 ) | ( ~n6344 & n13362 ) | ( n13361 & n13362 ) ;
  assign n13364 = ( n3179 & n4970 ) | ( n3179 & ~n13363 ) | ( n4970 & ~n13363 ) ;
  assign n13365 = ( ~n1524 & n3999 ) | ( ~n1524 & n11212 ) | ( n3999 & n11212 ) ;
  assign n13366 = n9947 ^ n4894 ^ n204 ;
  assign n13367 = n4545 | n13366 ;
  assign n13368 = ( n1118 & n6529 ) | ( n1118 & n13367 ) | ( n6529 & n13367 ) ;
  assign n13369 = ( n1075 & n2663 ) | ( n1075 & n13368 ) | ( n2663 & n13368 ) ;
  assign n13370 = n5800 & n8261 ;
  assign n13371 = n3683 ^ n3092 ^ 1'b0 ;
  assign n13373 = ( n771 & ~n2383 ) | ( n771 & n5307 ) | ( ~n2383 & n5307 ) ;
  assign n13372 = ( n298 & ~n5419 ) | ( n298 & n7429 ) | ( ~n5419 & n7429 ) ;
  assign n13374 = n13373 ^ n13372 ^ 1'b0 ;
  assign n13375 = n8328 | n13374 ;
  assign n13376 = n13371 & ~n13375 ;
  assign n13377 = n870 & ~n5397 ;
  assign n13378 = ~n3139 & n13377 ;
  assign n13379 = n6681 ^ n1575 ^ 1'b0 ;
  assign n13380 = n7561 | n13379 ;
  assign n13381 = n4093 ^ n3142 ^ n2386 ;
  assign n13382 = n2680 ^ n1675 ^ 1'b0 ;
  assign n13383 = ~n2404 & n12306 ;
  assign n13384 = ~n923 & n13383 ;
  assign n13385 = ( n5629 & n13382 ) | ( n5629 & n13384 ) | ( n13382 & n13384 ) ;
  assign n13386 = n13381 | n13385 ;
  assign n13387 = n9206 ^ n3950 ^ 1'b0 ;
  assign n13388 = ~n449 & n2034 ;
  assign n13389 = n13388 ^ n3038 ^ 1'b0 ;
  assign n13390 = ( n950 & ~n1547 ) | ( n950 & n13389 ) | ( ~n1547 & n13389 ) ;
  assign n13391 = n13390 ^ n5162 ^ 1'b0 ;
  assign n13392 = n13391 ^ n11852 ^ n8743 ;
  assign n13393 = n13392 ^ n6474 ^ 1'b0 ;
  assign n13394 = ~n1283 & n13393 ;
  assign n13396 = n775 & n9259 ;
  assign n13397 = n6002 & n13396 ;
  assign n13395 = ( n1527 & n2656 ) | ( n1527 & n10788 ) | ( n2656 & n10788 ) ;
  assign n13398 = n13397 ^ n13395 ^ n3689 ;
  assign n13399 = n5873 ^ n4394 ^ n4246 ;
  assign n13400 = ( ~n937 & n1732 ) | ( ~n937 & n13399 ) | ( n1732 & n13399 ) ;
  assign n13401 = ( n7063 & n8043 ) | ( n7063 & n13400 ) | ( n8043 & n13400 ) ;
  assign n13402 = n8343 ^ x94 ^ 1'b0 ;
  assign n13403 = n3486 | n13402 ;
  assign n13404 = n6998 ^ n5986 ^ 1'b0 ;
  assign n13405 = ( n995 & ~n8628 ) | ( n995 & n13404 ) | ( ~n8628 & n13404 ) ;
  assign n13406 = n1570 ^ n1353 ^ n1226 ;
  assign n13407 = n2372 & ~n13406 ;
  assign n13408 = n2832 & ~n11850 ;
  assign n13409 = ~n13407 & n13408 ;
  assign n13410 = ( n1512 & ~n2606 ) | ( n1512 & n4634 ) | ( ~n2606 & n4634 ) ;
  assign n13411 = n13410 ^ n4267 ^ n3551 ;
  assign n13412 = ( n708 & ~n8490 ) | ( n708 & n10104 ) | ( ~n8490 & n10104 ) ;
  assign n13413 = n5329 ^ n2080 ^ n2018 ;
  assign n13414 = n8785 ^ n5347 ^ n3843 ;
  assign n13415 = ( n2719 & n6885 ) | ( n2719 & n13414 ) | ( n6885 & n13414 ) ;
  assign n13416 = n10307 ^ n5843 ^ 1'b0 ;
  assign n13417 = ( ~n13413 & n13415 ) | ( ~n13413 & n13416 ) | ( n13415 & n13416 ) ;
  assign n13423 = n2474 | n9845 ;
  assign n13418 = n2303 | n2916 ;
  assign n13419 = n13418 ^ n4408 ^ 1'b0 ;
  assign n13420 = n13031 | n13419 ;
  assign n13421 = n959 & ~n13420 ;
  assign n13422 = n13421 ^ n12263 ^ x78 ;
  assign n13424 = n13423 ^ n13422 ^ n10199 ;
  assign n13425 = ( n346 & n4236 ) | ( n346 & ~n13334 ) | ( n4236 & ~n13334 ) ;
  assign n13426 = n10560 ^ n7016 ^ 1'b0 ;
  assign n13427 = ( ~n486 & n5842 ) | ( ~n486 & n10900 ) | ( n5842 & n10900 ) ;
  assign n13430 = ( n1020 & n1519 ) | ( n1020 & n11883 ) | ( n1519 & n11883 ) ;
  assign n13431 = n13430 ^ n1600 ^ n589 ;
  assign n13432 = n671 & ~n1287 ;
  assign n13433 = ~n13431 & n13432 ;
  assign n13428 = n1266 ^ n1048 ^ 1'b0 ;
  assign n13429 = n13428 ^ n8111 ^ n3924 ;
  assign n13434 = n13433 ^ n13429 ^ n6250 ;
  assign n13435 = ( n1437 & n3237 ) | ( n1437 & ~n8033 ) | ( n3237 & ~n8033 ) ;
  assign n13436 = n13435 ^ n1915 ^ 1'b0 ;
  assign n13437 = n4104 | n13436 ;
  assign n13438 = n4311 | n4345 ;
  assign n13439 = n13438 ^ n4191 ^ 1'b0 ;
  assign n13440 = ( n3764 & ~n9244 ) | ( n3764 & n13439 ) | ( ~n9244 & n13439 ) ;
  assign n13441 = ( n746 & n13437 ) | ( n746 & ~n13440 ) | ( n13437 & ~n13440 ) ;
  assign n13442 = n13441 ^ n2994 ^ 1'b0 ;
  assign n13444 = n3773 ^ n409 ^ 1'b0 ;
  assign n13445 = ( n1376 & n5725 ) | ( n1376 & ~n13444 ) | ( n5725 & ~n13444 ) ;
  assign n13443 = n3495 & n7284 ;
  assign n13446 = n13445 ^ n13443 ^ 1'b0 ;
  assign n13455 = ( n854 & n5408 ) | ( n854 & n8404 ) | ( n5408 & n8404 ) ;
  assign n13456 = n13455 ^ n11718 ^ n1758 ;
  assign n13449 = ( ~n783 & n1159 ) | ( ~n783 & n3223 ) | ( n1159 & n3223 ) ;
  assign n13447 = n9105 ^ n3251 ^ 1'b0 ;
  assign n13448 = ~n8839 & n13447 ;
  assign n13450 = n13449 ^ n13448 ^ 1'b0 ;
  assign n13451 = ~n11922 & n12024 ;
  assign n13452 = ( n6012 & ~n13450 ) | ( n6012 & n13451 ) | ( ~n13450 & n13451 ) ;
  assign n13453 = n4392 ^ n350 ^ 1'b0 ;
  assign n13454 = ~n13452 & n13453 ;
  assign n13457 = n13456 ^ n13454 ^ 1'b0 ;
  assign n13462 = n12892 ^ n10380 ^ 1'b0 ;
  assign n13463 = n13462 ^ n901 ^ 1'b0 ;
  assign n13464 = n13463 ^ n5125 ^ 1'b0 ;
  assign n13465 = n12545 | n13464 ;
  assign n13458 = n2156 ^ n1963 ^ n190 ;
  assign n13459 = n6246 | n13458 ;
  assign n13460 = n3166 | n13459 ;
  assign n13461 = ( ~n3295 & n6606 ) | ( ~n3295 & n13460 ) | ( n6606 & n13460 ) ;
  assign n13466 = n13465 ^ n13461 ^ n6251 ;
  assign n13467 = n8965 ^ n266 ^ 1'b0 ;
  assign n13468 = n13466 | n13467 ;
  assign n13469 = ( n11585 & n13457 ) | ( n11585 & n13468 ) | ( n13457 & n13468 ) ;
  assign n13470 = n5170 ^ n1099 ^ 1'b0 ;
  assign n13471 = ( ~n4239 & n8251 ) | ( ~n4239 & n10552 ) | ( n8251 & n10552 ) ;
  assign n13472 = n498 & n6083 ;
  assign n13473 = ~n1314 & n13472 ;
  assign n13474 = n13473 ^ n5411 ^ 1'b0 ;
  assign n13475 = n9219 ^ n4492 ^ x11 ;
  assign n13476 = ~n5501 & n13475 ;
  assign n13477 = ~n12593 & n13476 ;
  assign n13478 = n13477 ^ n6250 ^ n6247 ;
  assign n13479 = n13478 ^ n6063 ^ 1'b0 ;
  assign n13480 = n6845 ^ n5906 ^ n5015 ;
  assign n13481 = n9250 & n9666 ;
  assign n13482 = ~n13480 & n13481 ;
  assign n13483 = ( ~n636 & n2804 ) | ( ~n636 & n8641 ) | ( n2804 & n8641 ) ;
  assign n13484 = n1610 | n8024 ;
  assign n13485 = n13484 ^ n3454 ^ 1'b0 ;
  assign n13486 = n13485 ^ n7868 ^ 1'b0 ;
  assign n13487 = n1929 & n13486 ;
  assign n13488 = n13487 ^ n2981 ^ 1'b0 ;
  assign n13489 = n1532 & ~n13488 ;
  assign n13490 = ( n1037 & n13483 ) | ( n1037 & n13489 ) | ( n13483 & n13489 ) ;
  assign n13491 = ~n975 & n4401 ;
  assign n13492 = n5272 & n13491 ;
  assign n13493 = n12715 | n13492 ;
  assign n13494 = n13490 | n13493 ;
  assign n13495 = n4532 | n6379 ;
  assign n13496 = n4905 & ~n13495 ;
  assign n13497 = ( n1571 & n4130 ) | ( n1571 & n13496 ) | ( n4130 & n13496 ) ;
  assign n13498 = n13451 ^ n10400 ^ n5439 ;
  assign n13499 = n2596 & ~n6465 ;
  assign n13500 = n7568 & n13499 ;
  assign n13501 = n13500 ^ n12999 ^ 1'b0 ;
  assign n13502 = ~x34 & n476 ;
  assign n13503 = n13502 ^ n3617 ^ n1591 ;
  assign n13504 = ( ~n6899 & n11605 ) | ( ~n6899 & n12315 ) | ( n11605 & n12315 ) ;
  assign n13505 = n13504 ^ n2897 ^ n2022 ;
  assign n13506 = ( n1606 & n3631 ) | ( n1606 & n6768 ) | ( n3631 & n6768 ) ;
  assign n13508 = n12413 ^ n3905 ^ n1868 ;
  assign n13507 = ( ~n4257 & n8306 ) | ( ~n4257 & n9409 ) | ( n8306 & n9409 ) ;
  assign n13509 = n13508 ^ n13507 ^ n3889 ;
  assign n13510 = n13506 & n13509 ;
  assign n13511 = ~n4744 & n13510 ;
  assign n13512 = ( n4017 & ~n5019 ) | ( n4017 & n8033 ) | ( ~n5019 & n8033 ) ;
  assign n13513 = n2873 | n13512 ;
  assign n13514 = n10736 & ~n13513 ;
  assign n13515 = n11830 ^ n3063 ^ 1'b0 ;
  assign n13516 = n10193 ^ n2789 ^ 1'b0 ;
  assign n13517 = ( ~n2430 & n3446 ) | ( ~n2430 & n13516 ) | ( n3446 & n13516 ) ;
  assign n13518 = ( ~n1880 & n5758 ) | ( ~n1880 & n7902 ) | ( n5758 & n7902 ) ;
  assign n13519 = ( n1942 & n13517 ) | ( n1942 & ~n13518 ) | ( n13517 & ~n13518 ) ;
  assign n13520 = ( n3074 & ~n13515 ) | ( n3074 & n13519 ) | ( ~n13515 & n13519 ) ;
  assign n13521 = n8162 | n12475 ;
  assign n13522 = ( ~n2743 & n5322 ) | ( ~n2743 & n13521 ) | ( n5322 & n13521 ) ;
  assign n13524 = n6138 ^ n2098 ^ 1'b0 ;
  assign n13525 = ( n160 & n3110 ) | ( n160 & n13524 ) | ( n3110 & n13524 ) ;
  assign n13526 = n13525 ^ n2517 ^ 1'b0 ;
  assign n13527 = ~n6116 & n13526 ;
  assign n13528 = ~n4365 & n13527 ;
  assign n13529 = n8764 & n13528 ;
  assign n13530 = n13529 ^ n480 ^ 1'b0 ;
  assign n13531 = n5771 & ~n13530 ;
  assign n13532 = ( ~n2069 & n10509 ) | ( ~n2069 & n13531 ) | ( n10509 & n13531 ) ;
  assign n13523 = n591 & n2158 ;
  assign n13533 = n13532 ^ n13523 ^ 1'b0 ;
  assign n13534 = n2825 ^ n1954 ^ 1'b0 ;
  assign n13535 = n4149 & n13534 ;
  assign n13536 = n13535 ^ n4574 ^ 1'b0 ;
  assign n13537 = n10997 ^ n4642 ^ 1'b0 ;
  assign n13538 = n4300 & ~n9440 ;
  assign n13539 = n11838 | n13538 ;
  assign n13540 = n8864 ^ n5870 ^ n1242 ;
  assign n13541 = ( ~n2882 & n3589 ) | ( ~n2882 & n9296 ) | ( n3589 & n9296 ) ;
  assign n13542 = n448 | n13541 ;
  assign n13543 = n295 & ~n13542 ;
  assign n13544 = n5987 ^ n2348 ^ n216 ;
  assign n13545 = n13544 ^ n9257 ^ 1'b0 ;
  assign n13546 = n13545 ^ n11317 ^ n9762 ;
  assign n13547 = ( n5696 & ~n10662 ) | ( n5696 & n13546 ) | ( ~n10662 & n13546 ) ;
  assign n13548 = n3474 & ~n13547 ;
  assign n13549 = n435 & n13548 ;
  assign n13551 = n6199 ^ n4302 ^ n1130 ;
  assign n13552 = ( n2426 & ~n4813 ) | ( n2426 & n13551 ) | ( ~n4813 & n13551 ) ;
  assign n13553 = n13552 ^ n7871 ^ 1'b0 ;
  assign n13554 = n1962 | n13553 ;
  assign n13550 = ( n3574 & n5487 ) | ( n3574 & n6210 ) | ( n5487 & n6210 ) ;
  assign n13555 = n13554 ^ n13550 ^ x123 ;
  assign n13556 = n7757 ^ n3246 ^ 1'b0 ;
  assign n13557 = n13556 ^ n11390 ^ n4181 ;
  assign n13558 = n9389 ^ n5862 ^ n4213 ;
  assign n13559 = n2198 & n4147 ;
  assign n13560 = n3418 & n13559 ;
  assign n13561 = ( n2293 & ~n7934 ) | ( n2293 & n13560 ) | ( ~n7934 & n13560 ) ;
  assign n13562 = ( n1376 & n7739 ) | ( n1376 & n10566 ) | ( n7739 & n10566 ) ;
  assign n13563 = ( n6365 & n13219 ) | ( n6365 & n13562 ) | ( n13219 & n13562 ) ;
  assign n13569 = ~n3197 & n13290 ;
  assign n13570 = n13569 ^ n178 ^ 1'b0 ;
  assign n13571 = n423 & n4398 ;
  assign n13572 = n13570 & n13571 ;
  assign n13567 = ( n1197 & ~n1644 ) | ( n1197 & n3236 ) | ( ~n1644 & n3236 ) ;
  assign n13568 = n1860 & n13567 ;
  assign n13573 = n13572 ^ n13568 ^ 1'b0 ;
  assign n13564 = n12158 ^ n9600 ^ n3690 ;
  assign n13565 = ( n4270 & ~n11106 ) | ( n4270 & n13564 ) | ( ~n11106 & n13564 ) ;
  assign n13566 = n3964 | n13565 ;
  assign n13574 = n13573 ^ n13566 ^ 1'b0 ;
  assign n13575 = n4240 ^ n3862 ^ 1'b0 ;
  assign n13576 = ( ~n4553 & n11738 ) | ( ~n4553 & n13575 ) | ( n11738 & n13575 ) ;
  assign n13577 = n10083 & ~n12983 ;
  assign n13580 = ( n1013 & n4964 ) | ( n1013 & n6346 ) | ( n4964 & n6346 ) ;
  assign n13578 = ( n6580 & n7405 ) | ( n6580 & ~n10758 ) | ( n7405 & ~n10758 ) ;
  assign n13579 = n6159 | n13578 ;
  assign n13581 = n13580 ^ n13579 ^ n3973 ;
  assign n13582 = n429 & ~n6816 ;
  assign n13583 = n13582 ^ n1744 ^ 1'b0 ;
  assign n13584 = n13583 ^ n9006 ^ n1987 ;
  assign n13585 = n13584 ^ n8630 ^ n4025 ;
  assign n13586 = n8577 & n8815 ;
  assign n13587 = ~n13585 & n13586 ;
  assign n13588 = n13587 ^ n7313 ^ n630 ;
  assign n13589 = ( n1559 & n4271 ) | ( n1559 & ~n11080 ) | ( n4271 & ~n11080 ) ;
  assign n13590 = ( n4968 & n6786 ) | ( n4968 & n13589 ) | ( n6786 & n13589 ) ;
  assign n13592 = n6658 ^ x88 ^ 1'b0 ;
  assign n13593 = ~n5110 & n13592 ;
  assign n13594 = ( n1188 & n3390 ) | ( n1188 & n13593 ) | ( n3390 & n13593 ) ;
  assign n13591 = ( n1149 & n3783 ) | ( n1149 & ~n6976 ) | ( n3783 & ~n6976 ) ;
  assign n13595 = n13594 ^ n13591 ^ n12670 ;
  assign n13596 = ~x53 & n12328 ;
  assign n13601 = ~n11616 & n11925 ;
  assign n13597 = n8002 ^ n2740 ^ 1'b0 ;
  assign n13598 = ~n1495 & n13597 ;
  assign n13599 = ~n2389 & n13598 ;
  assign n13600 = n1573 & n13599 ;
  assign n13602 = n13601 ^ n13600 ^ 1'b0 ;
  assign n13603 = n8943 ^ n5318 ^ n1478 ;
  assign n13604 = n12323 & ~n13603 ;
  assign n13605 = ( n7473 & ~n7724 ) | ( n7473 & n10660 ) | ( ~n7724 & n10660 ) ;
  assign n13606 = n13605 ^ n4906 ^ n4343 ;
  assign n13607 = ( n6617 & n11564 ) | ( n6617 & ~n13492 ) | ( n11564 & ~n13492 ) ;
  assign n13608 = n10380 ^ n5283 ^ n4673 ;
  assign n13609 = n13608 ^ n1413 ^ 1'b0 ;
  assign n13610 = ( ~n721 & n12958 ) | ( ~n721 & n13609 ) | ( n12958 & n13609 ) ;
  assign n13611 = ( n1893 & ~n13181 ) | ( n1893 & n13610 ) | ( ~n13181 & n13610 ) ;
  assign n13612 = n3055 & n5376 ;
  assign n13613 = n9701 ^ n3147 ^ 1'b0 ;
  assign n13614 = n2959 & ~n13613 ;
  assign n13615 = n5141 & ~n13614 ;
  assign n13616 = ( n627 & n1254 ) | ( n627 & n12792 ) | ( n1254 & n12792 ) ;
  assign n13617 = ( ~n11540 & n13615 ) | ( ~n11540 & n13616 ) | ( n13615 & n13616 ) ;
  assign n13618 = ( x115 & ~n137 ) | ( x115 & n5813 ) | ( ~n137 & n5813 ) ;
  assign n13622 = ( ~n683 & n1268 ) | ( ~n683 & n2370 ) | ( n1268 & n2370 ) ;
  assign n13619 = n2622 & n5915 ;
  assign n13620 = n13619 ^ n5289 ^ 1'b0 ;
  assign n13621 = n13620 ^ n7072 ^ 1'b0 ;
  assign n13623 = n13622 ^ n13621 ^ n12458 ;
  assign n13624 = ( n3238 & ~n6483 ) | ( n3238 & n6860 ) | ( ~n6483 & n6860 ) ;
  assign n13625 = n1441 & ~n4608 ;
  assign n13626 = n10659 | n13625 ;
  assign n13627 = n4590 | n13626 ;
  assign n13628 = ~n13624 & n13627 ;
  assign n13629 = n8082 ^ n8023 ^ 1'b0 ;
  assign n13630 = ~n9317 & n13629 ;
  assign n13631 = n1584 & n13630 ;
  assign n13632 = ( n3297 & n13628 ) | ( n3297 & ~n13631 ) | ( n13628 & ~n13631 ) ;
  assign n13633 = ~n2033 & n3575 ;
  assign n13634 = ( n6028 & n6623 ) | ( n6028 & ~n13633 ) | ( n6623 & ~n13633 ) ;
  assign n13635 = ~n6596 & n10210 ;
  assign n13636 = ~n13634 & n13635 ;
  assign n13637 = ( n4420 & n11897 ) | ( n4420 & ~n13636 ) | ( n11897 & ~n13636 ) ;
  assign n13646 = ( n8316 & n8376 ) | ( n8316 & ~n9352 ) | ( n8376 & ~n9352 ) ;
  assign n13644 = n11346 & ~n11563 ;
  assign n13645 = n13644 ^ n11544 ^ 1'b0 ;
  assign n13640 = n2732 & ~n3298 ;
  assign n13641 = n13640 ^ n4557 ^ 1'b0 ;
  assign n13638 = n3969 | n12398 ;
  assign n13639 = n13638 ^ n9508 ^ 1'b0 ;
  assign n13642 = n13641 ^ n13639 ^ n5545 ;
  assign n13643 = n13642 ^ n6567 ^ 1'b0 ;
  assign n13647 = n13646 ^ n13645 ^ n13643 ;
  assign n13648 = n10096 ^ n4811 ^ 1'b0 ;
  assign n13649 = n10858 & n13648 ;
  assign n13650 = n2251 ^ n1728 ^ 1'b0 ;
  assign n13651 = n2053 ^ n1339 ^ 1'b0 ;
  assign n13652 = n758 & n3902 ;
  assign n13653 = n8965 & n13652 ;
  assign n13654 = n13651 | n13653 ;
  assign n13655 = n13650 | n13654 ;
  assign n13656 = n2101 ^ n1522 ^ n904 ;
  assign n13657 = n1559 & n13656 ;
  assign n13658 = ~n5466 & n13657 ;
  assign n13660 = n2902 | n6649 ;
  assign n13659 = n10437 ^ n1778 ^ 1'b0 ;
  assign n13661 = n13660 ^ n13659 ^ 1'b0 ;
  assign n13662 = ( n5155 & n5866 ) | ( n5155 & ~n7831 ) | ( n5866 & ~n7831 ) ;
  assign n13663 = n13662 ^ n12517 ^ n1301 ;
  assign n13664 = n5658 ^ n3023 ^ n2060 ;
  assign n13665 = ( n2101 & ~n4352 ) | ( n2101 & n4481 ) | ( ~n4352 & n4481 ) ;
  assign n13666 = n13664 & n13665 ;
  assign n13667 = n13666 ^ n5371 ^ 1'b0 ;
  assign n13668 = n3520 & ~n13667 ;
  assign n13669 = ~n6738 & n10978 ;
  assign n13670 = n13668 | n13669 ;
  assign n13671 = n13670 ^ n8919 ^ 1'b0 ;
  assign n13672 = n12735 ^ n5470 ^ n1097 ;
  assign n13673 = ( n1040 & n3922 ) | ( n1040 & ~n8812 ) | ( n3922 & ~n8812 ) ;
  assign n13674 = ( n4151 & n7003 ) | ( n4151 & ~n9805 ) | ( n7003 & ~n9805 ) ;
  assign n13675 = n13674 ^ n8143 ^ 1'b0 ;
  assign n13676 = ( n1058 & ~n13673 ) | ( n1058 & n13675 ) | ( ~n13673 & n13675 ) ;
  assign n13677 = n13676 ^ n5346 ^ n2790 ;
  assign n13678 = n9128 ^ n7567 ^ n3592 ;
  assign n13679 = n5009 ^ n3902 ^ 1'b0 ;
  assign n13680 = ( ~n3883 & n11090 ) | ( ~n3883 & n12029 ) | ( n11090 & n12029 ) ;
  assign n13681 = n13679 | n13680 ;
  assign n13682 = n8377 ^ n4353 ^ 1'b0 ;
  assign n13683 = n1706 | n13682 ;
  assign n13684 = n12190 ^ n11463 ^ n2925 ;
  assign n13685 = n13684 ^ n7309 ^ n2552 ;
  assign n13686 = n8644 ^ n2968 ^ n854 ;
  assign n13687 = ~n4611 & n6650 ;
  assign n13688 = ( n2819 & n13157 ) | ( n2819 & ~n13687 ) | ( n13157 & ~n13687 ) ;
  assign n13689 = ( ~n4677 & n13686 ) | ( ~n4677 & n13688 ) | ( n13686 & n13688 ) ;
  assign n13690 = n13689 ^ n6189 ^ n1854 ;
  assign n13692 = ( ~n1300 & n3053 ) | ( ~n1300 & n7407 ) | ( n3053 & n7407 ) ;
  assign n13691 = n3975 & n5777 ;
  assign n13693 = n13692 ^ n13691 ^ 1'b0 ;
  assign n13694 = ~n5254 & n7806 ;
  assign n13695 = n13694 ^ n3441 ^ 1'b0 ;
  assign n13696 = n13695 ^ n4883 ^ n460 ;
  assign n13697 = n9637 ^ n5833 ^ n675 ;
  assign n13698 = n13697 ^ n8958 ^ n1081 ;
  assign n13700 = n13345 ^ n4590 ^ n200 ;
  assign n13701 = n13700 ^ n469 ^ 1'b0 ;
  assign n13699 = ~n3377 & n11869 ;
  assign n13702 = n13701 ^ n13699 ^ 1'b0 ;
  assign n13704 = n3136 ^ n2296 ^ n738 ;
  assign n13705 = n13704 ^ n8806 ^ 1'b0 ;
  assign n13703 = n4145 & ~n12959 ;
  assign n13706 = n13705 ^ n13703 ^ 1'b0 ;
  assign n13709 = ~n7350 & n10595 ;
  assign n13707 = n771 | n11029 ;
  assign n13708 = ~n3319 & n13707 ;
  assign n13710 = n13709 ^ n13708 ^ 1'b0 ;
  assign n13711 = n8811 & ~n11760 ;
  assign n13714 = n917 & ~n1769 ;
  assign n13712 = ( n1416 & ~n5168 ) | ( n1416 & n6404 ) | ( ~n5168 & n6404 ) ;
  assign n13713 = n13712 ^ n3790 ^ n168 ;
  assign n13715 = n13714 ^ n13713 ^ n8054 ;
  assign n13716 = n13715 ^ n9178 ^ 1'b0 ;
  assign n13717 = n8178 | n9628 ;
  assign n13718 = n13716 & n13717 ;
  assign n13719 = n13711 & n13718 ;
  assign n13721 = ( n5638 & ~n13423 ) | ( n5638 & n13715 ) | ( ~n13423 & n13715 ) ;
  assign n13720 = n9586 & ~n11280 ;
  assign n13722 = n13721 ^ n13720 ^ 1'b0 ;
  assign n13723 = n2043 & n2125 ;
  assign n13724 = n13723 ^ n7480 ^ 1'b0 ;
  assign n13725 = n3361 & ~n13724 ;
  assign n13726 = n13722 & ~n13725 ;
  assign n13729 = ( n3211 & n4311 ) | ( n3211 & ~n8966 ) | ( n4311 & ~n8966 ) ;
  assign n13730 = ~n2146 & n7268 ;
  assign n13731 = n13730 ^ n4019 ^ n1936 ;
  assign n13732 = ( n1318 & n13729 ) | ( n1318 & n13731 ) | ( n13729 & n13731 ) ;
  assign n13727 = ~n9314 & n11329 ;
  assign n13728 = ( n5391 & ~n8533 ) | ( n5391 & n13727 ) | ( ~n8533 & n13727 ) ;
  assign n13733 = n13732 ^ n13728 ^ n13419 ;
  assign n13740 = n4926 | n12727 ;
  assign n13741 = ( n4615 & n4717 ) | ( n4615 & ~n5043 ) | ( n4717 & ~n5043 ) ;
  assign n13742 = ( n9508 & n13584 ) | ( n9508 & n13741 ) | ( n13584 & n13741 ) ;
  assign n13743 = n13742 ^ n13011 ^ n2097 ;
  assign n13744 = ( n9696 & ~n13740 ) | ( n9696 & n13743 ) | ( ~n13740 & n13743 ) ;
  assign n13734 = n852 & ~n6828 ;
  assign n13735 = ~n778 & n13734 ;
  assign n13736 = ( ~n445 & n1351 ) | ( ~n445 & n5623 ) | ( n1351 & n5623 ) ;
  assign n13737 = n13736 ^ n3061 ^ 1'b0 ;
  assign n13738 = ~n2903 & n13737 ;
  assign n13739 = ( n11957 & ~n13735 ) | ( n11957 & n13738 ) | ( ~n13735 & n13738 ) ;
  assign n13745 = n13744 ^ n13739 ^ n13295 ;
  assign n13746 = n864 & ~n1322 ;
  assign n13747 = n5316 ^ n4612 ^ 1'b0 ;
  assign n13748 = ~n13746 & n13747 ;
  assign n13753 = n3571 ^ n3416 ^ n2779 ;
  assign n13750 = n3324 & ~n3840 ;
  assign n13751 = n13750 ^ n9144 ^ 1'b0 ;
  assign n13752 = n13751 ^ n13688 ^ n10284 ;
  assign n13754 = n13753 ^ n13752 ^ 1'b0 ;
  assign n13749 = n4507 & ~n11833 ;
  assign n13755 = n13754 ^ n13749 ^ 1'b0 ;
  assign n13759 = ( n779 & n9640 ) | ( n779 & ~n11779 ) | ( n9640 & ~n11779 ) ;
  assign n13756 = n13036 ^ n3699 ^ n1822 ;
  assign n13757 = ( n679 & n11528 ) | ( n679 & ~n13756 ) | ( n11528 & ~n13756 ) ;
  assign n13758 = n241 & n13757 ;
  assign n13760 = n13759 ^ n13758 ^ n2398 ;
  assign n13761 = n9095 ^ n3822 ^ n2727 ;
  assign n13762 = n13761 ^ n12505 ^ n3833 ;
  assign n13763 = n13562 ^ n3236 ^ n1537 ;
  assign n13764 = n13763 ^ n10718 ^ 1'b0 ;
  assign n13765 = n13762 | n13764 ;
  assign n13766 = ( ~n4735 & n5554 ) | ( ~n4735 & n10522 ) | ( n5554 & n10522 ) ;
  assign n13767 = ( n2449 & n2810 ) | ( n2449 & ~n4893 ) | ( n2810 & ~n4893 ) ;
  assign n13768 = ~n4971 & n13767 ;
  assign n13769 = n13768 ^ n2970 ^ n791 ;
  assign n13770 = ( n8740 & ~n13766 ) | ( n8740 & n13769 ) | ( ~n13766 & n13769 ) ;
  assign n13771 = n13770 ^ n12200 ^ 1'b0 ;
  assign n13772 = n11957 ^ n3393 ^ n588 ;
  assign n13773 = n13772 ^ n9727 ^ 1'b0 ;
  assign n13774 = n13773 ^ n6208 ^ 1'b0 ;
  assign n13775 = n13608 ^ n11662 ^ n2508 ;
  assign n13776 = n10691 ^ n4869 ^ n3707 ;
  assign n13777 = ( n2565 & n4496 ) | ( n2565 & ~n12124 ) | ( n4496 & ~n12124 ) ;
  assign n13778 = n13777 ^ n9081 ^ 1'b0 ;
  assign n13779 = ( ~n334 & n12976 ) | ( ~n334 & n13778 ) | ( n12976 & n13778 ) ;
  assign n13780 = n8705 ^ n7953 ^ 1'b0 ;
  assign n13781 = n13780 ^ n5780 ^ n4858 ;
  assign n13782 = n9937 | n13546 ;
  assign n13783 = n1696 | n6421 ;
  assign n13784 = n9967 ^ n7749 ^ n1326 ;
  assign n13785 = n13784 ^ n11218 ^ n4970 ;
  assign n13786 = ( n2003 & ~n13783 ) | ( n2003 & n13785 ) | ( ~n13783 & n13785 ) ;
  assign n13787 = ( n994 & n3631 ) | ( n994 & ~n6660 ) | ( n3631 & ~n6660 ) ;
  assign n13788 = ~n521 & n1982 ;
  assign n13789 = n4680 | n5786 ;
  assign n13790 = n7277 & ~n13789 ;
  assign n13791 = n1981 | n8822 ;
  assign n13792 = ( n13788 & n13790 ) | ( n13788 & ~n13791 ) | ( n13790 & ~n13791 ) ;
  assign n13793 = n135 & n9073 ;
  assign n13797 = n7766 ^ n7602 ^ 1'b0 ;
  assign n13794 = ~n8399 & n8439 ;
  assign n13795 = ( x45 & ~n11957 ) | ( x45 & n13794 ) | ( ~n11957 & n13794 ) ;
  assign n13796 = n13795 ^ n6402 ^ 1'b0 ;
  assign n13798 = n13797 ^ n13796 ^ n4939 ;
  assign n13804 = n4608 & n7317 ;
  assign n13800 = ( n5128 & ~n8161 ) | ( n5128 & n10988 ) | ( ~n8161 & n10988 ) ;
  assign n13801 = n4002 & n13800 ;
  assign n13802 = ~n10028 & n13801 ;
  assign n13803 = n13802 ^ n8244 ^ n5313 ;
  assign n13799 = n12072 ^ n10465 ^ 1'b0 ;
  assign n13805 = n13804 ^ n13803 ^ n13799 ;
  assign n13806 = n6325 & ~n13805 ;
  assign n13812 = ( n571 & n3513 ) | ( n571 & n6343 ) | ( n3513 & n6343 ) ;
  assign n13808 = n9067 ^ n4110 ^ 1'b0 ;
  assign n13809 = n2997 & n13808 ;
  assign n13807 = n5647 | n6937 ;
  assign n13810 = n13809 ^ n13807 ^ 1'b0 ;
  assign n13811 = n13810 ^ n9068 ^ n7962 ;
  assign n13813 = n13812 ^ n13811 ^ n4640 ;
  assign n13814 = ( n199 & n258 ) | ( n199 & ~n4645 ) | ( n258 & ~n4645 ) ;
  assign n13815 = ( n3788 & n12973 ) | ( n3788 & n13814 ) | ( n12973 & n13814 ) ;
  assign n13816 = n13815 ^ n4261 ^ 1'b0 ;
  assign n13817 = n13813 & n13816 ;
  assign n13818 = n13817 ^ n7512 ^ n7419 ;
  assign n13819 = ( n1925 & n2281 ) | ( n1925 & ~n10627 ) | ( n2281 & ~n10627 ) ;
  assign n13820 = n2471 | n13819 ;
  assign n13821 = n6879 | n13820 ;
  assign n13827 = ( n4647 & ~n5531 ) | ( n4647 & n11235 ) | ( ~n5531 & n11235 ) ;
  assign n13822 = n4785 ^ n4442 ^ n2990 ;
  assign n13823 = n924 | n6120 ;
  assign n13824 = n13822 | n13823 ;
  assign n13825 = n13824 ^ n5932 ^ n2079 ;
  assign n13826 = ( ~n395 & n1362 ) | ( ~n395 & n13825 ) | ( n1362 & n13825 ) ;
  assign n13828 = n13827 ^ n13826 ^ 1'b0 ;
  assign n13829 = n13821 & n13828 ;
  assign n13830 = ( n1668 & n1839 ) | ( n1668 & ~n2002 ) | ( n1839 & ~n2002 ) ;
  assign n13831 = ~n6783 & n13830 ;
  assign n13832 = n6454 & ~n11349 ;
  assign n13833 = ( ~n907 & n13831 ) | ( ~n907 & n13832 ) | ( n13831 & n13832 ) ;
  assign n13834 = ( ~n5526 & n5916 ) | ( ~n5526 & n13833 ) | ( n5916 & n13833 ) ;
  assign n13835 = ( n3035 & n12643 ) | ( n3035 & n13834 ) | ( n12643 & n13834 ) ;
  assign n13836 = n13835 ^ n4891 ^ n339 ;
  assign n13837 = ( n3592 & n13829 ) | ( n3592 & ~n13836 ) | ( n13829 & ~n13836 ) ;
  assign n13838 = n13837 ^ n10350 ^ n8590 ;
  assign n13844 = n10178 ^ n4236 ^ n1935 ;
  assign n13843 = n3268 & n10358 ;
  assign n13845 = n13844 ^ n13843 ^ n12552 ;
  assign n13839 = n2484 & ~n3604 ;
  assign n13840 = n13839 ^ n5883 ^ 1'b0 ;
  assign n13841 = ~n5810 & n13840 ;
  assign n13842 = n7994 & n13841 ;
  assign n13846 = n13845 ^ n13842 ^ 1'b0 ;
  assign n13847 = ( n1795 & n3671 ) | ( n1795 & n11878 ) | ( n3671 & n11878 ) ;
  assign n13848 = n5862 ^ n3875 ^ n186 ;
  assign n13849 = n8029 & n13848 ;
  assign n13850 = n13847 & n13849 ;
  assign n13851 = ( n7351 & n10447 ) | ( n7351 & ~n13417 ) | ( n10447 & ~n13417 ) ;
  assign n13852 = ( n880 & n2529 ) | ( n880 & ~n6446 ) | ( n2529 & ~n6446 ) ;
  assign n13853 = n13852 ^ n6408 ^ n1158 ;
  assign n13854 = n12788 ^ n12702 ^ n4406 ;
  assign n13855 = ( n6228 & ~n10480 ) | ( n6228 & n13854 ) | ( ~n10480 & n13854 ) ;
  assign n13856 = n8073 ^ n2391 ^ 1'b0 ;
  assign n13857 = n7040 & n13856 ;
  assign n13858 = ( ~n1702 & n5714 ) | ( ~n1702 & n13857 ) | ( n5714 & n13857 ) ;
  assign n13859 = n4030 & n6664 ;
  assign n13860 = n6692 ^ n3360 ^ 1'b0 ;
  assign n13861 = ~n12104 & n13860 ;
  assign n13862 = n607 & ~n5178 ;
  assign n13863 = n13862 ^ n377 ^ 1'b0 ;
  assign n13864 = n8920 | n13863 ;
  assign n13865 = n3994 & ~n13864 ;
  assign n13866 = n1420 & ~n6869 ;
  assign n13867 = n9411 | n13866 ;
  assign n13868 = n13867 ^ n6004 ^ n1673 ;
  assign n13869 = ( n3541 & n13865 ) | ( n3541 & n13868 ) | ( n13865 & n13868 ) ;
  assign n13870 = n2517 & ~n13869 ;
  assign n13871 = n13870 ^ n12193 ^ n4941 ;
  assign n13872 = n8422 ^ n5586 ^ n278 ;
  assign n13873 = n13872 ^ n1408 ^ 1'b0 ;
  assign n13874 = n5591 & ~n13873 ;
  assign n13875 = n2990 | n12923 ;
  assign n13876 = n13875 ^ n1767 ^ n1538 ;
  assign n13877 = n528 & ~n2877 ;
  assign n13878 = n13877 ^ n5428 ^ 1'b0 ;
  assign n13881 = ( ~x31 & n1440 ) | ( ~x31 & n2762 ) | ( n1440 & n2762 ) ;
  assign n13879 = n6032 ^ n5939 ^ n3892 ;
  assign n13880 = n13879 ^ n10030 ^ n3574 ;
  assign n13882 = n13881 ^ n13880 ^ n13660 ;
  assign n13883 = n13878 & ~n13882 ;
  assign n13884 = n13876 & n13883 ;
  assign n13885 = n743 & ~n10451 ;
  assign n13886 = ( n2038 & ~n3380 ) | ( n2038 & n6483 ) | ( ~n3380 & n6483 ) ;
  assign n13887 = n13886 ^ n8270 ^ n4551 ;
  assign n13888 = n13887 ^ n12910 ^ n12752 ;
  assign n13889 = n5527 ^ n3370 ^ n1997 ;
  assign n13890 = n13889 ^ n7736 ^ n4431 ;
  assign n13891 = n1809 & n3335 ;
  assign n13892 = n5140 ^ n460 ^ 1'b0 ;
  assign n13893 = n13891 & ~n13892 ;
  assign n13894 = n4834 ^ n4290 ^ n1699 ;
  assign n13895 = ( n4271 & ~n13893 ) | ( n4271 & n13894 ) | ( ~n13893 & n13894 ) ;
  assign n13896 = n13895 ^ n9555 ^ n877 ;
  assign n13897 = x105 & n13078 ;
  assign n13898 = n13897 ^ n12172 ^ n6063 ;
  assign n13899 = n8691 ^ n8630 ^ n5252 ;
  assign n13900 = ( n5634 & ~n7246 ) | ( n5634 & n13899 ) | ( ~n7246 & n13899 ) ;
  assign n13901 = n6680 | n13900 ;
  assign n13902 = n13636 & ~n13901 ;
  assign n13903 = ( ~n670 & n4341 ) | ( ~n670 & n5501 ) | ( n4341 & n5501 ) ;
  assign n13904 = ( n238 & n3931 ) | ( n238 & ~n12583 ) | ( n3931 & ~n12583 ) ;
  assign n13905 = n13903 & ~n13904 ;
  assign n13906 = ( n1325 & n5601 ) | ( n1325 & n9524 ) | ( n5601 & n9524 ) ;
  assign n13907 = ( n3187 & ~n6320 ) | ( n3187 & n13906 ) | ( ~n6320 & n13906 ) ;
  assign n13908 = n324 & ~n1625 ;
  assign n13909 = n13386 ^ n3999 ^ 1'b0 ;
  assign n13910 = n13908 & ~n13909 ;
  assign n13911 = n11269 ^ x27 ^ 1'b0 ;
  assign n13912 = n12674 | n13911 ;
  assign n13913 = ~n369 & n865 ;
  assign n13914 = n430 & n13913 ;
  assign n13915 = n13914 ^ n6437 ^ n5559 ;
  assign n13916 = n13915 ^ n5621 ^ n4632 ;
  assign n13917 = ( n4378 & n5428 ) | ( n4378 & n13916 ) | ( n5428 & n13916 ) ;
  assign n13918 = n1227 & n4082 ;
  assign n13919 = n4448 & n13918 ;
  assign n13920 = n2529 | n13919 ;
  assign n13921 = n3186 & n7530 ;
  assign n13922 = n13921 ^ n4239 ^ 1'b0 ;
  assign n13923 = n13920 & ~n13922 ;
  assign n13924 = ( n4560 & ~n13917 ) | ( n4560 & n13923 ) | ( ~n13917 & n13923 ) ;
  assign n13925 = ( n2343 & ~n3982 ) | ( n2343 & n4913 ) | ( ~n3982 & n4913 ) ;
  assign n13926 = n2222 & ~n7735 ;
  assign n13927 = n13926 ^ n6590 ^ 1'b0 ;
  assign n13928 = ( n1650 & ~n2081 ) | ( n1650 & n13927 ) | ( ~n2081 & n13927 ) ;
  assign n13929 = n13928 ^ n13551 ^ n4014 ;
  assign n13930 = ~n7058 & n13929 ;
  assign n13935 = n130 & ~n5858 ;
  assign n13936 = n13935 ^ n4553 ^ 1'b0 ;
  assign n13931 = n3511 ^ n410 ^ 1'b0 ;
  assign n13932 = ~n6711 & n13931 ;
  assign n13933 = n13932 ^ n10601 ^ n6929 ;
  assign n13934 = ~n2767 & n13933 ;
  assign n13937 = n13936 ^ n13934 ^ 1'b0 ;
  assign n13938 = n13428 ^ n2611 ^ x42 ;
  assign n13939 = n1184 & ~n13938 ;
  assign n13940 = ~n3834 & n13939 ;
  assign n13941 = n6253 | n10571 ;
  assign n13942 = n13941 ^ n5022 ^ n635 ;
  assign n13943 = n13942 ^ n9068 ^ n2348 ;
  assign n13944 = ( n6294 & n7404 ) | ( n6294 & ~n9597 ) | ( n7404 & ~n9597 ) ;
  assign n13947 = n5916 ^ n1263 ^ 1'b0 ;
  assign n13945 = n12016 ^ n1703 ^ 1'b0 ;
  assign n13946 = n5117 & ~n13945 ;
  assign n13948 = n13947 ^ n13946 ^ 1'b0 ;
  assign n13949 = n8797 & ~n13948 ;
  assign n13950 = n10819 ^ n2702 ^ n549 ;
  assign n13951 = n1538 & ~n13950 ;
  assign n13952 = ~n10582 & n13951 ;
  assign n13953 = n8651 & ~n10707 ;
  assign n13954 = ( ~n5802 & n10118 ) | ( ~n5802 & n13953 ) | ( n10118 & n13953 ) ;
  assign n13955 = n3809 ^ n1567 ^ 1'b0 ;
  assign n13956 = n8135 ^ n6603 ^ n352 ;
  assign n13957 = n13955 | n13956 ;
  assign n13958 = n6823 | n13957 ;
  assign n13960 = n12504 ^ n9382 ^ n6318 ;
  assign n13961 = x74 & n13960 ;
  assign n13962 = ~n13608 & n13961 ;
  assign n13959 = n10611 ^ n1445 ^ n453 ;
  assign n13963 = n13962 ^ n13959 ^ n3520 ;
  assign n13967 = x21 | n3108 ;
  assign n13968 = n13967 ^ n3421 ^ n2377 ;
  assign n13969 = ( ~n6485 & n6532 ) | ( ~n6485 & n13968 ) | ( n6532 & n13968 ) ;
  assign n13970 = n13969 ^ n10228 ^ 1'b0 ;
  assign n13971 = ~n4338 & n13970 ;
  assign n13972 = n7270 ^ n6106 ^ n278 ;
  assign n13973 = ( n768 & ~n13971 ) | ( n768 & n13972 ) | ( ~n13971 & n13972 ) ;
  assign n13964 = ( n3272 & ~n3853 ) | ( n3272 & n4420 ) | ( ~n3853 & n4420 ) ;
  assign n13965 = n10405 | n13964 ;
  assign n13966 = ( n6094 & ~n6183 ) | ( n6094 & n13965 ) | ( ~n6183 & n13965 ) ;
  assign n13974 = n13973 ^ n13966 ^ n5119 ;
  assign n13978 = n167 | n8042 ;
  assign n13979 = n13978 ^ n617 ^ 1'b0 ;
  assign n13977 = n10276 ^ n6995 ^ 1'b0 ;
  assign n13975 = n7882 ^ n3862 ^ n1341 ;
  assign n13976 = n13975 ^ n2292 ^ n921 ;
  assign n13980 = n13979 ^ n13977 ^ n13976 ;
  assign n13981 = n12360 ^ n4345 ^ n1755 ;
  assign n13982 = ( n2283 & ~n7382 ) | ( n2283 & n13981 ) | ( ~n7382 & n13981 ) ;
  assign n13983 = ( n3043 & ~n6361 ) | ( n3043 & n13982 ) | ( ~n6361 & n13982 ) ;
  assign n13984 = ~n1541 & n13983 ;
  assign n13985 = n7170 & n13984 ;
  assign n13986 = ~n1800 & n6159 ;
  assign n13987 = n6442 | n9468 ;
  assign n13988 = n2136 ^ n2124 ^ 1'b0 ;
  assign n13989 = ( ~n1376 & n5489 ) | ( ~n1376 & n6363 ) | ( n5489 & n6363 ) ;
  assign n13990 = n12259 ^ n5554 ^ 1'b0 ;
  assign n13991 = ( ~n8819 & n13989 ) | ( ~n8819 & n13990 ) | ( n13989 & n13990 ) ;
  assign n13992 = n7221 & n13991 ;
  assign n13993 = n1822 & ~n2837 ;
  assign n13994 = n1443 & ~n13993 ;
  assign n13995 = ~n3250 & n3418 ;
  assign n13996 = ( n1535 & n2036 ) | ( n1535 & n12634 ) | ( n2036 & n12634 ) ;
  assign n13997 = ( n8885 & n13995 ) | ( n8885 & ~n13996 ) | ( n13995 & ~n13996 ) ;
  assign n13998 = n13997 ^ n12864 ^ n12347 ;
  assign n13999 = n6200 ^ n5578 ^ n4545 ;
  assign n14000 = n1374 ^ n1129 ^ 1'b0 ;
  assign n14001 = n13999 & n14000 ;
  assign n14002 = n14001 ^ n10318 ^ n2538 ;
  assign n14006 = ( n6045 & ~n9029 ) | ( n6045 & n13309 ) | ( ~n9029 & n13309 ) ;
  assign n14007 = n6446 ^ n5620 ^ n5340 ;
  assign n14008 = ( n1240 & n14006 ) | ( n1240 & ~n14007 ) | ( n14006 & ~n14007 ) ;
  assign n14004 = n8248 & n10539 ;
  assign n14005 = n14004 ^ n1967 ^ 1'b0 ;
  assign n14003 = ( n6621 & ~n7911 ) | ( n6621 & n8812 ) | ( ~n7911 & n8812 ) ;
  assign n14009 = n14008 ^ n14005 ^ n14003 ;
  assign n14010 = ( ~n4940 & n7954 ) | ( ~n4940 & n13665 ) | ( n7954 & n13665 ) ;
  assign n14013 = ( n225 & n1899 ) | ( n225 & ~n7857 ) | ( n1899 & ~n7857 ) ;
  assign n14011 = n5254 ^ n3495 ^ 1'b0 ;
  assign n14012 = n5778 | n14011 ;
  assign n14014 = n14013 ^ n14012 ^ 1'b0 ;
  assign n14015 = n13609 ^ n1890 ^ n1317 ;
  assign n14016 = ( n2031 & n5373 ) | ( n2031 & n14015 ) | ( n5373 & n14015 ) ;
  assign n14017 = n9517 & n14016 ;
  assign n14018 = n14017 ^ n7884 ^ 1'b0 ;
  assign n14019 = n9064 ^ n8005 ^ 1'b0 ;
  assign n14020 = n5310 & n14019 ;
  assign n14021 = n14020 ^ n8659 ^ 1'b0 ;
  assign n14022 = n2506 & n14021 ;
  assign n14023 = n14022 ^ n7538 ^ n706 ;
  assign n14025 = n10377 ^ n5496 ^ 1'b0 ;
  assign n14026 = n2917 | n4167 ;
  assign n14027 = n14025 | n14026 ;
  assign n14028 = ( n4412 & ~n8475 ) | ( n4412 & n14027 ) | ( ~n8475 & n14027 ) ;
  assign n14024 = ( n5678 & n7445 ) | ( n5678 & ~n9802 ) | ( n7445 & ~n9802 ) ;
  assign n14029 = n14028 ^ n14024 ^ n9757 ;
  assign n14030 = ( n1869 & n2260 ) | ( n1869 & ~n4972 ) | ( n2260 & ~n4972 ) ;
  assign n14031 = ( n3653 & ~n5485 ) | ( n3653 & n14030 ) | ( ~n5485 & n14030 ) ;
  assign n14032 = ( ~n2896 & n7778 ) | ( ~n2896 & n14031 ) | ( n7778 & n14031 ) ;
  assign n14033 = ( n3788 & n6963 ) | ( n3788 & n10639 ) | ( n6963 & n10639 ) ;
  assign n14034 = n14033 ^ n5897 ^ 1'b0 ;
  assign n14035 = n6956 | n14034 ;
  assign n14036 = n14035 ^ n13531 ^ 1'b0 ;
  assign n14037 = ( n7800 & ~n13136 ) | ( n7800 & n14036 ) | ( ~n13136 & n14036 ) ;
  assign n14038 = n10670 ^ n7086 ^ 1'b0 ;
  assign n14047 = n1152 & ~n3840 ;
  assign n14048 = n2474 | n14047 ;
  assign n14049 = n14048 ^ n585 ^ 1'b0 ;
  assign n14040 = n9936 ^ n3453 ^ n2230 ;
  assign n14041 = ~n289 & n14040 ;
  assign n14039 = n12249 ^ n7947 ^ n2015 ;
  assign n14042 = n14041 ^ n14039 ^ n6713 ;
  assign n14043 = n1741 ^ n977 ^ 1'b0 ;
  assign n14044 = n2650 & n14043 ;
  assign n14045 = ( n268 & n14042 ) | ( n268 & n14044 ) | ( n14042 & n14044 ) ;
  assign n14046 = n14045 ^ n11328 ^ 1'b0 ;
  assign n14050 = n14049 ^ n14046 ^ n4869 ;
  assign n14051 = n9833 ^ n7809 ^ n2882 ;
  assign n14052 = n1055 & n14051 ;
  assign n14053 = n14052 ^ n1966 ^ 1'b0 ;
  assign n14054 = n14053 ^ n3238 ^ 1'b0 ;
  assign n14055 = n6876 ^ n4422 ^ n4184 ;
  assign n14056 = n14055 ^ n9917 ^ n699 ;
  assign n14057 = ( n2237 & ~n10937 ) | ( n2237 & n14056 ) | ( ~n10937 & n14056 ) ;
  assign n14058 = n231 | n6258 ;
  assign n14059 = ( n1764 & n10818 ) | ( n1764 & ~n14058 ) | ( n10818 & ~n14058 ) ;
  assign n14060 = n4654 ^ n2825 ^ 1'b0 ;
  assign n14061 = ~n6238 & n14060 ;
  assign n14062 = ~n14059 & n14061 ;
  assign n14065 = ( n4830 & ~n7373 ) | ( n4830 & n9696 ) | ( ~n7373 & n9696 ) ;
  assign n14063 = n1380 ^ n182 ^ 1'b0 ;
  assign n14064 = n2235 & ~n14063 ;
  assign n14066 = n14065 ^ n14064 ^ 1'b0 ;
  assign n14067 = n4388 ^ n1667 ^ 1'b0 ;
  assign n14068 = n1599 & n14067 ;
  assign n14069 = n13989 ^ n12068 ^ n11706 ;
  assign n14070 = n8146 ^ n1989 ^ n591 ;
  assign n14071 = ( n880 & n14069 ) | ( n880 & n14070 ) | ( n14069 & n14070 ) ;
  assign n14072 = ( n5972 & n14068 ) | ( n5972 & ~n14071 ) | ( n14068 & ~n14071 ) ;
  assign n14073 = n467 & ~n1100 ;
  assign n14074 = n4968 & n14073 ;
  assign n14075 = ~n4044 & n14074 ;
  assign n14076 = n7420 | n8161 ;
  assign n14077 = n14076 ^ x44 ^ 1'b0 ;
  assign n14078 = n7628 ^ n3141 ^ x28 ;
  assign n14079 = n14078 ^ n10023 ^ 1'b0 ;
  assign n14080 = n14077 & ~n14079 ;
  assign n14081 = n13614 ^ n11007 ^ n5978 ;
  assign n14082 = n12844 ^ n4199 ^ 1'b0 ;
  assign n14083 = n7105 ^ n6246 ^ n3730 ;
  assign n14084 = ( n8560 & ~n8739 ) | ( n8560 & n14083 ) | ( ~n8739 & n14083 ) ;
  assign n14086 = n4905 ^ n3868 ^ n2206 ;
  assign n14085 = n7475 ^ n5613 ^ n4207 ;
  assign n14087 = n14086 ^ n14085 ^ n9361 ;
  assign n14088 = n3384 | n4774 ;
  assign n14089 = n1047 | n4468 ;
  assign n14090 = n1836 & ~n14089 ;
  assign n14091 = ( ~n10351 & n14088 ) | ( ~n10351 & n14090 ) | ( n14088 & n14090 ) ;
  assign n14092 = ( ~n827 & n1204 ) | ( ~n827 & n8390 ) | ( n1204 & n8390 ) ;
  assign n14093 = n8007 | n14092 ;
  assign n14094 = n5916 ^ n1736 ^ n1545 ;
  assign n14095 = n14094 ^ n8440 ^ 1'b0 ;
  assign n14104 = n8996 ^ n7064 ^ n2281 ;
  assign n14096 = n7514 ^ n5916 ^ 1'b0 ;
  assign n14099 = n2885 | n4273 ;
  assign n14100 = n14099 ^ n1467 ^ 1'b0 ;
  assign n14097 = n1028 | n1112 ;
  assign n14098 = n1466 | n14097 ;
  assign n14101 = n14100 ^ n14098 ^ n1688 ;
  assign n14102 = ( n3197 & n5183 ) | ( n3197 & n14101 ) | ( n5183 & n14101 ) ;
  assign n14103 = n14096 | n14102 ;
  assign n14105 = n14104 ^ n14103 ^ 1'b0 ;
  assign n14106 = n12626 ^ n4909 ^ 1'b0 ;
  assign n14107 = n4528 & ~n14106 ;
  assign n14108 = n11075 ^ n917 ^ x32 ;
  assign n14109 = ( n3739 & n9007 ) | ( n3739 & n14108 ) | ( n9007 & n14108 ) ;
  assign n14110 = n3994 & ~n14109 ;
  assign n14111 = n14110 ^ n11211 ^ n6129 ;
  assign n14112 = n3856 | n4316 ;
  assign n14113 = n14112 ^ n2568 ^ 1'b0 ;
  assign n14114 = n14113 ^ n13614 ^ n7351 ;
  assign n14115 = ( n1603 & n5018 ) | ( n1603 & n7703 ) | ( n5018 & n7703 ) ;
  assign n14116 = n4936 | n14115 ;
  assign n14117 = n14116 ^ n12909 ^ n5817 ;
  assign n14118 = n14117 ^ n2377 ^ n1363 ;
  assign n14119 = ( n10140 & n13589 ) | ( n10140 & ~n14118 ) | ( n13589 & ~n14118 ) ;
  assign n14120 = n6566 ^ n3392 ^ n423 ;
  assign n14121 = n5054 & ~n9119 ;
  assign n14122 = ~n1751 & n14121 ;
  assign n14125 = n6498 ^ n405 ^ 1'b0 ;
  assign n14123 = n10306 ^ n7449 ^ n4659 ;
  assign n14124 = n394 | n14123 ;
  assign n14126 = n14125 ^ n14124 ^ 1'b0 ;
  assign n14127 = n3234 ^ x21 ^ 1'b0 ;
  assign n14128 = n5741 & n14127 ;
  assign n14129 = ( n699 & ~n7977 ) | ( n699 & n14128 ) | ( ~n7977 & n14128 ) ;
  assign n14130 = n10056 ^ n5219 ^ 1'b0 ;
  assign n14131 = n14129 & ~n14130 ;
  assign n14132 = n1573 & n14131 ;
  assign n14133 = n6474 ^ n2366 ^ 1'b0 ;
  assign n14134 = ~n9237 & n14133 ;
  assign n14135 = ( n706 & n8156 ) | ( n706 & ~n11651 ) | ( n8156 & ~n11651 ) ;
  assign n14136 = n14135 ^ n2191 ^ n1335 ;
  assign n14137 = ( n10916 & n14134 ) | ( n10916 & n14136 ) | ( n14134 & n14136 ) ;
  assign n14138 = ( n1242 & ~n1566 ) | ( n1242 & n4950 ) | ( ~n1566 & n4950 ) ;
  assign n14139 = n13712 ^ n9678 ^ 1'b0 ;
  assign n14140 = n14139 ^ n9144 ^ n3559 ;
  assign n14141 = ~n6173 & n7066 ;
  assign n14142 = n1038 & n14141 ;
  assign n14143 = ~n3766 & n10251 ;
  assign n14144 = ~n7955 & n14143 ;
  assign n14145 = n14144 ^ n4770 ^ n4067 ;
  assign n14146 = ~n12534 & n14145 ;
  assign n14147 = n816 | n5578 ;
  assign n14148 = n14147 ^ n3831 ^ 1'b0 ;
  assign n14149 = n6949 | n9409 ;
  assign n14150 = ( n4061 & n14148 ) | ( n4061 & ~n14149 ) | ( n14148 & ~n14149 ) ;
  assign n14151 = ( n1929 & n2324 ) | ( n1929 & n14150 ) | ( n2324 & n14150 ) ;
  assign n14152 = ( n10641 & n14146 ) | ( n10641 & n14151 ) | ( n14146 & n14151 ) ;
  assign n14158 = ~n6138 & n8241 ;
  assign n14159 = n14158 ^ n3515 ^ 1'b0 ;
  assign n14154 = n4201 ^ n1919 ^ 1'b0 ;
  assign n14155 = n7337 & ~n14154 ;
  assign n14153 = n1496 & n5116 ;
  assign n14156 = n14155 ^ n14153 ^ 1'b0 ;
  assign n14157 = n12994 | n14156 ;
  assign n14160 = n14159 ^ n14157 ^ 1'b0 ;
  assign n14161 = n1044 & ~n4711 ;
  assign n14162 = n14161 ^ n10767 ^ n3368 ;
  assign n14163 = ~n7370 & n8511 ;
  assign n14164 = n4800 ^ n870 ^ 1'b0 ;
  assign n14165 = n6209 ^ n4338 ^ x24 ;
  assign n14166 = ( n1148 & n6911 ) | ( n1148 & ~n14165 ) | ( n6911 & ~n14165 ) ;
  assign n14167 = n5699 & n8541 ;
  assign n14168 = n14167 ^ n3058 ^ 1'b0 ;
  assign n14169 = n2582 | n14168 ;
  assign n14170 = n5087 & ~n8240 ;
  assign n14171 = n14170 ^ n718 ^ 1'b0 ;
  assign n14172 = n10323 ^ n3375 ^ 1'b0 ;
  assign n14173 = n6403 ^ n4765 ^ n510 ;
  assign n14174 = n2611 & ~n14173 ;
  assign n14175 = n14174 ^ n6937 ^ 1'b0 ;
  assign n14176 = n2909 ^ n2716 ^ 1'b0 ;
  assign n14177 = ( n2253 & ~n2787 ) | ( n2253 & n10100 ) | ( ~n2787 & n10100 ) ;
  assign n14178 = n14177 ^ n8319 ^ n7678 ;
  assign n14179 = n14178 ^ n12046 ^ n9616 ;
  assign n14180 = n9386 ^ n5589 ^ 1'b0 ;
  assign n14181 = n2978 & n14180 ;
  assign n14182 = n14181 ^ n13269 ^ n9331 ;
  assign n14183 = ( n5525 & n10319 ) | ( n5525 & ~n14182 ) | ( n10319 & ~n14182 ) ;
  assign n14184 = ( n751 & ~n11567 ) | ( n751 & n14183 ) | ( ~n11567 & n14183 ) ;
  assign n14185 = n14184 ^ n7171 ^ 1'b0 ;
  assign n14186 = ~n1617 & n14185 ;
  assign n14188 = ( ~n1900 & n2216 ) | ( ~n1900 & n3165 ) | ( n2216 & n3165 ) ;
  assign n14187 = ( n1467 & n3039 ) | ( n1467 & n9486 ) | ( n3039 & n9486 ) ;
  assign n14189 = n14188 ^ n14187 ^ 1'b0 ;
  assign n14190 = ~n3952 & n14189 ;
  assign n14196 = ( n2135 & n5225 ) | ( n2135 & n9132 ) | ( n5225 & n9132 ) ;
  assign n14191 = n2682 | n6586 ;
  assign n14192 = n11271 ^ n9301 ^ n5746 ;
  assign n14193 = n14192 ^ n5862 ^ n1696 ;
  assign n14194 = ( n12619 & n14191 ) | ( n12619 & n14193 ) | ( n14191 & n14193 ) ;
  assign n14195 = n10796 & n14194 ;
  assign n14197 = n14196 ^ n14195 ^ n317 ;
  assign n14198 = ( n4383 & n8292 ) | ( n4383 & n14197 ) | ( n8292 & n14197 ) ;
  assign n14199 = ( ~n5727 & n14190 ) | ( ~n5727 & n14198 ) | ( n14190 & n14198 ) ;
  assign n14200 = n7353 ^ n5649 ^ n3305 ;
  assign n14201 = n2510 ^ n130 ^ 1'b0 ;
  assign n14202 = n4375 | n14201 ;
  assign n14203 = n3244 ^ n2367 ^ n1060 ;
  assign n14204 = n11687 & n14203 ;
  assign n14205 = ~n1436 & n1976 ;
  assign n14206 = ~n5032 & n14205 ;
  assign n14207 = n14206 ^ n1404 ^ 1'b0 ;
  assign n14208 = ( n813 & ~n3621 ) | ( n813 & n12743 ) | ( ~n3621 & n12743 ) ;
  assign n14209 = n14208 ^ n291 ^ n284 ;
  assign n14210 = n14209 ^ n11984 ^ n7548 ;
  assign n14211 = n3165 & n8032 ;
  assign n14212 = ~n6760 & n14211 ;
  assign n14213 = ( ~n6399 & n14210 ) | ( ~n6399 & n14212 ) | ( n14210 & n14212 ) ;
  assign n14214 = n6454 ^ n4126 ^ n1847 ;
  assign n14215 = n13453 ^ n9019 ^ n2960 ;
  assign n14216 = n14215 ^ n1426 ^ n1136 ;
  assign n14217 = n14214 & n14216 ;
  assign n14222 = n4706 ^ n4418 ^ 1'b0 ;
  assign n14223 = n14222 ^ n2013 ^ 1'b0 ;
  assign n14224 = n10532 & ~n14223 ;
  assign n14218 = ( ~n6603 & n7891 ) | ( ~n6603 & n8995 ) | ( n7891 & n8995 ) ;
  assign n14219 = n10696 ^ n133 ^ 1'b0 ;
  assign n14220 = ~n14218 & n14219 ;
  assign n14221 = n2145 & n14220 ;
  assign n14225 = n14224 ^ n14221 ^ 1'b0 ;
  assign n14226 = ( n823 & ~n7367 ) | ( n823 & n9120 ) | ( ~n7367 & n9120 ) ;
  assign n14227 = n14226 ^ n6562 ^ n4343 ;
  assign n14228 = ( n7578 & ~n9235 ) | ( n7578 & n14227 ) | ( ~n9235 & n14227 ) ;
  assign n14229 = ~n14225 & n14228 ;
  assign n14230 = n14229 ^ n6562 ^ 1'b0 ;
  assign n14233 = n2343 ^ n1391 ^ n1109 ;
  assign n14231 = n8806 ^ n4425 ^ 1'b0 ;
  assign n14232 = ~n12968 & n14231 ;
  assign n14234 = n14233 ^ n14232 ^ n4354 ;
  assign n14235 = n5918 ^ n5044 ^ 1'b0 ;
  assign n14236 = n14235 ^ n4080 ^ 1'b0 ;
  assign n14237 = ( n3285 & ~n6443 ) | ( n3285 & n11695 ) | ( ~n6443 & n11695 ) ;
  assign n14238 = n7444 & n14237 ;
  assign n14239 = n3157 ^ n2739 ^ n1714 ;
  assign n14240 = ( n4611 & ~n13391 ) | ( n4611 & n14239 ) | ( ~n13391 & n14239 ) ;
  assign n14241 = n11204 & ~n14240 ;
  assign n14242 = ( n3723 & n10222 ) | ( n3723 & n14241 ) | ( n10222 & n14241 ) ;
  assign n14243 = ~n5181 & n7084 ;
  assign n14244 = n14243 ^ n4007 ^ 1'b0 ;
  assign n14245 = n6752 | n12356 ;
  assign n14246 = n14245 ^ n1912 ^ 1'b0 ;
  assign n14247 = ( n10183 & ~n14244 ) | ( n10183 & n14246 ) | ( ~n14244 & n14246 ) ;
  assign n14248 = n5487 ^ n1152 ^ n324 ;
  assign n14249 = n10806 ^ n4212 ^ 1'b0 ;
  assign n14250 = n1347 & ~n14249 ;
  assign n14251 = ( n5855 & ~n7685 ) | ( n5855 & n12352 ) | ( ~n7685 & n12352 ) ;
  assign n14252 = ( n11530 & n14250 ) | ( n11530 & ~n14251 ) | ( n14250 & ~n14251 ) ;
  assign n14253 = ~n889 & n1393 ;
  assign n14254 = n7194 & n14253 ;
  assign n14255 = n14254 ^ n10786 ^ n9741 ;
  assign n14256 = n2953 | n7837 ;
  assign n14257 = n14255 | n14256 ;
  assign n14258 = ( ~n4270 & n6004 ) | ( ~n4270 & n13465 ) | ( n6004 & n13465 ) ;
  assign n14259 = ( ~n2449 & n13439 ) | ( ~n2449 & n14258 ) | ( n13439 & n14258 ) ;
  assign n14260 = n3203 ^ n1796 ^ 1'b0 ;
  assign n14261 = ( n1795 & n9173 ) | ( n1795 & n9850 ) | ( n9173 & n9850 ) ;
  assign n14262 = ( n258 & n14260 ) | ( n258 & n14261 ) | ( n14260 & n14261 ) ;
  assign n14263 = ( n3285 & n4924 ) | ( n3285 & ~n10761 ) | ( n4924 & ~n10761 ) ;
  assign n14264 = n8811 ^ n650 ^ n583 ;
  assign n14265 = n13072 ^ n6135 ^ 1'b0 ;
  assign n14266 = n7233 & ~n14265 ;
  assign n14267 = n10328 ^ n9206 ^ 1'b0 ;
  assign n14268 = n14266 & n14267 ;
  assign n14269 = n14264 & n14268 ;
  assign n14270 = n14269 ^ n7414 ^ n5013 ;
  assign n14272 = ( n1263 & n4903 ) | ( n1263 & ~n10582 ) | ( n4903 & ~n10582 ) ;
  assign n14271 = n3450 ^ x34 ^ 1'b0 ;
  assign n14273 = n14272 ^ n14271 ^ n13527 ;
  assign n14274 = ~n8104 & n14273 ;
  assign n14275 = n14274 ^ n347 ^ 1'b0 ;
  assign n14276 = n1220 & n2692 ;
  assign n14277 = n773 & n14276 ;
  assign n14278 = n14277 ^ n4848 ^ n1668 ;
  assign n14279 = n4490 & ~n7372 ;
  assign n14280 = n14278 & n14279 ;
  assign n14281 = n1767 & n3068 ;
  assign n14282 = n8312 & n14281 ;
  assign n14283 = ( n3157 & ~n6098 ) | ( n3157 & n14282 ) | ( ~n6098 & n14282 ) ;
  assign n14284 = n4188 ^ n1434 ^ 1'b0 ;
  assign n14285 = n14284 ^ n7180 ^ n5481 ;
  assign n14291 = n11271 ^ n3782 ^ n1353 ;
  assign n14292 = n5174 ^ n2962 ^ n2774 ;
  assign n14293 = ~n3069 & n14292 ;
  assign n14294 = ~n14291 & n14293 ;
  assign n14286 = n2990 ^ n1945 ^ n1912 ;
  assign n14287 = n14286 ^ n12922 ^ n2455 ;
  assign n14288 = n14287 ^ n1095 ^ 1'b0 ;
  assign n14289 = n5510 & ~n14288 ;
  assign n14290 = n8021 | n14289 ;
  assign n14295 = n14294 ^ n14290 ^ n10979 ;
  assign n14296 = n6954 ^ n275 ^ 1'b0 ;
  assign n14297 = n11106 ^ n8822 ^ n921 ;
  assign n14298 = ~n6130 & n9247 ;
  assign n14299 = n9736 & n14298 ;
  assign n14300 = n14299 ^ n12577 ^ n1417 ;
  assign n14301 = ( n4465 & n11450 ) | ( n4465 & ~n14300 ) | ( n11450 & ~n14300 ) ;
  assign n14302 = ( n2120 & n14297 ) | ( n2120 & n14301 ) | ( n14297 & n14301 ) ;
  assign n14303 = n8655 ^ n1318 ^ 1'b0 ;
  assign n14304 = n6189 & ~n10784 ;
  assign n14305 = ( ~n9050 & n14303 ) | ( ~n9050 & n14304 ) | ( n14303 & n14304 ) ;
  assign n14306 = ( n2025 & ~n4659 ) | ( n2025 & n10669 ) | ( ~n4659 & n10669 ) ;
  assign n14307 = ( n2868 & n6978 ) | ( n2868 & n14306 ) | ( n6978 & n14306 ) ;
  assign n14308 = n13975 ^ n13269 ^ n7420 ;
  assign n14309 = n4651 & ~n14308 ;
  assign n14310 = n6365 & ~n10616 ;
  assign n14311 = n5108 ^ n1736 ^ n303 ;
  assign n14312 = ( ~n2070 & n4702 ) | ( ~n2070 & n14311 ) | ( n4702 & n14311 ) ;
  assign n14313 = n1193 & n14312 ;
  assign n14314 = n10759 ^ x80 ^ 1'b0 ;
  assign n14315 = ~n14313 & n14314 ;
  assign n14316 = n2973 & ~n4860 ;
  assign n14317 = n14316 ^ n1948 ^ 1'b0 ;
  assign n14319 = n7657 ^ n7290 ^ n869 ;
  assign n14318 = n13272 ^ n908 ^ 1'b0 ;
  assign n14320 = n14319 ^ n14318 ^ 1'b0 ;
  assign n14321 = ~n14317 & n14320 ;
  assign n14322 = ( n4689 & ~n6098 ) | ( n4689 & n10445 ) | ( ~n6098 & n10445 ) ;
  assign n14323 = n12010 ^ n2733 ^ n846 ;
  assign n14324 = n9883 ^ n2785 ^ 1'b0 ;
  assign n14325 = ( n387 & ~n1572 ) | ( n387 & n13166 ) | ( ~n1572 & n13166 ) ;
  assign n14326 = ( n703 & n2486 ) | ( n703 & ~n13036 ) | ( n2486 & ~n13036 ) ;
  assign n14327 = ( n6679 & n10493 ) | ( n6679 & ~n14326 ) | ( n10493 & ~n14326 ) ;
  assign n14328 = n6172 ^ n2043 ^ 1'b0 ;
  assign n14329 = n1101 | n14328 ;
  assign n14330 = n11598 & ~n14329 ;
  assign n14333 = ( ~n5490 & n6109 ) | ( ~n5490 & n7741 ) | ( n6109 & n7741 ) ;
  assign n14331 = n12944 ^ n3205 ^ n2299 ;
  assign n14332 = ( n964 & ~n7721 ) | ( n964 & n14331 ) | ( ~n7721 & n14331 ) ;
  assign n14334 = n14333 ^ n14332 ^ n3049 ;
  assign n14335 = n13585 & ~n14334 ;
  assign n14336 = ( n2078 & ~n5922 ) | ( n2078 & n6020 ) | ( ~n5922 & n6020 ) ;
  assign n14337 = n225 & ~n14336 ;
  assign n14338 = n14337 ^ n11698 ^ 1'b0 ;
  assign n14339 = n1533 & n8333 ;
  assign n14340 = n14339 ^ n3391 ^ 1'b0 ;
  assign n14341 = n14340 ^ n9087 ^ n3840 ;
  assign n14342 = n5663 ^ n1727 ^ n1282 ;
  assign n14343 = n14342 ^ n7952 ^ n6676 ;
  assign n14344 = n2120 | n7821 ;
  assign n14345 = n14344 ^ n3073 ^ 1'b0 ;
  assign n14346 = n2552 ^ n1257 ^ 1'b0 ;
  assign n14347 = n934 | n5101 ;
  assign n14348 = n11769 | n14347 ;
  assign n14349 = ( ~n7120 & n14346 ) | ( ~n7120 & n14348 ) | ( n14346 & n14348 ) ;
  assign n14350 = n13997 ^ n8998 ^ n4794 ;
  assign n14351 = ( n1822 & n3420 ) | ( n1822 & n10262 ) | ( n3420 & n10262 ) ;
  assign n14352 = n10588 ^ n8166 ^ 1'b0 ;
  assign n14353 = n11788 | n14352 ;
  assign n14354 = n4494 ^ n2778 ^ n1474 ;
  assign n14355 = ( x66 & n4913 ) | ( x66 & n14354 ) | ( n4913 & n14354 ) ;
  assign n14356 = ~n7522 & n14355 ;
  assign n14357 = n9144 ^ n3997 ^ 1'b0 ;
  assign n14358 = n8270 ^ n8085 ^ 1'b0 ;
  assign n14359 = ~n14144 & n14358 ;
  assign n14360 = ( n1012 & n7818 ) | ( n1012 & n7906 ) | ( n7818 & n7906 ) ;
  assign n14361 = n10580 ^ n2928 ^ 1'b0 ;
  assign n14362 = n14360 & ~n14361 ;
  assign n14363 = ( ~n457 & n14359 ) | ( ~n457 & n14362 ) | ( n14359 & n14362 ) ;
  assign n14364 = ( n4467 & n14357 ) | ( n4467 & n14363 ) | ( n14357 & n14363 ) ;
  assign n14365 = n6358 ^ n802 ^ 1'b0 ;
  assign n14366 = ( ~n2686 & n3870 ) | ( ~n2686 & n11236 ) | ( n3870 & n11236 ) ;
  assign n14367 = n12524 ^ n6363 ^ n4290 ;
  assign n14368 = n5213 ^ n746 ^ n594 ;
  assign n14369 = ( n3783 & n11651 ) | ( n3783 & n14368 ) | ( n11651 & n14368 ) ;
  assign n14370 = n2055 & n13434 ;
  assign n14371 = n14370 ^ n5604 ^ 1'b0 ;
  assign n14372 = n785 | n5068 ;
  assign n14373 = n2225 & ~n14372 ;
  assign n14374 = ( n8434 & ~n10031 ) | ( n8434 & n14373 ) | ( ~n10031 & n14373 ) ;
  assign n14375 = n6102 ^ n4675 ^ 1'b0 ;
  assign n14376 = ( ~n9930 & n12097 ) | ( ~n9930 & n12747 ) | ( n12097 & n12747 ) ;
  assign n14377 = n14376 ^ n10083 ^ 1'b0 ;
  assign n14380 = n164 | n8313 ;
  assign n14378 = ( n969 & ~n3630 ) | ( n969 & n12703 ) | ( ~n3630 & n12703 ) ;
  assign n14379 = ( n2132 & n14155 ) | ( n2132 & ~n14378 ) | ( n14155 & ~n14378 ) ;
  assign n14381 = n14380 ^ n14379 ^ 1'b0 ;
  assign n14382 = n9048 & n10480 ;
  assign n14383 = n6407 & n14382 ;
  assign n14384 = ~n2652 & n5266 ;
  assign n14385 = n14384 ^ n4132 ^ 1'b0 ;
  assign n14386 = ( n13057 & ~n14332 ) | ( n13057 & n14385 ) | ( ~n14332 & n14385 ) ;
  assign n14389 = ( n784 & ~n3315 ) | ( n784 & n5214 ) | ( ~n3315 & n5214 ) ;
  assign n14387 = n4657 & n9898 ;
  assign n14388 = n14387 ^ n9402 ^ 1'b0 ;
  assign n14390 = n14389 ^ n14388 ^ 1'b0 ;
  assign n14391 = ~n14386 & n14390 ;
  assign n14392 = n12139 ^ n10745 ^ n6272 ;
  assign n14393 = n14392 ^ n7715 ^ 1'b0 ;
  assign n14394 = n5311 ^ n4627 ^ 1'b0 ;
  assign n14395 = n14393 & n14394 ;
  assign n14396 = n12100 ^ n6299 ^ n5921 ;
  assign n14397 = n7341 ^ n6895 ^ x9 ;
  assign n14398 = n3147 | n5502 ;
  assign n14399 = n14397 & ~n14398 ;
  assign n14400 = n2005 | n5199 ;
  assign n14401 = n14400 ^ n9699 ^ 1'b0 ;
  assign n14402 = n2663 & ~n9364 ;
  assign n14403 = n14402 ^ n1906 ^ 1'b0 ;
  assign n14404 = n14401 & n14403 ;
  assign n14405 = n408 & n4011 ;
  assign n14406 = ~n3892 & n10351 ;
  assign n14407 = ~n14405 & n14406 ;
  assign n14408 = ( n3700 & n6953 ) | ( n3700 & ~n11174 ) | ( n6953 & ~n11174 ) ;
  assign n14409 = n4451 | n14360 ;
  assign n14410 = n11669 ^ n6555 ^ 1'b0 ;
  assign n14411 = n14409 & n14410 ;
  assign n14412 = ( n5198 & n14408 ) | ( n5198 & n14411 ) | ( n14408 & n14411 ) ;
  assign n14414 = n5087 | n9400 ;
  assign n14415 = n6900 ^ n3698 ^ 1'b0 ;
  assign n14416 = ~n13524 & n14415 ;
  assign n14417 = ( n13889 & n14414 ) | ( n13889 & ~n14416 ) | ( n14414 & ~n14416 ) ;
  assign n14413 = ~n3623 & n7463 ;
  assign n14418 = n14417 ^ n14413 ^ 1'b0 ;
  assign n14419 = n14418 ^ n6290 ^ n3812 ;
  assign n14420 = n3600 ^ n1139 ^ 1'b0 ;
  assign n14421 = ( n6368 & ~n10313 ) | ( n6368 & n14420 ) | ( ~n10313 & n14420 ) ;
  assign n14424 = ( n1306 & ~n1889 ) | ( n1306 & n4333 ) | ( ~n1889 & n4333 ) ;
  assign n14425 = n14424 ^ n8581 ^ n2504 ;
  assign n14422 = ( n3077 & n5875 ) | ( n3077 & ~n10582 ) | ( n5875 & ~n10582 ) ;
  assign n14423 = n14422 ^ n1193 ^ 1'b0 ;
  assign n14426 = n14425 ^ n14423 ^ n2578 ;
  assign n14427 = ( n1488 & ~n14421 ) | ( n1488 & n14426 ) | ( ~n14421 & n14426 ) ;
  assign n14428 = n4503 ^ x10 ^ 1'b0 ;
  assign n14429 = ~n8966 & n14428 ;
  assign n14430 = ( n6337 & n13421 ) | ( n6337 & n14429 ) | ( n13421 & n14429 ) ;
  assign n14431 = n10460 ^ n6344 ^ 1'b0 ;
  assign n14432 = n11528 | n14431 ;
  assign n14433 = ( n573 & n10702 ) | ( n573 & ~n14432 ) | ( n10702 & ~n14432 ) ;
  assign n14434 = n1343 & n2074 ;
  assign n14435 = n14434 ^ n4289 ^ 1'b0 ;
  assign n14436 = n14435 ^ n4508 ^ 1'b0 ;
  assign n14437 = n10283 | n14436 ;
  assign n14438 = n14437 ^ n4739 ^ n4319 ;
  assign n14439 = ( n8760 & ~n14424 ) | ( n8760 & n14438 ) | ( ~n14424 & n14438 ) ;
  assign n14440 = n12143 ^ n9753 ^ n7968 ;
  assign n14443 = ( n1719 & n5197 ) | ( n1719 & n6585 ) | ( n5197 & n6585 ) ;
  assign n14441 = ~n265 & n10764 ;
  assign n14442 = n3471 & n14441 ;
  assign n14444 = n14443 ^ n14442 ^ n3345 ;
  assign n14445 = n2607 | n14444 ;
  assign n14446 = n345 | n14445 ;
  assign n14452 = n5383 & n7515 ;
  assign n14453 = n14452 ^ n11080 ^ 1'b0 ;
  assign n14449 = n4910 ^ n2057 ^ 1'b0 ;
  assign n14450 = n4833 | n14449 ;
  assign n14451 = n14450 ^ n7013 ^ n4821 ;
  assign n14447 = n3101 & ~n7836 ;
  assign n14448 = ( n630 & ~n11239 ) | ( n630 & n14447 ) | ( ~n11239 & n14447 ) ;
  assign n14454 = n14453 ^ n14451 ^ n14448 ;
  assign n14455 = ( n252 & n3138 ) | ( n252 & ~n7627 ) | ( n3138 & ~n7627 ) ;
  assign n14456 = n726 | n3194 ;
  assign n14457 = n3772 & ~n14456 ;
  assign n14458 = x94 | n2605 ;
  assign n14459 = n9987 ^ n5868 ^ n3529 ;
  assign n14460 = ( n2801 & n9917 ) | ( n2801 & n14459 ) | ( n9917 & n14459 ) ;
  assign n14461 = n14460 ^ n11024 ^ 1'b0 ;
  assign n14462 = n1687 | n6607 ;
  assign n14463 = n14462 ^ n4292 ^ 1'b0 ;
  assign n14464 = ~n3392 & n7749 ;
  assign n14465 = n9093 & ~n14464 ;
  assign n14466 = ~n14463 & n14465 ;
  assign n14467 = n12903 ^ x54 ^ 1'b0 ;
  assign n14468 = n3227 & ~n14467 ;
  assign n14469 = ~n5559 & n7163 ;
  assign n14470 = n9328 & n14469 ;
  assign n14471 = n14470 ^ n9652 ^ 1'b0 ;
  assign n14472 = n9659 & n14471 ;
  assign n14473 = n2019 ^ n1845 ^ n1728 ;
  assign n14476 = ( n1472 & n3330 ) | ( n1472 & n4901 ) | ( n3330 & n4901 ) ;
  assign n14474 = n9143 ^ n2452 ^ n1252 ;
  assign n14475 = ~n8403 & n14474 ;
  assign n14477 = n14476 ^ n14475 ^ 1'b0 ;
  assign n14478 = n7367 ^ n1824 ^ 1'b0 ;
  assign n14479 = n238 & ~n14478 ;
  assign n14480 = ( ~n812 & n3544 ) | ( ~n812 & n9905 ) | ( n3544 & n9905 ) ;
  assign n14481 = ( n10234 & n14479 ) | ( n10234 & ~n14480 ) | ( n14479 & ~n14480 ) ;
  assign n14482 = n9010 ^ n4453 ^ 1'b0 ;
  assign n14483 = n9079 ^ n6508 ^ 1'b0 ;
  assign n14484 = ( n2417 & n4697 ) | ( n2417 & n5152 ) | ( n4697 & n5152 ) ;
  assign n14485 = ( n1184 & ~n3243 ) | ( n1184 & n9032 ) | ( ~n3243 & n9032 ) ;
  assign n14486 = ( n3879 & n14484 ) | ( n3879 & ~n14485 ) | ( n14484 & ~n14485 ) ;
  assign n14487 = n6835 & n14486 ;
  assign n14488 = n14487 ^ n7908 ^ n2592 ;
  assign n14489 = ( n1138 & n3848 ) | ( n1138 & n4115 ) | ( n3848 & n4115 ) ;
  assign n14490 = n14489 ^ n1655 ^ 1'b0 ;
  assign n14491 = n14490 ^ n3622 ^ 1'b0 ;
  assign n14492 = ~n478 & n14491 ;
  assign n14493 = ( n4742 & n10122 ) | ( n4742 & ~n14492 ) | ( n10122 & ~n14492 ) ;
  assign n14499 = n2235 & n8295 ;
  assign n14500 = n14499 ^ n3710 ^ 1'b0 ;
  assign n14501 = n14500 ^ n11984 ^ n1667 ;
  assign n14497 = n9803 ^ n3565 ^ n1440 ;
  assign n14496 = ~n2126 & n2473 ;
  assign n14498 = n14497 ^ n14496 ^ 1'b0 ;
  assign n14494 = n10582 & ~n10636 ;
  assign n14495 = n6690 & n14494 ;
  assign n14502 = n14501 ^ n14498 ^ n14495 ;
  assign n14503 = n5622 ^ n3384 ^ n3175 ;
  assign n14504 = ~n5223 & n6507 ;
  assign n14505 = n14504 ^ n4837 ^ 1'b0 ;
  assign n14506 = ( n6999 & n14503 ) | ( n6999 & n14505 ) | ( n14503 & n14505 ) ;
  assign n14507 = ( n2600 & ~n3111 ) | ( n2600 & n10377 ) | ( ~n3111 & n10377 ) ;
  assign n14508 = ( ~n9559 & n9728 ) | ( ~n9559 & n14507 ) | ( n9728 & n14507 ) ;
  assign n14509 = n4279 ^ n4117 ^ 1'b0 ;
  assign n14510 = ~n8343 & n14509 ;
  assign n14511 = ( n11792 & n14508 ) | ( n11792 & n14510 ) | ( n14508 & n14510 ) ;
  assign n14512 = n13772 ^ n2500 ^ 1'b0 ;
  assign n14513 = n14512 ^ n4697 ^ n3746 ;
  assign n14521 = ( ~n1129 & n2080 ) | ( ~n1129 & n2791 ) | ( n2080 & n2791 ) ;
  assign n14522 = n6181 | n11756 ;
  assign n14523 = n14521 | n14522 ;
  assign n14517 = ( n1812 & n8625 ) | ( n1812 & ~n9913 ) | ( n8625 & ~n9913 ) ;
  assign n14514 = n10441 ^ n4103 ^ 1'b0 ;
  assign n14515 = n5854 & ~n14514 ;
  assign n14516 = n14515 ^ n9455 ^ n7067 ;
  assign n14518 = n14517 ^ n14516 ^ n11275 ;
  assign n14519 = n14518 ^ n3472 ^ 1'b0 ;
  assign n14520 = ( x44 & n12048 ) | ( x44 & n14519 ) | ( n12048 & n14519 ) ;
  assign n14524 = n14523 ^ n14520 ^ n2724 ;
  assign n14525 = n14524 ^ n2622 ^ 1'b0 ;
  assign n14526 = n12455 ^ n2539 ^ 1'b0 ;
  assign n14527 = n779 | n4000 ;
  assign n14528 = n14527 ^ n1981 ^ 1'b0 ;
  assign n14529 = ~n1863 & n5329 ;
  assign n14530 = ~n8443 & n14529 ;
  assign n14531 = ( ~x34 & n14065 ) | ( ~x34 & n14530 ) | ( n14065 & n14530 ) ;
  assign n14532 = n14531 ^ n8956 ^ n7991 ;
  assign n14533 = n12646 ^ n6416 ^ n2755 ;
  assign n14534 = ~n6637 & n12118 ;
  assign n14535 = n14534 ^ n7905 ^ 1'b0 ;
  assign n14536 = n1940 | n2902 ;
  assign n14537 = n14536 ^ n3853 ^ 1'b0 ;
  assign n14538 = n14537 ^ n9904 ^ 1'b0 ;
  assign n14539 = n6447 ^ n4784 ^ 1'b0 ;
  assign n14540 = n10513 & ~n14539 ;
  assign n14541 = n14540 ^ n3190 ^ 1'b0 ;
  assign n14542 = n2835 | n14541 ;
  assign n14543 = n5276 ^ n649 ^ 1'b0 ;
  assign n14544 = n14542 | n14543 ;
  assign n14545 = n11080 ^ n7552 ^ n4242 ;
  assign n14546 = ( x28 & n14507 ) | ( x28 & ~n14545 ) | ( n14507 & ~n14545 ) ;
  assign n14547 = ( n5962 & ~n6336 ) | ( n5962 & n6555 ) | ( ~n6336 & n6555 ) ;
  assign n14548 = ( ~x55 & n9380 ) | ( ~x55 & n14547 ) | ( n9380 & n14547 ) ;
  assign n14549 = n1832 | n2899 ;
  assign n14550 = x113 & ~n3417 ;
  assign n14551 = n14550 ^ n10358 ^ 1'b0 ;
  assign n14553 = ( ~n1528 & n5935 ) | ( ~n1528 & n9871 ) | ( n5935 & n9871 ) ;
  assign n14552 = ~n5899 & n11727 ;
  assign n14554 = n14553 ^ n14552 ^ 1'b0 ;
  assign n14555 = n14554 ^ n12149 ^ n8611 ;
  assign n14556 = ( ~n14549 & n14551 ) | ( ~n14549 & n14555 ) | ( n14551 & n14555 ) ;
  assign n14557 = n1677 & ~n2550 ;
  assign n14558 = n14557 ^ n14220 ^ n9640 ;
  assign n14559 = n14558 ^ n4374 ^ x16 ;
  assign n14560 = n5865 & ~n10559 ;
  assign n14561 = n12151 & n13429 ;
  assign n14562 = ( n9258 & n14560 ) | ( n9258 & ~n14561 ) | ( n14560 & ~n14561 ) ;
  assign n14563 = n14562 ^ n13880 ^ 1'b0 ;
  assign n14568 = n2918 ^ n173 ^ 1'b0 ;
  assign n14564 = n4427 ^ n2319 ^ n335 ;
  assign n14565 = n5960 | n7743 ;
  assign n14566 = n14564 | n14565 ;
  assign n14567 = ( x108 & n1514 ) | ( x108 & ~n14566 ) | ( n1514 & ~n14566 ) ;
  assign n14569 = n14568 ^ n14567 ^ n8309 ;
  assign n14570 = ( ~n5735 & n6511 ) | ( ~n5735 & n8885 ) | ( n6511 & n8885 ) ;
  assign n14571 = n2975 & n3683 ;
  assign n14572 = n4339 & ~n14571 ;
  assign n14573 = ~n4493 & n14572 ;
  assign n14574 = n3179 & n3305 ;
  assign n14575 = n14574 ^ n14490 ^ 1'b0 ;
  assign n14576 = n14575 ^ n11810 ^ n3989 ;
  assign n14577 = n1986 | n14576 ;
  assign n14578 = n14577 ^ n2560 ^ 1'b0 ;
  assign n14579 = n11861 ^ n4683 ^ 1'b0 ;
  assign n14580 = ( n1696 & n3252 ) | ( n1696 & n12392 ) | ( n3252 & n12392 ) ;
  assign n14581 = ( n11065 & ~n12164 ) | ( n11065 & n14580 ) | ( ~n12164 & n14580 ) ;
  assign n14582 = n4778 ^ n1767 ^ n517 ;
  assign n14583 = n7568 ^ n458 ^ n226 ;
  assign n14584 = n6601 ^ n6342 ^ 1'b0 ;
  assign n14585 = ( n9966 & n14583 ) | ( n9966 & n14584 ) | ( n14583 & n14584 ) ;
  assign n14586 = n5139 ^ n2341 ^ n1663 ;
  assign n14587 = ( n7697 & n10133 ) | ( n7697 & n12108 ) | ( n10133 & n12108 ) ;
  assign n14588 = n4507 & ~n6876 ;
  assign n14589 = n14588 ^ n10971 ^ 1'b0 ;
  assign n14590 = n10210 ^ n8590 ^ n738 ;
  assign n14591 = n14590 ^ n2292 ^ 1'b0 ;
  assign n14592 = n14589 & n14591 ;
  assign n14595 = ~n1206 & n5468 ;
  assign n14593 = ~n1655 & n9359 ;
  assign n14594 = n14593 ^ n4389 ^ n1759 ;
  assign n14596 = n14595 ^ n14594 ^ n7903 ;
  assign n14597 = n14596 ^ n14297 ^ n3252 ;
  assign n14598 = n850 & n4877 ;
  assign n14599 = n4930 | n14598 ;
  assign n14602 = n4139 & n8696 ;
  assign n14603 = n3592 & n14602 ;
  assign n14600 = n7475 ^ n5581 ^ n1544 ;
  assign n14601 = n11970 | n14600 ;
  assign n14604 = n14603 ^ n14601 ^ 1'b0 ;
  assign n14605 = n4112 ^ n2978 ^ n857 ;
  assign n14606 = n2582 ^ n1616 ^ n1418 ;
  assign n14607 = n14606 ^ n4505 ^ 1'b0 ;
  assign n14608 = n13579 & n14607 ;
  assign n14609 = ( ~n10725 & n14605 ) | ( ~n10725 & n14608 ) | ( n14605 & n14608 ) ;
  assign n14615 = ~n1790 & n9769 ;
  assign n14616 = n9382 & n14615 ;
  assign n14613 = n10488 ^ n2031 ^ 1'b0 ;
  assign n14614 = n14613 ^ n1430 ^ 1'b0 ;
  assign n14610 = n4055 | n11589 ;
  assign n14611 = n14610 ^ n10339 ^ 1'b0 ;
  assign n14612 = ( n822 & n5950 ) | ( n822 & ~n14611 ) | ( n5950 & ~n14611 ) ;
  assign n14617 = n14616 ^ n14614 ^ n14612 ;
  assign n14618 = ( n613 & ~n3384 ) | ( n613 & n5289 ) | ( ~n3384 & n5289 ) ;
  assign n14619 = ( n3488 & n8313 ) | ( n3488 & n14618 ) | ( n8313 & n14618 ) ;
  assign n14620 = n9761 | n12650 ;
  assign n14621 = ( n8069 & ~n14619 ) | ( n8069 & n14620 ) | ( ~n14619 & n14620 ) ;
  assign n14622 = ( n10691 & n12096 ) | ( n10691 & n13014 ) | ( n12096 & n13014 ) ;
  assign n14623 = ( n2406 & n13844 ) | ( n2406 & ~n14622 ) | ( n13844 & ~n14622 ) ;
  assign n14624 = ( n6273 & n6975 ) | ( n6273 & n12475 ) | ( n6975 & n12475 ) ;
  assign n14626 = n3416 ^ n2656 ^ 1'b0 ;
  assign n14627 = n4405 | n14626 ;
  assign n14625 = n10251 ^ n9421 ^ 1'b0 ;
  assign n14628 = n14627 ^ n14625 ^ 1'b0 ;
  assign n14629 = n14624 & n14628 ;
  assign n14630 = n4575 & n8717 ;
  assign n14631 = n14630 ^ n9048 ^ 1'b0 ;
  assign n14632 = n3223 | n14631 ;
  assign n14633 = n10557 & ~n14632 ;
  assign n14634 = ( n213 & n9124 ) | ( n213 & n14633 ) | ( n9124 & n14633 ) ;
  assign n14635 = n11819 ^ n9644 ^ n3657 ;
  assign n14640 = n6731 ^ n4317 ^ n2108 ;
  assign n14636 = ~n3348 & n7412 ;
  assign n14637 = ~n1632 & n14636 ;
  assign n14638 = n4857 & n10116 ;
  assign n14639 = n14637 & n14638 ;
  assign n14641 = n14640 ^ n14639 ^ n8630 ;
  assign n14642 = n14641 ^ n4896 ^ 1'b0 ;
  assign n14643 = n14239 & ~n14642 ;
  assign n14644 = n4474 ^ n1652 ^ 1'b0 ;
  assign n14645 = ~n2653 & n13736 ;
  assign n14646 = n5287 & n14645 ;
  assign n14647 = ( n6181 & n14644 ) | ( n6181 & n14646 ) | ( n14644 & n14646 ) ;
  assign n14648 = n12653 & ~n14647 ;
  assign n14649 = n14648 ^ n3222 ^ 1'b0 ;
  assign n14650 = n14649 ^ n13912 ^ n6732 ;
  assign n14651 = ( ~n2206 & n9806 ) | ( ~n2206 & n10146 ) | ( n9806 & n10146 ) ;
  assign n14652 = n14651 ^ n6850 ^ 1'b0 ;
  assign n14653 = n14652 ^ n9059 ^ n5549 ;
  assign n14654 = ( n742 & n10662 ) | ( n742 & n14653 ) | ( n10662 & n14653 ) ;
  assign n14655 = ( n5967 & n9762 ) | ( n5967 & ~n14654 ) | ( n9762 & ~n14654 ) ;
  assign n14656 = ~n3737 & n7947 ;
  assign n14657 = n14656 ^ n9424 ^ n2305 ;
  assign n14658 = ( n11646 & n12096 ) | ( n11646 & n14657 ) | ( n12096 & n14657 ) ;
  assign n14663 = ( n195 & n3340 ) | ( n195 & ~n5316 ) | ( n3340 & ~n5316 ) ;
  assign n14662 = ( n7977 & ~n9729 ) | ( n7977 & n10349 ) | ( ~n9729 & n10349 ) ;
  assign n14659 = n1671 | n2448 ;
  assign n14660 = n7853 | n14659 ;
  assign n14661 = ( ~n3839 & n14451 ) | ( ~n3839 & n14660 ) | ( n14451 & n14660 ) ;
  assign n14664 = n14663 ^ n14662 ^ n14661 ;
  assign n14665 = n8376 | n11443 ;
  assign n14666 = n14664 & ~n14665 ;
  assign n14667 = n11472 ^ n5429 ^ n3223 ;
  assign n14668 = n11139 ^ n9254 ^ n4902 ;
  assign n14669 = ( n5535 & n9149 ) | ( n5535 & n14668 ) | ( n9149 & n14668 ) ;
  assign n14670 = n4740 ^ n2271 ^ 1'b0 ;
  assign n14671 = n14669 | n14670 ;
  assign n14678 = n12653 ^ n3049 ^ n542 ;
  assign n14675 = n11853 ^ n5437 ^ 1'b0 ;
  assign n14676 = ~n3025 & n14675 ;
  assign n14672 = n1405 & n2083 ;
  assign n14673 = n14672 ^ n4410 ^ 1'b0 ;
  assign n14674 = ( n789 & n7692 ) | ( n789 & n14673 ) | ( n7692 & n14673 ) ;
  assign n14677 = n14676 ^ n14674 ^ n2732 ;
  assign n14679 = n14678 ^ n14677 ^ n1914 ;
  assign n14680 = ( n8950 & n14671 ) | ( n8950 & n14679 ) | ( n14671 & n14679 ) ;
  assign n14681 = n8651 ^ n5374 ^ n582 ;
  assign n14682 = ( x37 & ~n2630 ) | ( x37 & n10916 ) | ( ~n2630 & n10916 ) ;
  assign n14683 = ( n3947 & n14671 ) | ( n3947 & ~n14682 ) | ( n14671 & ~n14682 ) ;
  assign n14684 = n11686 ^ n3345 ^ 1'b0 ;
  assign n14687 = ( ~n2329 & n3174 ) | ( ~n2329 & n4303 ) | ( n3174 & n4303 ) ;
  assign n14688 = ( n7708 & n10505 ) | ( n7708 & n14687 ) | ( n10505 & n14687 ) ;
  assign n14685 = ( n2903 & n6568 ) | ( n2903 & n8552 ) | ( n6568 & n8552 ) ;
  assign n14686 = ~n9561 & n14685 ;
  assign n14689 = n14688 ^ n14686 ^ 1'b0 ;
  assign n14690 = n3402 | n3629 ;
  assign n14691 = n14689 & ~n14690 ;
  assign n14692 = n6785 ^ n4878 ^ n4412 ;
  assign n14693 = n2224 & n14692 ;
  assign n14694 = n14693 ^ n13606 ^ 1'b0 ;
  assign n14696 = x56 & ~n3648 ;
  assign n14695 = ( n2798 & n3111 ) | ( n2798 & n11243 ) | ( n3111 & n11243 ) ;
  assign n14697 = n14696 ^ n14695 ^ n12134 ;
  assign n14698 = n11821 ^ n3396 ^ 1'b0 ;
  assign n14699 = ( ~n1704 & n3689 ) | ( ~n1704 & n12024 ) | ( n3689 & n12024 ) ;
  assign n14700 = ( n5068 & n7061 ) | ( n5068 & n11199 ) | ( n7061 & n11199 ) ;
  assign n14701 = ( n13057 & n14699 ) | ( n13057 & n14700 ) | ( n14699 & n14700 ) ;
  assign n14702 = n2575 ^ n1555 ^ 1'b0 ;
  assign n14703 = n14702 ^ n13042 ^ n3902 ;
  assign n14704 = n2853 ^ n331 ^ 1'b0 ;
  assign n14705 = ~n8059 & n14704 ;
  assign n14706 = n14705 ^ n2469 ^ 1'b0 ;
  assign n14707 = n14706 ^ n2479 ^ n742 ;
  assign n14708 = n7169 & n7809 ;
  assign n14709 = ~n1932 & n14708 ;
  assign n14710 = n4539 & ~n5444 ;
  assign n14711 = n13011 ^ n4906 ^ n1732 ;
  assign n14712 = n7375 | n8314 ;
  assign n14713 = n14712 ^ n2927 ^ 1'b0 ;
  assign n14720 = n13686 ^ n5609 ^ 1'b0 ;
  assign n14714 = ( n1379 & ~n2570 ) | ( n1379 & n7133 ) | ( ~n2570 & n7133 ) ;
  assign n14715 = ( n2113 & n7903 ) | ( n2113 & n14714 ) | ( n7903 & n14714 ) ;
  assign n14716 = ( ~n5149 & n5665 ) | ( ~n5149 & n7152 ) | ( n5665 & n7152 ) ;
  assign n14717 = ( n840 & ~n5279 ) | ( n840 & n7582 ) | ( ~n5279 & n7582 ) ;
  assign n14718 = ( n14715 & n14716 ) | ( n14715 & ~n14717 ) | ( n14716 & ~n14717 ) ;
  assign n14719 = n3247 | n14718 ;
  assign n14721 = n14720 ^ n14719 ^ 1'b0 ;
  assign n14722 = ( n14711 & ~n14713 ) | ( n14711 & n14721 ) | ( ~n14713 & n14721 ) ;
  assign n14723 = n12150 ^ n4281 ^ 1'b0 ;
  assign n14724 = n6422 | n14723 ;
  assign n14725 = n14724 ^ n12364 ^ n4148 ;
  assign n14726 = ~n7662 & n14725 ;
  assign n14727 = n1193 | n14726 ;
  assign n14728 = n11927 & n14727 ;
  assign n14729 = ( n2394 & n3698 ) | ( n2394 & ~n5132 ) | ( n3698 & ~n5132 ) ;
  assign n14730 = n3271 & ~n11292 ;
  assign n14731 = n14729 & n14730 ;
  assign n14732 = ( n6222 & ~n12552 ) | ( n6222 & n14731 ) | ( ~n12552 & n14731 ) ;
  assign n14733 = ( n3570 & ~n5793 ) | ( n3570 & n14732 ) | ( ~n5793 & n14732 ) ;
  assign n14734 = ( ~n2049 & n8028 ) | ( ~n2049 & n12314 ) | ( n8028 & n12314 ) ;
  assign n14735 = ( n2744 & n3573 ) | ( n2744 & ~n14734 ) | ( n3573 & ~n14734 ) ;
  assign n14736 = ( ~n4539 & n10445 ) | ( ~n4539 & n12060 ) | ( n10445 & n12060 ) ;
  assign n14737 = ( n4779 & ~n14735 ) | ( n4779 & n14736 ) | ( ~n14735 & n14736 ) ;
  assign n14738 = n10152 ^ n2209 ^ n1241 ;
  assign n14741 = n2528 ^ n1581 ^ 1'b0 ;
  assign n14739 = n275 | n4547 ;
  assign n14740 = n14739 ^ n622 ^ 1'b0 ;
  assign n14742 = n14741 ^ n14740 ^ n9101 ;
  assign n14743 = n10200 ^ n6610 ^ 1'b0 ;
  assign n14744 = n9466 & n14743 ;
  assign n14745 = n5074 ^ n165 ^ 1'b0 ;
  assign n14746 = ( n7976 & n11316 ) | ( n7976 & n14745 ) | ( n11316 & n14745 ) ;
  assign n14747 = ( n2188 & ~n5162 ) | ( n2188 & n10157 ) | ( ~n5162 & n10157 ) ;
  assign n14748 = n6904 ^ n3840 ^ n1904 ;
  assign n14749 = n14748 ^ n7702 ^ 1'b0 ;
  assign n14750 = ~n1354 & n14749 ;
  assign n14751 = ( ~n3790 & n10294 ) | ( ~n3790 & n14750 ) | ( n10294 & n14750 ) ;
  assign n14752 = n8519 ^ n5633 ^ n4086 ;
  assign n14753 = n11815 ^ x53 ^ 1'b0 ;
  assign n14754 = n14753 ^ n4845 ^ n2172 ;
  assign n14755 = ( n2519 & ~n14752 ) | ( n2519 & n14754 ) | ( ~n14752 & n14754 ) ;
  assign n14756 = ( n1876 & ~n4019 ) | ( n1876 & n8602 ) | ( ~n4019 & n8602 ) ;
  assign n14757 = n14756 ^ n2502 ^ n693 ;
  assign n14758 = ( n1152 & ~n14755 ) | ( n1152 & n14757 ) | ( ~n14755 & n14757 ) ;
  assign n14759 = n8391 & ~n12148 ;
  assign n14761 = ( n261 & n1121 ) | ( n261 & n10669 ) | ( n1121 & n10669 ) ;
  assign n14760 = n10497 ^ n4532 ^ n2558 ;
  assign n14762 = n14761 ^ n14760 ^ n7334 ;
  assign n14763 = n14759 & n14762 ;
  assign n14764 = ~n11916 & n14763 ;
  assign n14765 = n564 & n5132 ;
  assign n14766 = n14765 ^ x72 ^ 1'b0 ;
  assign n14767 = ( n1679 & n6198 ) | ( n1679 & ~n10760 ) | ( n6198 & ~n10760 ) ;
  assign n14768 = n1534 & n14767 ;
  assign n14769 = n14766 & n14768 ;
  assign n14770 = ~n12619 & n14769 ;
  assign n14771 = ~n3402 & n8603 ;
  assign n14772 = n14771 ^ n227 ^ 1'b0 ;
  assign n14773 = n5775 | n9397 ;
  assign n14774 = n14772 & ~n14773 ;
  assign n14775 = ( ~n1357 & n3891 ) | ( ~n1357 & n10276 ) | ( n3891 & n10276 ) ;
  assign n14779 = n6008 ^ n662 ^ 1'b0 ;
  assign n14780 = ~n2115 & n14779 ;
  assign n14781 = n860 & n14780 ;
  assign n14782 = n14781 ^ n6278 ^ 1'b0 ;
  assign n14776 = n918 & n4874 ;
  assign n14777 = n6384 & n14776 ;
  assign n14778 = n4024 & n14777 ;
  assign n14783 = n14782 ^ n14778 ^ n13751 ;
  assign n14784 = ~n14775 & n14783 ;
  assign n14786 = n3271 ^ n3138 ^ n372 ;
  assign n14787 = ~n1747 & n2483 ;
  assign n14788 = ~n14786 & n14787 ;
  assign n14785 = n7233 ^ n6714 ^ 1'b0 ;
  assign n14789 = n14788 ^ n14785 ^ n10551 ;
  assign n14790 = n2994 ^ n405 ^ 1'b0 ;
  assign n14791 = n6414 | n14790 ;
  assign n14792 = ( n1721 & n2611 ) | ( n1721 & n14791 ) | ( n2611 & n14791 ) ;
  assign n14793 = n4767 | n9325 ;
  assign n14794 = n9734 & ~n14793 ;
  assign n14795 = ( n4872 & ~n14792 ) | ( n4872 & n14794 ) | ( ~n14792 & n14794 ) ;
  assign n14796 = n2386 ^ n1635 ^ 1'b0 ;
  assign n14797 = n12881 & ~n14796 ;
  assign n14798 = ~n5078 & n14797 ;
  assign n14799 = n13333 ^ n2639 ^ 1'b0 ;
  assign n14800 = n2779 & ~n14799 ;
  assign n14801 = n13821 & n14800 ;
  assign n14802 = ~n5871 & n14801 ;
  assign n14803 = ( n2136 & n14798 ) | ( n2136 & n14802 ) | ( n14798 & n14802 ) ;
  assign n14804 = ~n13468 & n14803 ;
  assign n14805 = n14678 ^ n3782 ^ n896 ;
  assign n14806 = n14471 | n14805 ;
  assign n14807 = n14806 ^ n1194 ^ 1'b0 ;
  assign n14808 = ~n1413 & n8632 ;
  assign n14809 = n14808 ^ n12140 ^ 1'b0 ;
  assign n14810 = n494 | n3142 ;
  assign n14811 = ( ~n2439 & n14604 ) | ( ~n2439 & n14810 ) | ( n14604 & n14810 ) ;
  assign n14812 = n14486 ^ n11277 ^ 1'b0 ;
  assign n14813 = n14812 ^ n11645 ^ 1'b0 ;
  assign n14814 = n4221 | n7465 ;
  assign n14815 = n8428 | n14814 ;
  assign n14816 = ( n5556 & n12602 ) | ( n5556 & ~n14815 ) | ( n12602 & ~n14815 ) ;
  assign n14817 = ( n11470 & ~n12935 ) | ( n11470 & n14816 ) | ( ~n12935 & n14816 ) ;
  assign n14822 = n2858 | n6547 ;
  assign n14823 = n14822 ^ n914 ^ 1'b0 ;
  assign n14818 = ~n342 & n1078 ;
  assign n14819 = n14818 ^ n4762 ^ 1'b0 ;
  assign n14820 = ( ~n509 & n1146 ) | ( ~n509 & n2676 ) | ( n1146 & n2676 ) ;
  assign n14821 = ~n14819 & n14820 ;
  assign n14824 = n14823 ^ n14821 ^ n8802 ;
  assign n14825 = ( ~n6954 & n9202 ) | ( ~n6954 & n14824 ) | ( n9202 & n14824 ) ;
  assign n14827 = n6838 ^ n294 ^ 1'b0 ;
  assign n14828 = n2038 & ~n14827 ;
  assign n14829 = ~n10368 & n14828 ;
  assign n14826 = ~n8033 & n13501 ;
  assign n14830 = n14829 ^ n14826 ^ 1'b0 ;
  assign n14831 = n3683 ^ n783 ^ n746 ;
  assign n14832 = n6678 & n14831 ;
  assign n14833 = n3823 | n14832 ;
  assign n14834 = n6883 | n9248 ;
  assign n14835 = n129 | n14834 ;
  assign n14836 = n10719 | n14835 ;
  assign n14837 = n2747 & ~n12643 ;
  assign n14838 = ( ~n6716 & n6915 ) | ( ~n6716 & n8049 ) | ( n6915 & n8049 ) ;
  assign n14839 = n6466 ^ n2768 ^ 1'b0 ;
  assign n14840 = ( n373 & n14838 ) | ( n373 & ~n14839 ) | ( n14838 & ~n14839 ) ;
  assign n14841 = n14840 ^ n2809 ^ n1856 ;
  assign n14842 = ~n14558 & n14841 ;
  assign n14848 = ( n774 & n5442 ) | ( n774 & n6282 ) | ( n5442 & n6282 ) ;
  assign n14843 = ~n2363 & n3852 ;
  assign n14844 = n14843 ^ n5116 ^ 1'b0 ;
  assign n14845 = n2631 | n14844 ;
  assign n14846 = n12944 & ~n14845 ;
  assign n14847 = n14846 ^ n3241 ^ 1'b0 ;
  assign n14849 = n14848 ^ n14847 ^ n2545 ;
  assign n14850 = n14849 ^ n10056 ^ n6886 ;
  assign n14851 = ~n5559 & n14850 ;
  assign n14852 = ( n156 & n6385 ) | ( n156 & ~n12544 ) | ( n6385 & ~n12544 ) ;
  assign n14853 = n14852 ^ n5027 ^ n1561 ;
  assign n14854 = ( n1594 & n4157 ) | ( n1594 & n9800 ) | ( n4157 & n9800 ) ;
  assign n14855 = n6524 ^ n5077 ^ n3284 ;
  assign n14856 = ( n369 & n4058 ) | ( n369 & n14855 ) | ( n4058 & n14855 ) ;
  assign n14857 = ( n1982 & n14854 ) | ( n1982 & ~n14856 ) | ( n14854 & ~n14856 ) ;
  assign n14860 = n4560 ^ n4003 ^ n861 ;
  assign n14858 = ( x57 & n4905 ) | ( x57 & ~n5333 ) | ( n4905 & ~n5333 ) ;
  assign n14859 = n14858 ^ n7135 ^ n3717 ;
  assign n14861 = n14860 ^ n14859 ^ 1'b0 ;
  assign n14862 = n9769 ^ n555 ^ 1'b0 ;
  assign n14863 = ( n3759 & n11906 ) | ( n3759 & ~n14862 ) | ( n11906 & ~n14862 ) ;
  assign n14864 = ( n4607 & ~n12101 ) | ( n4607 & n13968 ) | ( ~n12101 & n13968 ) ;
  assign n14865 = ( n6743 & ~n11620 ) | ( n6743 & n12663 ) | ( ~n11620 & n12663 ) ;
  assign n14866 = n8809 | n13914 ;
  assign n14867 = n828 & ~n1290 ;
  assign n14868 = ~n9880 & n14867 ;
  assign n14869 = n5704 & n14868 ;
  assign n14870 = n14869 ^ n6622 ^ 1'b0 ;
  assign n14871 = ( ~n1931 & n6679 ) | ( ~n1931 & n9643 ) | ( n6679 & n9643 ) ;
  assign n14876 = n9549 ^ n4828 ^ 1'b0 ;
  assign n14877 = n813 & ~n14876 ;
  assign n14872 = n3932 & n14588 ;
  assign n14873 = ~n7416 & n14872 ;
  assign n14874 = n14873 ^ n923 ^ 1'b0 ;
  assign n14875 = n14874 ^ n11255 ^ 1'b0 ;
  assign n14878 = n14877 ^ n14875 ^ n7894 ;
  assign n14879 = n3899 | n14878 ;
  assign n14880 = ( n7282 & ~n7874 ) | ( n7282 & n13551 ) | ( ~n7874 & n13551 ) ;
  assign n14881 = ( n6057 & n11949 ) | ( n6057 & n14880 ) | ( n11949 & n14880 ) ;
  assign n14882 = ( n131 & n3108 ) | ( n131 & ~n7468 ) | ( n3108 & ~n7468 ) ;
  assign n14883 = ( ~n5683 & n6697 ) | ( ~n5683 & n14882 ) | ( n6697 & n14882 ) ;
  assign n14884 = n14883 ^ n9647 ^ n9238 ;
  assign n14885 = ( ~n6242 & n11086 ) | ( ~n6242 & n12312 ) | ( n11086 & n12312 ) ;
  assign n14886 = ~n2767 & n7424 ;
  assign n14887 = ( ~n8255 & n14885 ) | ( ~n8255 & n14886 ) | ( n14885 & n14886 ) ;
  assign n14888 = n1472 & n3883 ;
  assign n14889 = n13661 ^ n12770 ^ 1'b0 ;
  assign n14890 = n11966 & n14889 ;
  assign n14891 = ( n5848 & n6669 ) | ( n5848 & n12654 ) | ( n6669 & n12654 ) ;
  assign n14892 = ( n4696 & n5025 ) | ( n4696 & n14891 ) | ( n5025 & n14891 ) ;
  assign n14893 = ~n6514 & n14521 ;
  assign n14894 = n14892 & n14893 ;
  assign n14897 = n2771 ^ n1647 ^ n926 ;
  assign n14895 = n7595 ^ n3807 ^ 1'b0 ;
  assign n14896 = ~n10919 & n14895 ;
  assign n14898 = n14897 ^ n14896 ^ n3735 ;
  assign n14900 = n6572 ^ n602 ^ 1'b0 ;
  assign n14899 = n12095 ^ n9696 ^ 1'b0 ;
  assign n14901 = n14900 ^ n14899 ^ n6639 ;
  assign n14902 = ( n3536 & n4738 ) | ( n3536 & ~n11489 ) | ( n4738 & ~n11489 ) ;
  assign n14903 = ( n3508 & ~n8851 ) | ( n3508 & n14902 ) | ( ~n8851 & n14902 ) ;
  assign n14904 = ~n3351 & n14903 ;
  assign n14905 = ~n9117 & n14904 ;
  assign n14906 = n5307 ^ n3833 ^ n2338 ;
  assign n14907 = ~n5068 & n7858 ;
  assign n14908 = ( n13833 & n14750 ) | ( n13833 & ~n14907 ) | ( n14750 & ~n14907 ) ;
  assign n14909 = n14908 ^ n6691 ^ 1'b0 ;
  assign n14910 = n456 & ~n14909 ;
  assign n14911 = n4017 & n14910 ;
  assign n14912 = n14911 ^ n4349 ^ 1'b0 ;
  assign n14913 = n14912 ^ n7319 ^ 1'b0 ;
  assign n14914 = n14906 | n14913 ;
  assign n14915 = n10694 & ~n14914 ;
  assign n14916 = n14915 ^ n6133 ^ 1'b0 ;
  assign n14917 = n13905 ^ n11607 ^ n10449 ;
  assign n14918 = n2744 | n6145 ;
  assign n14919 = n14918 ^ n4314 ^ 1'b0 ;
  assign n14920 = n10696 | n14919 ;
  assign n14922 = ( n1127 & ~n3845 ) | ( n1127 & n9137 ) | ( ~n3845 & n9137 ) ;
  assign n14923 = n11373 & n14922 ;
  assign n14924 = n14923 ^ n11008 ^ 1'b0 ;
  assign n14925 = n10662 & ~n14924 ;
  assign n14921 = ~n8007 & n10073 ;
  assign n14926 = n14925 ^ n14921 ^ n7749 ;
  assign n14927 = n9647 ^ n4628 ^ n1058 ;
  assign n14928 = n7977 & n14927 ;
  assign n14929 = ~n3496 & n14928 ;
  assign n14930 = n12478 ^ n12356 ^ n2178 ;
  assign n14931 = ( n5207 & ~n11803 ) | ( n5207 & n14930 ) | ( ~n11803 & n14930 ) ;
  assign n14932 = ( n1778 & ~n11907 ) | ( n1778 & n14840 ) | ( ~n11907 & n14840 ) ;
  assign n14933 = n14932 ^ n10745 ^ 1'b0 ;
  assign n14934 = n14931 & ~n14933 ;
  assign n14935 = n409 & ~n5601 ;
  assign n14936 = n3157 & ~n6826 ;
  assign n14937 = n2034 & ~n8235 ;
  assign n14938 = ( x88 & ~n424 ) | ( x88 & n2372 ) | ( ~n424 & n2372 ) ;
  assign n14939 = ( n14936 & ~n14937 ) | ( n14936 & n14938 ) | ( ~n14937 & n14938 ) ;
  assign n14940 = n5372 & n14939 ;
  assign n14941 = ( n4259 & ~n4752 ) | ( n4259 & n11827 ) | ( ~n4752 & n11827 ) ;
  assign n14942 = n14941 ^ n3147 ^ 1'b0 ;
  assign n14943 = n14942 ^ n9805 ^ n151 ;
  assign n14949 = ~n5397 & n8853 ;
  assign n14950 = ~n1531 & n14949 ;
  assign n14944 = n1333 & ~n2713 ;
  assign n14945 = n1997 & ~n7854 ;
  assign n14946 = n14945 ^ n6898 ^ 1'b0 ;
  assign n14947 = ( n1145 & n1666 ) | ( n1145 & ~n14946 ) | ( n1666 & ~n14946 ) ;
  assign n14948 = ( n14033 & n14944 ) | ( n14033 & ~n14947 ) | ( n14944 & ~n14947 ) ;
  assign n14951 = n14950 ^ n14948 ^ 1'b0 ;
  assign n14952 = n4424 & n14951 ;
  assign n14953 = ( n11640 & n14943 ) | ( n11640 & ~n14952 ) | ( n14943 & ~n14952 ) ;
  assign n14954 = ( n1550 & n11074 ) | ( n1550 & ~n13002 ) | ( n11074 & ~n13002 ) ;
  assign n14960 = n4072 ^ n2269 ^ 1'b0 ;
  assign n14955 = n10283 ^ n2025 ^ x119 ;
  assign n14956 = n14955 ^ n3599 ^ n1220 ;
  assign n14957 = n14956 ^ n14015 ^ n1399 ;
  assign n14958 = n14957 ^ n13352 ^ 1'b0 ;
  assign n14959 = n4056 & n14958 ;
  assign n14961 = n14960 ^ n14959 ^ n10944 ;
  assign n14962 = n12340 | n14961 ;
  assign n14963 = n8694 ^ n6963 ^ 1'b0 ;
  assign n14965 = ~n414 & n715 ;
  assign n14964 = n7530 ^ n2656 ^ 1'b0 ;
  assign n14966 = n14965 ^ n14964 ^ n11903 ;
  assign n14967 = ( n2282 & ~n14963 ) | ( n2282 & n14966 ) | ( ~n14963 & n14966 ) ;
  assign n14968 = n1028 & ~n7821 ;
  assign n14969 = ( n1749 & n3408 ) | ( n1749 & n5101 ) | ( n3408 & n5101 ) ;
  assign n14970 = n14969 ^ n7959 ^ 1'b0 ;
  assign n14971 = n12888 ^ n12141 ^ n3643 ;
  assign n14973 = ( x75 & n726 ) | ( x75 & n992 ) | ( n726 & n992 ) ;
  assign n14974 = n14973 ^ n2270 ^ 1'b0 ;
  assign n14975 = n14974 ^ n6639 ^ 1'b0 ;
  assign n14972 = n5715 ^ n3889 ^ 1'b0 ;
  assign n14976 = n14975 ^ n14972 ^ n10829 ;
  assign n14977 = n1027 | n1266 ;
  assign n14978 = n13788 | n14977 ;
  assign n14979 = n13496 ^ n6216 ^ n255 ;
  assign n14980 = ( x92 & n5569 ) | ( x92 & ~n14979 ) | ( n5569 & ~n14979 ) ;
  assign n14981 = ( ~n3736 & n5443 ) | ( ~n3736 & n9227 ) | ( n5443 & n9227 ) ;
  assign n14982 = n14487 | n14981 ;
  assign n14983 = n4028 & n6172 ;
  assign n14984 = ( n4062 & n14334 ) | ( n4062 & ~n14983 ) | ( n14334 & ~n14983 ) ;
  assign n14986 = n6330 ^ n2563 ^ x102 ;
  assign n14987 = n14986 ^ n4521 ^ 1'b0 ;
  assign n14988 = n6178 | n14987 ;
  assign n14985 = n4139 & n11780 ;
  assign n14989 = n14988 ^ n14985 ^ 1'b0 ;
  assign n14991 = ( n285 & n4077 ) | ( n285 & n4784 ) | ( n4077 & n4784 ) ;
  assign n14990 = n11589 | n14418 ;
  assign n14992 = n14991 ^ n14990 ^ 1'b0 ;
  assign n14993 = n3238 ^ n2320 ^ 1'b0 ;
  assign n14994 = ~n2547 & n14993 ;
  assign n14995 = n3822 ^ n3009 ^ 1'b0 ;
  assign n14996 = n8904 & n14995 ;
  assign n14997 = n14996 ^ n9826 ^ 1'b0 ;
  assign n14998 = ( ~n2631 & n9984 ) | ( ~n2631 & n14997 ) | ( n9984 & n14997 ) ;
  assign n14999 = ( n3916 & n6432 ) | ( n3916 & ~n14998 ) | ( n6432 & ~n14998 ) ;
  assign n15000 = n8434 ^ n3524 ^ n912 ;
  assign n15001 = ~n2086 & n11868 ;
  assign n15002 = n7895 ^ n6352 ^ 1'b0 ;
  assign n15003 = n6832 & n15002 ;
  assign n15004 = ( n8416 & ~n15001 ) | ( n8416 & n15003 ) | ( ~n15001 & n15003 ) ;
  assign n15005 = n15004 ^ n9769 ^ n1764 ;
  assign n15006 = n11325 ^ n10429 ^ n578 ;
  assign n15007 = n5723 ^ n2426 ^ 1'b0 ;
  assign n15008 = n15007 ^ n6782 ^ 1'b0 ;
  assign n15009 = n2112 ^ n203 ^ 1'b0 ;
  assign n15010 = n2627 & n15009 ;
  assign n15011 = n10963 & n15010 ;
  assign n15012 = n14854 & n15011 ;
  assign n15013 = n4074 & ~n15012 ;
  assign n15014 = ~n2258 & n15013 ;
  assign n15015 = ( n8074 & ~n15008 ) | ( n8074 & n15014 ) | ( ~n15008 & n15014 ) ;
  assign n15016 = ( n2202 & ~n4387 ) | ( n2202 & n11219 ) | ( ~n4387 & n11219 ) ;
  assign n15017 = n15016 ^ n2930 ^ n2509 ;
  assign n15018 = n15017 ^ n2599 ^ 1'b0 ;
  assign n15019 = n1801 | n15018 ;
  assign n15020 = n2142 & n9443 ;
  assign n15021 = n15020 ^ n8878 ^ 1'b0 ;
  assign n15022 = n1410 & n15021 ;
  assign n15026 = n3174 & ~n3654 ;
  assign n15023 = n3951 | n10875 ;
  assign n15024 = n2747 & ~n15023 ;
  assign n15025 = n7548 | n15024 ;
  assign n15027 = n15026 ^ n15025 ^ 1'b0 ;
  assign n15029 = ( ~x44 & n10145 ) | ( ~x44 & n11496 ) | ( n10145 & n11496 ) ;
  assign n15028 = n9012 ^ n8469 ^ n144 ;
  assign n15030 = n15029 ^ n15028 ^ n10788 ;
  assign n15031 = n12001 ^ n8886 ^ n780 ;
  assign n15032 = n15031 ^ n13485 ^ n4176 ;
  assign n15036 = ( n11705 & n12700 ) | ( n11705 & n14354 ) | ( n12700 & n14354 ) ;
  assign n15037 = n15036 ^ n11785 ^ n4930 ;
  assign n15033 = n4406 | n7424 ;
  assign n15034 = n7164 | n12864 ;
  assign n15035 = n15033 & n15034 ;
  assign n15038 = n15037 ^ n15035 ^ 1'b0 ;
  assign n15043 = n3491 | n7285 ;
  assign n15039 = n8793 ^ n4642 ^ 1'b0 ;
  assign n15040 = n2851 | n15039 ;
  assign n15041 = n5826 ^ n721 ^ 1'b0 ;
  assign n15042 = n15040 | n15041 ;
  assign n15044 = n15043 ^ n15042 ^ n8677 ;
  assign n15045 = n4690 | n13258 ;
  assign n15046 = ( n3559 & n6923 ) | ( n3559 & ~n11757 ) | ( n6923 & ~n11757 ) ;
  assign n15047 = ~n5468 & n15046 ;
  assign n15048 = n3596 | n3788 ;
  assign n15049 = n5265 | n15048 ;
  assign n15050 = n15049 ^ n8676 ^ 1'b0 ;
  assign n15051 = n15050 ^ n11325 ^ n5371 ;
  assign n15052 = n11349 & n15051 ;
  assign n15053 = ( x23 & n10355 ) | ( x23 & ~n11005 ) | ( n10355 & ~n11005 ) ;
  assign n15054 = n15053 ^ n11979 ^ 1'b0 ;
  assign n15055 = n3741 ^ n2169 ^ 1'b0 ;
  assign n15056 = n1695 & n2293 ;
  assign n15057 = n15056 ^ n8654 ^ 1'b0 ;
  assign n15058 = n14335 & n15057 ;
  assign n15061 = ( x110 & n507 ) | ( x110 & ~n6555 ) | ( n507 & ~n6555 ) ;
  assign n15059 = n4800 | n5778 ;
  assign n15060 = n15059 ^ n4232 ^ 1'b0 ;
  assign n15062 = n15061 ^ n15060 ^ n5196 ;
  assign n15063 = n11623 ^ n11207 ^ 1'b0 ;
  assign n15064 = n3787 & ~n15063 ;
  assign n15065 = ~n2063 & n15064 ;
  assign n15066 = n15065 ^ n13534 ^ n4326 ;
  assign n15067 = ( n10898 & ~n11658 ) | ( n10898 & n15066 ) | ( ~n11658 & n15066 ) ;
  assign n15068 = n15062 | n15067 ;
  assign n15069 = ( ~n165 & n2900 ) | ( ~n165 & n12090 ) | ( n2900 & n12090 ) ;
  assign n15070 = n15069 ^ n11068 ^ n3304 ;
  assign n15071 = n2075 & n4657 ;
  assign n15072 = n15071 ^ n4104 ^ 1'b0 ;
  assign n15073 = n3268 & n15072 ;
  assign n15074 = n13393 ^ n1317 ^ 1'b0 ;
  assign n15075 = n12980 & ~n15074 ;
  assign n15076 = n7242 ^ n314 ^ 1'b0 ;
  assign n15077 = n5295 & n15076 ;
  assign n15078 = n5539 ^ n4677 ^ n2580 ;
  assign n15079 = n15078 ^ n14039 ^ n3261 ;
  assign n15080 = ( ~n7266 & n15077 ) | ( ~n7266 & n15079 ) | ( n15077 & n15079 ) ;
  assign n15081 = ( n3721 & n14600 ) | ( n3721 & n15080 ) | ( n14600 & n15080 ) ;
  assign n15082 = n8916 ^ n5327 ^ 1'b0 ;
  assign n15083 = n926 & ~n5865 ;
  assign n15084 = n15083 ^ n5958 ^ 1'b0 ;
  assign n15085 = ( n2322 & n4517 ) | ( n2322 & ~n5918 ) | ( n4517 & ~n5918 ) ;
  assign n15086 = n15085 ^ n10919 ^ n9267 ;
  assign n15087 = n15086 ^ n1158 ^ 1'b0 ;
  assign n15088 = n15087 ^ n2074 ^ n568 ;
  assign n15089 = ( n4189 & n15084 ) | ( n4189 & n15088 ) | ( n15084 & n15088 ) ;
  assign n15091 = n9640 ^ n6494 ^ n2517 ;
  assign n15090 = n8662 & n13371 ;
  assign n15092 = n15091 ^ n15090 ^ n497 ;
  assign n15093 = ( x68 & n3129 ) | ( x68 & n8923 ) | ( n3129 & n8923 ) ;
  assign n15097 = ( n1211 & n4545 ) | ( n1211 & n9413 ) | ( n4545 & n9413 ) ;
  assign n15094 = ( n3536 & n4748 ) | ( n3536 & n11805 ) | ( n4748 & n11805 ) ;
  assign n15095 = n12177 | n15094 ;
  assign n15096 = n2963 | n15095 ;
  assign n15098 = n15097 ^ n15096 ^ 1'b0 ;
  assign n15099 = ( n1571 & n7121 ) | ( n1571 & n8620 ) | ( n7121 & n8620 ) ;
  assign n15100 = n8315 & n15099 ;
  assign n15101 = n2596 & n3878 ;
  assign n15102 = n15101 ^ n7842 ^ n1712 ;
  assign n15103 = n2109 & ~n8394 ;
  assign n15104 = ( n1853 & ~n8698 ) | ( n1853 & n13722 ) | ( ~n8698 & n13722 ) ;
  assign n15105 = ( n5375 & n7485 ) | ( n5375 & ~n14651 ) | ( n7485 & ~n14651 ) ;
  assign n15106 = n15105 ^ n4524 ^ 1'b0 ;
  assign n15107 = ( n1262 & n6314 ) | ( n1262 & n7369 ) | ( n6314 & n7369 ) ;
  assign n15108 = ~n2033 & n2818 ;
  assign n15109 = n15108 ^ n11891 ^ 1'b0 ;
  assign n15110 = n11616 ^ n11067 ^ n2047 ;
  assign n15111 = ( n203 & ~n4320 ) | ( n203 & n14676 ) | ( ~n4320 & n14676 ) ;
  assign n15112 = n15111 ^ n4901 ^ n4720 ;
  assign n15113 = ( n5107 & n15110 ) | ( n5107 & n15112 ) | ( n15110 & n15112 ) ;
  assign n15114 = n15113 ^ n1573 ^ 1'b0 ;
  assign n15115 = ~n8789 & n15114 ;
  assign n15116 = n15115 ^ n4375 ^ 1'b0 ;
  assign n15117 = n14220 & ~n15116 ;
  assign n15118 = n10397 ^ n3553 ^ 1'b0 ;
  assign n15119 = n2953 | n15118 ;
  assign n15120 = n12918 ^ n12742 ^ n3712 ;
  assign n15121 = n2068 & ~n7117 ;
  assign n15122 = ( n7351 & n13164 ) | ( n7351 & n15121 ) | ( n13164 & n15121 ) ;
  assign n15123 = n944 | n2215 ;
  assign n15124 = n15123 ^ n5468 ^ n2796 ;
  assign n15125 = ( n5032 & n13257 ) | ( n5032 & ~n15124 ) | ( n13257 & ~n15124 ) ;
  assign n15126 = n15125 ^ n8539 ^ n1399 ;
  assign n15127 = n2097 | n13228 ;
  assign n15128 = n15127 ^ n5035 ^ 1'b0 ;
  assign n15129 = n15128 ^ n14273 ^ n3243 ;
  assign n15130 = n1871 & ~n6584 ;
  assign n15131 = n1125 | n6872 ;
  assign n15132 = n9533 ^ n6251 ^ 1'b0 ;
  assign n15133 = n9010 & ~n15132 ;
  assign n15134 = n13186 ^ n10624 ^ 1'b0 ;
  assign n15135 = ( n11906 & n15133 ) | ( n11906 & n15134 ) | ( n15133 & n15134 ) ;
  assign n15136 = ~n2654 & n13916 ;
  assign n15137 = n15136 ^ n6864 ^ 1'b0 ;
  assign n15138 = n1925 | n8080 ;
  assign n15139 = ( n1261 & n3941 ) | ( n1261 & ~n8111 ) | ( n3941 & ~n8111 ) ;
  assign n15140 = n3292 & n5521 ;
  assign n15141 = n15140 ^ n11756 ^ 1'b0 ;
  assign n15142 = ~n9787 & n15141 ;
  assign n15143 = n15142 ^ n6327 ^ 1'b0 ;
  assign n15144 = n9647 ^ n6900 ^ n1074 ;
  assign n15145 = n4986 | n6404 ;
  assign n15146 = n15144 | n15145 ;
  assign n15147 = n15146 ^ n13178 ^ 1'b0 ;
  assign n15148 = ( n9441 & ~n15143 ) | ( n9441 & n15147 ) | ( ~n15143 & n15147 ) ;
  assign n15149 = n13162 & n15148 ;
  assign n15150 = n15139 & n15149 ;
  assign n15151 = ( ~n3510 & n3754 ) | ( ~n3510 & n7575 ) | ( n3754 & n7575 ) ;
  assign n15152 = ( n6783 & ~n6797 ) | ( n6783 & n15151 ) | ( ~n6797 & n15151 ) ;
  assign n15153 = n15152 ^ n2372 ^ n831 ;
  assign n15154 = n6011 & ~n6352 ;
  assign n15155 = n15154 ^ n1108 ^ 1'b0 ;
  assign n15156 = n15155 ^ n5735 ^ n3318 ;
  assign n15157 = n15156 ^ n5701 ^ n3079 ;
  assign n15158 = n15157 ^ n5787 ^ n2759 ;
  assign n15159 = ( n273 & n1940 ) | ( n273 & ~n5962 ) | ( n1940 & ~n5962 ) ;
  assign n15160 = n15159 ^ n7567 ^ n2868 ;
  assign n15161 = ( n3640 & ~n6420 ) | ( n3640 & n6872 ) | ( ~n6420 & n6872 ) ;
  assign n15162 = ( n520 & n1997 ) | ( n520 & n2671 ) | ( n1997 & n2671 ) ;
  assign n15163 = n15162 ^ n4581 ^ 1'b0 ;
  assign n15164 = ~n4619 & n15163 ;
  assign n15169 = ~n2358 & n6404 ;
  assign n15170 = n15169 ^ n3651 ^ 1'b0 ;
  assign n15166 = n13162 ^ n4600 ^ n2166 ;
  assign n15165 = ( ~n783 & n6604 ) | ( ~n783 & n12144 ) | ( n6604 & n12144 ) ;
  assign n15167 = n15166 ^ n15165 ^ n4833 ;
  assign n15168 = n15167 ^ n3227 ^ n644 ;
  assign n15171 = n15170 ^ n15168 ^ n2439 ;
  assign n15172 = ( n7130 & n15164 ) | ( n7130 & n15171 ) | ( n15164 & n15171 ) ;
  assign n15173 = ( n10465 & ~n15161 ) | ( n10465 & n15172 ) | ( ~n15161 & n15172 ) ;
  assign n15174 = n15173 ^ n9769 ^ n3353 ;
  assign n15179 = n6430 ^ n1890 ^ 1'b0 ;
  assign n15175 = n5349 & ~n7912 ;
  assign n15176 = ~n4855 & n15175 ;
  assign n15177 = n665 | n15176 ;
  assign n15178 = n15177 ^ n3551 ^ 1'b0 ;
  assign n15180 = n15179 ^ n15178 ^ n1437 ;
  assign n15181 = n4129 ^ n2411 ^ x126 ;
  assign n15182 = n15181 ^ n4505 ^ 1'b0 ;
  assign n15183 = x65 ^ x50 ^ 1'b0 ;
  assign n15184 = ~n2124 & n15183 ;
  assign n15185 = ( n2678 & n5294 ) | ( n2678 & ~n15184 ) | ( n5294 & ~n15184 ) ;
  assign n15186 = ( ~n1929 & n6134 ) | ( ~n1929 & n8194 ) | ( n6134 & n8194 ) ;
  assign n15187 = ( n2267 & n6360 ) | ( n2267 & n6413 ) | ( n6360 & n6413 ) ;
  assign n15188 = n15187 ^ x115 ^ 1'b0 ;
  assign n15189 = n15186 | n15188 ;
  assign n15190 = n12934 ^ n7787 ^ n4223 ;
  assign n15191 = ( n641 & n1797 ) | ( n641 & ~n5562 ) | ( n1797 & ~n5562 ) ;
  assign n15192 = n15191 ^ n6175 ^ 1'b0 ;
  assign n15193 = n6992 & ~n13444 ;
  assign n15194 = n3622 & n15193 ;
  assign n15195 = n15194 ^ n4946 ^ 1'b0 ;
  assign n15196 = ~n10133 & n15195 ;
  assign n15197 = n15196 ^ n11540 ^ n642 ;
  assign n15198 = ( n6156 & n6859 ) | ( n6156 & n11362 ) | ( n6859 & n11362 ) ;
  assign n15199 = ~n1259 & n5630 ;
  assign n15200 = n15199 ^ n5589 ^ 1'b0 ;
  assign n15201 = n15200 ^ n8308 ^ n578 ;
  assign n15202 = n3991 & ~n10436 ;
  assign n15203 = ~n8921 & n15202 ;
  assign n15204 = n15203 ^ n11346 ^ n4418 ;
  assign n15205 = ( n3783 & n12361 ) | ( n3783 & n15204 ) | ( n12361 & n15204 ) ;
  assign n15206 = ( n1236 & ~n5723 ) | ( n1236 & n7230 ) | ( ~n5723 & n7230 ) ;
  assign n15207 = ( n3886 & n14487 ) | ( n3886 & ~n15206 ) | ( n14487 & ~n15206 ) ;
  assign n15211 = n11927 ^ n4650 ^ n2727 ;
  assign n15212 = n15061 & ~n15211 ;
  assign n15213 = n6357 & n15212 ;
  assign n15208 = n1575 & n1840 ;
  assign n15209 = n13352 ^ n6203 ^ 1'b0 ;
  assign n15210 = n15208 | n15209 ;
  assign n15214 = n15213 ^ n15210 ^ 1'b0 ;
  assign n15215 = n1212 & n15214 ;
  assign n15216 = n12888 ^ n4492 ^ n3973 ;
  assign n15217 = ( n5108 & ~n6148 ) | ( n5108 & n9809 ) | ( ~n6148 & n9809 ) ;
  assign n15218 = ( n6561 & ~n10689 ) | ( n6561 & n15217 ) | ( ~n10689 & n15217 ) ;
  assign n15219 = ( n4404 & n13332 ) | ( n4404 & n15218 ) | ( n13332 & n15218 ) ;
  assign n15221 = ( n1672 & n5451 ) | ( n1672 & n7601 ) | ( n5451 & n7601 ) ;
  assign n15220 = n12457 ^ n6749 ^ 1'b0 ;
  assign n15222 = n15221 ^ n15220 ^ n12263 ;
  assign n15223 = n1555 & ~n8413 ;
  assign n15224 = n9190 ^ n4330 ^ 1'b0 ;
  assign n15225 = n2261 | n15224 ;
  assign n15226 = ~n4497 & n10868 ;
  assign n15227 = n15226 ^ n3382 ^ 1'b0 ;
  assign n15228 = n3296 ^ n1741 ^ n645 ;
  assign n15229 = n15228 ^ n8696 ^ n7043 ;
  assign n15232 = ( n1532 & n4329 ) | ( n1532 & n4640 ) | ( n4329 & n4640 ) ;
  assign n15230 = ~n780 & n12161 ;
  assign n15231 = n15230 ^ n12471 ^ 1'b0 ;
  assign n15233 = n15232 ^ n15231 ^ n10002 ;
  assign n15234 = ( n6401 & n7505 ) | ( n6401 & n7854 ) | ( n7505 & n7854 ) ;
  assign n15235 = n15234 ^ n14230 ^ n13228 ;
  assign n15239 = n6056 ^ n393 ^ 1'b0 ;
  assign n15236 = n1772 & ~n8358 ;
  assign n15237 = ~n7844 & n15236 ;
  assign n15238 = n15237 ^ n13715 ^ 1'b0 ;
  assign n15240 = n15239 ^ n15238 ^ n6001 ;
  assign n15241 = n6084 ^ n1347 ^ 1'b0 ;
  assign n15242 = ~n3050 & n15241 ;
  assign n15243 = ~n10244 & n15242 ;
  assign n15244 = n7202 ^ n1363 ^ n290 ;
  assign n15245 = ~n5778 & n15244 ;
  assign n15250 = x61 & ~n5305 ;
  assign n15251 = n15250 ^ n12493 ^ n7465 ;
  assign n15246 = ( n3043 & ~n4690 ) | ( n3043 & n6184 ) | ( ~n4690 & n6184 ) ;
  assign n15247 = n15246 ^ n3034 ^ 1'b0 ;
  assign n15248 = ( ~n3769 & n7715 ) | ( ~n3769 & n15247 ) | ( n7715 & n15247 ) ;
  assign n15249 = n15248 ^ n9362 ^ n6180 ;
  assign n15252 = n15251 ^ n15249 ^ n11405 ;
  assign n15253 = n3651 & ~n11795 ;
  assign n15254 = n5424 & n15253 ;
  assign n15255 = ( n6346 & n8242 ) | ( n6346 & ~n15254 ) | ( n8242 & ~n15254 ) ;
  assign n15256 = n13094 & n15255 ;
  assign n15257 = n15256 ^ n13178 ^ n484 ;
  assign n15258 = ( n3146 & n4126 ) | ( n3146 & n4945 ) | ( n4126 & n4945 ) ;
  assign n15259 = n15258 ^ n8863 ^ n4702 ;
  assign n15261 = n5682 ^ n5407 ^ n611 ;
  assign n15260 = n7803 ^ n6033 ^ n5778 ;
  assign n15262 = n15261 ^ n15260 ^ n7475 ;
  assign n15263 = n2029 & ~n15262 ;
  assign n15264 = n13532 & n15263 ;
  assign n15265 = n737 | n15264 ;
  assign n15266 = n15259 & ~n15265 ;
  assign n15274 = n2324 ^ n1809 ^ n184 ;
  assign n15267 = ( ~n2445 & n4756 ) | ( ~n2445 & n8315 ) | ( n4756 & n8315 ) ;
  assign n15270 = n14858 ^ n1544 ^ n1376 ;
  assign n15271 = ( n1500 & ~n4752 ) | ( n1500 & n15270 ) | ( ~n4752 & n15270 ) ;
  assign n15268 = n14674 ^ n12513 ^ 1'b0 ;
  assign n15269 = ~n924 & n15268 ;
  assign n15272 = n15271 ^ n15269 ^ n212 ;
  assign n15273 = n15267 | n15272 ;
  assign n15275 = n15274 ^ n15273 ^ 1'b0 ;
  assign n15276 = ( x42 & n3872 ) | ( x42 & n4568 ) | ( n3872 & n4568 ) ;
  assign n15277 = n15276 ^ n4292 ^ 1'b0 ;
  assign n15278 = n15277 ^ n10930 ^ n2560 ;
  assign n15279 = ( n2825 & n4743 ) | ( n2825 & n15278 ) | ( n4743 & n15278 ) ;
  assign n15280 = n921 & n8704 ;
  assign n15281 = n5184 ^ n2768 ^ 1'b0 ;
  assign n15282 = n384 | n15281 ;
  assign n15283 = n6569 & ~n15282 ;
  assign n15284 = n3240 & n15283 ;
  assign n15285 = n4442 & ~n6997 ;
  assign n15286 = n15285 ^ n1277 ^ 1'b0 ;
  assign n15287 = n6937 ^ n3801 ^ 1'b0 ;
  assign n15288 = n1113 & n15287 ;
  assign n15289 = ( n771 & n7163 ) | ( n771 & ~n15288 ) | ( n7163 & ~n15288 ) ;
  assign n15290 = ~n6953 & n15289 ;
  assign n15291 = n8700 ^ n5439 ^ n2770 ;
  assign n15292 = ( n1140 & ~n10858 ) | ( n1140 & n15291 ) | ( ~n10858 & n15291 ) ;
  assign n15293 = ( ~n787 & n9407 ) | ( ~n787 & n14389 ) | ( n9407 & n14389 ) ;
  assign n15294 = n15293 ^ n4015 ^ n3631 ;
  assign n15295 = n10707 ^ n445 ^ 1'b0 ;
  assign n15296 = n589 | n15295 ;
  assign n15297 = n15296 ^ n7090 ^ n2034 ;
  assign n15298 = n1459 & ~n6434 ;
  assign n15299 = ~n10037 & n15298 ;
  assign n15300 = n2356 ^ n748 ^ 1'b0 ;
  assign n15301 = n15300 ^ n10136 ^ n5591 ;
  assign n15302 = n10872 | n15301 ;
  assign n15303 = n15228 ^ n10386 ^ 1'b0 ;
  assign n15304 = n15303 ^ n1259 ^ 1'b0 ;
  assign n15305 = ( n5421 & n12085 ) | ( n5421 & n15304 ) | ( n12085 & n15304 ) ;
  assign n15307 = n10210 ^ n3898 ^ 1'b0 ;
  assign n15306 = n10974 ^ n10595 ^ n6939 ;
  assign n15308 = n15307 ^ n15306 ^ 1'b0 ;
  assign n15309 = n2821 & n11002 ;
  assign n15310 = n15309 ^ n8855 ^ 1'b0 ;
  assign n15311 = ~n7922 & n15310 ;
  assign n15312 = ( n6328 & n9484 ) | ( n6328 & ~n15311 ) | ( n9484 & ~n15311 ) ;
  assign n15313 = n15312 ^ n14170 ^ n13148 ;
  assign n15314 = ( n197 & ~n4611 ) | ( n197 & n6401 ) | ( ~n4611 & n6401 ) ;
  assign n15315 = n15314 ^ n12754 ^ n7948 ;
  assign n15316 = ( n1966 & n3300 ) | ( n1966 & n13122 ) | ( n3300 & n13122 ) ;
  assign n15317 = n15316 ^ n443 ^ 1'b0 ;
  assign n15326 = ~n4187 & n5220 ;
  assign n15327 = ~n6760 & n15326 ;
  assign n15328 = n15327 ^ n11045 ^ n7422 ;
  assign n15321 = n15159 ^ n7287 ^ 1'b0 ;
  assign n15322 = n14930 & ~n15321 ;
  assign n15323 = n3434 ^ n3385 ^ 1'b0 ;
  assign n15324 = n15322 & ~n15323 ;
  assign n15325 = n15324 ^ n11632 ^ n10115 ;
  assign n15318 = ( n2486 & n3850 ) | ( n2486 & ~n10276 ) | ( n3850 & ~n10276 ) ;
  assign n15319 = n15318 ^ n3792 ^ n2044 ;
  assign n15320 = n13589 | n15319 ;
  assign n15329 = n15328 ^ n15325 ^ n15320 ;
  assign n15337 = n14193 ^ n2136 ^ 1'b0 ;
  assign n15338 = ~n6489 & n15337 ;
  assign n15330 = ( ~n2849 & n3095 ) | ( ~n2849 & n4626 ) | ( n3095 & n4626 ) ;
  assign n15331 = n6384 ^ x114 ^ 1'b0 ;
  assign n15332 = n15331 ^ n9089 ^ n6816 ;
  assign n15333 = n15330 | n15332 ;
  assign n15334 = n8566 & n9419 ;
  assign n15335 = n15334 ^ n10403 ^ 1'b0 ;
  assign n15336 = ( ~n5917 & n15333 ) | ( ~n5917 & n15335 ) | ( n15333 & n15335 ) ;
  assign n15339 = n15338 ^ n15336 ^ n12456 ;
  assign n15340 = n10181 ^ n5093 ^ 1'b0 ;
  assign n15341 = n12140 ^ n9688 ^ n6352 ;
  assign n15342 = n9339 | n15341 ;
  assign n15343 = n13419 ^ n10364 ^ n386 ;
  assign n15345 = ~n2776 & n5050 ;
  assign n15344 = ( n738 & ~n1466 ) | ( n738 & n9059 ) | ( ~n1466 & n9059 ) ;
  assign n15346 = n15345 ^ n15344 ^ 1'b0 ;
  assign n15347 = n5135 & n9016 ;
  assign n15348 = n15347 ^ n7505 ^ x102 ;
  assign n15349 = n13056 ^ n2940 ^ 1'b0 ;
  assign n15350 = n7052 | n10715 ;
  assign n15351 = ( n14254 & n15349 ) | ( n14254 & n15350 ) | ( n15349 & n15350 ) ;
  assign n15352 = n6325 ^ n5269 ^ n143 ;
  assign n15353 = n2910 & n15352 ;
  assign n15354 = n15351 & n15353 ;
  assign n15355 = n4004 ^ n3181 ^ 1'b0 ;
  assign n15356 = ( ~n931 & n4416 ) | ( ~n931 & n10002 ) | ( n4416 & n10002 ) ;
  assign n15357 = n15356 ^ n8544 ^ 1'b0 ;
  assign n15358 = n10942 ^ n7290 ^ 1'b0 ;
  assign n15359 = n1136 | n15358 ;
  assign n15360 = n9048 ^ n4417 ^ n1833 ;
  assign n15361 = n15359 | n15360 ;
  assign n15362 = n13906 ^ n13391 ^ n5721 ;
  assign n15363 = n15361 | n15362 ;
  assign n15364 = n11883 & n15363 ;
  assign n15365 = n15364 ^ n8261 ^ 1'b0 ;
  assign n15366 = ( n8341 & ~n15357 ) | ( n8341 & n15365 ) | ( ~n15357 & n15365 ) ;
  assign n15367 = n1575 & n2724 ;
  assign n15368 = ( n2729 & n8658 ) | ( n2729 & n15367 ) | ( n8658 & n15367 ) ;
  assign n15369 = n15368 ^ n9640 ^ n829 ;
  assign n15370 = ( n5686 & n9395 ) | ( n5686 & ~n15369 ) | ( n9395 & ~n15369 ) ;
  assign n15371 = n6149 | n15370 ;
  assign n15372 = n11614 ^ n2689 ^ n441 ;
  assign n15373 = ( n2015 & n6556 ) | ( n2015 & n11748 ) | ( n6556 & n11748 ) ;
  assign n15377 = n1394 & n2479 ;
  assign n15378 = n4944 & n13656 ;
  assign n15379 = ( n1017 & n15377 ) | ( n1017 & ~n15378 ) | ( n15377 & ~n15378 ) ;
  assign n15374 = n1632 & n7233 ;
  assign n15375 = ~n8385 & n15374 ;
  assign n15376 = n15375 ^ n4583 ^ n3133 ;
  assign n15380 = n15379 ^ n15376 ^ n5682 ;
  assign n15381 = n8470 ^ n3775 ^ 1'b0 ;
  assign n15382 = ~n7522 & n15381 ;
  assign n15383 = ( n4227 & n15380 ) | ( n4227 & ~n15382 ) | ( n15380 & ~n15382 ) ;
  assign n15384 = n3967 ^ n3366 ^ n2529 ;
  assign n15385 = n12973 | n15384 ;
  assign n15386 = n4871 & n6636 ;
  assign n15387 = ~n3271 & n15386 ;
  assign n15388 = n11430 & n12360 ;
  assign n15389 = n15387 & n15388 ;
  assign n15390 = ~n3860 & n12576 ;
  assign n15391 = n15390 ^ n4429 ^ x56 ;
  assign n15392 = n5073 | n14846 ;
  assign n15393 = n15391 & ~n15392 ;
  assign n15399 = ( ~n6471 & n13414 ) | ( ~n6471 & n13429 ) | ( n13414 & n13429 ) ;
  assign n15394 = n4102 | n13078 ;
  assign n15395 = n15394 ^ n666 ^ 1'b0 ;
  assign n15396 = ~n6388 & n15395 ;
  assign n15397 = ( x43 & ~n3297 ) | ( x43 & n15396 ) | ( ~n3297 & n15396 ) ;
  assign n15398 = ( n5556 & n8166 ) | ( n5556 & ~n15397 ) | ( n8166 & ~n15397 ) ;
  assign n15400 = n15399 ^ n15398 ^ n13123 ;
  assign n15401 = ( n6777 & ~n9123 ) | ( n6777 & n10948 ) | ( ~n9123 & n10948 ) ;
  assign n15402 = n15401 ^ n7202 ^ n1222 ;
  assign n15403 = n11427 ^ n7512 ^ n7223 ;
  assign n15404 = ( n9550 & n15053 ) | ( n9550 & ~n15403 ) | ( n15053 & ~n15403 ) ;
  assign n15410 = ~n3753 & n3960 ;
  assign n15405 = n1496 ^ x45 ^ 1'b0 ;
  assign n15407 = n11584 ^ n8917 ^ n671 ;
  assign n15406 = n4043 | n6933 ;
  assign n15408 = n15407 ^ n15406 ^ n647 ;
  assign n15409 = ( ~n4683 & n15405 ) | ( ~n4683 & n15408 ) | ( n15405 & n15408 ) ;
  assign n15411 = n15410 ^ n15409 ^ 1'b0 ;
  assign n15412 = n7103 ^ n2170 ^ n1071 ;
  assign n15413 = n334 | n15412 ;
  assign n15414 = n8988 & ~n15413 ;
  assign n15415 = n14061 ^ n8920 ^ n3985 ;
  assign n15416 = ~n2663 & n8540 ;
  assign n15417 = ~n15415 & n15416 ;
  assign n15418 = n1433 & ~n2676 ;
  assign n15419 = n10555 ^ n229 ^ x22 ;
  assign n15420 = n15327 ^ n5734 ^ n1208 ;
  assign n15421 = ( n4525 & n12576 ) | ( n4525 & ~n15420 ) | ( n12576 & ~n15420 ) ;
  assign n15422 = ( ~n15418 & n15419 ) | ( ~n15418 & n15421 ) | ( n15419 & n15421 ) ;
  assign n15423 = n9812 ^ n7130 ^ n4699 ;
  assign n15424 = n9532 ^ n6185 ^ n5562 ;
  assign n15425 = n7680 & ~n15424 ;
  assign n15426 = n15423 & n15425 ;
  assign n15427 = ( n6216 & n10778 ) | ( n6216 & ~n15426 ) | ( n10778 & ~n15426 ) ;
  assign n15428 = n1483 & n10298 ;
  assign n15429 = n15428 ^ n970 ^ 1'b0 ;
  assign n15430 = n5637 | n15429 ;
  assign n15431 = n15430 ^ n12276 ^ 1'b0 ;
  assign n15432 = n4794 ^ n1685 ^ 1'b0 ;
  assign n15433 = n1681 | n15432 ;
  assign n15434 = n163 & ~n13768 ;
  assign n15435 = n6346 | n15434 ;
  assign n15436 = ( n7135 & n15433 ) | ( n7135 & n15435 ) | ( n15433 & n15435 ) ;
  assign n15437 = n14489 ^ n11086 ^ n3630 ;
  assign n15438 = n7810 ^ n2760 ^ x80 ;
  assign n15439 = n11180 ^ n9872 ^ n7759 ;
  assign n15440 = n1638 | n12095 ;
  assign n15441 = n15439 & ~n15440 ;
  assign n15442 = n15441 ^ n10567 ^ n5213 ;
  assign n15443 = ~n4717 & n7367 ;
  assign n15444 = n15443 ^ n11012 ^ n2489 ;
  assign n15445 = n15444 ^ n14045 ^ n2043 ;
  assign n15446 = n2360 | n4988 ;
  assign n15447 = n15446 ^ n7218 ^ 1'b0 ;
  assign n15451 = ( ~n3123 & n9352 ) | ( ~n3123 & n11873 ) | ( n9352 & n11873 ) ;
  assign n15448 = n2683 & ~n3155 ;
  assign n15449 = n9167 | n14673 ;
  assign n15450 = n15448 & n15449 ;
  assign n15452 = n15451 ^ n15450 ^ 1'b0 ;
  assign n15453 = ( n1542 & n2219 ) | ( n1542 & n3050 ) | ( n2219 & n3050 ) ;
  assign n15454 = n15453 ^ n7035 ^ n4548 ;
  assign n15455 = ( ~n8097 & n9110 ) | ( ~n8097 & n15454 ) | ( n9110 & n15454 ) ;
  assign n15456 = n15452 | n15455 ;
  assign n15457 = n11111 & ~n15456 ;
  assign n15458 = n4891 ^ n4064 ^ 1'b0 ;
  assign n15459 = n4717 & ~n15458 ;
  assign n15460 = ( n1158 & n9935 ) | ( n1158 & n15459 ) | ( n9935 & n15459 ) ;
  assign n15461 = ~n5248 & n6900 ;
  assign n15462 = n15460 & n15461 ;
  assign n15463 = ~n13552 & n15462 ;
  assign n15464 = ( n1638 & ~n4932 ) | ( n1638 & n7530 ) | ( ~n4932 & n7530 ) ;
  assign n15465 = n760 & n15464 ;
  assign n15466 = ( ~n7453 & n10114 ) | ( ~n7453 & n15465 ) | ( n10114 & n15465 ) ;
  assign n15468 = n12618 ^ n4072 ^ 1'b0 ;
  assign n15469 = n15468 ^ n11486 ^ 1'b0 ;
  assign n15470 = n4148 & n15469 ;
  assign n15467 = ( n1095 & ~n5036 ) | ( n1095 & n12513 ) | ( ~n5036 & n12513 ) ;
  assign n15471 = n15470 ^ n15467 ^ 1'b0 ;
  assign n15472 = n5620 ^ n4461 ^ n3730 ;
  assign n15473 = n1514 ^ n1250 ^ n613 ;
  assign n15474 = ( n5469 & ~n13863 ) | ( n5469 & n15473 ) | ( ~n13863 & n15473 ) ;
  assign n15475 = ~n1555 & n15474 ;
  assign n15476 = n15472 & n15475 ;
  assign n15477 = n15476 ^ n1583 ^ 1'b0 ;
  assign n15478 = ~n1258 & n15477 ;
  assign n15479 = ~n3176 & n3237 ;
  assign n15480 = n4045 ^ n1462 ^ 1'b0 ;
  assign n15481 = n15479 & ~n15480 ;
  assign n15482 = n13956 ^ n11990 ^ n1554 ;
  assign n15483 = n4701 ^ n3944 ^ n2679 ;
  assign n15484 = n15483 ^ n5916 ^ n489 ;
  assign n15485 = ( n5589 & n7246 ) | ( n5589 & n12648 ) | ( n7246 & n12648 ) ;
  assign n15486 = n8475 ^ n8198 ^ n1954 ;
  assign n15487 = ( ~n913 & n11292 ) | ( ~n913 & n15486 ) | ( n11292 & n15486 ) ;
  assign n15488 = n1734 | n15487 ;
  assign n15489 = n15485 | n15488 ;
  assign n15490 = ( n4584 & ~n15484 ) | ( n4584 & n15489 ) | ( ~n15484 & n15489 ) ;
  assign n15491 = ( ~n1203 & n14555 ) | ( ~n1203 & n14627 ) | ( n14555 & n14627 ) ;
  assign n15492 = n7168 | n10049 ;
  assign n15493 = ( ~n2592 & n6142 ) | ( ~n2592 & n6881 ) | ( n6142 & n6881 ) ;
  assign n15494 = n6250 & n15493 ;
  assign n15495 = n6869 & n15494 ;
  assign n15496 = n15495 ^ n9317 ^ n6394 ;
  assign n15500 = n6975 ^ n4918 ^ n2753 ;
  assign n15497 = n7913 ^ n1228 ^ 1'b0 ;
  assign n15498 = n5317 & ~n15497 ;
  assign n15499 = n10963 & n15498 ;
  assign n15501 = n15500 ^ n15499 ^ 1'b0 ;
  assign n15502 = ( n11552 & n15496 ) | ( n11552 & ~n15501 ) | ( n15496 & ~n15501 ) ;
  assign n15503 = n7922 | n14306 ;
  assign n15504 = n15503 ^ n13886 ^ 1'b0 ;
  assign n15505 = n13277 & n15504 ;
  assign n15506 = n15502 & n15505 ;
  assign n15511 = n2175 ^ n969 ^ n664 ;
  assign n15512 = n15511 ^ n3736 ^ n3382 ;
  assign n15513 = ( n5285 & n8019 ) | ( n5285 & n15512 ) | ( n8019 & n15512 ) ;
  assign n15507 = ( n2091 & n4043 ) | ( n2091 & n15140 ) | ( n4043 & n15140 ) ;
  assign n15508 = ( n5982 & ~n12075 ) | ( n5982 & n15507 ) | ( ~n12075 & n15507 ) ;
  assign n15509 = n15228 | n15508 ;
  assign n15510 = n11412 & ~n15509 ;
  assign n15514 = n15513 ^ n15510 ^ 1'b0 ;
  assign n15515 = ( n9790 & ~n11047 ) | ( n9790 & n11414 ) | ( ~n11047 & n11414 ) ;
  assign n15516 = n15515 ^ n4105 ^ 1'b0 ;
  assign n15517 = ( n2434 & ~n5063 ) | ( n2434 & n6173 ) | ( ~n5063 & n6173 ) ;
  assign n15521 = n8986 ^ n3209 ^ n909 ;
  assign n15519 = n8033 ^ n2154 ^ 1'b0 ;
  assign n15520 = n11584 | n15519 ;
  assign n15522 = n15521 ^ n15520 ^ n9682 ;
  assign n15523 = n7141 & n11060 ;
  assign n15524 = n15522 & n15523 ;
  assign n15518 = n273 & ~n3703 ;
  assign n15525 = n15524 ^ n15518 ^ 1'b0 ;
  assign n15526 = ~n3469 & n15525 ;
  assign n15527 = n15526 ^ n1793 ^ 1'b0 ;
  assign n15528 = n14233 ^ x21 ^ 1'b0 ;
  assign n15529 = n15528 ^ n6697 ^ n4825 ;
  assign n15530 = n8020 | n11154 ;
  assign n15531 = n15529 & ~n15530 ;
  assign n15532 = n6218 ^ n4798 ^ n1492 ;
  assign n15533 = n15532 ^ n7515 ^ n169 ;
  assign n15534 = ( ~n1362 & n12089 ) | ( ~n1362 & n15533 ) | ( n12089 & n15533 ) ;
  assign n15535 = x12 & ~n12063 ;
  assign n15536 = ~n2500 & n15535 ;
  assign n15540 = n12967 ^ n6987 ^ 1'b0 ;
  assign n15541 = n6721 & ~n15540 ;
  assign n15542 = ( n10312 & n11345 ) | ( n10312 & ~n15541 ) | ( n11345 & ~n15541 ) ;
  assign n15537 = n10333 ^ n7567 ^ n1288 ;
  assign n15538 = n8291 ^ n4294 ^ n2038 ;
  assign n15539 = ( n1748 & ~n15537 ) | ( n1748 & n15538 ) | ( ~n15537 & n15538 ) ;
  assign n15543 = n15542 ^ n15539 ^ n7595 ;
  assign n15544 = n7268 ^ n3860 ^ 1'b0 ;
  assign n15545 = n15544 ^ n2349 ^ 1'b0 ;
  assign n15546 = n15543 & n15545 ;
  assign n15547 = n13707 ^ n6813 ^ n6530 ;
  assign n15548 = n252 | n6446 ;
  assign n15549 = n737 & ~n15548 ;
  assign n15550 = ( n900 & ~n3925 ) | ( n900 & n15549 ) | ( ~n3925 & n15549 ) ;
  assign n15551 = ( n3574 & n13716 ) | ( n3574 & n15550 ) | ( n13716 & n15550 ) ;
  assign n15552 = n4278 ^ n2775 ^ n2423 ;
  assign n15553 = n8446 & ~n15552 ;
  assign n15555 = n9730 ^ n8384 ^ n2613 ;
  assign n15554 = n4790 ^ n3708 ^ n3043 ;
  assign n15556 = n15555 ^ n15554 ^ 1'b0 ;
  assign n15557 = ~n15553 & n15556 ;
  assign n15558 = n9249 & n14022 ;
  assign n15559 = n663 & ~n4984 ;
  assign n15560 = n15559 ^ n10696 ^ n7514 ;
  assign n15561 = n15560 ^ n4721 ^ n2805 ;
  assign n15562 = ( n9504 & n10459 ) | ( n9504 & ~n11508 ) | ( n10459 & ~n11508 ) ;
  assign n15563 = ( ~n2934 & n4879 ) | ( ~n2934 & n8781 ) | ( n4879 & n8781 ) ;
  assign n15565 = n12346 ^ n6072 ^ n4641 ;
  assign n15566 = n15565 ^ n9952 ^ 1'b0 ;
  assign n15567 = ~n7702 & n15566 ;
  assign n15564 = ( ~n926 & n5125 ) | ( ~n926 & n14226 ) | ( n5125 & n14226 ) ;
  assign n15568 = n15567 ^ n15564 ^ n8915 ;
  assign n15569 = n15563 & ~n15568 ;
  assign n15570 = ( n1883 & n3285 ) | ( n1883 & ~n6396 ) | ( n3285 & ~n6396 ) ;
  assign n15571 = n2059 ^ n1455 ^ 1'b0 ;
  assign n15572 = n15571 ^ n7756 ^ n2280 ;
  assign n15573 = ( n4247 & n8934 ) | ( n4247 & n15572 ) | ( n8934 & n15572 ) ;
  assign n15574 = ( n1797 & ~n15570 ) | ( n1797 & n15573 ) | ( ~n15570 & n15573 ) ;
  assign n15575 = ~n3470 & n15574 ;
  assign n15576 = n8531 ^ n3543 ^ n810 ;
  assign n15577 = n15576 ^ n4612 ^ 1'b0 ;
  assign n15578 = n14098 ^ n9619 ^ n5756 ;
  assign n15579 = n15578 ^ n5281 ^ 1'b0 ;
  assign n15580 = n15579 ^ n11325 ^ 1'b0 ;
  assign n15581 = ~n2816 & n9617 ;
  assign n15582 = n4195 ^ n2234 ^ 1'b0 ;
  assign n15583 = x106 & n15582 ;
  assign n15584 = n15583 ^ n5409 ^ n5359 ;
  assign n15585 = n15584 ^ n11276 ^ 1'b0 ;
  assign n15586 = ( n1341 & n15581 ) | ( n1341 & ~n15585 ) | ( n15581 & ~n15585 ) ;
  assign n15587 = n5626 | n9116 ;
  assign n15588 = n15587 ^ n860 ^ 1'b0 ;
  assign n15589 = n9064 | n15588 ;
  assign n15590 = ( ~n3920 & n3959 ) | ( ~n3920 & n15589 ) | ( n3959 & n15589 ) ;
  assign n15591 = n6375 ^ n3462 ^ 1'b0 ;
  assign n15592 = ~n10311 & n15591 ;
  assign n15594 = ~n1223 & n8758 ;
  assign n15595 = n2672 & n15594 ;
  assign n15593 = n2925 ^ n2839 ^ 1'b0 ;
  assign n15596 = n15595 ^ n15593 ^ 1'b0 ;
  assign n15597 = n6514 | n15596 ;
  assign n15598 = ( n1873 & n2289 ) | ( n1873 & ~n9506 ) | ( n2289 & ~n9506 ) ;
  assign n15599 = n11796 & n11970 ;
  assign n15600 = ~n13404 & n15599 ;
  assign n15601 = ( n7427 & n11448 ) | ( n7427 & ~n15600 ) | ( n11448 & ~n15600 ) ;
  assign n15602 = n15601 ^ n1459 ^ n841 ;
  assign n15603 = n15550 ^ n2251 ^ 1'b0 ;
  assign n15604 = n15603 ^ n4083 ^ n2164 ;
  assign n15605 = ( n10592 & n12057 ) | ( n10592 & n15604 ) | ( n12057 & n15604 ) ;
  assign n15607 = n15565 ^ n471 ^ 1'b0 ;
  assign n15606 = ( n397 & n2743 ) | ( n397 & n15571 ) | ( n2743 & n15571 ) ;
  assign n15608 = n15607 ^ n15606 ^ 1'b0 ;
  assign n15609 = ( n1723 & ~n7595 ) | ( n1723 & n13342 ) | ( ~n7595 & n13342 ) ;
  assign n15610 = n5464 ^ n1562 ^ n899 ;
  assign n15611 = ( x100 & n7160 ) | ( x100 & ~n15610 ) | ( n7160 & ~n15610 ) ;
  assign n15612 = n10101 ^ n8299 ^ n2423 ;
  assign n15613 = ( n1003 & n1582 ) | ( n1003 & ~n7634 ) | ( n1582 & ~n7634 ) ;
  assign n15614 = ~n12198 & n15613 ;
  assign n15615 = n15614 ^ n7178 ^ 1'b0 ;
  assign n15616 = n15612 & ~n15615 ;
  assign n15617 = n7667 ^ n6156 ^ n5279 ;
  assign n15618 = n15617 ^ n14575 ^ n8485 ;
  assign n15619 = n7284 ^ n2788 ^ 1'b0 ;
  assign n15620 = ~n3688 & n15619 ;
  assign n15621 = n2923 ^ n726 ^ n558 ;
  assign n15623 = ( n4915 & n10825 ) | ( n4915 & ~n11270 ) | ( n10825 & ~n11270 ) ;
  assign n15624 = ~n3199 & n4352 ;
  assign n15625 = n15623 & n15624 ;
  assign n15626 = n15625 ^ n3505 ^ n1755 ;
  assign n15622 = n10537 & n15420 ;
  assign n15627 = n15626 ^ n15622 ^ n8742 ;
  assign n15628 = n762 & n1024 ;
  assign n15629 = ( n347 & n3449 ) | ( n347 & n15628 ) | ( n3449 & n15628 ) ;
  assign n15633 = ( n2185 & n3789 ) | ( n2185 & n9676 ) | ( n3789 & n9676 ) ;
  assign n15632 = n7583 ^ n1428 ^ 1'b0 ;
  assign n15634 = n15633 ^ n15632 ^ n8057 ;
  assign n15635 = ( n172 & ~n8177 ) | ( n172 & n15634 ) | ( ~n8177 & n15634 ) ;
  assign n15630 = n5331 | n11010 ;
  assign n15631 = n15630 ^ n223 ^ 1'b0 ;
  assign n15636 = n15635 ^ n15631 ^ n14197 ;
  assign n15637 = n2792 | n11814 ;
  assign n15638 = n3623 & ~n15637 ;
  assign n15639 = ~n5872 & n12171 ;
  assign n15640 = n7198 & n15639 ;
  assign n15641 = ( n9880 & n12227 ) | ( n9880 & ~n15640 ) | ( n12227 & ~n15640 ) ;
  assign n15642 = ~n1323 & n1480 ;
  assign n15643 = n15641 & n15642 ;
  assign n15644 = ( ~n11047 & n15638 ) | ( ~n11047 & n15643 ) | ( n15638 & n15643 ) ;
  assign n15645 = n15644 ^ n14460 ^ n567 ;
  assign n15647 = n14936 ^ n6561 ^ n5462 ;
  assign n15646 = ( n715 & n1235 ) | ( n715 & ~n3100 ) | ( n1235 & ~n3100 ) ;
  assign n15648 = n15647 ^ n15646 ^ n12342 ;
  assign n15649 = n10585 ^ n1864 ^ 1'b0 ;
  assign n15650 = n1418 & ~n15649 ;
  assign n15651 = ( n204 & n2431 ) | ( n204 & ~n4469 ) | ( n2431 & ~n4469 ) ;
  assign n15652 = n1809 & n15651 ;
  assign n15653 = n2097 & n2942 ;
  assign n15654 = n7494 ^ n755 ^ 1'b0 ;
  assign n15655 = ~n15653 & n15654 ;
  assign n15656 = ( n4907 & n7268 ) | ( n4907 & n15655 ) | ( n7268 & n15655 ) ;
  assign n15657 = n7199 ^ n3666 ^ n991 ;
  assign n15659 = n858 | n4804 ;
  assign n15658 = ~n7881 & n8650 ;
  assign n15660 = n15659 ^ n15658 ^ 1'b0 ;
  assign n15661 = n15660 ^ n8572 ^ 1'b0 ;
  assign n15662 = ~n6236 & n15661 ;
  assign n15663 = ( n1560 & n15657 ) | ( n1560 & n15662 ) | ( n15657 & n15662 ) ;
  assign n15665 = x105 & n8577 ;
  assign n15666 = n10116 ^ n9782 ^ 1'b0 ;
  assign n15667 = n15665 & n15666 ;
  assign n15664 = n10523 | n11830 ;
  assign n15668 = n15667 ^ n15664 ^ n4367 ;
  assign n15669 = n7702 ^ n5560 ^ n4939 ;
  assign n15670 = n3016 | n15669 ;
  assign n15671 = n3043 & ~n15670 ;
  assign n15672 = n3701 & n11244 ;
  assign n15673 = n15671 & n15672 ;
  assign n15676 = n8753 ^ n5516 ^ 1'b0 ;
  assign n15675 = n770 & ~n1283 ;
  assign n15677 = n15676 ^ n15675 ^ 1'b0 ;
  assign n15678 = ( x60 & ~n8581 ) | ( x60 & n15677 ) | ( ~n8581 & n15677 ) ;
  assign n15674 = ( n1155 & ~n1265 ) | ( n1155 & n2796 ) | ( ~n1265 & n2796 ) ;
  assign n15679 = n15678 ^ n15674 ^ n13109 ;
  assign n15680 = n13063 ^ n7000 ^ 1'b0 ;
  assign n15681 = n8385 & ~n15680 ;
  assign n15682 = ( n4902 & n14669 ) | ( n4902 & n15681 ) | ( n14669 & n15681 ) ;
  assign n15683 = n5284 ^ x71 ^ 1'b0 ;
  assign n15684 = n6648 | n15683 ;
  assign n15685 = n15684 ^ n9446 ^ 1'b0 ;
  assign n15686 = n11148 | n15685 ;
  assign n15687 = n5356 & ~n15686 ;
  assign n15689 = n2450 & n2891 ;
  assign n15690 = n6073 & n15689 ;
  assign n15691 = n15690 ^ n1917 ^ n1652 ;
  assign n15688 = ~n3784 & n6201 ;
  assign n15692 = n15691 ^ n15688 ^ 1'b0 ;
  assign n15693 = n8929 ^ n8211 ^ 1'b0 ;
  assign n15694 = n5754 & ~n15693 ;
  assign n15695 = n15694 ^ n11635 ^ n3473 ;
  assign n15700 = ~n5438 & n12632 ;
  assign n15701 = ~n14025 & n15700 ;
  assign n15702 = n15701 ^ n8124 ^ n647 ;
  assign n15696 = n12932 ^ n8035 ^ n1708 ;
  assign n15697 = n2572 ^ n2036 ^ 1'b0 ;
  assign n15698 = ( n459 & n9689 ) | ( n459 & n15697 ) | ( n9689 & n15697 ) ;
  assign n15699 = n15696 | n15698 ;
  assign n15703 = n15702 ^ n15699 ^ n10866 ;
  assign n15704 = n6034 & ~n15703 ;
  assign n15705 = n15704 ^ n2455 ^ 1'b0 ;
  assign n15707 = ( n1688 & n2712 ) | ( n1688 & ~n7421 ) | ( n2712 & ~n7421 ) ;
  assign n15708 = ( ~n9558 & n13297 ) | ( ~n9558 & n15707 ) | ( n13297 & n15707 ) ;
  assign n15706 = n3008 & ~n12407 ;
  assign n15709 = n15708 ^ n15706 ^ 1'b0 ;
  assign n15711 = ( n5655 & ~n8295 ) | ( n5655 & n10070 ) | ( ~n8295 & n10070 ) ;
  assign n15710 = ( n1377 & ~n2159 ) | ( n1377 & n8220 ) | ( ~n2159 & n8220 ) ;
  assign n15712 = n15711 ^ n15710 ^ n5232 ;
  assign n15713 = n6939 & n12311 ;
  assign n15714 = n675 ^ n650 ^ 1'b0 ;
  assign n15715 = n7066 & n15714 ;
  assign n15723 = ( ~n581 & n6736 ) | ( ~n581 & n9725 ) | ( n6736 & n9725 ) ;
  assign n15716 = n2488 ^ n690 ^ n655 ;
  assign n15717 = n11957 ^ n3083 ^ 1'b0 ;
  assign n15718 = n1580 & n3544 ;
  assign n15719 = ~n1424 & n15718 ;
  assign n15720 = n15719 ^ n1619 ^ n525 ;
  assign n15721 = ( ~n15716 & n15717 ) | ( ~n15716 & n15720 ) | ( n15717 & n15720 ) ;
  assign n15722 = ( n6341 & n14027 ) | ( n6341 & n15721 ) | ( n14027 & n15721 ) ;
  assign n15724 = n15723 ^ n15722 ^ n5827 ;
  assign n15730 = n10185 ^ n9478 ^ 1'b0 ;
  assign n15731 = n15730 ^ n3257 ^ 1'b0 ;
  assign n15728 = n8839 ^ n8514 ^ n3525 ;
  assign n15729 = ( n6927 & ~n7350 ) | ( n6927 & n15728 ) | ( ~n7350 & n15728 ) ;
  assign n15725 = n7086 ^ n1952 ^ n436 ;
  assign n15726 = n15725 ^ n8156 ^ n1829 ;
  assign n15727 = n15726 ^ n15112 ^ n5786 ;
  assign n15732 = n15731 ^ n15729 ^ n15727 ;
  assign n15733 = n6759 ^ n1924 ^ 1'b0 ;
  assign n15734 = n1342 | n15733 ;
  assign n15735 = n15734 ^ n1301 ^ 1'b0 ;
  assign n15736 = n15735 ^ x116 ^ 1'b0 ;
  assign n15737 = n15736 ^ n472 ^ 1'b0 ;
  assign n15739 = n2055 & n4713 ;
  assign n15740 = n15739 ^ n12506 ^ 1'b0 ;
  assign n15738 = n3397 & n9572 ;
  assign n15741 = n15740 ^ n15738 ^ 1'b0 ;
  assign n15742 = ~n196 & n15741 ;
  assign n15743 = n5596 & n15742 ;
  assign n15744 = ( ~n359 & n2246 ) | ( ~n359 & n5753 ) | ( n2246 & n5753 ) ;
  assign n15745 = n15744 ^ n3885 ^ 1'b0 ;
  assign n15746 = n14101 & ~n15745 ;
  assign n15747 = n15746 ^ n3510 ^ n397 ;
  assign n15748 = n7630 ^ n6820 ^ 1'b0 ;
  assign n15749 = ~n15396 & n15748 ;
  assign n15750 = n15749 ^ n6569 ^ 1'b0 ;
  assign n15751 = ~n10772 & n15750 ;
  assign n15752 = ( n2968 & ~n9439 ) | ( n2968 & n15186 ) | ( ~n9439 & n15186 ) ;
  assign n15753 = n15752 ^ n4717 ^ n3063 ;
  assign n15754 = ( ~n4601 & n10083 ) | ( ~n4601 & n14964 ) | ( n10083 & n14964 ) ;
  assign n15755 = n15754 ^ n5949 ^ n2222 ;
  assign n15756 = ~n8442 & n15755 ;
  assign n15759 = n13593 ^ n4348 ^ n2038 ;
  assign n15757 = n10264 ^ n9966 ^ 1'b0 ;
  assign n15758 = n14129 & ~n15757 ;
  assign n15760 = n15759 ^ n15758 ^ 1'b0 ;
  assign n15761 = n14215 ^ n8509 ^ n6750 ;
  assign n15762 = n2142 & n15761 ;
  assign n15763 = ~n15016 & n15660 ;
  assign n15764 = n13246 & n15763 ;
  assign n15765 = ( n482 & ~n9073 ) | ( n482 & n9392 ) | ( ~n9073 & n9392 ) ;
  assign n15769 = n1376 | n2772 ;
  assign n15770 = ( n616 & ~n2559 ) | ( n616 & n11120 ) | ( ~n2559 & n11120 ) ;
  assign n15771 = n15770 ^ n2937 ^ n2896 ;
  assign n15772 = ( n4893 & ~n15769 ) | ( n4893 & n15771 ) | ( ~n15769 & n15771 ) ;
  assign n15773 = ( n2915 & n7161 ) | ( n2915 & ~n15772 ) | ( n7161 & ~n15772 ) ;
  assign n15766 = n7700 ^ n3775 ^ n1843 ;
  assign n15767 = n6072 & ~n8633 ;
  assign n15768 = n15766 & n15767 ;
  assign n15774 = n15773 ^ n15768 ^ 1'b0 ;
  assign n15775 = ~n15765 & n15774 ;
  assign n15776 = ( n1981 & n2105 ) | ( n1981 & ~n4792 ) | ( n2105 & ~n4792 ) ;
  assign n15777 = n1571 & n1820 ;
  assign n15778 = n15777 ^ n8705 ^ n2580 ;
  assign n15779 = ~n15776 & n15778 ;
  assign n15780 = ( ~n1557 & n11789 ) | ( ~n1557 & n14906 ) | ( n11789 & n14906 ) ;
  assign n15789 = ~n6837 & n7117 ;
  assign n15790 = n3391 & ~n15789 ;
  assign n15791 = n2526 & n15790 ;
  assign n15784 = n14854 ^ n7471 ^ n7216 ;
  assign n15785 = ( ~n3524 & n15633 ) | ( ~n3524 & n15784 ) | ( n15633 & n15784 ) ;
  assign n15782 = ~n1579 & n3786 ;
  assign n15783 = n15782 ^ n11234 ^ 1'b0 ;
  assign n15786 = n15785 ^ n15783 ^ n8040 ;
  assign n15787 = ( n2394 & n8728 ) | ( n2394 & n15786 ) | ( n8728 & n15786 ) ;
  assign n15781 = n4789 & n8946 ;
  assign n15788 = n15787 ^ n15781 ^ 1'b0 ;
  assign n15792 = n15791 ^ n15788 ^ n13688 ;
  assign n15793 = ~n10049 & n11465 ;
  assign n15794 = ~n1763 & n15793 ;
  assign n15795 = n5530 & n15046 ;
  assign n15796 = n15794 & n15795 ;
  assign n15797 = n10778 ^ n1071 ^ 1'b0 ;
  assign n15798 = n322 & ~n15797 ;
  assign n15799 = ~n8642 & n15798 ;
  assign n15803 = ( n913 & ~n4234 ) | ( n913 & n11579 ) | ( ~n4234 & n11579 ) ;
  assign n15800 = n4600 & n4651 ;
  assign n15801 = n15800 ^ n13462 ^ 1'b0 ;
  assign n15802 = ( n2103 & ~n6812 ) | ( n2103 & n15801 ) | ( ~n6812 & n15801 ) ;
  assign n15804 = n15803 ^ n15802 ^ n13342 ;
  assign n15805 = ( n2842 & n3902 ) | ( n2842 & n14100 ) | ( n3902 & n14100 ) ;
  assign n15806 = ( x8 & n5053 ) | ( x8 & n5681 ) | ( n5053 & n5681 ) ;
  assign n15807 = n15806 ^ n5496 ^ 1'b0 ;
  assign n15808 = n15805 & ~n15807 ;
  assign n15809 = ( n2234 & n15804 ) | ( n2234 & n15808 ) | ( n15804 & n15808 ) ;
  assign n15810 = n15809 ^ x104 ^ 1'b0 ;
  assign n15811 = ( n3133 & ~n5218 ) | ( n3133 & n10995 ) | ( ~n5218 & n10995 ) ;
  assign n15812 = n10358 & ~n13217 ;
  assign n15813 = ~n15811 & n15812 ;
  assign n15816 = n7913 ^ n2703 ^ n844 ;
  assign n15817 = n3558 & ~n15816 ;
  assign n15814 = n2935 & ~n5156 ;
  assign n15815 = n15814 ^ n8651 ^ 1'b0 ;
  assign n15818 = n15817 ^ n15815 ^ n974 ;
  assign n15819 = ( n260 & n5586 ) | ( n260 & n15818 ) | ( n5586 & n15818 ) ;
  assign n15820 = n10534 & ~n15819 ;
  assign n15821 = n15813 & n15820 ;
  assign n15822 = n8160 & ~n10199 ;
  assign n15823 = n15822 ^ n7090 ^ 1'b0 ;
  assign n15824 = n4030 ^ n1695 ^ 1'b0 ;
  assign n15825 = n342 | n2724 ;
  assign n15826 = ~n15824 & n15825 ;
  assign n15827 = n15826 ^ n6466 ^ 1'b0 ;
  assign n15828 = n15827 ^ n1912 ^ 1'b0 ;
  assign n15829 = n3941 | n15828 ;
  assign n15830 = n12700 ^ n5582 ^ n541 ;
  assign n15831 = n15830 ^ n10691 ^ 1'b0 ;
  assign n15832 = ( n15823 & n15829 ) | ( n15823 & ~n15831 ) | ( n15829 & ~n15831 ) ;
  assign n15833 = n3926 ^ n1138 ^ 1'b0 ;
  assign n15834 = n14471 ^ n4828 ^ 1'b0 ;
  assign n15835 = ( n1912 & ~n2172 ) | ( n1912 & n4974 ) | ( ~n2172 & n4974 ) ;
  assign n15836 = ( n5796 & ~n7113 ) | ( n5796 & n14420 ) | ( ~n7113 & n14420 ) ;
  assign n15837 = ( n488 & n2408 ) | ( n488 & ~n15836 ) | ( n2408 & ~n15836 ) ;
  assign n15843 = ~n2837 & n8015 ;
  assign n15838 = n2059 | n11882 ;
  assign n15839 = n15838 ^ n2770 ^ 1'b0 ;
  assign n15840 = n15839 ^ n5397 ^ n650 ;
  assign n15841 = n2998 & ~n15840 ;
  assign n15842 = n15841 ^ n14798 ^ 1'b0 ;
  assign n15844 = n15843 ^ n15842 ^ n5993 ;
  assign n15846 = ( n3751 & ~n5195 ) | ( n3751 & n7497 ) | ( ~n5195 & n7497 ) ;
  assign n15847 = n15846 ^ n6874 ^ n6494 ;
  assign n15845 = ( n1635 & ~n2136 ) | ( n1635 & n8128 ) | ( ~n2136 & n8128 ) ;
  assign n15848 = n15847 ^ n15845 ^ n6692 ;
  assign n15849 = n1159 | n11406 ;
  assign n15850 = n5041 | n15849 ;
  assign n15851 = n9098 & n15850 ;
  assign n15852 = n15851 ^ n7944 ^ 1'b0 ;
  assign n15853 = ~n5162 & n7977 ;
  assign n15854 = n15853 ^ n5181 ^ 1'b0 ;
  assign n15855 = n9052 ^ n8359 ^ 1'b0 ;
  assign n15856 = n15854 & n15855 ;
  assign n15857 = n6027 ^ n460 ^ 1'b0 ;
  assign n15858 = n15857 ^ n7906 ^ n4798 ;
  assign n15859 = ( n13863 & ~n15856 ) | ( n13863 & n15858 ) | ( ~n15856 & n15858 ) ;
  assign n15860 = n15859 ^ n7330 ^ n3675 ;
  assign n15861 = ( n4873 & n11405 ) | ( n4873 & n14688 ) | ( n11405 & n14688 ) ;
  assign n15862 = n15861 ^ n13184 ^ 1'b0 ;
  assign n15863 = ~n2922 & n11227 ;
  assign n15864 = ~n3158 & n15863 ;
  assign n15865 = ( n4693 & n14266 ) | ( n4693 & n15864 ) | ( n14266 & n15864 ) ;
  assign n15866 = ( n11344 & n11597 ) | ( n11344 & n15865 ) | ( n11597 & n15865 ) ;
  assign n15867 = n5604 | n15866 ;
  assign n15868 = ( ~n4544 & n4817 ) | ( ~n4544 & n8152 ) | ( n4817 & n8152 ) ;
  assign n15869 = n11794 ^ n1246 ^ 1'b0 ;
  assign n15870 = ( n5672 & n14038 ) | ( n5672 & n15869 ) | ( n14038 & n15869 ) ;
  assign n15871 = ~n2085 & n4487 ;
  assign n15872 = n15870 & n15871 ;
  assign n15873 = n1201 & ~n3506 ;
  assign n15874 = n15873 ^ n12693 ^ n8853 ;
  assign n15875 = x102 & n4884 ;
  assign n15876 = ~n2660 & n15875 ;
  assign n15877 = n15874 | n15876 ;
  assign n15878 = ( n11496 & n13797 ) | ( n11496 & n15877 ) | ( n13797 & n15877 ) ;
  assign n15879 = ( ~n3592 & n6337 ) | ( ~n3592 & n9367 ) | ( n6337 & n9367 ) ;
  assign n15880 = ( ~n6543 & n12360 ) | ( ~n6543 & n15879 ) | ( n12360 & n15879 ) ;
  assign n15881 = n15880 ^ n15495 ^ n13593 ;
  assign n15882 = n5868 | n7230 ;
  assign n15883 = n1954 & ~n15882 ;
  assign n15884 = n15883 ^ n705 ^ 1'b0 ;
  assign n15885 = ( n1136 & ~n1138 ) | ( n1136 & n1818 ) | ( ~n1138 & n1818 ) ;
  assign n15886 = n11894 ^ n4083 ^ n359 ;
  assign n15887 = n9632 & ~n15886 ;
  assign n15888 = n15885 & n15887 ;
  assign n15889 = n3533 & ~n15888 ;
  assign n15890 = n15889 ^ n12830 ^ 1'b0 ;
  assign n15891 = n14024 & ~n15890 ;
  assign n15892 = n9070 & n15891 ;
  assign n15893 = ( ~n1907 & n4322 ) | ( ~n1907 & n6352 ) | ( n4322 & n6352 ) ;
  assign n15894 = ( n1901 & n6971 ) | ( n1901 & ~n14271 ) | ( n6971 & ~n14271 ) ;
  assign n15895 = n15893 | n15894 ;
  assign n15896 = ( ~n543 & n1003 ) | ( ~n543 & n7829 ) | ( n1003 & n7829 ) ;
  assign n15897 = n15896 ^ n12798 ^ n10575 ;
  assign n15898 = n15801 ^ n3019 ^ 1'b0 ;
  assign n15899 = ( n2944 & ~n14070 ) | ( n2944 & n15898 ) | ( ~n14070 & n15898 ) ;
  assign n15900 = n205 & ~n713 ;
  assign n15901 = ( ~n6611 & n10522 ) | ( ~n6611 & n15900 ) | ( n10522 & n15900 ) ;
  assign n15902 = n2942 & n15901 ;
  assign n15906 = n2412 & n2839 ;
  assign n15907 = n15906 ^ n587 ^ 1'b0 ;
  assign n15908 = n15907 ^ n7984 ^ n2894 ;
  assign n15903 = n13832 ^ n12316 ^ n760 ;
  assign n15904 = ~n8033 & n11616 ;
  assign n15905 = n15903 & n15904 ;
  assign n15909 = n15908 ^ n15905 ^ n11105 ;
  assign n15910 = n15909 ^ n4408 ^ 1'b0 ;
  assign n15911 = ~n9347 & n15910 ;
  assign n15912 = ~n12695 & n15911 ;
  assign n15913 = n15912 ^ n596 ^ 1'b0 ;
  assign n15914 = ( n1745 & n2267 ) | ( n1745 & n4292 ) | ( n2267 & n4292 ) ;
  assign n15915 = ~n6243 & n15914 ;
  assign n15916 = ~n6956 & n12517 ;
  assign n15917 = ~n1908 & n15916 ;
  assign n15918 = ( n2663 & n3888 ) | ( n2663 & n15917 ) | ( n3888 & n15917 ) ;
  assign n15919 = n1422 & ~n11584 ;
  assign n15920 = n4010 & n15919 ;
  assign n15921 = n15920 ^ n14923 ^ 1'b0 ;
  assign n15922 = n3959 ^ n245 ^ 1'b0 ;
  assign n15923 = n3456 & ~n3988 ;
  assign n15924 = n6996 ^ n5189 ^ 1'b0 ;
  assign n15928 = n2729 ^ n1293 ^ n510 ;
  assign n15929 = n12903 ^ n4732 ^ 1'b0 ;
  assign n15930 = n15928 | n15929 ;
  assign n15926 = ~n2788 & n6088 ;
  assign n15927 = n15926 ^ n15121 ^ n1142 ;
  assign n15925 = n10946 ^ n10713 ^ n2436 ;
  assign n15931 = n15930 ^ n15927 ^ n15925 ;
  assign n15932 = ( n1725 & ~n8885 ) | ( n1725 & n12548 ) | ( ~n8885 & n12548 ) ;
  assign n15933 = n8037 ^ x0 ^ 1'b0 ;
  assign n15934 = ( n6738 & n7348 ) | ( n6738 & n15933 ) | ( n7348 & n15933 ) ;
  assign n15935 = ( n3356 & ~n4227 ) | ( n3356 & n15934 ) | ( ~n4227 & n15934 ) ;
  assign n15936 = ( n13746 & n15932 ) | ( n13746 & ~n15935 ) | ( n15932 & ~n15935 ) ;
  assign n15937 = n8254 ^ n626 ^ 1'b0 ;
  assign n15938 = n10820 ^ n5269 ^ n2863 ;
  assign n15939 = n10302 | n15938 ;
  assign n15940 = n15939 ^ n8534 ^ 1'b0 ;
  assign n15941 = ( ~n9176 & n10034 ) | ( ~n9176 & n15940 ) | ( n10034 & n15940 ) ;
  assign n15942 = n3490 & n8667 ;
  assign n15943 = n10266 ^ n7383 ^ n6700 ;
  assign n15944 = n15435 ^ n4303 ^ 1'b0 ;
  assign n15945 = n15839 & ~n15944 ;
  assign n15946 = n15945 ^ n7270 ^ 1'b0 ;
  assign n15947 = n1594 & n15659 ;
  assign n15948 = n3014 | n15947 ;
  assign n15949 = n15948 ^ n15777 ^ n7545 ;
  assign n15950 = ( n1096 & ~n4257 ) | ( n1096 & n15949 ) | ( ~n4257 & n15949 ) ;
  assign n15951 = n11023 ^ n640 ^ 1'b0 ;
  assign n15952 = n15950 & ~n15951 ;
  assign n15953 = ( n508 & ~n1680 ) | ( n508 & n3456 ) | ( ~n1680 & n3456 ) ;
  assign n15954 = n14735 & ~n15953 ;
  assign n15959 = n4575 ^ n1665 ^ 1'b0 ;
  assign n15960 = ( n11883 & n13381 ) | ( n11883 & ~n15959 ) | ( n13381 & ~n15959 ) ;
  assign n15961 = n9363 & ~n15960 ;
  assign n15962 = n15961 ^ n1027 ^ 1'b0 ;
  assign n15958 = ( n2650 & ~n4064 ) | ( n2650 & n11837 ) | ( ~n4064 & n11837 ) ;
  assign n15963 = n15962 ^ n15958 ^ 1'b0 ;
  assign n15956 = n13941 ^ n7986 ^ 1'b0 ;
  assign n15957 = n4819 & n15956 ;
  assign n15955 = ( n1912 & n2579 ) | ( n1912 & ~n12911 ) | ( n2579 & ~n12911 ) ;
  assign n15964 = n15963 ^ n15957 ^ n15955 ;
  assign n15965 = n15964 ^ n6578 ^ 1'b0 ;
  assign n15966 = n15843 & n15965 ;
  assign n15967 = ( n1404 & ~n3783 ) | ( n1404 & n10727 ) | ( ~n3783 & n10727 ) ;
  assign n15968 = n11234 ^ n6064 ^ 1'b0 ;
  assign n15969 = ~n10104 & n15968 ;
  assign n15970 = ( n7644 & n9034 ) | ( n7644 & ~n15969 ) | ( n9034 & ~n15969 ) ;
  assign n15971 = n15970 ^ n5942 ^ 1'b0 ;
  assign n15972 = ~n287 & n15971 ;
  assign n15973 = n15972 ^ n5898 ^ n3191 ;
  assign n15974 = ~n4831 & n4964 ;
  assign n15975 = ~n6233 & n15974 ;
  assign n15976 = x123 | n15975 ;
  assign n15977 = ~n1899 & n10718 ;
  assign n15978 = n15977 ^ n5714 ^ 1'b0 ;
  assign n15979 = n15978 ^ n4214 ^ 1'b0 ;
  assign n15982 = n3111 ^ n1172 ^ n880 ;
  assign n15980 = ( n3809 & n5507 ) | ( n3809 & ~n9173 ) | ( n5507 & ~n9173 ) ;
  assign n15981 = n15980 ^ n15351 ^ 1'b0 ;
  assign n15983 = n15982 ^ n15981 ^ n11982 ;
  assign n15984 = n4386 | n15983 ;
  assign n15985 = n15979 & ~n15984 ;
  assign n15986 = n7568 ^ n170 ^ 1'b0 ;
  assign n15988 = ( n1445 & n3654 ) | ( n1445 & n7644 ) | ( n3654 & n7644 ) ;
  assign n15989 = n15988 ^ n10448 ^ n6522 ;
  assign n15990 = ( n3966 & ~n4320 ) | ( n3966 & n15989 ) | ( ~n4320 & n15989 ) ;
  assign n15987 = ~n1927 & n11346 ;
  assign n15991 = n15990 ^ n15987 ^ 1'b0 ;
  assign n15992 = n15986 & ~n15991 ;
  assign n15993 = n4290 ^ n2295 ^ n312 ;
  assign n15994 = n9093 & ~n15908 ;
  assign n15995 = n15994 ^ n14125 ^ 1'b0 ;
  assign n15996 = ( ~n8764 & n15993 ) | ( ~n8764 & n15995 ) | ( n15993 & n15995 ) ;
  assign n15997 = n7189 ^ n1914 ^ 1'b0 ;
  assign n15998 = n15997 ^ n3336 ^ 1'b0 ;
  assign n15999 = n6534 | n14817 ;
  assign n16000 = n15999 ^ n2265 ^ 1'b0 ;
  assign n16001 = ( n2800 & ~n10028 ) | ( n2800 & n16000 ) | ( ~n10028 & n16000 ) ;
  assign n16002 = n8248 & n13729 ;
  assign n16003 = n16002 ^ n15026 ^ 1'b0 ;
  assign n16004 = n16003 ^ n14755 ^ 1'b0 ;
  assign n16005 = ( n3744 & n9674 ) | ( n3744 & ~n12257 ) | ( n9674 & ~n12257 ) ;
  assign n16006 = ( ~n9528 & n11935 ) | ( ~n9528 & n16005 ) | ( n11935 & n16005 ) ;
  assign n16007 = ( n1441 & n6253 ) | ( n1441 & n11079 ) | ( n6253 & n11079 ) ;
  assign n16008 = n13133 ^ n12502 ^ n6215 ;
  assign n16009 = n16008 ^ n5581 ^ 1'b0 ;
  assign n16010 = ~n16007 & n16009 ;
  assign n16011 = ~n706 & n5013 ;
  assign n16012 = n3220 & n16011 ;
  assign n16013 = ( n894 & n2790 ) | ( n894 & ~n16012 ) | ( n2790 & ~n16012 ) ;
  assign n16014 = n4392 ^ n2550 ^ n2113 ;
  assign n16015 = n8990 ^ n7994 ^ n3843 ;
  assign n16016 = n3380 | n15433 ;
  assign n16017 = n16016 ^ n8475 ^ 1'b0 ;
  assign n16018 = ( n16014 & n16015 ) | ( n16014 & n16017 ) | ( n16015 & n16017 ) ;
  assign n16019 = ~x91 & n1761 ;
  assign n16020 = n4606 ^ n702 ^ n131 ;
  assign n16021 = ( n3076 & ~n9451 ) | ( n3076 & n16020 ) | ( ~n9451 & n16020 ) ;
  assign n16022 = ( n3913 & n16019 ) | ( n3913 & n16021 ) | ( n16019 & n16021 ) ;
  assign n16023 = ( n619 & n3991 ) | ( n619 & n9848 ) | ( n3991 & n9848 ) ;
  assign n16024 = ( n2803 & n10784 ) | ( n2803 & ~n16023 ) | ( n10784 & ~n16023 ) ;
  assign n16025 = n16024 ^ n6785 ^ 1'b0 ;
  assign n16026 = n8102 ^ n3564 ^ 1'b0 ;
  assign n16027 = n395 & ~n16026 ;
  assign n16028 = n16027 ^ n11328 ^ 1'b0 ;
  assign n16031 = n15387 ^ n2724 ^ 1'b0 ;
  assign n16029 = n8319 | n12111 ;
  assign n16030 = n16029 ^ n7236 ^ 1'b0 ;
  assign n16032 = n16031 ^ n16030 ^ n4864 ;
  assign n16033 = n11671 ^ n1529 ^ 1'b0 ;
  assign n16034 = n16033 ^ n11909 ^ n1146 ;
  assign n16035 = n10419 ^ n1162 ^ 1'b0 ;
  assign n16036 = n7882 | n16035 ;
  assign n16037 = n7492 | n11012 ;
  assign n16038 = n9522 & ~n16037 ;
  assign n16039 = ( ~n8777 & n12008 ) | ( ~n8777 & n16038 ) | ( n12008 & n16038 ) ;
  assign n16040 = n16039 ^ n7421 ^ 1'b0 ;
  assign n16042 = ( ~n5470 & n7936 ) | ( ~n5470 & n8333 ) | ( n7936 & n8333 ) ;
  assign n16041 = n1361 & n5986 ;
  assign n16043 = n16042 ^ n16041 ^ n15882 ;
  assign n16051 = ~n5563 & n13872 ;
  assign n16052 = ~n6184 & n16051 ;
  assign n16044 = n1626 & n6756 ;
  assign n16045 = n7892 & n16044 ;
  assign n16046 = n16045 ^ n2642 ^ 1'b0 ;
  assign n16047 = n15804 | n16046 ;
  assign n16048 = n16047 ^ n4458 ^ 1'b0 ;
  assign n16049 = n16048 ^ n14086 ^ 1'b0 ;
  assign n16050 = n3309 | n16049 ;
  assign n16053 = n16052 ^ n16050 ^ n12513 ;
  assign n16054 = ~n12314 & n15356 ;
  assign n16055 = n16054 ^ x95 ^ 1'b0 ;
  assign n16056 = n16055 ^ n9561 ^ n319 ;
  assign n16057 = n16056 ^ n13596 ^ n5599 ;
  assign n16058 = n15698 ^ n5310 ^ n3905 ;
  assign n16059 = n6773 ^ n6153 ^ n5277 ;
  assign n16060 = n2910 & ~n3117 ;
  assign n16064 = n8442 & ~n9968 ;
  assign n16065 = n16064 ^ n13219 ^ 1'b0 ;
  assign n16061 = ~n4291 & n13190 ;
  assign n16062 = n16061 ^ n15740 ^ 1'b0 ;
  assign n16063 = ( ~n1613 & n1931 ) | ( ~n1613 & n16062 ) | ( n1931 & n16062 ) ;
  assign n16066 = n16065 ^ n16063 ^ n2832 ;
  assign n16067 = n16060 & n16066 ;
  assign n16068 = n16059 & n16067 ;
  assign n16070 = ( ~n862 & n4562 ) | ( ~n862 & n7240 ) | ( n4562 & n7240 ) ;
  assign n16071 = ( ~n11325 & n15007 ) | ( ~n11325 & n16070 ) | ( n15007 & n16070 ) ;
  assign n16069 = n5678 ^ n5123 ^ n3421 ;
  assign n16072 = n16071 ^ n16069 ^ 1'b0 ;
  assign n16073 = n9850 | n12215 ;
  assign n16074 = ~n423 & n1242 ;
  assign n16075 = ( n487 & n9883 ) | ( n487 & n16074 ) | ( n9883 & n16074 ) ;
  assign n16076 = n13991 ^ n12990 ^ n10421 ;
  assign n16077 = n6768 | n9247 ;
  assign n16078 = n13455 ^ n464 ^ 1'b0 ;
  assign n16079 = n15372 ^ n14897 ^ 1'b0 ;
  assign n16080 = ~n9004 & n16079 ;
  assign n16081 = n9363 ^ n623 ^ 1'b0 ;
  assign n16082 = n665 | n16081 ;
  assign n16083 = n4694 | n16082 ;
  assign n16084 = n16083 ^ n10297 ^ 1'b0 ;
  assign n16085 = n10791 ^ n5949 ^ 1'b0 ;
  assign n16086 = n2298 | n3450 ;
  assign n16087 = n16086 ^ n6898 ^ n2020 ;
  assign n16088 = n16087 ^ n7330 ^ n3353 ;
  assign n16089 = n9705 & n10468 ;
  assign n16090 = n6684 ^ n2340 ^ n2154 ;
  assign n16091 = n5127 ^ n680 ^ 1'b0 ;
  assign n16092 = n6929 ^ n4721 ^ 1'b0 ;
  assign n16093 = n16091 & ~n16092 ;
  assign n16094 = n1362 & ~n14209 ;
  assign n16095 = x115 & n8279 ;
  assign n16096 = n16095 ^ n9467 ^ 1'b0 ;
  assign n16097 = ( n677 & n3467 ) | ( n677 & n16096 ) | ( n3467 & n16096 ) ;
  assign n16098 = n12912 ^ n6742 ^ n6125 ;
  assign n16099 = ( n1976 & n4861 ) | ( n1976 & n11722 ) | ( n4861 & n11722 ) ;
  assign n16100 = ( n10758 & n16098 ) | ( n10758 & ~n16099 ) | ( n16098 & ~n16099 ) ;
  assign n16101 = n835 | n2212 ;
  assign n16102 = n14194 | n16101 ;
  assign n16103 = ( n7063 & ~n15587 ) | ( n7063 & n16102 ) | ( ~n15587 & n16102 ) ;
  assign n16104 = ~n11421 & n16103 ;
  assign n16105 = n16104 ^ n14357 ^ 1'b0 ;
  assign n16106 = n3122 | n11498 ;
  assign n16107 = n7226 & n9442 ;
  assign n16108 = ~n16106 & n16107 ;
  assign n16109 = n5150 | n9394 ;
  assign n16110 = n5035 & ~n16109 ;
  assign n16111 = n8155 | n16110 ;
  assign n16112 = n6469 & ~n16111 ;
  assign n16113 = n16112 ^ n9521 ^ 1'b0 ;
  assign n16114 = n10973 ^ n332 ^ 1'b0 ;
  assign n16115 = ( ~n2219 & n4017 ) | ( ~n2219 & n4202 ) | ( n4017 & n4202 ) ;
  assign n16118 = ~n4474 & n11799 ;
  assign n16116 = ( n1409 & ~n6082 ) | ( n1409 & n12315 ) | ( ~n6082 & n12315 ) ;
  assign n16117 = n9887 & ~n16116 ;
  assign n16119 = n16118 ^ n16117 ^ 1'b0 ;
  assign n16120 = n16119 ^ n7714 ^ n6594 ;
  assign n16121 = ( n16114 & n16115 ) | ( n16114 & ~n16120 ) | ( n16115 & ~n16120 ) ;
  assign n16124 = ( ~n4992 & n6084 ) | ( ~n4992 & n13217 ) | ( n6084 & n13217 ) ;
  assign n16125 = ( n3286 & ~n4801 ) | ( n3286 & n16124 ) | ( ~n4801 & n16124 ) ;
  assign n16122 = n2385 & ~n5248 ;
  assign n16123 = n1085 & n16122 ;
  assign n16126 = n16125 ^ n16123 ^ n7175 ;
  assign n16127 = ( n9244 & n14564 ) | ( n9244 & n16126 ) | ( n14564 & n16126 ) ;
  assign n16128 = n16127 ^ n14745 ^ n6240 ;
  assign n16129 = ~n15005 & n16128 ;
  assign n16130 = n14084 ^ n9405 ^ 1'b0 ;
  assign n16131 = n7743 ^ n4634 ^ n1739 ;
  assign n16132 = n12757 & n16131 ;
  assign n16133 = n3344 & ~n7878 ;
  assign n16136 = n5259 ^ n2359 ^ 1'b0 ;
  assign n16134 = ( ~n7661 & n14443 ) | ( ~n7661 & n14944 ) | ( n14443 & n14944 ) ;
  assign n16135 = n5241 & ~n16134 ;
  assign n16137 = n16136 ^ n16135 ^ 1'b0 ;
  assign n16138 = n13642 & ~n16137 ;
  assign n16139 = ( ~n4342 & n5241 ) | ( ~n4342 & n9039 ) | ( n5241 & n9039 ) ;
  assign n16140 = n16139 ^ n2129 ^ n459 ;
  assign n16141 = n16140 ^ n7950 ^ n3132 ;
  assign n16142 = n2652 | n7364 ;
  assign n16143 = n14627 & ~n16142 ;
  assign n16144 = ( n4607 & n13784 ) | ( n4607 & n16143 ) | ( n13784 & n16143 ) ;
  assign n16145 = n6656 & n9721 ;
  assign n16146 = n6464 & n16145 ;
  assign n16151 = ( n3211 & n5518 ) | ( n3211 & ~n10714 ) | ( n5518 & ~n10714 ) ;
  assign n16148 = n4464 ^ n4008 ^ n852 ;
  assign n16149 = n16148 ^ n6983 ^ 1'b0 ;
  assign n16150 = ~n3975 & n16149 ;
  assign n16152 = n16151 ^ n16150 ^ n8846 ;
  assign n16147 = n11731 ^ n1496 ^ n416 ;
  assign n16153 = n16152 ^ n16147 ^ n4394 ;
  assign n16154 = n2426 & n4990 ;
  assign n16155 = n16154 ^ n7163 ^ 1'b0 ;
  assign n16156 = ( x10 & n568 ) | ( x10 & ~n993 ) | ( n568 & ~n993 ) ;
  assign n16157 = ( n395 & n6601 ) | ( n395 & ~n16156 ) | ( n6601 & ~n16156 ) ;
  assign n16158 = n1987 | n16157 ;
  assign n16159 = n16158 ^ n371 ^ 1'b0 ;
  assign n16160 = n16159 ^ n175 ^ x71 ;
  assign n16161 = ( ~n1910 & n16155 ) | ( ~n1910 & n16160 ) | ( n16155 & n16160 ) ;
  assign n16162 = ( n2506 & ~n7644 ) | ( n2506 & n10125 ) | ( ~n7644 & n10125 ) ;
  assign n16168 = n370 | n8827 ;
  assign n16163 = n581 ^ n397 ^ n275 ;
  assign n16164 = ( n5142 & n7494 ) | ( n5142 & ~n16163 ) | ( n7494 & ~n16163 ) ;
  assign n16165 = ( n1040 & ~n1268 ) | ( n1040 & n16164 ) | ( ~n1268 & n16164 ) ;
  assign n16166 = ( n6745 & ~n14726 ) | ( n6745 & n16165 ) | ( ~n14726 & n16165 ) ;
  assign n16167 = n1628 | n16166 ;
  assign n16169 = n16168 ^ n16167 ^ 1'b0 ;
  assign n16170 = ~n1908 & n11515 ;
  assign n16171 = ( n410 & n9451 ) | ( n410 & ~n16170 ) | ( n9451 & ~n16170 ) ;
  assign n16172 = n16048 ^ n13465 ^ n1460 ;
  assign n16177 = n10229 | n13572 ;
  assign n16173 = n8466 ^ n5028 ^ n649 ;
  assign n16174 = n16173 ^ n7256 ^ n6004 ;
  assign n16175 = n16174 ^ n11917 ^ 1'b0 ;
  assign n16176 = n5919 | n16175 ;
  assign n16178 = n16177 ^ n16176 ^ 1'b0 ;
  assign n16179 = n13038 ^ n8629 ^ n3725 ;
  assign n16180 = n2586 & ~n13072 ;
  assign n16181 = n13206 ^ n690 ^ 1'b0 ;
  assign n16182 = n13639 & ~n16181 ;
  assign n16183 = n9395 ^ n4775 ^ n1177 ;
  assign n16184 = n15708 ^ n7842 ^ n3132 ;
  assign n16185 = ( n4102 & n4756 ) | ( n4102 & n16184 ) | ( n4756 & n16184 ) ;
  assign n16187 = ( n2992 & n3327 ) | ( n2992 & ~n6051 ) | ( n3327 & ~n6051 ) ;
  assign n16188 = n7254 ^ n4685 ^ n778 ;
  assign n16189 = n10324 | n16188 ;
  assign n16190 = ( n1133 & n16187 ) | ( n1133 & n16189 ) | ( n16187 & n16189 ) ;
  assign n16186 = n10940 ^ n4128 ^ n1421 ;
  assign n16191 = n16190 ^ n16186 ^ n5714 ;
  assign n16192 = n353 ^ x115 ^ 1'b0 ;
  assign n16194 = n11797 ^ n597 ^ n555 ;
  assign n16193 = n9569 ^ n7177 ^ n3095 ;
  assign n16195 = n16194 ^ n16193 ^ 1'b0 ;
  assign n16196 = n16195 ^ n8694 ^ n405 ;
  assign n16197 = ( n4660 & n14520 ) | ( n4660 & ~n16196 ) | ( n14520 & ~n16196 ) ;
  assign n16198 = n4062 ^ n3762 ^ n2511 ;
  assign n16199 = n12556 | n16198 ;
  assign n16200 = n6264 ^ n5322 ^ n4879 ;
  assign n16201 = n16200 ^ n5695 ^ 1'b0 ;
  assign n16202 = n6818 | n16201 ;
  assign n16203 = n11090 ^ n5728 ^ 1'b0 ;
  assign n16204 = n6503 & n16203 ;
  assign n16205 = ( n1212 & n2790 ) | ( n1212 & n4241 ) | ( n2790 & n4241 ) ;
  assign n16206 = ( n2351 & n5451 ) | ( n2351 & ~n16205 ) | ( n5451 & ~n16205 ) ;
  assign n16207 = n584 & ~n3421 ;
  assign n16208 = n16207 ^ n393 ^ 1'b0 ;
  assign n16209 = n8989 ^ n1242 ^ 1'b0 ;
  assign n16210 = ( n3127 & n4770 ) | ( n3127 & n12205 ) | ( n4770 & n12205 ) ;
  assign n16211 = ( n16208 & n16209 ) | ( n16208 & n16210 ) | ( n16209 & n16210 ) ;
  assign n16212 = n16211 ^ n10880 ^ 1'b0 ;
  assign n16221 = ( x70 & n838 ) | ( x70 & n1501 ) | ( n838 & n1501 ) ;
  assign n16219 = ~n1843 & n5046 ;
  assign n16220 = ( n718 & n6182 ) | ( n718 & ~n16219 ) | ( n6182 & ~n16219 ) ;
  assign n16214 = ( n2269 & n4639 ) | ( n2269 & ~n13525 ) | ( n4639 & ~n13525 ) ;
  assign n16215 = n8912 & ~n16214 ;
  assign n16216 = n16215 ^ n440 ^ 1'b0 ;
  assign n16213 = n4241 ^ n1785 ^ 1'b0 ;
  assign n16217 = n16216 ^ n16213 ^ n5632 ;
  assign n16218 = n16217 ^ n2425 ^ 1'b0 ;
  assign n16222 = n16221 ^ n16220 ^ n16218 ;
  assign n16223 = n3295 ^ n3100 ^ 1'b0 ;
  assign n16228 = ( n499 & ~n10595 ) | ( n499 & n14936 ) | ( ~n10595 & n14936 ) ;
  assign n16229 = ( ~n715 & n4527 ) | ( ~n715 & n12188 ) | ( n4527 & n12188 ) ;
  assign n16230 = ( ~n324 & n2706 ) | ( ~n324 & n10627 ) | ( n2706 & n10627 ) ;
  assign n16231 = ( ~n1170 & n9670 ) | ( ~n1170 & n16230 ) | ( n9670 & n16230 ) ;
  assign n16232 = ( ~n16228 & n16229 ) | ( ~n16228 & n16231 ) | ( n16229 & n16231 ) ;
  assign n16224 = n4257 | n10365 ;
  assign n16225 = n12881 | n16224 ;
  assign n16226 = n10816 & n16225 ;
  assign n16227 = ~n15324 & n16226 ;
  assign n16233 = n16232 ^ n16227 ^ n7811 ;
  assign n16234 = ( ~n1099 & n7466 ) | ( ~n1099 & n8848 ) | ( n7466 & n8848 ) ;
  assign n16236 = n8109 ^ n2437 ^ 1'b0 ;
  assign n16237 = ( ~n5650 & n13772 ) | ( ~n5650 & n16236 ) | ( n13772 & n16236 ) ;
  assign n16235 = n7425 ^ n3997 ^ 1'b0 ;
  assign n16238 = n16237 ^ n16235 ^ n7353 ;
  assign n16239 = ( ~n8779 & n16234 ) | ( ~n8779 & n16238 ) | ( n16234 & n16238 ) ;
  assign n16240 = n5485 & ~n6610 ;
  assign n16241 = n2889 & n16240 ;
  assign n16242 = n16241 ^ n12845 ^ n8048 ;
  assign n16245 = ( ~n2022 & n4687 ) | ( ~n2022 & n4861 ) | ( n4687 & n4861 ) ;
  assign n16243 = n9572 ^ n6940 ^ 1'b0 ;
  assign n16244 = n6507 & n16243 ;
  assign n16246 = n16245 ^ n16244 ^ n15420 ;
  assign n16247 = n16242 | n16246 ;
  assign n16248 = ( ~n4982 & n5260 ) | ( ~n4982 & n8590 ) | ( n5260 & n8590 ) ;
  assign n16249 = n15123 ^ n1486 ^ n600 ;
  assign n16250 = n16249 ^ n3835 ^ 1'b0 ;
  assign n16251 = ~n14698 & n16250 ;
  assign n16252 = n6897 ^ n5862 ^ 1'b0 ;
  assign n16253 = n16252 ^ n537 ^ 1'b0 ;
  assign n16254 = ( n4855 & ~n10148 ) | ( n4855 & n16253 ) | ( ~n10148 & n16253 ) ;
  assign n16255 = n10415 ^ n9644 ^ n6997 ;
  assign n16256 = n2069 & n16255 ;
  assign n16257 = n16254 & n16256 ;
  assign n16258 = n3172 & n4145 ;
  assign n16259 = n8553 | n14785 ;
  assign n16260 = n16259 ^ n3045 ^ 1'b0 ;
  assign n16261 = n16260 ^ n3924 ^ 1'b0 ;
  assign n16262 = n7654 & n16261 ;
  assign n16263 = n16262 ^ n10883 ^ 1'b0 ;
  assign n16264 = n4553 ^ n1225 ^ n972 ;
  assign n16265 = n2079 & n2294 ;
  assign n16266 = n16265 ^ n5659 ^ 1'b0 ;
  assign n16267 = n16264 | n16266 ;
  assign n16268 = n4392 & ~n16267 ;
  assign n16269 = n14741 ^ n5336 ^ 1'b0 ;
  assign n16270 = n16269 ^ n9853 ^ n2741 ;
  assign n16271 = n16270 ^ n10178 ^ x63 ;
  assign n16272 = ( n3907 & ~n5699 ) | ( n3907 & n6617 ) | ( ~n5699 & n6617 ) ;
  assign n16273 = ( n3822 & n7229 ) | ( n3822 & ~n8394 ) | ( n7229 & ~n8394 ) ;
  assign n16274 = n10012 ^ n7415 ^ n7208 ;
  assign n16275 = ( n3960 & ~n16273 ) | ( n3960 & n16274 ) | ( ~n16273 & n16274 ) ;
  assign n16276 = ~n15086 & n16275 ;
  assign n16277 = n16272 & n16276 ;
  assign n16278 = n7656 & ~n16277 ;
  assign n16279 = n16278 ^ n16191 ^ 1'b0 ;
  assign n16285 = n6820 & ~n10559 ;
  assign n16286 = ~n491 & n16285 ;
  assign n16287 = ( n3582 & n5313 ) | ( n3582 & n16286 ) | ( n5313 & n16286 ) ;
  assign n16288 = n4579 ^ n2916 ^ n1176 ;
  assign n16289 = ( n2381 & n2837 ) | ( n2381 & n16288 ) | ( n2837 & n16288 ) ;
  assign n16290 = n16289 ^ n6846 ^ n1633 ;
  assign n16291 = ( ~n1783 & n2964 ) | ( ~n1783 & n16290 ) | ( n2964 & n16290 ) ;
  assign n16292 = n16287 & ~n16291 ;
  assign n16293 = ~n1273 & n16292 ;
  assign n16280 = n3428 & ~n3693 ;
  assign n16281 = n8203 ^ n1480 ^ 1'b0 ;
  assign n16282 = ( n2184 & n16280 ) | ( n2184 & ~n16281 ) | ( n16280 & ~n16281 ) ;
  assign n16283 = n16282 ^ n15016 ^ 1'b0 ;
  assign n16284 = n3600 & n16283 ;
  assign n16294 = n16293 ^ n16284 ^ 1'b0 ;
  assign n16295 = ( ~n3967 & n4566 ) | ( ~n3967 & n11870 ) | ( n4566 & n11870 ) ;
  assign n16296 = n6256 ^ n435 ^ 1'b0 ;
  assign n16297 = n16295 | n16296 ;
  assign n16298 = ( n2198 & ~n2295 ) | ( n2198 & n13344 ) | ( ~n2295 & n13344 ) ;
  assign n16299 = ( n3437 & ~n16297 ) | ( n3437 & n16298 ) | ( ~n16297 & n16298 ) ;
  assign n16300 = ~n1151 & n3306 ;
  assign n16301 = n3454 & n16300 ;
  assign n16302 = n4515 | n16301 ;
  assign n16303 = n16299 | n16302 ;
  assign n16304 = n3941 & n4504 ;
  assign n16305 = n16304 ^ n3301 ^ 1'b0 ;
  assign n16306 = n13150 ^ n12545 ^ n7559 ;
  assign n16307 = n2003 & n16306 ;
  assign n16308 = n16305 & n16307 ;
  assign n16309 = n4690 & ~n15982 ;
  assign n16310 = ~n16308 & n16309 ;
  assign n16313 = n5381 & ~n5817 ;
  assign n16314 = n3157 & n16313 ;
  assign n16311 = ( n1750 & ~n2126 ) | ( n1750 & n6189 ) | ( ~n2126 & n6189 ) ;
  assign n16312 = n16311 ^ n14554 ^ n9412 ;
  assign n16315 = n16314 ^ n16312 ^ n14055 ;
  assign n16316 = ( n13615 & n16310 ) | ( n13615 & ~n16315 ) | ( n16310 & ~n16315 ) ;
  assign n16317 = ( n2780 & ~n6886 ) | ( n2780 & n7829 ) | ( ~n6886 & n7829 ) ;
  assign n16318 = ( n12342 & ~n13011 ) | ( n12342 & n16317 ) | ( ~n13011 & n16317 ) ;
  assign n16319 = n14633 ^ n5423 ^ n1421 ;
  assign n16321 = ~n5949 & n6187 ;
  assign n16320 = n13172 ^ n10533 ^ n1993 ;
  assign n16322 = n16321 ^ n16320 ^ 1'b0 ;
  assign n16323 = ~n11040 & n16322 ;
  assign n16324 = ( ~n16318 & n16319 ) | ( ~n16318 & n16323 ) | ( n16319 & n16323 ) ;
  assign n16325 = n9312 ^ n6088 ^ 1'b0 ;
  assign n16327 = n679 & ~n10133 ;
  assign n16326 = n7202 & n11496 ;
  assign n16328 = n16327 ^ n16326 ^ 1'b0 ;
  assign n16329 = n10405 ^ n5000 ^ 1'b0 ;
  assign n16330 = n11074 & ~n16329 ;
  assign n16331 = ( n241 & ~n4967 ) | ( n241 & n6739 ) | ( ~n4967 & n6739 ) ;
  assign n16332 = ( ~n6552 & n8103 ) | ( ~n6552 & n16331 ) | ( n8103 & n16331 ) ;
  assign n16333 = n13021 ^ n4515 ^ 1'b0 ;
  assign n16334 = ( n1623 & ~n4336 ) | ( n1623 & n5624 ) | ( ~n4336 & n5624 ) ;
  assign n16339 = n14435 ^ n10142 ^ n959 ;
  assign n16335 = n2073 & ~n4932 ;
  assign n16336 = n16335 ^ n5905 ^ 1'b0 ;
  assign n16337 = ~n11563 & n16336 ;
  assign n16338 = n16337 ^ n3513 ^ 1'b0 ;
  assign n16340 = n16339 ^ n16338 ^ n4664 ;
  assign n16341 = ( n13135 & n16334 ) | ( n13135 & ~n16340 ) | ( n16334 & ~n16340 ) ;
  assign n16342 = n7299 ^ n6397 ^ 1'b0 ;
  assign n16343 = n5723 | n16342 ;
  assign n16344 = n9279 ^ n5855 ^ n3000 ;
  assign n16345 = ~n3503 & n13627 ;
  assign n16346 = ( ~n3334 & n6992 ) | ( ~n3334 & n14051 ) | ( n6992 & n14051 ) ;
  assign n16347 = n16345 & n16346 ;
  assign n16348 = ~n16344 & n16347 ;
  assign n16350 = ~n900 & n5651 ;
  assign n16351 = n16350 ^ n3061 ^ 1'b0 ;
  assign n16349 = ~n5061 & n8498 ;
  assign n16352 = n16351 ^ n16349 ^ 1'b0 ;
  assign n16353 = ~n4114 & n16352 ;
  assign n16354 = n729 & n16353 ;
  assign n16355 = ( ~n1447 & n11545 ) | ( ~n1447 & n16354 ) | ( n11545 & n16354 ) ;
  assign n16356 = n5371 ^ n804 ^ 1'b0 ;
  assign n16357 = n4374 ^ n3602 ^ n639 ;
  assign n16358 = ( n1647 & n5629 ) | ( n1647 & n16357 ) | ( n5629 & n16357 ) ;
  assign n16359 = ( n6910 & n9850 ) | ( n6910 & n16358 ) | ( n9850 & n16358 ) ;
  assign n16360 = n16359 ^ n3309 ^ 1'b0 ;
  assign n16361 = n9467 ^ n4061 ^ 1'b0 ;
  assign n16362 = n2524 & n16361 ;
  assign n16363 = n2592 | n9703 ;
  assign n16364 = x11 & n16363 ;
  assign n16365 = ~n4569 & n16364 ;
  assign n16366 = n11511 & n16365 ;
  assign n16367 = n13414 ^ n12418 ^ n10848 ;
  assign n16368 = n3609 & n10623 ;
  assign n16369 = n16368 ^ n11321 ^ 1'b0 ;
  assign n16370 = n16369 ^ n4085 ^ n3293 ;
  assign n16371 = n8851 ^ n7481 ^ n7311 ;
  assign n16372 = n16371 ^ n13269 ^ n12905 ;
  assign n16373 = n15228 ^ n462 ^ 1'b0 ;
  assign n16374 = n2611 & n16373 ;
  assign n16375 = n543 & n16374 ;
  assign n16376 = n2022 | n9608 ;
  assign n16377 = n16376 ^ n754 ^ 1'b0 ;
  assign n16378 = n16377 ^ n6813 ^ n3971 ;
  assign n16379 = n7490 & ~n16378 ;
  assign n16380 = ( n10512 & n16375 ) | ( n10512 & ~n16379 ) | ( n16375 & ~n16379 ) ;
  assign n16381 = n13697 ^ n5774 ^ n1230 ;
  assign n16382 = n9067 ^ n2425 ^ n285 ;
  assign n16383 = ~n13620 & n16382 ;
  assign n16384 = ~n4261 & n6113 ;
  assign n16385 = n16384 ^ n11026 ^ 1'b0 ;
  assign n16386 = n13899 & ~n16385 ;
  assign n16387 = n16386 ^ n12748 ^ 1'b0 ;
  assign n16390 = n5967 ^ n3851 ^ n2364 ;
  assign n16388 = ( n1066 & ~n10368 ) | ( n1066 & n11146 ) | ( ~n10368 & n11146 ) ;
  assign n16389 = ( n6569 & ~n7245 ) | ( n6569 & n16388 ) | ( ~n7245 & n16388 ) ;
  assign n16391 = n16390 ^ n16389 ^ 1'b0 ;
  assign n16392 = n16391 ^ n8771 ^ n6508 ;
  assign n16393 = ~n2686 & n16392 ;
  assign n16394 = n15721 & n16393 ;
  assign n16395 = n2738 ^ n264 ^ 1'b0 ;
  assign n16396 = n13165 & n14908 ;
  assign n16397 = n8820 & ~n15564 ;
  assign n16398 = n16397 ^ n10488 ^ 1'b0 ;
  assign n16399 = ~n5899 & n10343 ;
  assign n16400 = n16399 ^ n4850 ^ n1117 ;
  assign n16401 = n16400 ^ n15690 ^ 1'b0 ;
  assign n16402 = n13777 ^ n11118 ^ 1'b0 ;
  assign n16403 = ( n1665 & n10123 ) | ( n1665 & n11363 ) | ( n10123 & n11363 ) ;
  assign n16404 = n16403 ^ n12703 ^ n5073 ;
  assign n16405 = n9649 ^ n2443 ^ n2363 ;
  assign n16406 = n16030 & n16405 ;
  assign n16407 = n16404 | n16406 ;
  assign n16408 = n16019 ^ n6538 ^ n1893 ;
  assign n16409 = ( n7834 & n13693 ) | ( n7834 & n16408 ) | ( n13693 & n16408 ) ;
  assign n16410 = n9013 ^ n7175 ^ 1'b0 ;
  assign n16411 = n2232 & n16410 ;
  assign n16412 = n2789 & ~n10837 ;
  assign n16413 = n4200 & ~n11463 ;
  assign n16414 = n16413 ^ n10623 ^ 1'b0 ;
  assign n16415 = ( n6388 & n10058 ) | ( n6388 & n10502 ) | ( n10058 & n10502 ) ;
  assign n16416 = ~n10976 & n13971 ;
  assign n16417 = n16415 & n16416 ;
  assign n16418 = n16417 ^ n10011 ^ 1'b0 ;
  assign n16421 = n8140 & ~n8195 ;
  assign n16419 = ( n3125 & n3747 ) | ( n3125 & n5004 ) | ( n3747 & n5004 ) ;
  assign n16420 = ( n3080 & n9298 ) | ( n3080 & ~n16419 ) | ( n9298 & ~n16419 ) ;
  assign n16422 = n16421 ^ n16420 ^ n7280 ;
  assign n16423 = ( n3731 & n7389 ) | ( n3731 & ~n9031 ) | ( n7389 & ~n9031 ) ;
  assign n16424 = n15186 ^ n671 ^ 1'b0 ;
  assign n16425 = n569 & ~n16424 ;
  assign n16426 = ( n830 & n1938 ) | ( n830 & n11472 ) | ( n1938 & n11472 ) ;
  assign n16427 = ( n1527 & n3125 ) | ( n1527 & n8928 ) | ( n3125 & n8928 ) ;
  assign n16428 = ~n16426 & n16427 ;
  assign n16429 = n7868 & n16428 ;
  assign n16430 = n16425 & ~n16429 ;
  assign n16431 = ~n9865 & n16430 ;
  assign n16432 = ( ~n2739 & n4545 ) | ( ~n2739 & n11915 ) | ( n4545 & n11915 ) ;
  assign n16433 = ( n3574 & n14399 ) | ( n3574 & n15628 ) | ( n14399 & n15628 ) ;
  assign n16436 = n3682 ^ n3038 ^ n2971 ;
  assign n16437 = n9597 ^ n5718 ^ n2190 ;
  assign n16438 = n6448 & ~n16437 ;
  assign n16439 = ( n9614 & n16436 ) | ( n9614 & ~n16438 ) | ( n16436 & ~n16438 ) ;
  assign n16434 = n3866 | n9682 ;
  assign n16435 = n16434 ^ n541 ^ 1'b0 ;
  assign n16440 = n16439 ^ n16435 ^ 1'b0 ;
  assign n16441 = n16440 ^ n14094 ^ n5428 ;
  assign n16442 = n16441 ^ n2940 ^ n773 ;
  assign n16443 = n8710 & ~n15565 ;
  assign n16444 = n16443 ^ n16042 ^ 1'b0 ;
  assign n16445 = n16444 ^ n3134 ^ 1'b0 ;
  assign n16446 = n13803 & ~n16445 ;
  assign n16447 = n3466 | n13210 ;
  assign n16448 = n16447 ^ n10397 ^ 1'b0 ;
  assign n16449 = n5837 ^ n2678 ^ 1'b0 ;
  assign n16450 = n8473 | n16449 ;
  assign n16451 = n3574 & n16450 ;
  assign n16452 = n9907 ^ n234 ^ 1'b0 ;
  assign n16453 = ~n16451 & n16452 ;
  assign n16454 = n16453 ^ n14266 ^ 1'b0 ;
  assign n16455 = n11160 ^ n11121 ^ n10060 ;
  assign n16456 = n6209 | n8588 ;
  assign n16457 = n16456 ^ n6228 ^ 1'b0 ;
  assign n16458 = ( n4751 & n7080 ) | ( n4751 & ~n16457 ) | ( n7080 & ~n16457 ) ;
  assign n16459 = n620 | n16458 ;
  assign n16460 = n15818 ^ n13357 ^ n4891 ;
  assign n16461 = ( n1952 & n7230 ) | ( n1952 & ~n15221 ) | ( n7230 & ~n15221 ) ;
  assign n16462 = ( ~n7844 & n16238 ) | ( ~n7844 & n16461 ) | ( n16238 & n16461 ) ;
  assign n16463 = n16462 ^ n5303 ^ n4761 ;
  assign n16464 = ( ~n9538 & n10869 ) | ( ~n9538 & n16463 ) | ( n10869 & n16463 ) ;
  assign n16465 = ( n6197 & n15152 ) | ( n6197 & ~n16464 ) | ( n15152 & ~n16464 ) ;
  assign n16466 = ( n201 & n1978 ) | ( n201 & ~n5311 ) | ( n1978 & ~n5311 ) ;
  assign n16467 = n16466 ^ n13389 ^ 1'b0 ;
  assign n16468 = n4591 & ~n16467 ;
  assign n16469 = n6033 & n16468 ;
  assign n16470 = n10912 ^ n6742 ^ x100 ;
  assign n16471 = ( n4649 & n5230 ) | ( n4649 & ~n8255 ) | ( n5230 & ~n8255 ) ;
  assign n16472 = n16471 ^ n3409 ^ n2388 ;
  assign n16473 = ( n5138 & n6823 ) | ( n5138 & ~n9717 ) | ( n6823 & ~n9717 ) ;
  assign n16474 = n16473 ^ n15677 ^ 1'b0 ;
  assign n16475 = n11341 ^ n4159 ^ 1'b0 ;
  assign n16476 = ~n4012 & n16475 ;
  assign n16477 = x41 & ~n16476 ;
  assign n16478 = n7143 ^ n332 ^ 1'b0 ;
  assign n16479 = ~n16477 & n16478 ;
  assign n16480 = ( n5468 & n16365 ) | ( n5468 & n16479 ) | ( n16365 & n16479 ) ;
  assign n16481 = ( n3686 & n8954 ) | ( n3686 & ~n15538 ) | ( n8954 & ~n15538 ) ;
  assign n16482 = n2995 | n6355 ;
  assign n16483 = n16482 ^ n15246 ^ 1'b0 ;
  assign n16484 = n16481 & ~n16483 ;
  assign n16485 = n2631 ^ n1992 ^ 1'b0 ;
  assign n16486 = n1914 & n16485 ;
  assign n16487 = n6386 ^ n1898 ^ 1'b0 ;
  assign n16488 = n15542 | n16487 ;
  assign n16489 = ( n3556 & n11541 ) | ( n3556 & ~n16488 ) | ( n11541 & ~n16488 ) ;
  assign n16490 = n4543 | n7520 ;
  assign n16491 = n16490 ^ n2592 ^ 1'b0 ;
  assign n16492 = n16491 ^ n15111 ^ x48 ;
  assign n16493 = n2962 & ~n8744 ;
  assign n16494 = n9883 & n16493 ;
  assign n16495 = n6759 ^ n1009 ^ 1'b0 ;
  assign n16496 = n16495 ^ n1326 ^ n627 ;
  assign n16497 = n16496 ^ n3217 ^ 1'b0 ;
  assign n16498 = n16494 | n16497 ;
  assign n16499 = n3731 | n11474 ;
  assign n16500 = n16499 ^ n4749 ^ 1'b0 ;
  assign n16501 = ~n9672 & n12074 ;
  assign n16502 = n16501 ^ n8175 ^ 1'b0 ;
  assign n16503 = ( n12960 & n16500 ) | ( n12960 & ~n16502 ) | ( n16500 & ~n16502 ) ;
  assign n16504 = ( n9158 & n13088 ) | ( n9158 & ~n16503 ) | ( n13088 & ~n16503 ) ;
  assign n16505 = n13979 ^ n1987 ^ 1'b0 ;
  assign n16506 = n11349 ^ n10584 ^ 1'b0 ;
  assign n16507 = n4590 & n16506 ;
  assign n16508 = n16507 ^ n13431 ^ n3093 ;
  assign n16509 = n8496 ^ n4066 ^ n3408 ;
  assign n16510 = n16509 ^ n5218 ^ 1'b0 ;
  assign n16511 = ( n2524 & ~n16508 ) | ( n2524 & n16510 ) | ( ~n16508 & n16510 ) ;
  assign n16512 = n8966 | n9171 ;
  assign n16513 = n6566 ^ n713 ^ 1'b0 ;
  assign n16514 = ~n16512 & n16513 ;
  assign n16515 = ( n517 & ~n7275 ) | ( n517 & n8764 ) | ( ~n7275 & n8764 ) ;
  assign n16516 = n11698 ^ n9057 ^ 1'b0 ;
  assign n16517 = ( n4762 & n16220 ) | ( n4762 & ~n16516 ) | ( n16220 & ~n16516 ) ;
  assign n16518 = ( n11157 & n16515 ) | ( n11157 & n16517 ) | ( n16515 & n16517 ) ;
  assign n16519 = ( n4253 & n16514 ) | ( n4253 & ~n16518 ) | ( n16514 & ~n16518 ) ;
  assign n16520 = ( n6353 & n8636 ) | ( n6353 & n11772 ) | ( n8636 & n11772 ) ;
  assign n16521 = ( n13335 & ~n15553 ) | ( n13335 & n16520 ) | ( ~n15553 & n16520 ) ;
  assign n16522 = n16521 ^ n13465 ^ n7425 ;
  assign n16524 = ( n4304 & n9771 ) | ( n4304 & n12654 ) | ( n9771 & n12654 ) ;
  assign n16523 = n544 & ~n6363 ;
  assign n16525 = n16524 ^ n16523 ^ 1'b0 ;
  assign n16526 = ~n335 & n9622 ;
  assign n16527 = ~n4090 & n16526 ;
  assign n16528 = n16527 ^ n8618 ^ n7940 ;
  assign n16529 = n16528 ^ n15501 ^ n9592 ;
  assign n16530 = ~n253 & n8354 ;
  assign n16531 = ( n3032 & n6542 ) | ( n3032 & n16281 ) | ( n6542 & n16281 ) ;
  assign n16532 = ( n2859 & ~n5981 ) | ( n2859 & n16531 ) | ( ~n5981 & n16531 ) ;
  assign n16533 = n14498 ^ n6886 ^ 1'b0 ;
  assign n16534 = n16533 ^ n14215 ^ n644 ;
  assign n16535 = n16534 ^ n4034 ^ n1876 ;
  assign n16536 = ( ~n16530 & n16532 ) | ( ~n16530 & n16535 ) | ( n16532 & n16535 ) ;
  assign n16537 = ( n5438 & n5841 ) | ( n5438 & ~n9237 ) | ( n5841 & ~n9237 ) ;
  assign n16538 = ( ~n3498 & n13780 ) | ( ~n3498 & n16537 ) | ( n13780 & n16537 ) ;
  assign n16539 = ( ~n272 & n4567 ) | ( ~n272 & n16538 ) | ( n4567 & n16538 ) ;
  assign n16540 = ( n7059 & ~n13021 ) | ( n7059 & n13601 ) | ( ~n13021 & n13601 ) ;
  assign n16541 = n15155 ^ n12234 ^ 1'b0 ;
  assign n16542 = ( ~n8717 & n12707 ) | ( ~n8717 & n16541 ) | ( n12707 & n16541 ) ;
  assign n16548 = ( n3320 & ~n8280 ) | ( n3320 & n12787 ) | ( ~n8280 & n12787 ) ;
  assign n16545 = ~n1216 & n3677 ;
  assign n16546 = ~n425 & n16545 ;
  assign n16547 = n4164 & ~n16546 ;
  assign n16549 = n16548 ^ n16547 ^ 1'b0 ;
  assign n16543 = n3916 ^ n1417 ^ n719 ;
  assign n16544 = n16543 ^ n15655 ^ n6109 ;
  assign n16550 = n16549 ^ n16544 ^ 1'b0 ;
  assign n16551 = ( ~n5836 & n8759 ) | ( ~n5836 & n16550 ) | ( n8759 & n16550 ) ;
  assign n16555 = ( n3113 & n4645 ) | ( n3113 & ~n8343 ) | ( n4645 & ~n8343 ) ;
  assign n16552 = ( n6256 & n8781 ) | ( n6256 & n16229 ) | ( n8781 & n16229 ) ;
  assign n16553 = ( n8256 & ~n13264 ) | ( n8256 & n16552 ) | ( ~n13264 & n16552 ) ;
  assign n16554 = ~n13052 & n16553 ;
  assign n16556 = n16555 ^ n16554 ^ n13272 ;
  assign n16557 = ( ~n2482 & n4622 ) | ( ~n2482 & n6825 ) | ( n4622 & n6825 ) ;
  assign n16558 = ( n247 & n4752 ) | ( n247 & ~n16557 ) | ( n4752 & ~n16557 ) ;
  assign n16559 = n2697 & n13104 ;
  assign n16560 = n16558 & n16559 ;
  assign n16561 = ( x26 & ~n8967 ) | ( x26 & n16560 ) | ( ~n8967 & n16560 ) ;
  assign n16564 = n7202 ^ n3292 ^ n1462 ;
  assign n16565 = n16564 ^ n9120 ^ 1'b0 ;
  assign n16562 = n5494 ^ n2071 ^ 1'b0 ;
  assign n16563 = n16562 ^ n12154 ^ n2500 ;
  assign n16566 = n16565 ^ n16563 ^ 1'b0 ;
  assign n16567 = ( n637 & ~n748 ) | ( n637 & n2393 ) | ( ~n748 & n2393 ) ;
  assign n16568 = n16567 ^ n16118 ^ n12740 ;
  assign n16575 = ~n220 & n860 ;
  assign n16576 = n16575 ^ n10666 ^ 1'b0 ;
  assign n16577 = n3737 & n16576 ;
  assign n16573 = ( n1172 & ~n5761 ) | ( n1172 & n12249 ) | ( ~n5761 & n12249 ) ;
  assign n16571 = n7726 ^ n1620 ^ 1'b0 ;
  assign n16569 = n1227 & n3470 ;
  assign n16570 = n15893 & n16569 ;
  assign n16572 = n16571 ^ n16570 ^ 1'b0 ;
  assign n16574 = n16573 ^ n16572 ^ n3068 ;
  assign n16578 = n16577 ^ n16574 ^ n5715 ;
  assign n16579 = ( n5430 & ~n6352 ) | ( n5430 & n12054 ) | ( ~n6352 & n12054 ) ;
  assign n16580 = ( n2386 & n4388 ) | ( n2386 & n4899 ) | ( n4388 & n4899 ) ;
  assign n16581 = n16580 ^ n11247 ^ 1'b0 ;
  assign n16582 = n10251 ^ n5065 ^ n1947 ;
  assign n16583 = ~n9400 & n16582 ;
  assign n16584 = n16583 ^ n11769 ^ n1323 ;
  assign n16585 = n16584 ^ n15031 ^ n12583 ;
  assign n16586 = n15289 ^ n4064 ^ 1'b0 ;
  assign n16587 = n1307 & n16586 ;
  assign n16588 = ( n4431 & n13876 ) | ( n4431 & n16587 ) | ( n13876 & n16587 ) ;
  assign n16589 = n13440 ^ n3421 ^ n2548 ;
  assign n16597 = n4396 | n10768 ;
  assign n16598 = n16597 ^ n5609 ^ 1'b0 ;
  assign n16595 = ( n845 & ~n3799 ) | ( n845 & n7063 ) | ( ~n3799 & n7063 ) ;
  assign n16593 = ( n1859 & n4346 ) | ( n1859 & n12259 ) | ( n4346 & n12259 ) ;
  assign n16590 = ( ~n1686 & n2511 ) | ( ~n1686 & n8205 ) | ( n2511 & n8205 ) ;
  assign n16591 = n16590 ^ n4353 ^ n239 ;
  assign n16592 = n10575 & ~n16591 ;
  assign n16594 = n16593 ^ n16592 ^ 1'b0 ;
  assign n16596 = n16595 ^ n16594 ^ n14942 ;
  assign n16599 = n16598 ^ n16596 ^ n4470 ;
  assign n16600 = ( n445 & ~n7576 ) | ( n445 & n16599 ) | ( ~n7576 & n16599 ) ;
  assign n16601 = n7104 & ~n16600 ;
  assign n16602 = n4947 | n13960 ;
  assign n16603 = n11641 ^ n8630 ^ n805 ;
  assign n16604 = ( n1143 & n3845 ) | ( n1143 & n7463 ) | ( n3845 & n7463 ) ;
  assign n16605 = n16604 ^ n10568 ^ n8308 ;
  assign n16606 = ~n5525 & n9973 ;
  assign n16607 = n16606 ^ n13463 ^ 1'b0 ;
  assign n16608 = ~n5699 & n16607 ;
  assign n16609 = ( n5359 & n16425 ) | ( n5359 & ~n16608 ) | ( n16425 & ~n16608 ) ;
  assign n16610 = n3200 & n8230 ;
  assign n16611 = n16610 ^ n15969 ^ 1'b0 ;
  assign n16612 = ( n11767 & n13373 ) | ( n11767 & ~n16611 ) | ( n13373 & ~n16611 ) ;
  assign n16613 = n9445 ^ n2488 ^ 1'b0 ;
  assign n16614 = n4507 & ~n16613 ;
  assign n16615 = n8775 & n16614 ;
  assign n16616 = ~n16612 & n16615 ;
  assign n16617 = n16616 ^ n9043 ^ 1'b0 ;
  assign n16618 = n5541 & ~n8533 ;
  assign n16619 = n9848 ^ n2788 ^ n1677 ;
  assign n16620 = ( n3879 & n4946 ) | ( n3879 & n6521 ) | ( n4946 & n6521 ) ;
  assign n16621 = ~n4676 & n4697 ;
  assign n16622 = n16620 & n16621 ;
  assign n16623 = ( n12043 & n16619 ) | ( n12043 & ~n16622 ) | ( n16619 & ~n16622 ) ;
  assign n16624 = n14342 ^ n10652 ^ n129 ;
  assign n16625 = n16624 ^ n11735 ^ 1'b0 ;
  assign n16626 = n2942 & ~n16625 ;
  assign n16627 = n16626 ^ n15864 ^ n5802 ;
  assign n16628 = n8781 ^ n7502 ^ n7313 ;
  assign n16629 = n7700 ^ n6589 ^ n424 ;
  assign n16630 = ( n1327 & n7976 ) | ( n1327 & ~n16629 ) | ( n7976 & ~n16629 ) ;
  assign n16631 = n1965 | n5910 ;
  assign n16632 = n13134 | n16631 ;
  assign n16633 = n16632 ^ n1492 ^ 1'b0 ;
  assign n16634 = n6532 & n16633 ;
  assign n16635 = n13827 ^ n10597 ^ n5771 ;
  assign n16636 = n16635 ^ n13813 ^ 1'b0 ;
  assign n16637 = n13675 & ~n16636 ;
  assign n16638 = n16637 ^ n12094 ^ n2137 ;
  assign n16639 = n8103 ^ n3411 ^ n1543 ;
  assign n16640 = n16639 ^ n6861 ^ 1'b0 ;
  assign n16641 = n1437 | n2031 ;
  assign n16642 = n11794 & ~n16641 ;
  assign n16643 = n16642 ^ n13824 ^ n8241 ;
  assign n16644 = n16643 ^ n13707 ^ n4970 ;
  assign n16645 = ~n1075 & n16235 ;
  assign n16646 = n9363 ^ n6394 ^ n4758 ;
  assign n16647 = n2892 | n16646 ;
  assign n16649 = n3057 & n5234 ;
  assign n16650 = n4702 & n16649 ;
  assign n16648 = n9705 ^ n5160 ^ n1744 ;
  assign n16651 = n16650 ^ n16648 ^ n9573 ;
  assign n16652 = ~n2363 & n4028 ;
  assign n16653 = n16652 ^ n3575 ^ n639 ;
  assign n16654 = ( ~n2960 & n6199 ) | ( ~n2960 & n8966 ) | ( n6199 & n8966 ) ;
  assign n16655 = n16654 ^ n15986 ^ 1'b0 ;
  assign n16656 = n16653 & ~n16655 ;
  assign n16657 = ( n9475 & n11847 ) | ( n9475 & n16656 ) | ( n11847 & n16656 ) ;
  assign n16658 = n467 & ~n5235 ;
  assign n16659 = n7193 & ~n13310 ;
  assign n16660 = ~n16658 & n16659 ;
  assign n16662 = ( ~n745 & n1151 ) | ( ~n745 & n8191 ) | ( n1151 & n8191 ) ;
  assign n16661 = ~n4956 & n15460 ;
  assign n16663 = n16662 ^ n16661 ^ 1'b0 ;
  assign n16664 = n11914 ^ n5297 ^ 1'b0 ;
  assign n16665 = ~n303 & n16664 ;
  assign n16666 = ( n331 & n3184 ) | ( n331 & ~n16665 ) | ( n3184 & ~n16665 ) ;
  assign n16667 = n13997 ^ n1953 ^ n533 ;
  assign n16668 = ( ~n13088 & n15453 ) | ( ~n13088 & n16667 ) | ( n15453 & n16667 ) ;
  assign n16669 = n9231 | n14726 ;
  assign n16670 = n7178 ^ n1635 ^ n1116 ;
  assign n16671 = ( n1250 & n10114 ) | ( n1250 & ~n16670 ) | ( n10114 & ~n16670 ) ;
  assign n16672 = n5336 ^ n2702 ^ n362 ;
  assign n16673 = n3039 ^ n2961 ^ n1695 ;
  assign n16674 = ~n4798 & n16673 ;
  assign n16675 = ~n16672 & n16674 ;
  assign n16676 = n9248 ^ n4331 ^ n659 ;
  assign n16677 = ( n2281 & n5470 ) | ( n2281 & n16676 ) | ( n5470 & n16676 ) ;
  assign n16678 = ~n1775 & n16677 ;
  assign n16679 = ~n16675 & n16678 ;
  assign n16680 = n15699 ^ n15206 ^ n3593 ;
  assign n16681 = ( n3528 & n3660 ) | ( n3528 & n5657 ) | ( n3660 & n5657 ) ;
  assign n16682 = ( n13297 & n13502 ) | ( n13297 & ~n16681 ) | ( n13502 & ~n16681 ) ;
  assign n16683 = ( ~n11769 & n14065 ) | ( ~n11769 & n14618 ) | ( n14065 & n14618 ) ;
  assign n16684 = n865 & ~n16683 ;
  assign n16685 = n3530 & n16684 ;
  assign n16687 = ( n1746 & n3365 ) | ( n1746 & ~n4624 ) | ( n3365 & ~n4624 ) ;
  assign n16686 = ~n5186 & n8856 ;
  assign n16688 = n16687 ^ n16686 ^ x113 ;
  assign n16689 = ( n2565 & ~n3139 ) | ( n2565 & n11669 ) | ( ~n3139 & n11669 ) ;
  assign n16690 = n9384 | n16689 ;
  assign n16691 = n11881 ^ n2225 ^ 1'b0 ;
  assign n16692 = n5652 & n13614 ;
  assign n16693 = n16691 & n16692 ;
  assign n16694 = ( ~n962 & n3257 ) | ( ~n962 & n16693 ) | ( n3257 & n16693 ) ;
  assign n16695 = ( ~n216 & n1192 ) | ( ~n216 & n16694 ) | ( n1192 & n16694 ) ;
  assign n16696 = ( x73 & ~n2467 ) | ( x73 & n2918 ) | ( ~n2467 & n2918 ) ;
  assign n16697 = ( n2287 & ~n5108 ) | ( n2287 & n16696 ) | ( ~n5108 & n16696 ) ;
  assign n16698 = n16697 ^ n6811 ^ n3080 ;
  assign n16699 = n6975 & ~n16628 ;
  assign n16700 = n7878 & n16699 ;
  assign n16701 = ( n467 & ~n8092 ) | ( n467 & n14692 ) | ( ~n8092 & n14692 ) ;
  assign n16702 = n4030 ^ n1977 ^ 1'b0 ;
  assign n16703 = n7912 & ~n12218 ;
  assign n16704 = n16702 & n16703 ;
  assign n16705 = n16704 ^ n5324 ^ 1'b0 ;
  assign n16706 = n16701 | n16705 ;
  assign n16707 = n6943 ^ n5877 ^ n4284 ;
  assign n16708 = n10232 & n11153 ;
  assign n16709 = n16708 ^ n3536 ^ 1'b0 ;
  assign n16710 = n16709 ^ n6091 ^ n2581 ;
  assign n16711 = n1001 & ~n4195 ;
  assign n16712 = n16711 ^ n6210 ^ 1'b0 ;
  assign n16713 = n4760 ^ n566 ^ 1'b0 ;
  assign n16714 = n2454 & n16713 ;
  assign n16715 = n16126 ^ n14844 ^ n8611 ;
  assign n16716 = ( ~n4750 & n16714 ) | ( ~n4750 & n16715 ) | ( n16714 & n16715 ) ;
  assign n16717 = n6487 ^ n6055 ^ n1060 ;
  assign n16724 = n3754 ^ n3675 ^ n3056 ;
  assign n16725 = n6153 | n16724 ;
  assign n16726 = n16725 ^ n4791 ^ 1'b0 ;
  assign n16718 = n9195 ^ n1515 ^ 1'b0 ;
  assign n16719 = n13684 & ~n16718 ;
  assign n16720 = ( n611 & n4801 ) | ( n611 & n10528 ) | ( n4801 & n10528 ) ;
  assign n16721 = ~n9658 & n16720 ;
  assign n16722 = ~n16719 & n16721 ;
  assign n16723 = n685 & ~n16722 ;
  assign n16727 = n16726 ^ n16723 ^ 1'b0 ;
  assign n16728 = n16727 ^ n8414 ^ n6042 ;
  assign n16729 = n1269 & n7621 ;
  assign n16730 = n360 | n10053 ;
  assign n16731 = n16729 | n16730 ;
  assign n16732 = ( n16717 & ~n16728 ) | ( n16717 & n16731 ) | ( ~n16728 & n16731 ) ;
  assign n16733 = n202 & ~n14639 ;
  assign n16734 = ~n4378 & n16733 ;
  assign n16735 = ( n2212 & n5089 ) | ( n2212 & n8581 ) | ( n5089 & n8581 ) ;
  assign n16736 = ~n4848 & n10528 ;
  assign n16737 = n16735 & n16736 ;
  assign n16738 = n14244 ^ n11069 ^ 1'b0 ;
  assign n16739 = ~n6336 & n16363 ;
  assign n16740 = n16738 & n16739 ;
  assign n16741 = n1379 ^ n598 ^ 1'b0 ;
  assign n16742 = ( n7636 & n16740 ) | ( n7636 & ~n16741 ) | ( n16740 & ~n16741 ) ;
  assign n16751 = ( n3999 & ~n6277 ) | ( n3999 & n9853 ) | ( ~n6277 & n9853 ) ;
  assign n16749 = n2358 | n2498 ;
  assign n16745 = n6238 | n14729 ;
  assign n16746 = n1273 | n16745 ;
  assign n16744 = n9909 ^ n1050 ^ n667 ;
  assign n16743 = ( ~n648 & n875 ) | ( ~n648 & n6658 ) | ( n875 & n6658 ) ;
  assign n16747 = n16746 ^ n16744 ^ n16743 ;
  assign n16748 = n16747 ^ n3952 ^ 1'b0 ;
  assign n16750 = n16749 ^ n16748 ^ 1'b0 ;
  assign n16752 = n16751 ^ n16750 ^ n15963 ;
  assign n16759 = ( x68 & n1360 ) | ( x68 & ~n3350 ) | ( n1360 & ~n3350 ) ;
  assign n16760 = ( ~n1212 & n1472 ) | ( ~n1212 & n13608 ) | ( n1472 & n13608 ) ;
  assign n16761 = n16759 | n16760 ;
  assign n16762 = n16761 ^ n13865 ^ n3762 ;
  assign n16753 = ( n3047 & n5496 ) | ( n3047 & n5665 ) | ( n5496 & n5665 ) ;
  assign n16755 = n16334 ^ n10318 ^ n8995 ;
  assign n16754 = n9346 ^ n7429 ^ n5279 ;
  assign n16756 = n16755 ^ n16754 ^ n4873 ;
  assign n16757 = n16756 ^ n6754 ^ n1802 ;
  assign n16758 = ~n16753 & n16757 ;
  assign n16763 = n16762 ^ n16758 ^ 1'b0 ;
  assign n16764 = ~n645 & n6676 ;
  assign n16765 = n16764 ^ n2188 ^ 1'b0 ;
  assign n16767 = ~n2470 & n5117 ;
  assign n16768 = n16767 ^ n4732 ^ 1'b0 ;
  assign n16766 = ( ~n5406 & n6948 ) | ( ~n5406 & n12407 ) | ( n6948 & n12407 ) ;
  assign n16769 = n16768 ^ n16766 ^ n3208 ;
  assign n16770 = n4994 | n15933 ;
  assign n16771 = n16770 ^ n14877 ^ n13631 ;
  assign n16772 = ( n7726 & n10153 ) | ( n7726 & n14692 ) | ( n10153 & n14692 ) ;
  assign n16773 = ~n6732 & n15521 ;
  assign n16774 = n7913 ^ n2125 ^ 1'b0 ;
  assign n16780 = ( n2852 & n5078 ) | ( n2852 & n10772 ) | ( n5078 & n10772 ) ;
  assign n16781 = ( n4604 & n10583 ) | ( n4604 & n16780 ) | ( n10583 & n16780 ) ;
  assign n16775 = n2252 & ~n8015 ;
  assign n16776 = ( n2794 & n6513 ) | ( n2794 & n16775 ) | ( n6513 & n16775 ) ;
  assign n16777 = ~n15304 & n15421 ;
  assign n16778 = n16777 ^ n7674 ^ 1'b0 ;
  assign n16779 = n16776 | n16778 ;
  assign n16782 = n16781 ^ n16779 ^ 1'b0 ;
  assign n16783 = ( ~n3242 & n7697 ) | ( ~n3242 & n10200 ) | ( n7697 & n10200 ) ;
  assign n16784 = n4562 & n5435 ;
  assign n16785 = n4294 & n12271 ;
  assign n16786 = ~n16784 & n16785 ;
  assign n16787 = n7801 ^ n4112 ^ n2814 ;
  assign n16788 = ( n16783 & n16786 ) | ( n16783 & ~n16787 ) | ( n16786 & ~n16787 ) ;
  assign n16789 = n6972 ^ n6893 ^ 1'b0 ;
  assign n16790 = n762 & n7461 ;
  assign n16791 = ( n9739 & n16789 ) | ( n9739 & ~n16790 ) | ( n16789 & ~n16790 ) ;
  assign n16792 = n16791 ^ n7495 ^ n4813 ;
  assign n16793 = n14010 ^ n12983 ^ n5822 ;
  assign n16794 = n2302 & n15288 ;
  assign n16795 = n16794 ^ n13333 ^ 1'b0 ;
  assign n16796 = ~n3190 & n3315 ;
  assign n16797 = n16796 ^ n13309 ^ n2813 ;
  assign n16798 = n16797 ^ n16480 ^ 1'b0 ;
  assign n16799 = n170 | n3854 ;
  assign n16800 = n16799 ^ n9790 ^ 1'b0 ;
  assign n16801 = ( n1990 & ~n16213 ) | ( n1990 & n16800 ) | ( ~n16213 & n16800 ) ;
  assign n16802 = n14901 ^ n13715 ^ n4417 ;
  assign n16803 = ( ~n1123 & n12334 ) | ( ~n1123 & n14042 ) | ( n12334 & n14042 ) ;
  assign n16804 = ( n5892 & ~n6279 ) | ( n5892 & n16803 ) | ( ~n6279 & n16803 ) ;
  assign n16805 = n1212 & n3861 ;
  assign n16806 = n9589 & ~n15259 ;
  assign n16807 = n16806 ^ n10191 ^ 1'b0 ;
  assign n16808 = n13073 ^ n9786 ^ n9147 ;
  assign n16809 = n16808 ^ n13179 ^ n7510 ;
  assign n16810 = n5686 | n13766 ;
  assign n16811 = n2454 & n12676 ;
  assign n16812 = ( n189 & ~n10254 ) | ( n189 & n16811 ) | ( ~n10254 & n16811 ) ;
  assign n16813 = n16812 ^ n8553 ^ 1'b0 ;
  assign n16814 = n6861 ^ n5734 ^ n859 ;
  assign n16815 = n1869 & n16814 ;
  assign n16819 = ( n4107 & ~n4872 ) | ( n4107 & n13914 ) | ( ~n4872 & n13914 ) ;
  assign n16820 = n16819 ^ n1942 ^ 1'b0 ;
  assign n16817 = x8 & ~n12312 ;
  assign n16816 = ( n7519 & ~n7935 ) | ( n7519 & n9713 ) | ( ~n7935 & n9713 ) ;
  assign n16818 = n16817 ^ n16816 ^ n1002 ;
  assign n16821 = n16820 ^ n16818 ^ 1'b0 ;
  assign n16822 = ( n8831 & ~n13521 ) | ( n8831 & n16821 ) | ( ~n13521 & n16821 ) ;
  assign n16823 = ( n1651 & n5829 ) | ( n1651 & ~n11402 ) | ( n5829 & ~n11402 ) ;
  assign n16824 = n2140 & ~n6574 ;
  assign n16825 = n11321 & n16824 ;
  assign n16826 = ( ~n1227 & n1862 ) | ( ~n1227 & n8354 ) | ( n1862 & n8354 ) ;
  assign n16827 = ( ~n3985 & n13794 ) | ( ~n3985 & n16826 ) | ( n13794 & n16826 ) ;
  assign n16828 = n2921 & ~n12297 ;
  assign n16829 = n7198 & n16828 ;
  assign n16830 = n2510 | n16829 ;
  assign n16831 = n16827 & ~n16830 ;
  assign n16835 = ( n979 & n2854 ) | ( n979 & ~n3807 ) | ( n2854 & ~n3807 ) ;
  assign n16832 = n3967 ^ n3462 ^ 1'b0 ;
  assign n16833 = n15576 & n16832 ;
  assign n16834 = ( n2670 & n8095 ) | ( n2670 & n16833 ) | ( n8095 & n16833 ) ;
  assign n16836 = n16835 ^ n16834 ^ 1'b0 ;
  assign n16837 = ( ~n1054 & n9561 ) | ( ~n1054 & n16836 ) | ( n9561 & n16836 ) ;
  assign n16838 = n5303 ^ n3662 ^ n623 ;
  assign n16839 = ( n4757 & n8676 ) | ( n4757 & n16838 ) | ( n8676 & n16838 ) ;
  assign n16840 = n5178 ^ n393 ^ 1'b0 ;
  assign n16841 = ( n449 & ~n6633 ) | ( n449 & n16840 ) | ( ~n6633 & n16840 ) ;
  assign n16842 = n13447 ^ n13276 ^ 1'b0 ;
  assign n16843 = n11653 & ~n16842 ;
  assign n16844 = ( n2003 & n3580 ) | ( n2003 & n12798 ) | ( n3580 & n12798 ) ;
  assign n16845 = n16844 ^ n16747 ^ n1834 ;
  assign n16846 = ( n357 & n2159 ) | ( n357 & ~n2675 ) | ( n2159 & ~n2675 ) ;
  assign n16847 = ~n1801 & n4999 ;
  assign n16848 = ~n16846 & n16847 ;
  assign n16849 = n16848 ^ n15241 ^ n9752 ;
  assign n16850 = ~n4015 & n10804 ;
  assign n16851 = n3444 ^ n2120 ^ n194 ;
  assign n16852 = n16851 ^ n11079 ^ n3069 ;
  assign n16853 = n16654 ^ n8336 ^ n3848 ;
  assign n16854 = n16853 ^ n7888 ^ 1'b0 ;
  assign n16855 = n308 | n16854 ;
  assign n16856 = n9216 ^ n182 ^ x47 ;
  assign n16857 = n16856 ^ n9880 ^ n6457 ;
  assign n16858 = n16855 | n16857 ;
  assign n16859 = ~n2878 & n7716 ;
  assign n16860 = n9832 & n16859 ;
  assign n16861 = ( n4306 & ~n4584 ) | ( n4306 & n12876 ) | ( ~n4584 & n12876 ) ;
  assign n16862 = n11941 ^ n2642 ^ 1'b0 ;
  assign n16863 = n16862 ^ n4744 ^ 1'b0 ;
  assign n16864 = n16861 & ~n16863 ;
  assign n16867 = n11535 ^ n5080 ^ n2759 ;
  assign n16868 = n16867 ^ n1865 ^ n1528 ;
  assign n16865 = n8679 ^ n5616 ^ 1'b0 ;
  assign n16866 = n16865 ^ n12937 ^ 1'b0 ;
  assign n16869 = n16868 ^ n16866 ^ n14984 ;
  assign n16870 = ( n9506 & n10845 ) | ( n9506 & n12512 ) | ( n10845 & n12512 ) ;
  assign n16871 = ( n7330 & n14724 ) | ( n7330 & n16870 ) | ( n14724 & n16870 ) ;
  assign n16872 = n6604 ^ n3268 ^ n1834 ;
  assign n16873 = ( ~n277 & n1126 ) | ( ~n277 & n7280 ) | ( n1126 & n7280 ) ;
  assign n16874 = n16873 ^ n14687 ^ n13634 ;
  assign n16875 = ( n8028 & ~n14051 ) | ( n8028 & n16874 ) | ( ~n14051 & n16874 ) ;
  assign n16877 = ( n1326 & ~n3506 ) | ( n1326 & n3676 ) | ( ~n3506 & n3676 ) ;
  assign n16876 = ~n2425 & n7399 ;
  assign n16878 = n16877 ^ n16876 ^ 1'b0 ;
  assign n16879 = n6431 | n13979 ;
  assign n16880 = ( ~n1113 & n2891 ) | ( ~n1113 & n4761 ) | ( n2891 & n4761 ) ;
  assign n16881 = n7533 & ~n10513 ;
  assign n16882 = n16881 ^ n4696 ^ n2810 ;
  assign n16883 = n4601 & n16882 ;
  assign n16884 = ~n16880 & n16883 ;
  assign n16885 = n8674 | n16884 ;
  assign n16886 = n13570 ^ n12166 ^ n1246 ;
  assign n16887 = ( n1534 & ~n3463 ) | ( n1534 & n8121 ) | ( ~n3463 & n8121 ) ;
  assign n16888 = n10996 ^ n8133 ^ n1912 ;
  assign n16889 = ~n1795 & n16218 ;
  assign n16890 = n16888 & n16889 ;
  assign n16891 = n440 & n5518 ;
  assign n16892 = n16891 ^ n1751 ^ 1'b0 ;
  assign n16893 = n16892 ^ n9996 ^ n5602 ;
  assign n16894 = n5432 & ~n11157 ;
  assign n16895 = n16894 ^ n5091 ^ 1'b0 ;
  assign n16896 = ( ~n9624 & n16893 ) | ( ~n9624 & n16895 ) | ( n16893 & n16895 ) ;
  assign n16897 = ( n16887 & ~n16890 ) | ( n16887 & n16896 ) | ( ~n16890 & n16896 ) ;
  assign n16899 = n2656 ^ n1428 ^ 1'b0 ;
  assign n16898 = n5644 | n6186 ;
  assign n16900 = n16899 ^ n16898 ^ 1'b0 ;
  assign n16901 = n13847 ^ n4451 ^ 1'b0 ;
  assign n16902 = ( n2279 & n16900 ) | ( n2279 & n16901 ) | ( n16900 & n16901 ) ;
  assign n16903 = ( n16886 & n16897 ) | ( n16886 & ~n16902 ) | ( n16897 & ~n16902 ) ;
  assign n16904 = ( ~n1785 & n4175 ) | ( ~n1785 & n6524 ) | ( n4175 & n6524 ) ;
  assign n16905 = n16904 ^ n2002 ^ n597 ;
  assign n16906 = n16905 ^ n11735 ^ n3484 ;
  assign n16907 = n15838 ^ n11561 ^ n2002 ;
  assign n16908 = ( ~n1552 & n2916 ) | ( ~n1552 & n4483 ) | ( n2916 & n4483 ) ;
  assign n16909 = ( n4742 & n7316 ) | ( n4742 & ~n16908 ) | ( n7316 & ~n16908 ) ;
  assign n16910 = n11369 ^ n8851 ^ n8338 ;
  assign n16911 = ( n4343 & n4587 ) | ( n4343 & ~n16910 ) | ( n4587 & ~n16910 ) ;
  assign n16912 = n16911 ^ n10006 ^ n1059 ;
  assign n16920 = n11815 ^ n1079 ^ 1'b0 ;
  assign n16921 = n6764 & ~n16920 ;
  assign n16915 = n1804 | n5125 ;
  assign n16916 = n15947 ^ n1848 ^ 1'b0 ;
  assign n16917 = ~n4252 & n16916 ;
  assign n16918 = ( n11383 & ~n16915 ) | ( n11383 & n16917 ) | ( ~n16915 & n16917 ) ;
  assign n16913 = n2369 ^ n2044 ^ n1341 ;
  assign n16914 = n16913 ^ n7453 ^ n596 ;
  assign n16919 = n16918 ^ n16914 ^ 1'b0 ;
  assign n16922 = n16921 ^ n16919 ^ n13068 ;
  assign n16923 = n9739 ^ n5133 ^ n3622 ;
  assign n16924 = n16923 ^ n3474 ^ n1496 ;
  assign n16925 = n16924 ^ n13632 ^ n5307 ;
  assign n16926 = n7918 ^ n2224 ^ 1'b0 ;
  assign n16927 = ~n8320 & n16926 ;
  assign n16928 = n16927 ^ n11304 ^ n3849 ;
  assign n16929 = n15829 ^ n13074 ^ n10233 ;
  assign n16930 = n5950 ^ n5533 ^ n4149 ;
  assign n16931 = n12526 & ~n13331 ;
  assign n16932 = n8950 & n16931 ;
  assign n16933 = n12604 | n16932 ;
  assign n16934 = ( n16570 & ~n16930 ) | ( n16570 & n16933 ) | ( ~n16930 & n16933 ) ;
  assign n16935 = n3707 ^ n2476 ^ 1'b0 ;
  assign n16936 = ( n3869 & n11080 ) | ( n3869 & n16935 ) | ( n11080 & n16935 ) ;
  assign n16937 = ( n9727 & n14640 ) | ( n9727 & n16936 ) | ( n14640 & n16936 ) ;
  assign n16938 = ~n5471 & n16937 ;
  assign n16939 = n10067 ^ n5780 ^ 1'b0 ;
  assign n16940 = n1307 & n16939 ;
  assign n16941 = n15270 ^ n1911 ^ 1'b0 ;
  assign n16942 = ~n16855 & n16941 ;
  assign n16944 = n7489 ^ n3744 ^ n1033 ;
  assign n16943 = ( n265 & n5018 ) | ( n265 & ~n8631 ) | ( n5018 & ~n8631 ) ;
  assign n16945 = n16944 ^ n16943 ^ 1'b0 ;
  assign n16946 = n1463 & n16945 ;
  assign n16947 = n5805 ^ n5754 ^ 1'b0 ;
  assign n16948 = ( n1580 & n4417 ) | ( n1580 & n12794 ) | ( n4417 & n12794 ) ;
  assign n16949 = ( n1780 & n7427 ) | ( n1780 & n16948 ) | ( n7427 & n16948 ) ;
  assign n16950 = ( n1919 & n12541 ) | ( n1919 & ~n14732 ) | ( n12541 & ~n14732 ) ;
  assign n16951 = n8749 ^ n2103 ^ 1'b0 ;
  assign n16952 = ~n3765 & n16951 ;
  assign n16953 = ( n3869 & n12501 ) | ( n3869 & ~n16188 ) | ( n12501 & ~n16188 ) ;
  assign n16954 = ( ~n5063 & n8021 ) | ( ~n5063 & n16953 ) | ( n8021 & n16953 ) ;
  assign n16955 = n3973 & n16954 ;
  assign n16956 = n6547 & n16955 ;
  assign n16957 = n8227 ^ n5235 ^ n4767 ;
  assign n16958 = n3658 | n16957 ;
  assign n16959 = n14116 & ~n16958 ;
  assign n16960 = n12577 ^ n9440 ^ n514 ;
  assign n16961 = ( n3093 & n12835 ) | ( n3093 & ~n15989 ) | ( n12835 & ~n15989 ) ;
  assign n16962 = n10140 ^ n7589 ^ x108 ;
  assign n16963 = n16962 ^ n9460 ^ n8233 ;
  assign n16972 = n2454 & n7066 ;
  assign n16973 = n2526 & n16972 ;
  assign n16974 = n7871 | n16973 ;
  assign n16975 = n6078 | n16974 ;
  assign n16964 = n3730 | n7837 ;
  assign n16965 = n16964 ^ n14096 ^ 1'b0 ;
  assign n16966 = ( n4357 & n7494 ) | ( n4357 & ~n10582 ) | ( n7494 & ~n10582 ) ;
  assign n16967 = n4007 ^ n2781 ^ 1'b0 ;
  assign n16968 = ( n1964 & n12351 ) | ( n1964 & ~n16967 ) | ( n12351 & ~n16967 ) ;
  assign n16969 = n16968 ^ n9945 ^ n7335 ;
  assign n16970 = n16966 & n16969 ;
  assign n16971 = n16965 & n16970 ;
  assign n16976 = n16975 ^ n16971 ^ n4097 ;
  assign n16977 = n7662 ^ n3880 ^ 1'b0 ;
  assign n16978 = n14128 ^ n8956 ^ n5225 ;
  assign n16979 = n12796 ^ n10446 ^ n8198 ;
  assign n16980 = n16979 ^ n4404 ^ n3380 ;
  assign n16981 = ( ~n563 & n12695 ) | ( ~n563 & n16980 ) | ( n12695 & n16980 ) ;
  assign n16982 = n10665 ^ n9026 ^ n6946 ;
  assign n16983 = n3734 & n3795 ;
  assign n16984 = n16983 ^ n3144 ^ 1'b0 ;
  assign n16989 = ( n3188 & ~n6406 ) | ( n3188 & n8751 ) | ( ~n6406 & n8751 ) ;
  assign n16985 = n3673 | n4568 ;
  assign n16986 = n16985 ^ n777 ^ 1'b0 ;
  assign n16987 = n5099 & ~n9084 ;
  assign n16988 = n16986 & n16987 ;
  assign n16990 = n16989 ^ n16988 ^ 1'b0 ;
  assign n16991 = n16984 | n16990 ;
  assign n16992 = n2779 ^ n2210 ^ 1'b0 ;
  assign n16993 = ~n2375 & n16992 ;
  assign n16994 = n16993 ^ n6299 ^ 1'b0 ;
  assign n16995 = n12618 | n16994 ;
  assign n16996 = ~n6935 & n14547 ;
  assign n16997 = n16996 ^ n12346 ^ 1'b0 ;
  assign n16998 = n8012 & n16997 ;
  assign n16999 = n16995 | n16998 ;
  assign n17000 = n5539 ^ n1947 ^ 1'b0 ;
  assign n17001 = n17000 ^ n13580 ^ n3601 ;
  assign n17002 = ( n622 & n1219 ) | ( n622 & ~n17001 ) | ( n1219 & ~n17001 ) ;
  assign n17003 = ( n442 & n12574 ) | ( n442 & ~n17002 ) | ( n12574 & ~n17002 ) ;
  assign n17004 = ( n4137 & n9302 ) | ( n4137 & ~n11169 ) | ( n9302 & ~n11169 ) ;
  assign n17005 = ( n310 & n322 ) | ( n310 & n345 ) | ( n322 & n345 ) ;
  assign n17006 = n17005 ^ n10931 ^ 1'b0 ;
  assign n17010 = ~n587 & n13222 ;
  assign n17007 = n15449 ^ n1662 ^ 1'b0 ;
  assign n17008 = n13387 ^ n443 ^ 1'b0 ;
  assign n17009 = n17007 | n17008 ;
  assign n17011 = n17010 ^ n17009 ^ 1'b0 ;
  assign n17012 = n5245 ^ n1900 ^ n585 ;
  assign n17013 = n16219 ^ n8941 ^ n6161 ;
  assign n17014 = n17013 ^ n12966 ^ 1'b0 ;
  assign n17015 = n17014 ^ n1159 ^ 1'b0 ;
  assign n17016 = ~n17012 & n17015 ;
  assign n17017 = ( n5900 & n15096 ) | ( n5900 & ~n17016 ) | ( n15096 & ~n17016 ) ;
  assign n17018 = ( ~n607 & n2369 ) | ( ~n607 & n12679 ) | ( n2369 & n12679 ) ;
  assign n17019 = n5452 ^ n5249 ^ n3292 ;
  assign n17020 = ( n2771 & ~n2889 ) | ( n2771 & n17019 ) | ( ~n2889 & n17019 ) ;
  assign n17021 = ( n4650 & ~n17018 ) | ( n4650 & n17020 ) | ( ~n17018 & n17020 ) ;
  assign n17022 = ( ~n1619 & n5825 ) | ( ~n1619 & n17021 ) | ( n5825 & n17021 ) ;
  assign n17023 = n14515 ^ n5340 ^ 1'b0 ;
  assign n17024 = n1025 & ~n2972 ;
  assign n17026 = ( n3201 & ~n6565 ) | ( n3201 & n6773 ) | ( ~n6565 & n6773 ) ;
  assign n17025 = n10064 ^ n4587 ^ n1629 ;
  assign n17027 = n17026 ^ n17025 ^ n6489 ;
  assign n17028 = n3321 ^ n264 ^ 1'b0 ;
  assign n17029 = ( n828 & n9237 ) | ( n828 & ~n17028 ) | ( n9237 & ~n17028 ) ;
  assign n17030 = n1248 & n7282 ;
  assign n17031 = n10892 ^ n10058 ^ n3622 ;
  assign n17032 = ( n3860 & ~n11025 ) | ( n3860 & n17031 ) | ( ~n11025 & n17031 ) ;
  assign n17033 = n8078 | n17032 ;
  assign n17034 = n17033 ^ n11238 ^ 1'b0 ;
  assign n17035 = n11373 & ~n13077 ;
  assign n17036 = ( ~n461 & n5135 ) | ( ~n461 & n5793 ) | ( n5135 & n5793 ) ;
  assign n17037 = n11957 & ~n17036 ;
  assign n17041 = n9277 ^ n6202 ^ n3385 ;
  assign n17038 = n14450 ^ n10824 ^ n2271 ;
  assign n17039 = n17038 ^ n15684 ^ 1'b0 ;
  assign n17040 = n12327 & n17039 ;
  assign n17042 = n17041 ^ n17040 ^ 1'b0 ;
  assign n17043 = ~n17037 & n17042 ;
  assign n17044 = ( n8059 & n8240 ) | ( n8059 & n16675 ) | ( n8240 & n16675 ) ;
  assign n17047 = n5465 ^ n3153 ^ n1048 ;
  assign n17045 = ~n4413 & n6374 ;
  assign n17046 = n17045 ^ n17012 ^ 1'b0 ;
  assign n17048 = n17047 ^ n17046 ^ n2355 ;
  assign n17049 = n7842 & ~n8166 ;
  assign n17050 = n4536 | n5733 ;
  assign n17051 = n1745 & ~n17050 ;
  assign n17052 = ( n1114 & n3703 ) | ( n1114 & n16851 ) | ( n3703 & n16851 ) ;
  assign n17053 = n636 & n12696 ;
  assign n17054 = n17052 & n17053 ;
  assign n17055 = ( ~n1069 & n6351 ) | ( ~n1069 & n7778 ) | ( n6351 & n7778 ) ;
  assign n17056 = n14617 | n17055 ;
  assign n17057 = n17056 ^ n5658 ^ 1'b0 ;
  assign n17058 = n2069 & n4891 ;
  assign n17059 = ~n651 & n17058 ;
  assign n17060 = n17059 ^ n11884 ^ n6520 ;
  assign n17063 = n9473 ^ n4022 ^ n132 ;
  assign n17061 = n16155 ^ n9405 ^ 1'b0 ;
  assign n17062 = ( n1045 & n15293 ) | ( n1045 & n17061 ) | ( n15293 & n17061 ) ;
  assign n17064 = n17063 ^ n17062 ^ n12198 ;
  assign n17065 = ( n2480 & n6081 ) | ( n2480 & ~n11202 ) | ( n6081 & ~n11202 ) ;
  assign n17066 = n2036 & n9199 ;
  assign n17067 = n17066 ^ n2309 ^ 1'b0 ;
  assign n17068 = n17067 ^ n14085 ^ n6414 ;
  assign n17069 = n2309 ^ n528 ^ x64 ;
  assign n17070 = ~n1330 & n17069 ;
  assign n17071 = n1690 & n17070 ;
  assign n17072 = ~n3339 & n10098 ;
  assign n17073 = n10547 & n17072 ;
  assign n17074 = n8884 ^ n4788 ^ n1710 ;
  assign n17075 = n7164 & n13417 ;
  assign n17076 = n17075 ^ n11681 ^ 1'b0 ;
  assign n17077 = n4044 & n17076 ;
  assign n17078 = n5439 & n10064 ;
  assign n17079 = n17078 ^ n6524 ^ 1'b0 ;
  assign n17080 = ( n4051 & n5965 ) | ( n4051 & ~n17079 ) | ( n5965 & ~n17079 ) ;
  assign n17081 = n15789 ^ n9771 ^ 1'b0 ;
  assign n17082 = ( x40 & ~n885 ) | ( x40 & n17081 ) | ( ~n885 & n17081 ) ;
  assign n17083 = ( ~n1541 & n2978 ) | ( ~n1541 & n17082 ) | ( n2978 & n17082 ) ;
  assign n17084 = ~n3904 & n9054 ;
  assign n17085 = ( ~n1339 & n3679 ) | ( ~n1339 & n17084 ) | ( n3679 & n17084 ) ;
  assign n17086 = n17085 ^ n1171 ^ 1'b0 ;
  assign n17087 = n13809 & ~n16264 ;
  assign n17088 = n14507 & n17087 ;
  assign n17089 = ( n2917 & n14396 ) | ( n2917 & ~n17088 ) | ( n14396 & ~n17088 ) ;
  assign n17090 = n1972 ^ n1373 ^ 1'b0 ;
  assign n17091 = n10133 & n15686 ;
  assign n17092 = ( ~n7408 & n7972 ) | ( ~n7408 & n17091 ) | ( n7972 & n17091 ) ;
  assign n17093 = n17092 ^ n12892 ^ n1915 ;
  assign n17094 = n17093 ^ n6320 ^ n5174 ;
  assign n17095 = ( n8695 & ~n17090 ) | ( n8695 & n17094 ) | ( ~n17090 & n17094 ) ;
  assign n17096 = n6222 ^ n3256 ^ 1'b0 ;
  assign n17097 = n7502 & n17096 ;
  assign n17098 = n10571 | n12841 ;
  assign n17099 = n17098 ^ n3588 ^ n642 ;
  assign n17100 = ( n4551 & ~n5113 ) | ( n4551 & n7700 ) | ( ~n5113 & n7700 ) ;
  assign n17101 = ~n6458 & n17100 ;
  assign n17102 = n13008 ^ n4844 ^ 1'b0 ;
  assign n17103 = n17102 ^ n8727 ^ n3326 ;
  assign n17108 = ( n2848 & n7332 ) | ( n2848 & ~n9172 ) | ( n7332 & ~n9172 ) ;
  assign n17104 = n8731 ^ n175 ^ 1'b0 ;
  assign n17105 = n1254 & n17104 ;
  assign n17106 = n17105 ^ n11825 ^ 1'b0 ;
  assign n17107 = ~n10170 & n17106 ;
  assign n17109 = n17108 ^ n17107 ^ 1'b0 ;
  assign n17110 = n3641 | n6253 ;
  assign n17111 = n17110 ^ n2452 ^ 1'b0 ;
  assign n17112 = n2573 & n7564 ;
  assign n17113 = ~n17111 & n17112 ;
  assign n17114 = ( n10884 & n13537 ) | ( n10884 & ~n17113 ) | ( n13537 & ~n17113 ) ;
  assign n17115 = n4130 & ~n9873 ;
  assign n17116 = n16681 ^ n13358 ^ 1'b0 ;
  assign n17117 = n904 | n17116 ;
  assign n17118 = n6653 & ~n17117 ;
  assign n17119 = n13857 ^ n5647 ^ 1'b0 ;
  assign n17120 = n4040 | n17119 ;
  assign n17121 = n8065 ^ n1534 ^ 1'b0 ;
  assign n17122 = ( ~n13068 & n17120 ) | ( ~n13068 & n17121 ) | ( n17120 & n17121 ) ;
  assign n17123 = n10246 | n17122 ;
  assign n17124 = n17123 ^ n13224 ^ 1'b0 ;
  assign n17125 = ~n3992 & n4053 ;
  assign n17126 = n9306 ^ n4422 ^ 1'b0 ;
  assign n17127 = ( n685 & n825 ) | ( n685 & n4684 ) | ( n825 & n4684 ) ;
  assign n17128 = n17127 ^ n4326 ^ n1208 ;
  assign n17129 = n13560 ^ n11653 ^ 1'b0 ;
  assign n17130 = n12424 ^ n9595 ^ n1955 ;
  assign n17131 = n17130 ^ n12248 ^ 1'b0 ;
  assign n17132 = n10332 & ~n17131 ;
  assign n17133 = ( ~n6908 & n17129 ) | ( ~n6908 & n17132 ) | ( n17129 & n17132 ) ;
  assign n17134 = n7565 ^ n6569 ^ n1927 ;
  assign n17135 = n3136 | n13772 ;
  assign n17136 = ( n11773 & n17134 ) | ( n11773 & ~n17135 ) | ( n17134 & ~n17135 ) ;
  assign n17138 = n6696 ^ n2061 ^ n192 ;
  assign n17139 = ( ~n12827 & n15020 ) | ( ~n12827 & n17138 ) | ( n15020 & n17138 ) ;
  assign n17137 = n6063 & n6970 ;
  assign n17140 = n17139 ^ n17137 ^ 1'b0 ;
  assign n17141 = n12562 ^ n5311 ^ n3395 ;
  assign n17143 = ~n1557 & n2097 ;
  assign n17144 = ~n5218 & n17143 ;
  assign n17145 = ( ~n6246 & n13651 ) | ( ~n6246 & n17144 ) | ( n13651 & n17144 ) ;
  assign n17142 = n7771 ^ n7415 ^ 1'b0 ;
  assign n17146 = n17145 ^ n17142 ^ 1'b0 ;
  assign n17147 = ( n2839 & n5887 ) | ( n2839 & n13058 ) | ( n5887 & n13058 ) ;
  assign n17148 = n6679 | n15542 ;
  assign n17149 = n17148 ^ n6826 ^ 1'b0 ;
  assign n17150 = x115 | n7633 ;
  assign n17151 = ( n1668 & ~n1728 ) | ( n1668 & n2495 ) | ( ~n1728 & n2495 ) ;
  assign n17152 = n17151 ^ n16595 ^ n13147 ;
  assign n17153 = n13035 ^ n3373 ^ n1942 ;
  assign n17154 = ~n5572 & n17153 ;
  assign n17155 = ~n16176 & n17154 ;
  assign n17156 = ( n5100 & n7468 ) | ( n5100 & ~n10772 ) | ( n7468 & ~n10772 ) ;
  assign n17157 = n11844 ^ n11221 ^ 1'b0 ;
  assign n17158 = n14612 & ~n17157 ;
  assign n17159 = ( n10692 & n17156 ) | ( n10692 & ~n17158 ) | ( n17156 & ~n17158 ) ;
  assign n17160 = ~n9530 & n13323 ;
  assign n17161 = ( ~n3357 & n5324 ) | ( ~n3357 & n5559 ) | ( n5324 & n5559 ) ;
  assign n17162 = n4585 | n9479 ;
  assign n17163 = n17161 | n17162 ;
  assign n17164 = n17160 | n17163 ;
  assign n17165 = n8604 ^ n8342 ^ 1'b0 ;
  assign n17166 = n5197 | n17165 ;
  assign n17167 = n17166 ^ n9550 ^ n1718 ;
  assign n17168 = n2498 ^ n2191 ^ 1'b0 ;
  assign n17169 = x121 & n17168 ;
  assign n17170 = ( n662 & n10835 ) | ( n662 & n17169 ) | ( n10835 & n17169 ) ;
  assign n17171 = ~n6899 & n14333 ;
  assign n17172 = n17076 & n17171 ;
  assign n17173 = ( n10439 & n10488 ) | ( n10439 & ~n15628 ) | ( n10488 & ~n15628 ) ;
  assign n17174 = ( n1766 & ~n3683 ) | ( n1766 & n8730 ) | ( ~n3683 & n8730 ) ;
  assign n17175 = n4252 ^ n840 ^ 1'b0 ;
  assign n17176 = ~n17174 & n17175 ;
  assign n17177 = n7994 & n17176 ;
  assign n17178 = n15978 ^ n1924 ^ n231 ;
  assign n17179 = ( n1765 & ~n6103 ) | ( n1765 & n12472 ) | ( ~n6103 & n12472 ) ;
  assign n17180 = n6344 | n17179 ;
  assign n17181 = n17178 & ~n17180 ;
  assign n17182 = ( n15716 & ~n16778 ) | ( n15716 & n17181 ) | ( ~n16778 & n17181 ) ;
  assign n17183 = n2353 ^ n1400 ^ 1'b0 ;
  assign n17184 = n16295 ^ n7749 ^ 1'b0 ;
  assign n17185 = n6145 | n17184 ;
  assign n17186 = n15406 ^ n4389 ^ 1'b0 ;
  assign n17187 = n17186 ^ n9796 ^ 1'b0 ;
  assign n17188 = n17185 | n17187 ;
  assign n17189 = n17188 ^ n6004 ^ 1'b0 ;
  assign n17190 = n10759 ^ n10349 ^ n8295 ;
  assign n17191 = n8363 & n14517 ;
  assign n17192 = n8431 ^ n2772 ^ n296 ;
  assign n17193 = n17192 ^ n16178 ^ 1'b0 ;
  assign n17194 = ~n11229 & n17193 ;
  assign n17195 = ( n1484 & ~n9769 ) | ( n1484 & n11169 ) | ( ~n9769 & n11169 ) ;
  assign n17196 = n5870 | n13063 ;
  assign n17197 = n17196 ^ n15050 ^ 1'b0 ;
  assign n17198 = n17197 ^ n7633 ^ 1'b0 ;
  assign n17199 = ~n17195 & n17198 ;
  assign n17200 = ( n1946 & ~n3392 ) | ( n1946 & n4491 ) | ( ~n3392 & n4491 ) ;
  assign n17201 = n17200 ^ n15390 ^ n5222 ;
  assign n17202 = ( ~n8491 & n17199 ) | ( ~n8491 & n17201 ) | ( n17199 & n17201 ) ;
  assign n17203 = n10022 | n14445 ;
  assign n17204 = n17202 & ~n17203 ;
  assign n17205 = ~n5864 & n9195 ;
  assign n17206 = ~n4307 & n17205 ;
  assign n17207 = ( n4541 & n4857 ) | ( n4541 & ~n17206 ) | ( n4857 & ~n17206 ) ;
  assign n17208 = ~n14235 & n17207 ;
  assign n17209 = n7083 & n17208 ;
  assign n17210 = n17209 ^ n5201 ^ 1'b0 ;
  assign n17211 = n9806 ^ n8574 ^ 1'b0 ;
  assign n17212 = n11317 ^ n4081 ^ n2074 ;
  assign n17213 = ( n432 & n16711 ) | ( n432 & ~n17212 ) | ( n16711 & ~n17212 ) ;
  assign n17214 = n10494 & n17213 ;
  assign n17215 = ~n17211 & n17214 ;
  assign n17216 = n9397 & ~n17215 ;
  assign n17217 = n17216 ^ n10463 ^ n5321 ;
  assign n17218 = n16125 ^ n136 ^ 1'b0 ;
  assign n17219 = n531 & ~n15444 ;
  assign n17220 = n15331 ^ n10080 ^ n3891 ;
  assign n17221 = n10941 ^ n7512 ^ n3117 ;
  assign n17222 = ~n16126 & n17221 ;
  assign n17223 = n17222 ^ n13908 ^ n5372 ;
  assign n17224 = n4195 ^ n2789 ^ n1908 ;
  assign n17225 = ( ~n1671 & n10646 ) | ( ~n1671 & n17224 ) | ( n10646 & n17224 ) ;
  assign n17226 = ~n1605 & n17225 ;
  assign n17227 = n17226 ^ n8609 ^ 1'b0 ;
  assign n17228 = n5215 | n17227 ;
  assign n17229 = n9705 & ~n17228 ;
  assign n17230 = ( ~n12515 & n14863 ) | ( ~n12515 & n15552 ) | ( n14863 & n15552 ) ;
  assign n17231 = ( n571 & n3174 ) | ( n571 & ~n4671 ) | ( n3174 & ~n4671 ) ;
  assign n17232 = ~n16670 & n17231 ;
  assign n17233 = n2227 ^ n2154 ^ 1'b0 ;
  assign n17234 = ( n921 & n8740 ) | ( n921 & ~n13945 ) | ( n8740 & ~n13945 ) ;
  assign n17235 = n8226 | n16168 ;
  assign n17236 = n17234 | n17235 ;
  assign n17237 = n4651 & ~n10241 ;
  assign n17238 = n2515 & n17237 ;
  assign n17239 = ( n10313 & ~n15806 ) | ( n10313 & n15840 ) | ( ~n15806 & n15840 ) ;
  assign n17240 = ( n5214 & n12201 ) | ( n5214 & ~n17239 ) | ( n12201 & ~n17239 ) ;
  assign n17241 = ( n2172 & n17238 ) | ( n2172 & n17240 ) | ( n17238 & n17240 ) ;
  assign n17242 = n2994 & ~n17241 ;
  assign n17243 = ~n5157 & n17242 ;
  assign n17244 = n15993 ^ n7270 ^ n1185 ;
  assign n17245 = n17244 ^ n6388 ^ n3402 ;
  assign n17246 = ( n3040 & ~n14831 ) | ( n3040 & n17245 ) | ( ~n14831 & n17245 ) ;
  assign n17247 = n10256 ^ n4751 ^ 1'b0 ;
  assign n17248 = ( n2007 & ~n7303 ) | ( n2007 & n8650 ) | ( ~n7303 & n8650 ) ;
  assign n17249 = ( ~n11161 & n17247 ) | ( ~n11161 & n17248 ) | ( n17247 & n17248 ) ;
  assign n17250 = n1686 & ~n4356 ;
  assign n17251 = n14557 & n17250 ;
  assign n17252 = ~n1876 & n16042 ;
  assign n17253 = n17251 & n17252 ;
  assign n17254 = ( n3256 & n13982 ) | ( n3256 & ~n17253 ) | ( n13982 & ~n17253 ) ;
  assign n17255 = ( n5859 & n17249 ) | ( n5859 & n17254 ) | ( n17249 & n17254 ) ;
  assign n17256 = n11871 ^ n11338 ^ n4681 ;
  assign n17257 = n10430 ^ n5142 ^ n4739 ;
  assign n17258 = n3957 ^ n3931 ^ n2926 ;
  assign n17259 = n7317 & n17258 ;
  assign n17260 = n10429 ^ n3205 ^ n919 ;
  assign n17269 = ( n8806 & n11589 ) | ( n8806 & ~n13766 ) | ( n11589 & ~n13766 ) ;
  assign n17263 = n2493 ^ n421 ^ 1'b0 ;
  assign n17264 = n17263 ^ n5699 ^ n2206 ;
  assign n17265 = n12611 & ~n17264 ;
  assign n17266 = n17265 ^ n3198 ^ n2043 ;
  assign n17267 = n14596 ^ n11032 ^ n2693 ;
  assign n17268 = ( n2339 & n17266 ) | ( n2339 & ~n17267 ) | ( n17266 & ~n17267 ) ;
  assign n17261 = n6408 ^ n3155 ^ 1'b0 ;
  assign n17262 = n3472 & n17261 ;
  assign n17270 = n17269 ^ n17268 ^ n17262 ;
  assign n17271 = n6118 ^ n3009 ^ 1'b0 ;
  assign n17272 = ( n1703 & n5080 ) | ( n1703 & ~n9050 ) | ( n5080 & ~n9050 ) ;
  assign n17273 = n17272 ^ n7765 ^ 1'b0 ;
  assign n17274 = ( n9112 & n17271 ) | ( n9112 & ~n17273 ) | ( n17271 & ~n17273 ) ;
  assign n17276 = n4874 ^ n4056 ^ n3270 ;
  assign n17277 = n17276 ^ n1486 ^ 1'b0 ;
  assign n17278 = n380 | n17277 ;
  assign n17279 = n6901 & ~n17278 ;
  assign n17280 = n17279 ^ n4403 ^ 1'b0 ;
  assign n17275 = ( n1339 & n2424 ) | ( n1339 & n7695 ) | ( n2424 & n7695 ) ;
  assign n17281 = n17280 ^ n17275 ^ n15585 ;
  assign n17282 = n12522 ^ n2523 ^ 1'b0 ;
  assign n17283 = n7935 & n17282 ;
  assign n17284 = n17283 ^ n10179 ^ n1934 ;
  assign n17285 = n1753 ^ n462 ^ 1'b0 ;
  assign n17286 = ~n17284 & n17285 ;
  assign n17287 = ~n1849 & n3525 ;
  assign n17288 = n4605 | n4770 ;
  assign n17289 = n17287 & n17288 ;
  assign n17290 = ~n16687 & n17289 ;
  assign n17291 = n7370 ^ n4649 ^ 1'b0 ;
  assign n17292 = ( n4592 & n16761 ) | ( n4592 & n17291 ) | ( n16761 & n17291 ) ;
  assign n17293 = n13848 ^ n5228 ^ 1'b0 ;
  assign n17294 = n7582 | n17293 ;
  assign n17295 = n17294 ^ n9952 ^ n5416 ;
  assign n17296 = ( n7578 & n10214 ) | ( n7578 & n17295 ) | ( n10214 & n17295 ) ;
  assign n17297 = n17296 ^ n8821 ^ n7613 ;
  assign n17298 = n413 | n9811 ;
  assign n17299 = n969 & ~n2634 ;
  assign n17300 = n4270 | n17299 ;
  assign n17301 = n2896 | n17300 ;
  assign n17302 = n7047 ^ n2134 ^ 1'b0 ;
  assign n17303 = n17301 & ~n17302 ;
  assign n17304 = ( ~n5898 & n7867 ) | ( ~n5898 & n8496 ) | ( n7867 & n8496 ) ;
  assign n17305 = n2448 ^ n664 ^ n383 ;
  assign n17306 = n1142 & n17305 ;
  assign n17307 = n17306 ^ n3862 ^ 1'b0 ;
  assign n17308 = ( n5149 & n17304 ) | ( n5149 & n17307 ) | ( n17304 & n17307 ) ;
  assign n17309 = ( ~n1751 & n1779 ) | ( ~n1751 & n3220 ) | ( n1779 & n3220 ) ;
  assign n17310 = n17309 ^ n9133 ^ 1'b0 ;
  assign n17311 = x125 & ~n12090 ;
  assign n17312 = n17311 ^ n12029 ^ 1'b0 ;
  assign n17313 = ( n324 & ~n3931 ) | ( n324 & n4674 ) | ( ~n3931 & n4674 ) ;
  assign n17314 = ( n2514 & ~n16260 ) | ( n2514 & n17313 ) | ( ~n16260 & n17313 ) ;
  assign n17315 = n14780 ^ n4987 ^ 1'b0 ;
  assign n17316 = ( n809 & n1213 ) | ( n809 & n17315 ) | ( n1213 & n17315 ) ;
  assign n17317 = n4480 & n12748 ;
  assign n17318 = n17317 ^ n15567 ^ 1'b0 ;
  assign n17319 = ~n17316 & n17318 ;
  assign n17320 = n17319 ^ n6635 ^ 1'b0 ;
  assign n17321 = n7000 & ~n17320 ;
  assign n17322 = n17321 ^ n14390 ^ 1'b0 ;
  assign n17323 = ( ~n558 & n6120 ) | ( ~n558 & n13955 ) | ( n6120 & n13955 ) ;
  assign n17324 = ( ~n3427 & n6750 ) | ( ~n3427 & n17323 ) | ( n6750 & n17323 ) ;
  assign n17325 = ( n8565 & n14028 ) | ( n8565 & ~n17324 ) | ( n14028 & ~n17324 ) ;
  assign n17326 = ~n1550 & n1948 ;
  assign n17327 = n17326 ^ n5487 ^ 1'b0 ;
  assign n17328 = ( n4623 & ~n5761 ) | ( n4623 & n17327 ) | ( ~n5761 & n17327 ) ;
  assign n17329 = n1515 & n3165 ;
  assign n17331 = ~n4143 & n4378 ;
  assign n17332 = n17331 ^ x14 ^ 1'b0 ;
  assign n17330 = ( n2377 & n3093 ) | ( n2377 & n13214 ) | ( n3093 & n13214 ) ;
  assign n17333 = n17332 ^ n17330 ^ n8015 ;
  assign n17341 = ( n1139 & n4541 ) | ( n1139 & n6222 ) | ( n4541 & n6222 ) ;
  assign n17337 = n5964 ^ x81 ^ 1'b0 ;
  assign n17338 = n1619 | n17337 ;
  assign n17339 = n17338 ^ n12551 ^ 1'b0 ;
  assign n17340 = n2498 | n17339 ;
  assign n17334 = x126 & ~n2222 ;
  assign n17335 = n17334 ^ n15997 ^ n6418 ;
  assign n17336 = n17335 ^ n15277 ^ n7002 ;
  assign n17342 = n17341 ^ n17340 ^ n17336 ;
  assign n17343 = n10866 | n16583 ;
  assign n17346 = n5703 & ~n10525 ;
  assign n17344 = n15368 ^ n4265 ^ n763 ;
  assign n17345 = n17344 ^ n14116 ^ 1'b0 ;
  assign n17347 = n17346 ^ n17345 ^ n1647 ;
  assign n17348 = n17347 ^ n10280 ^ n928 ;
  assign n17349 = ~n360 & n6726 ;
  assign n17350 = ~n3900 & n17349 ;
  assign n17351 = ( n3055 & n13770 ) | ( n3055 & ~n17350 ) | ( n13770 & ~n17350 ) ;
  assign n17352 = n7787 & n17351 ;
  assign n17353 = n17352 ^ x75 ^ 1'b0 ;
  assign n17355 = n4264 ^ n3044 ^ n2403 ;
  assign n17354 = n9160 ^ n7957 ^ 1'b0 ;
  assign n17356 = n17355 ^ n17354 ^ 1'b0 ;
  assign n17357 = ( n2708 & n12090 ) | ( n2708 & n12926 ) | ( n12090 & n12926 ) ;
  assign n17358 = n17357 ^ n12551 ^ n6593 ;
  assign n17359 = ( n7395 & n15818 ) | ( n7395 & ~n17358 ) | ( n15818 & ~n17358 ) ;
  assign n17360 = n4107 & n5139 ;
  assign n17361 = n16440 & n17360 ;
  assign n17362 = n11996 ^ n8958 ^ n187 ;
  assign n17363 = ~n2668 & n11080 ;
  assign n17364 = n1451 & n17363 ;
  assign n17365 = ( n3834 & ~n12227 ) | ( n3834 & n17364 ) | ( ~n12227 & n17364 ) ;
  assign n17366 = ~n3290 & n8934 ;
  assign n17367 = n17366 ^ n17357 ^ n12362 ;
  assign n17368 = n6738 | n12409 ;
  assign n17369 = n1958 | n17368 ;
  assign n17370 = n2282 & ~n12674 ;
  assign n17371 = n17370 ^ n8434 ^ 1'b0 ;
  assign n17372 = ( n5253 & n10145 ) | ( n5253 & ~n10595 ) | ( n10145 & ~n10595 ) ;
  assign n17373 = n17372 ^ n13239 ^ n11993 ;
  assign n17374 = ( n16155 & ~n16623 ) | ( n16155 & n17373 ) | ( ~n16623 & n17373 ) ;
  assign n17375 = n3032 ^ n2620 ^ 1'b0 ;
  assign n17376 = n1857 & n17375 ;
  assign n17377 = ( n6522 & n10267 ) | ( n6522 & n17376 ) | ( n10267 & n17376 ) ;
  assign n17378 = n5731 ^ n5270 ^ n149 ;
  assign n17379 = n17378 ^ n15839 ^ n14649 ;
  assign n17380 = ( n2156 & n17377 ) | ( n2156 & n17379 ) | ( n17377 & n17379 ) ;
  assign n17381 = ~n2191 & n11653 ;
  assign n17382 = n9128 & n17381 ;
  assign n17383 = n159 & ~n3032 ;
  assign n17384 = ( ~n9718 & n17382 ) | ( ~n9718 & n17383 ) | ( n17382 & n17383 ) ;
  assign n17385 = n13154 ^ n1861 ^ 1'b0 ;
  assign n17386 = ( n9880 & n15352 ) | ( n9880 & ~n16164 ) | ( n15352 & ~n16164 ) ;
  assign n17387 = ( ~n5451 & n12403 ) | ( ~n5451 & n14572 ) | ( n12403 & n14572 ) ;
  assign n17388 = n17387 ^ n4836 ^ n4581 ;
  assign n17389 = n17388 ^ n10666 ^ n8618 ;
  assign n17391 = ( ~n7406 & n8316 ) | ( ~n7406 & n13109 ) | ( n8316 & n13109 ) ;
  assign n17392 = n990 | n17391 ;
  assign n17393 = n4878 | n17392 ;
  assign n17394 = ( n4209 & n7710 ) | ( n4209 & n17393 ) | ( n7710 & n17393 ) ;
  assign n17390 = n6652 ^ n3570 ^ 1'b0 ;
  assign n17395 = n17394 ^ n17390 ^ n9458 ;
  assign n17396 = n17395 ^ n14065 ^ n4713 ;
  assign n17397 = ( n552 & n6839 ) | ( n552 & ~n14590 ) | ( n6839 & ~n14590 ) ;
  assign n17398 = n17397 ^ n2882 ^ 1'b0 ;
  assign n17404 = n17028 ^ n7844 ^ n3573 ;
  assign n17405 = ( n9519 & n12257 ) | ( n9519 & ~n17404 ) | ( n12257 & ~n17404 ) ;
  assign n17403 = n4999 & ~n13512 ;
  assign n17406 = n17405 ^ n17403 ^ 1'b0 ;
  assign n17407 = n7788 | n17406 ;
  assign n17402 = ( ~n1322 & n11323 ) | ( ~n1322 & n16567 ) | ( n11323 & n16567 ) ;
  assign n17408 = n17407 ^ n17402 ^ n782 ;
  assign n17401 = n5987 ^ n5244 ^ 1'b0 ;
  assign n17399 = n13700 ^ n7538 ^ 1'b0 ;
  assign n17400 = n17399 ^ n11174 ^ n9895 ;
  assign n17409 = n17408 ^ n17401 ^ n17400 ;
  assign n17410 = n5979 & ~n13996 ;
  assign n17411 = n17410 ^ n14935 ^ 1'b0 ;
  assign n17412 = n15241 ^ n1854 ^ 1'b0 ;
  assign n17413 = n3142 | n17412 ;
  assign n17414 = ( n2959 & ~n9190 ) | ( n2959 & n17413 ) | ( ~n9190 & n17413 ) ;
  assign n17415 = n11393 & ~n17414 ;
  assign n17416 = ~n17411 & n17415 ;
  assign n17417 = n11886 ^ n268 ^ 1'b0 ;
  assign n17419 = n1682 & ~n13273 ;
  assign n17420 = ~n1171 & n17419 ;
  assign n17418 = n7778 ^ n6419 ^ n3599 ;
  assign n17421 = n17420 ^ n17418 ^ n17081 ;
  assign n17422 = n2402 & ~n8548 ;
  assign n17423 = n17422 ^ n4959 ^ 1'b0 ;
  assign n17424 = n17423 ^ n8935 ^ n3534 ;
  assign n17425 = n1228 ^ n663 ^ 1'b0 ;
  assign n17426 = n927 & n17425 ;
  assign n17427 = ( ~n1929 & n13639 ) | ( ~n1929 & n17426 ) | ( n13639 & n17426 ) ;
  assign n17428 = n16291 ^ n14272 ^ n4256 ;
  assign n17431 = n4050 ^ n2572 ^ n345 ;
  assign n17432 = n811 & n6456 ;
  assign n17433 = ~n8949 & n17432 ;
  assign n17434 = ( n4030 & ~n16507 ) | ( n4030 & n17433 ) | ( ~n16507 & n17433 ) ;
  assign n17435 = ( n8711 & n17431 ) | ( n8711 & n17434 ) | ( n17431 & n17434 ) ;
  assign n17429 = x2 & ~n2398 ;
  assign n17430 = n17429 ^ n16835 ^ n13332 ;
  assign n17436 = n17435 ^ n17430 ^ 1'b0 ;
  assign n17437 = n2908 | n17436 ;
  assign n17439 = n11535 ^ n3682 ^ n2950 ;
  assign n17440 = n2429 & n5485 ;
  assign n17441 = ~n10448 & n17440 ;
  assign n17442 = n17441 ^ n4828 ^ n4338 ;
  assign n17443 = n17442 ^ n4738 ^ n840 ;
  assign n17444 = ( n7551 & n17439 ) | ( n7551 & ~n17443 ) | ( n17439 & ~n17443 ) ;
  assign n17438 = n646 & n9016 ;
  assign n17445 = n17444 ^ n17438 ^ 1'b0 ;
  assign n17446 = ~n1543 & n6325 ;
  assign n17447 = ( n5851 & ~n6912 ) | ( n5851 & n7986 ) | ( ~n6912 & n7986 ) ;
  assign n17448 = ( n3123 & n9800 ) | ( n3123 & n17447 ) | ( n9800 & n17447 ) ;
  assign n17449 = ( n3305 & ~n7243 ) | ( n3305 & n7265 ) | ( ~n7243 & n7265 ) ;
  assign n17450 = ( ~n4785 & n12165 ) | ( ~n4785 & n17449 ) | ( n12165 & n17449 ) ;
  assign n17451 = ( n5732 & n15719 ) | ( n5732 & n17450 ) | ( n15719 & n17450 ) ;
  assign n17452 = ( n4446 & n8421 ) | ( n4446 & n17451 ) | ( n8421 & n17451 ) ;
  assign n17453 = n17452 ^ n8207 ^ 1'b0 ;
  assign n17454 = n331 & ~n17453 ;
  assign n17455 = n17448 & n17454 ;
  assign n17456 = n17455 ^ n15304 ^ 1'b0 ;
  assign n17457 = n1764 & n6940 ;
  assign n17458 = ~n8571 & n12501 ;
  assign n17459 = n9264 | n17458 ;
  assign n17460 = x100 | n17459 ;
  assign n17461 = n17460 ^ n11445 ^ n2113 ;
  assign n17462 = ( ~n666 & n12300 ) | ( ~n666 & n15620 ) | ( n12300 & n15620 ) ;
  assign n17463 = n8718 ^ n7613 ^ n5689 ;
  assign n17464 = ( n2373 & ~n7141 ) | ( n2373 & n10309 ) | ( ~n7141 & n10309 ) ;
  assign n17465 = n5761 & ~n17464 ;
  assign n17466 = n17465 ^ n6546 ^ 1'b0 ;
  assign n17467 = n17463 & ~n17466 ;
  assign n17468 = n7306 ^ n6187 ^ n2077 ;
  assign n17469 = n2144 & ~n2495 ;
  assign n17470 = n17469 ^ n17156 ^ n13362 ;
  assign n17471 = n17470 ^ n1312 ^ 1'b0 ;
  assign n17472 = n17468 & n17471 ;
  assign n17473 = ( n409 & n2671 ) | ( n409 & ~n17200 ) | ( n2671 & ~n17200 ) ;
  assign n17474 = n7266 & ~n8852 ;
  assign n17475 = n17473 & n17474 ;
  assign n17476 = n17475 ^ n14170 ^ n8191 ;
  assign n17482 = n3577 & n5209 ;
  assign n17477 = n416 | n459 ;
  assign n17478 = n17477 ^ n2832 ^ 1'b0 ;
  assign n17479 = n17478 ^ n8855 ^ 1'b0 ;
  assign n17480 = ( ~n14761 & n14948 ) | ( ~n14761 & n17479 ) | ( n14948 & n17479 ) ;
  assign n17481 = n1738 & ~n17480 ;
  assign n17483 = n17482 ^ n17481 ^ n1096 ;
  assign n17484 = n17483 ^ n11942 ^ n1326 ;
  assign n17485 = n2204 & ~n17484 ;
  assign n17486 = ~n1507 & n6221 ;
  assign n17487 = n17486 ^ n5310 ^ 1'b0 ;
  assign n17488 = n3284 & ~n3976 ;
  assign n17489 = n2125 & ~n17488 ;
  assign n17490 = ( ~n2801 & n17487 ) | ( ~n2801 & n17489 ) | ( n17487 & n17489 ) ;
  assign n17494 = n1212 & n14319 ;
  assign n17495 = ~n8080 & n17494 ;
  assign n17496 = n17495 ^ n3981 ^ 1'b0 ;
  assign n17491 = n5629 & ~n15144 ;
  assign n17492 = ~n5510 & n17491 ;
  assign n17493 = ( ~n3782 & n16299 ) | ( ~n3782 & n17492 ) | ( n16299 & n17492 ) ;
  assign n17497 = n17496 ^ n17493 ^ n6487 ;
  assign n17498 = n16403 ^ n9776 ^ n6578 ;
  assign n17499 = n2079 & n6218 ;
  assign n17500 = n17499 ^ n1679 ^ 1'b0 ;
  assign n17501 = ( n4257 & n15036 ) | ( n4257 & n17500 ) | ( n15036 & n17500 ) ;
  assign n17502 = ( ~n3677 & n8369 ) | ( ~n3677 & n9215 ) | ( n8369 & n9215 ) ;
  assign n17503 = n17502 ^ n3354 ^ n619 ;
  assign n17504 = n9182 | n16436 ;
  assign n17505 = n6960 | n17504 ;
  assign n17506 = n10411 ^ n4164 ^ 1'b0 ;
  assign n17507 = n282 & ~n17506 ;
  assign n17508 = ~n6347 & n17507 ;
  assign n17510 = n6475 ^ n1882 ^ n1450 ;
  assign n17509 = n10429 ^ n8541 ^ n524 ;
  assign n17511 = n17510 ^ n17509 ^ n8029 ;
  assign n17512 = ( n4804 & ~n7475 ) | ( n4804 & n12523 ) | ( ~n7475 & n12523 ) ;
  assign n17513 = n17512 ^ n13509 ^ 1'b0 ;
  assign n17514 = ( ~n411 & n3254 ) | ( ~n411 & n3730 ) | ( n3254 & n3730 ) ;
  assign n17517 = n4587 | n9096 ;
  assign n17518 = n17517 ^ n2870 ^ 1'b0 ;
  assign n17516 = n3470 ^ n744 ^ 1'b0 ;
  assign n17515 = x45 & ~n5051 ;
  assign n17519 = n17518 ^ n17516 ^ n17515 ;
  assign n17520 = ~n17514 & n17519 ;
  assign n17521 = n14803 ^ n13832 ^ 1'b0 ;
  assign n17522 = n15791 ^ n11034 ^ 1'b0 ;
  assign n17523 = n5344 ^ n5220 ^ n4249 ;
  assign n17524 = n2895 | n17523 ;
  assign n17529 = n7439 ^ n3911 ^ n3464 ;
  assign n17530 = ( x41 & n2954 ) | ( x41 & n17529 ) | ( n2954 & n17529 ) ;
  assign n17531 = ( ~n319 & n6600 ) | ( ~n319 & n17530 ) | ( n6600 & n17530 ) ;
  assign n17525 = n10721 ^ n5313 ^ 1'b0 ;
  assign n17526 = n15361 ^ n600 ^ 1'b0 ;
  assign n17527 = ( n4566 & n17525 ) | ( n4566 & n17526 ) | ( n17525 & n17526 ) ;
  assign n17528 = n17527 ^ n13449 ^ 1'b0 ;
  assign n17532 = n17531 ^ n17528 ^ n15335 ;
  assign n17533 = ( x16 & n7909 ) | ( x16 & n14654 ) | ( n7909 & n14654 ) ;
  assign n17534 = n10673 ^ n4962 ^ 1'b0 ;
  assign n17535 = n15864 ^ n5738 ^ n5245 ;
  assign n17536 = n17535 ^ n14936 ^ n204 ;
  assign n17537 = ~n17534 & n17536 ;
  assign n17538 = ( n3422 & n6617 ) | ( n3422 & ~n10582 ) | ( n6617 & ~n10582 ) ;
  assign n17539 = n3518 ^ n2370 ^ 1'b0 ;
  assign n17540 = n11476 & ~n17539 ;
  assign n17541 = ( n3155 & n7953 ) | ( n3155 & n17540 ) | ( n7953 & n17540 ) ;
  assign n17545 = n5658 & n17276 ;
  assign n17542 = ( n3366 & ~n3955 ) | ( n3366 & n7628 ) | ( ~n3955 & n7628 ) ;
  assign n17543 = n17542 ^ n3454 ^ n2443 ;
  assign n17544 = n8483 & ~n17543 ;
  assign n17546 = n17545 ^ n17544 ^ n2237 ;
  assign n17547 = n17546 ^ x96 ^ 1'b0 ;
  assign n17548 = n17547 ^ n9524 ^ 1'b0 ;
  assign n17549 = n17541 | n17548 ;
  assign n17550 = n17538 & ~n17549 ;
  assign n17552 = ( n1440 & n9998 ) | ( n1440 & n14946 ) | ( n9998 & n14946 ) ;
  assign n17551 = ( n11398 & n11681 ) | ( n11398 & n11773 ) | ( n11681 & n11773 ) ;
  assign n17553 = n17552 ^ n17551 ^ n1141 ;
  assign n17554 = ( n1966 & ~n5696 ) | ( n1966 & n10359 ) | ( ~n5696 & n10359 ) ;
  assign n17555 = n5868 | n17554 ;
  assign n17556 = n1582 & ~n17555 ;
  assign n17557 = n17556 ^ n1703 ^ 1'b0 ;
  assign n17558 = n17557 ^ n6201 ^ n4490 ;
  assign n17559 = n17553 | n17558 ;
  assign n17560 = n15927 ^ n10767 ^ 1'b0 ;
  assign n17561 = n3811 | n3860 ;
  assign n17562 = n17561 ^ n7350 ^ 1'b0 ;
  assign n17563 = n17562 ^ n9402 ^ n2614 ;
  assign n17564 = n17563 ^ n7901 ^ n5698 ;
  assign n17565 = n4457 ^ n2762 ^ 1'b0 ;
  assign n17566 = n17565 ^ n16965 ^ n3188 ;
  assign n17567 = n7812 | n17413 ;
  assign n17568 = n5252 ^ n1246 ^ 1'b0 ;
  assign n17569 = n16136 & ~n17568 ;
  assign n17570 = n11828 ^ n11805 ^ 1'b0 ;
  assign n17571 = ( ~n8057 & n12834 ) | ( ~n8057 & n14233 ) | ( n12834 & n14233 ) ;
  assign n17572 = ( n2421 & n2513 ) | ( n2421 & n7986 ) | ( n2513 & n7986 ) ;
  assign n17573 = n5270 ^ n183 ^ 1'b0 ;
  assign n17574 = ~n15171 & n17573 ;
  assign n17575 = ( ~n5100 & n9300 ) | ( ~n5100 & n11078 ) | ( n9300 & n11078 ) ;
  assign n17576 = ( ~n1956 & n5368 ) | ( ~n1956 & n17575 ) | ( n5368 & n17575 ) ;
  assign n17577 = n10364 ^ n8215 ^ 1'b0 ;
  assign n17578 = ( n2951 & n10831 ) | ( n2951 & n17473 ) | ( n10831 & n17473 ) ;
  assign n17579 = ( n4760 & ~n8324 ) | ( n4760 & n9380 ) | ( ~n8324 & n9380 ) ;
  assign n17580 = n7878 | n17579 ;
  assign n17581 = n13886 ^ n8038 ^ n4390 ;
  assign n17582 = ( n1058 & n1755 ) | ( n1058 & ~n17581 ) | ( n1755 & ~n17581 ) ;
  assign n17583 = ~n2586 & n6018 ;
  assign n17584 = n17583 ^ n11719 ^ 1'b0 ;
  assign n17585 = ( ~n6314 & n17582 ) | ( ~n6314 & n17584 ) | ( n17582 & n17584 ) ;
  assign n17586 = ( n2190 & ~n2776 ) | ( n2190 & n6709 ) | ( ~n2776 & n6709 ) ;
  assign n17587 = n11093 & n17586 ;
  assign n17588 = n10178 & n17587 ;
  assign n17589 = n14832 ^ n10907 ^ 1'b0 ;
  assign n17590 = ( n5264 & ~n7015 ) | ( n5264 & n11120 ) | ( ~n7015 & n11120 ) ;
  assign n17591 = n17589 | n17590 ;
  assign n17592 = n17588 & ~n17591 ;
  assign n17593 = ( n1040 & ~n4957 ) | ( n1040 & n14125 ) | ( ~n4957 & n14125 ) ;
  assign n17594 = n7220 & n17593 ;
  assign n17595 = ~n919 & n17594 ;
  assign n17596 = n9064 | n11931 ;
  assign n17597 = n4771 & ~n17596 ;
  assign n17598 = n2554 & ~n4468 ;
  assign n17599 = ~n970 & n17598 ;
  assign n17600 = n17597 | n17599 ;
  assign n17601 = n10461 | n17600 ;
  assign n17602 = n17601 ^ n13546 ^ n9626 ;
  assign n17604 = ( n4502 & n9286 ) | ( n4502 & ~n15885 ) | ( n9286 & ~n15885 ) ;
  assign n17605 = ( n465 & n524 ) | ( n465 & ~n3198 ) | ( n524 & ~n3198 ) ;
  assign n17606 = ( n11058 & ~n17604 ) | ( n11058 & n17605 ) | ( ~n17604 & n17605 ) ;
  assign n17607 = n17606 ^ n11986 ^ n1348 ;
  assign n17608 = n2045 ^ n1235 ^ x21 ;
  assign n17609 = n11264 & ~n17608 ;
  assign n17610 = ( ~n13381 & n17607 ) | ( ~n13381 & n17609 ) | ( n17607 & n17609 ) ;
  assign n17603 = n13658 | n13940 ;
  assign n17611 = n17610 ^ n17603 ^ 1'b0 ;
  assign n17612 = n3938 ^ n1028 ^ 1'b0 ;
  assign n17613 = n4628 & n17612 ;
  assign n17614 = n17613 ^ n8688 ^ n3835 ;
  assign n17615 = n16351 ^ n4467 ^ 1'b0 ;
  assign n17616 = n7153 & ~n17615 ;
  assign n17617 = n17616 ^ n10632 ^ n5849 ;
  assign n17618 = ( n5305 & ~n5714 ) | ( n5305 & n6430 ) | ( ~n5714 & n6430 ) ;
  assign n17619 = n13732 & n17618 ;
  assign n17620 = ( n4179 & n11371 ) | ( n4179 & n17619 ) | ( n11371 & n17619 ) ;
  assign n17621 = n12307 ^ n1273 ^ 1'b0 ;
  assign n17622 = n3305 ^ n2775 ^ n516 ;
  assign n17623 = ( n5661 & ~n12792 ) | ( n5661 & n14459 ) | ( ~n12792 & n14459 ) ;
  assign n17624 = n5690 & n8868 ;
  assign n17625 = n6126 & ~n17624 ;
  assign n17626 = ~n17623 & n17625 ;
  assign n17627 = n12725 ^ n1216 ^ 1'b0 ;
  assign n17628 = n7427 ^ n1336 ^ 1'b0 ;
  assign n17629 = n5455 & n17628 ;
  assign n17630 = ~n11218 & n17629 ;
  assign n17631 = ~n7439 & n8081 ;
  assign n17632 = n17631 ^ n600 ^ 1'b0 ;
  assign n17633 = ( ~n14396 & n16216 ) | ( ~n14396 & n17632 ) | ( n16216 & n17632 ) ;
  assign n17634 = ( n8889 & n17630 ) | ( n8889 & n17633 ) | ( n17630 & n17633 ) ;
  assign n17635 = n5735 & n12944 ;
  assign n17636 = ( n6344 & n8156 ) | ( n6344 & n10959 ) | ( n8156 & n10959 ) ;
  assign n17637 = ~n17635 & n17636 ;
  assign n17638 = n17637 ^ n9238 ^ n6714 ;
  assign n17639 = ( n1934 & ~n10730 ) | ( n1934 & n15615 ) | ( ~n10730 & n15615 ) ;
  assign n17640 = ( ~n708 & n11705 ) | ( ~n708 & n11892 ) | ( n11705 & n11892 ) ;
  assign n17641 = n17640 ^ n11676 ^ n11238 ;
  assign n17642 = ~n315 & n377 ;
  assign n17643 = ( n4623 & n11623 ) | ( n4623 & n17642 ) | ( n11623 & n17642 ) ;
  assign n17644 = ( n3928 & ~n7560 ) | ( n3928 & n8170 ) | ( ~n7560 & n8170 ) ;
  assign n17645 = ( n6082 & n17643 ) | ( n6082 & n17644 ) | ( n17643 & n17644 ) ;
  assign n17646 = n4966 & ~n6099 ;
  assign n17647 = n17645 & n17646 ;
  assign n17648 = ( n2542 & n5554 ) | ( n2542 & n17647 ) | ( n5554 & n17647 ) ;
  assign n17649 = n17648 ^ n13665 ^ n4101 ;
  assign n17650 = n7036 ^ n4048 ^ 1'b0 ;
  assign n17651 = ( n975 & ~n10907 ) | ( n975 & n10938 ) | ( ~n10907 & n10938 ) ;
  assign n17652 = n10922 & ~n17651 ;
  assign n17653 = ~n17650 & n17652 ;
  assign n17654 = n10665 ^ n6426 ^ n754 ;
  assign n17657 = n7382 | n10377 ;
  assign n17655 = n8241 ^ n2209 ^ 1'b0 ;
  assign n17656 = n12544 | n17655 ;
  assign n17658 = n17657 ^ n17656 ^ 1'b0 ;
  assign n17659 = ~n17654 & n17658 ;
  assign n17660 = n14696 ^ n6004 ^ 1'b0 ;
  assign n17662 = ( ~n6635 & n9590 ) | ( ~n6635 & n11574 ) | ( n9590 & n11574 ) ;
  assign n17663 = n13435 & n17662 ;
  assign n17661 = ~n1983 & n5100 ;
  assign n17664 = n17663 ^ n17661 ^ n7115 ;
  assign n17666 = n8900 & ~n10336 ;
  assign n17667 = n17666 ^ n5849 ^ 1'b0 ;
  assign n17665 = ~n2353 & n10028 ;
  assign n17668 = n17667 ^ n17665 ^ n2366 ;
  assign n17670 = n11568 ^ n9544 ^ n7705 ;
  assign n17669 = n2800 | n10556 ;
  assign n17671 = n17670 ^ n17669 ^ 1'b0 ;
  assign n17672 = n5629 | n13719 ;
  assign n17673 = n17671 & ~n17672 ;
  assign n17678 = n6972 ^ n5369 ^ n2341 ;
  assign n17674 = n9767 ^ n2360 ^ n1486 ;
  assign n17675 = n8917 ^ n4883 ^ 1'b0 ;
  assign n17676 = n17674 & n17675 ;
  assign n17677 = ~n6282 & n17676 ;
  assign n17679 = n17678 ^ n17677 ^ 1'b0 ;
  assign n17682 = ( n3288 & n3843 ) | ( n3288 & n12922 ) | ( n3843 & n12922 ) ;
  assign n17680 = n3312 ^ n1294 ^ 1'b0 ;
  assign n17681 = ( n4775 & n13451 ) | ( n4775 & n17680 ) | ( n13451 & n17680 ) ;
  assign n17683 = n17682 ^ n17681 ^ n1005 ;
  assign n17684 = n12827 ^ n6355 ^ n5470 ;
  assign n17685 = n7240 & n9911 ;
  assign n17686 = n17685 ^ n15593 ^ 1'b0 ;
  assign n17687 = n17686 ^ n6549 ^ n947 ;
  assign n17688 = ~n2545 & n5009 ;
  assign n17689 = ( n9215 & ~n10654 ) | ( n9215 & n17688 ) | ( ~n10654 & n17688 ) ;
  assign n17690 = n8254 ^ n3057 ^ 1'b0 ;
  assign n17691 = n17690 ^ n9672 ^ n3579 ;
  assign n17692 = n8629 ^ n8383 ^ 1'b0 ;
  assign n17693 = ~n186 & n15061 ;
  assign n17694 = n2876 & n9530 ;
  assign n17695 = n2275 & n17694 ;
  assign n17696 = ( n5668 & n16371 ) | ( n5668 & n17695 ) | ( n16371 & n17695 ) ;
  assign n17697 = n13147 ^ n2771 ^ 1'b0 ;
  assign n17698 = n912 & n17697 ;
  assign n17699 = n8382 ^ n4279 ^ n2832 ;
  assign n17700 = n17699 ^ n3373 ^ 1'b0 ;
  assign n17701 = n2405 | n17700 ;
  assign n17702 = n9865 & ~n17701 ;
  assign n17703 = n901 & n17702 ;
  assign n17704 = n17698 & n17703 ;
  assign n17705 = n17704 ^ n14118 ^ n8686 ;
  assign n17706 = n5554 ^ n5383 ^ 1'b0 ;
  assign n17709 = n1911 & ~n7173 ;
  assign n17710 = ~n9404 & n17709 ;
  assign n17707 = n9029 ^ n3798 ^ n278 ;
  assign n17708 = ~n14046 & n17707 ;
  assign n17711 = n17710 ^ n17708 ^ 1'b0 ;
  assign n17712 = ( n1268 & n17706 ) | ( n1268 & ~n17711 ) | ( n17706 & ~n17711 ) ;
  assign n17713 = ( n1498 & n7437 ) | ( n1498 & ~n7471 ) | ( n7437 & ~n7471 ) ;
  assign n17714 = n17713 ^ n14128 ^ n13183 ;
  assign n17715 = n12635 ^ n3642 ^ n774 ;
  assign n17716 = ( n405 & n1345 ) | ( n405 & n17715 ) | ( n1345 & n17715 ) ;
  assign n17717 = ( ~n907 & n14961 ) | ( ~n907 & n17716 ) | ( n14961 & n17716 ) ;
  assign n17718 = n14429 & ~n16833 ;
  assign n17719 = n17718 ^ n8384 ^ n3942 ;
  assign n17720 = n12864 ^ n8033 ^ n1150 ;
  assign n17721 = n17720 ^ n13492 ^ n4862 ;
  assign n17722 = ( n838 & n2716 ) | ( n838 & ~n10423 ) | ( n2716 & ~n10423 ) ;
  assign n17723 = ~n6896 & n7641 ;
  assign n17724 = ~n3370 & n17723 ;
  assign n17725 = ( n4396 & n6598 ) | ( n4396 & ~n17724 ) | ( n6598 & ~n17724 ) ;
  assign n17726 = n2893 | n17725 ;
  assign n17727 = n17726 ^ x21 ^ 1'b0 ;
  assign n17728 = ( n1868 & n10293 ) | ( n1868 & ~n17727 ) | ( n10293 & ~n17727 ) ;
  assign n17729 = n17728 ^ n7046 ^ n7023 ;
  assign n17730 = n17729 ^ n15091 ^ n1071 ;
  assign n17731 = n4540 ^ n3402 ^ n1627 ;
  assign n17732 = n17731 ^ n11504 ^ n8136 ;
  assign n17733 = ( n2747 & ~n7992 ) | ( n2747 & n11222 ) | ( ~n7992 & n11222 ) ;
  assign n17734 = n17733 ^ n10294 ^ n805 ;
  assign n17735 = n2050 ^ n1967 ^ n1287 ;
  assign n17736 = n3773 ^ n2757 ^ 1'b0 ;
  assign n17737 = n17735 & ~n17736 ;
  assign n17738 = n8236 ^ n6092 ^ 1'b0 ;
  assign n17739 = n17738 ^ n8074 ^ n921 ;
  assign n17740 = ( ~n7519 & n17737 ) | ( ~n7519 & n17739 ) | ( n17737 & n17739 ) ;
  assign n17741 = n5414 ^ n2554 ^ n1276 ;
  assign n17742 = ( n5965 & ~n10652 ) | ( n5965 & n17542 ) | ( ~n10652 & n17542 ) ;
  assign n17743 = n8257 ^ n2388 ^ 1'b0 ;
  assign n17744 = n17742 & ~n17743 ;
  assign n17745 = n17744 ^ n7451 ^ 1'b0 ;
  assign n17746 = n2409 & n17745 ;
  assign n17747 = ( n7569 & ~n12576 ) | ( n7569 & n17746 ) | ( ~n12576 & n17746 ) ;
  assign n17748 = ( ~x68 & n2181 ) | ( ~x68 & n13567 ) | ( n2181 & n13567 ) ;
  assign n17749 = n4528 | n9119 ;
  assign n17750 = n17749 ^ n5602 ^ n2941 ;
  assign n17751 = n17738 ^ n6249 ^ 1'b0 ;
  assign n17752 = n14078 ^ n10803 ^ n6726 ;
  assign n17753 = n7153 & n13306 ;
  assign n17754 = ~n17752 & n17753 ;
  assign n17755 = ( n3926 & n8078 ) | ( n3926 & ~n17754 ) | ( n8078 & ~n17754 ) ;
  assign n17756 = n17755 ^ n739 ^ 1'b0 ;
  assign n17757 = n8592 & ~n17756 ;
  assign n17758 = ( n2198 & ~n5976 ) | ( n2198 & n11381 ) | ( ~n5976 & n11381 ) ;
  assign n17759 = n3616 ^ n1589 ^ x24 ;
  assign n17760 = n4889 | n9482 ;
  assign n17761 = n17759 | n17760 ;
  assign n17762 = n17761 ^ n11754 ^ n3861 ;
  assign n17763 = ( ~n7718 & n17758 ) | ( ~n7718 & n17762 ) | ( n17758 & n17762 ) ;
  assign n17764 = ( n9460 & ~n9824 ) | ( n9460 & n11111 ) | ( ~n9824 & n11111 ) ;
  assign n17771 = n2155 & ~n9869 ;
  assign n17765 = n582 & ~n12522 ;
  assign n17766 = n17765 ^ n4223 ^ 1'b0 ;
  assign n17767 = ( n5012 & ~n6850 ) | ( n5012 & n17766 ) | ( ~n6850 & n17766 ) ;
  assign n17768 = n17767 ^ n6893 ^ n6045 ;
  assign n17769 = n5659 & ~n17768 ;
  assign n17770 = ( ~n9462 & n13982 ) | ( ~n9462 & n17769 ) | ( n13982 & n17769 ) ;
  assign n17772 = n17771 ^ n17770 ^ 1'b0 ;
  assign n17773 = n4731 & n17772 ;
  assign n17774 = ~n6840 & n16590 ;
  assign n17778 = n13614 ^ n9382 ^ n6343 ;
  assign n17776 = ( n8398 & ~n9638 ) | ( n8398 & n13731 ) | ( ~n9638 & n13731 ) ;
  assign n17777 = n17776 ^ n4015 ^ n3032 ;
  assign n17775 = n10092 & n17510 ;
  assign n17779 = n17778 ^ n17777 ^ n17775 ;
  assign n17780 = ( n8637 & n11779 ) | ( n8637 & n16868 ) | ( n11779 & n16868 ) ;
  assign n17781 = n15276 ^ n13034 ^ n7481 ;
  assign n17782 = n17781 ^ n9354 ^ 1'b0 ;
  assign n17783 = n5236 | n12537 ;
  assign n17784 = n17783 ^ n15808 ^ 1'b0 ;
  assign n17785 = n9054 ^ n4724 ^ n3711 ;
  assign n17786 = n13372 ^ n1934 ^ n1413 ;
  assign n17787 = n17786 ^ n8061 ^ 1'b0 ;
  assign n17788 = ( ~n6347 & n9301 ) | ( ~n6347 & n17787 ) | ( n9301 & n17787 ) ;
  assign n17789 = ( n16619 & n17234 ) | ( n16619 & n17788 ) | ( n17234 & n17788 ) ;
  assign n17790 = ( n2914 & n17785 ) | ( n2914 & ~n17789 ) | ( n17785 & ~n17789 ) ;
  assign n17791 = n700 & ~n11405 ;
  assign n17792 = ( n12108 & n16426 ) | ( n12108 & n17791 ) | ( n16426 & n17791 ) ;
  assign n17793 = ( n8036 & n13769 ) | ( n8036 & ~n17792 ) | ( n13769 & ~n17792 ) ;
  assign n17794 = ~n6876 & n13667 ;
  assign n17795 = ( n531 & n3199 ) | ( n531 & ~n11583 ) | ( n3199 & ~n11583 ) ;
  assign n17796 = ( n1003 & n2772 ) | ( n1003 & ~n2922 ) | ( n2772 & ~n2922 ) ;
  assign n17797 = n5900 ^ n1863 ^ 1'b0 ;
  assign n17798 = n12357 & ~n17797 ;
  assign n17799 = n2302 & n17798 ;
  assign n17800 = ~n17796 & n17799 ;
  assign n17801 = ( n3946 & n17795 ) | ( n3946 & ~n17800 ) | ( n17795 & ~n17800 ) ;
  assign n17802 = n17801 ^ n10305 ^ 1'b0 ;
  assign n17803 = ~n5259 & n17802 ;
  assign n17804 = n17803 ^ n6221 ^ n4356 ;
  assign n17805 = ( n3094 & ~n10687 ) | ( n3094 & n16726 ) | ( ~n10687 & n16726 ) ;
  assign n17806 = n1973 | n16541 ;
  assign n17807 = ( ~n2931 & n3886 ) | ( ~n2931 & n4001 ) | ( n3886 & n4001 ) ;
  assign n17808 = n7721 ^ n5315 ^ n5149 ;
  assign n17809 = n9116 ^ n1606 ^ 1'b0 ;
  assign n17810 = n17808 | n17809 ;
  assign n17811 = n17807 | n17810 ;
  assign n17812 = n9173 | n17811 ;
  assign n17813 = ( n6890 & n15128 ) | ( n6890 & n15451 ) | ( n15128 & n15451 ) ;
  assign n17814 = n15347 ^ n9086 ^ 1'b0 ;
  assign n17815 = ( n2049 & n17813 ) | ( n2049 & ~n17814 ) | ( n17813 & ~n17814 ) ;
  assign n17817 = n2102 & ~n2800 ;
  assign n17816 = ( n6845 & n8790 ) | ( n6845 & ~n11196 ) | ( n8790 & ~n11196 ) ;
  assign n17818 = n17817 ^ n17816 ^ n3440 ;
  assign n17819 = n14333 ^ n7953 ^ 1'b0 ;
  assign n17820 = n17819 ^ n3624 ^ 1'b0 ;
  assign n17822 = n3986 ^ n2320 ^ n1822 ;
  assign n17821 = n10016 | n15594 ;
  assign n17823 = n17822 ^ n17821 ^ n17645 ;
  assign n17824 = ( n5434 & ~n16756 ) | ( n5434 & n17823 ) | ( ~n16756 & n17823 ) ;
  assign n17825 = ( n1701 & n2015 ) | ( n1701 & n2467 ) | ( n2015 & n2467 ) ;
  assign n17826 = ( ~n1004 & n4601 ) | ( ~n1004 & n5246 ) | ( n4601 & n5246 ) ;
  assign n17827 = ( n5295 & n10929 ) | ( n5295 & ~n17826 ) | ( n10929 & ~n17826 ) ;
  assign n17828 = ( n1129 & n17825 ) | ( n1129 & ~n17827 ) | ( n17825 & ~n17827 ) ;
  assign n17829 = n17828 ^ n12074 ^ n8033 ;
  assign n17830 = ( n1907 & n2771 ) | ( n1907 & ~n4668 ) | ( n2771 & ~n4668 ) ;
  assign n17831 = n17830 ^ n3413 ^ 1'b0 ;
  assign n17832 = x45 & ~n17831 ;
  assign n17833 = ( n6580 & n13300 ) | ( n6580 & ~n13430 ) | ( n13300 & ~n13430 ) ;
  assign n17834 = ( n10513 & ~n10986 ) | ( n10513 & n16435 ) | ( ~n10986 & n16435 ) ;
  assign n17835 = ( n10665 & n15318 ) | ( n10665 & n17834 ) | ( n15318 & n17834 ) ;
  assign n17836 = ~n14260 & n17835 ;
  assign n17837 = n17009 & n17836 ;
  assign n17838 = n17837 ^ n9534 ^ n2005 ;
  assign n17839 = ~n10256 & n15258 ;
  assign n17840 = ~n14065 & n17839 ;
  assign n17841 = n16775 ^ n8036 ^ n4675 ;
  assign n17842 = ( ~n1353 & n11702 ) | ( ~n1353 & n17841 ) | ( n11702 & n17841 ) ;
  assign n17843 = n685 & n8967 ;
  assign n17844 = n17843 ^ n14192 ^ 1'b0 ;
  assign n17845 = n17842 & n17844 ;
  assign n17846 = ~n5073 & n17845 ;
  assign n17847 = n17846 ^ n1129 ^ 1'b0 ;
  assign n17848 = ( n2800 & ~n4343 ) | ( n2800 & n12266 ) | ( ~n4343 & n12266 ) ;
  assign n17849 = n17584 ^ n10646 ^ n6000 ;
  assign n17850 = ( n988 & ~n4859 ) | ( n988 & n10930 ) | ( ~n4859 & n10930 ) ;
  assign n17851 = n8343 ^ n1993 ^ n1166 ;
  assign n17852 = n9751 ^ n3261 ^ n1732 ;
  assign n17853 = ( n9904 & n17851 ) | ( n9904 & ~n17852 ) | ( n17851 & ~n17852 ) ;
  assign n17854 = ( ~n13227 & n17850 ) | ( ~n13227 & n17853 ) | ( n17850 & n17853 ) ;
  assign n17855 = n5669 & ~n14883 ;
  assign n17856 = n17855 ^ n3969 ^ 1'b0 ;
  assign n17857 = n7160 & n17856 ;
  assign n17858 = n17854 & n17857 ;
  assign n17859 = n523 & ~n14812 ;
  assign n17860 = n17859 ^ n5524 ^ n3300 ;
  assign n17861 = n17860 ^ n4641 ^ 1'b0 ;
  assign n17862 = n12831 | n17861 ;
  assign n17863 = n3167 ^ n2915 ^ 1'b0 ;
  assign n17867 = ( ~n2159 & n2181 ) | ( ~n2159 & n2353 ) | ( n2181 & n2353 ) ;
  assign n17864 = ( n170 & n3850 ) | ( n170 & n6308 ) | ( n3850 & n6308 ) ;
  assign n17865 = ~n8567 & n17864 ;
  assign n17866 = n17865 ^ n4980 ^ 1'b0 ;
  assign n17868 = n17867 ^ n17866 ^ n5447 ;
  assign n17869 = ( n2650 & n17863 ) | ( n2650 & ~n17868 ) | ( n17863 & ~n17868 ) ;
  assign n17873 = ~n1799 & n5469 ;
  assign n17874 = n5613 & n17873 ;
  assign n17875 = ~n3437 & n17874 ;
  assign n17870 = n11712 ^ n3379 ^ 1'b0 ;
  assign n17871 = n897 & ~n8240 ;
  assign n17872 = ( n3766 & n17870 ) | ( n3766 & ~n17871 ) | ( n17870 & ~n17871 ) ;
  assign n17876 = n17875 ^ n17872 ^ 1'b0 ;
  assign n17877 = n6114 ^ n2579 ^ 1'b0 ;
  assign n17878 = n17877 ^ n8631 ^ n7398 ;
  assign n17879 = n11363 ^ n306 ^ 1'b0 ;
  assign n17880 = n7704 & ~n17879 ;
  assign n17881 = ~n17540 & n17880 ;
  assign n17884 = ( n159 & ~n4035 ) | ( n159 & n16245 ) | ( ~n4035 & n16245 ) ;
  assign n17882 = ~n4081 & n4738 ;
  assign n17883 = n17882 ^ n9559 ^ n7368 ;
  assign n17885 = n17884 ^ n17883 ^ n14644 ;
  assign n17889 = ( ~x47 & n1568 ) | ( ~x47 & n8981 ) | ( n1568 & n8981 ) ;
  assign n17887 = n12654 ^ n11885 ^ x59 ;
  assign n17886 = ( n2234 & n10146 ) | ( n2234 & n15170 ) | ( n10146 & n15170 ) ;
  assign n17888 = n17887 ^ n17886 ^ n2270 ;
  assign n17890 = n17889 ^ n17888 ^ n16253 ;
  assign n17891 = n4213 | n4786 ;
  assign n17892 = n15823 ^ n12314 ^ n8944 ;
  assign n17893 = ( n15247 & n17886 ) | ( n15247 & ~n17892 ) | ( n17886 & ~n17892 ) ;
  assign n17894 = ( n15648 & ~n17891 ) | ( n15648 & n17893 ) | ( ~n17891 & n17893 ) ;
  assign n17895 = n13756 ^ n1984 ^ 1'b0 ;
  assign n17896 = n15786 | n17895 ;
  assign n17897 = n1347 ^ n415 ^ 1'b0 ;
  assign n17898 = n17897 ^ n6693 ^ n4943 ;
  assign n17899 = n17898 ^ n16408 ^ 1'b0 ;
  assign n17900 = n12429 ^ n2880 ^ n2319 ;
  assign n17901 = n9234 & ~n17900 ;
  assign n17902 = n6253 & n17901 ;
  assign n17903 = ( n3768 & n4034 ) | ( n3768 & ~n15441 ) | ( n4034 & ~n15441 ) ;
  assign n17904 = ~n6765 & n11920 ;
  assign n17905 = ~n4363 & n17904 ;
  assign n17906 = n8346 & n17905 ;
  assign n17907 = ( x81 & ~n3148 ) | ( x81 & n13124 ) | ( ~n3148 & n13124 ) ;
  assign n17908 = ( n1521 & n9314 ) | ( n1521 & ~n13515 ) | ( n9314 & ~n13515 ) ;
  assign n17909 = n12040 | n12672 ;
  assign n17910 = ~n833 & n9717 ;
  assign n17911 = n17910 ^ n15349 ^ 1'b0 ;
  assign n17912 = n4431 | n17911 ;
  assign n17913 = n17912 ^ n2826 ^ 1'b0 ;
  assign n17914 = ~n835 & n10437 ;
  assign n17915 = ~n5122 & n17914 ;
  assign n17916 = n1955 & n6646 ;
  assign n17917 = n3942 & n17916 ;
  assign n17918 = n17917 ^ n5523 ^ 1'b0 ;
  assign n17919 = n3874 & n17918 ;
  assign n17920 = ~n3259 & n17919 ;
  assign n17921 = n8797 | n17920 ;
  assign n17922 = ( n3208 & ~n4179 ) | ( n3208 & n11283 ) | ( ~n4179 & n11283 ) ;
  assign n17923 = n17922 ^ n11807 ^ n7318 ;
  assign n17924 = ( n17915 & ~n17921 ) | ( n17915 & n17923 ) | ( ~n17921 & n17923 ) ;
  assign n17926 = n2482 ^ n1461 ^ x62 ;
  assign n17925 = n6979 ^ n3843 ^ n564 ;
  assign n17927 = n17926 ^ n17925 ^ n15111 ;
  assign n17928 = ( ~n3508 & n9708 ) | ( ~n3508 & n17729 ) | ( n9708 & n17729 ) ;
  assign n17929 = n17928 ^ n2463 ^ 1'b0 ;
  assign n17930 = n17929 ^ n3499 ^ 1'b0 ;
  assign n17936 = ( n5930 & ~n5932 ) | ( n5930 & n7396 ) | ( ~n5932 & n7396 ) ;
  assign n17937 = n13956 | n17936 ;
  assign n17932 = n13027 ^ n11199 ^ 1'b0 ;
  assign n17933 = n17932 ^ n16924 ^ n12323 ;
  assign n17931 = n4132 & ~n17185 ;
  assign n17934 = n17933 ^ n17931 ^ 1'b0 ;
  assign n17935 = ~n1710 & n17934 ;
  assign n17938 = n17937 ^ n17935 ^ 1'b0 ;
  assign n17939 = n4667 & ~n8214 ;
  assign n17940 = n17939 ^ n2146 ^ 1'b0 ;
  assign n17941 = n14867 ^ n13264 ^ 1'b0 ;
  assign n17942 = n17941 ^ n7626 ^ n3155 ;
  assign n17943 = n7138 ^ n6953 ^ n950 ;
  assign n17944 = n17943 ^ n17166 ^ n7204 ;
  assign n17945 = n10508 ^ n10299 ^ n7905 ;
  assign n17946 = ( ~n2653 & n11545 ) | ( ~n2653 & n17945 ) | ( n11545 & n17945 ) ;
  assign n17947 = n1153 | n8469 ;
  assign n17948 = n9118 | n16531 ;
  assign n17949 = n17947 & ~n17948 ;
  assign n17950 = n13905 ^ n11620 ^ n2389 ;
  assign n17951 = ~n17949 & n17950 ;
  assign n17952 = n17951 ^ n5436 ^ 1'b0 ;
  assign n17953 = ( n754 & n7714 ) | ( n754 & n10760 ) | ( n7714 & n10760 ) ;
  assign n17954 = n10374 ^ n3168 ^ n1100 ;
  assign n17955 = n17954 ^ n6096 ^ 1'b0 ;
  assign n17956 = n17953 | n17955 ;
  assign n17957 = n12096 ^ n3405 ^ n3146 ;
  assign n17958 = n9574 & n17957 ;
  assign n17959 = ( n1345 & n5711 ) | ( n1345 & ~n17958 ) | ( n5711 & ~n17958 ) ;
  assign n17960 = n17959 ^ n11850 ^ 1'b0 ;
  assign n17963 = n12980 ^ n2778 ^ n794 ;
  assign n17961 = ( n642 & n2267 ) | ( n642 & n3915 ) | ( n2267 & n3915 ) ;
  assign n17962 = ~n4946 & n17961 ;
  assign n17964 = n17963 ^ n17962 ^ x70 ;
  assign n17965 = ( n1704 & n4947 ) | ( n1704 & n11041 ) | ( n4947 & n11041 ) ;
  assign n17966 = n17965 ^ n2130 ^ 1'b0 ;
  assign n17967 = ~n282 & n17966 ;
  assign n17968 = n17967 ^ n15937 ^ n14897 ;
  assign n17969 = n9223 | n9937 ;
  assign n17970 = ( n15435 & n15794 ) | ( n15435 & n17969 ) | ( n15794 & n17969 ) ;
  assign n17972 = n2008 | n17473 ;
  assign n17973 = n17972 ^ n8391 ^ 1'b0 ;
  assign n17971 = ~n6537 & n15650 ;
  assign n17974 = n17973 ^ n17971 ^ 1'b0 ;
  assign n17975 = n12816 | n14038 ;
  assign n17976 = n6442 & ~n17975 ;
  assign n17977 = ( ~n7785 & n10316 ) | ( ~n7785 & n10886 ) | ( n10316 & n10886 ) ;
  assign n17978 = ~n8890 & n12793 ;
  assign n17979 = n17978 ^ n13391 ^ 1'b0 ;
  assign n17980 = n17977 & n17979 ;
  assign n17981 = n17397 ^ n9374 ^ n2986 ;
  assign n17982 = n7319 ^ n2630 ^ 1'b0 ;
  assign n17983 = ( n15813 & n16803 ) | ( n15813 & n17982 ) | ( n16803 & n17982 ) ;
  assign n17985 = n5622 & n10037 ;
  assign n17986 = n17985 ^ n5889 ^ 1'b0 ;
  assign n17984 = n6335 ^ n3934 ^ n1668 ;
  assign n17987 = n17986 ^ n17984 ^ n11839 ;
  assign n17988 = n6935 ^ n715 ^ 1'b0 ;
  assign n17989 = n17988 ^ n12371 ^ n5060 ;
  assign n17990 = n14474 ^ n10702 ^ n6350 ;
  assign n17991 = ( n816 & ~n3534 ) | ( n816 & n4845 ) | ( ~n3534 & n4845 ) ;
  assign n17992 = n17991 ^ n487 ^ 1'b0 ;
  assign n17993 = n8145 ^ n3060 ^ 1'b0 ;
  assign n17994 = n17992 & ~n17993 ;
  assign n17995 = ( n3788 & n17990 ) | ( n3788 & ~n17994 ) | ( n17990 & ~n17994 ) ;
  assign n17996 = n7716 & n8249 ;
  assign n17997 = n17996 ^ n6740 ^ 1'b0 ;
  assign n17998 = n17997 ^ n9129 ^ n5900 ;
  assign n17999 = ( n2957 & n10702 ) | ( n2957 & ~n15391 ) | ( n10702 & ~n15391 ) ;
  assign n18000 = n7332 ^ n6967 ^ 1'b0 ;
  assign n18001 = n4191 & ~n5112 ;
  assign n18002 = n18001 ^ n7864 ^ 1'b0 ;
  assign n18003 = n18000 & n18002 ;
  assign n18004 = ( ~n4103 & n7949 ) | ( ~n4103 & n18003 ) | ( n7949 & n18003 ) ;
  assign n18005 = n13323 ^ n7292 ^ n337 ;
  assign n18006 = n12359 & ~n18005 ;
  assign n18007 = n18006 ^ n6927 ^ 1'b0 ;
  assign n18008 = n4076 ^ n986 ^ 1'b0 ;
  assign n18009 = n17953 | n18008 ;
  assign n18010 = n2885 ^ n2115 ^ 1'b0 ;
  assign n18011 = n18010 ^ n15816 ^ n14523 ;
  assign n18012 = n18011 ^ n5557 ^ n636 ;
  assign n18013 = n11062 ^ n6279 ^ n3691 ;
  assign n18014 = n18013 ^ n4346 ^ x20 ;
  assign n18015 = n8234 ^ n6886 ^ 1'b0 ;
  assign n18016 = ( n7905 & n15741 ) | ( n7905 & ~n18015 ) | ( n15741 & ~n18015 ) ;
  assign n18017 = n18016 ^ n16760 ^ n7567 ;
  assign n18018 = n4041 & ~n4250 ;
  assign n18019 = n18018 ^ n16636 ^ n1394 ;
  assign n18020 = ( n139 & n3872 ) | ( n139 & ~n8541 ) | ( n3872 & ~n8541 ) ;
  assign n18021 = n2957 | n18020 ;
  assign n18022 = n18019 | n18021 ;
  assign n18023 = n18022 ^ n7974 ^ n5050 ;
  assign n18024 = n9790 ^ n1874 ^ 1'b0 ;
  assign n18025 = ~n3506 & n18024 ;
  assign n18026 = n18025 ^ n16783 ^ n1887 ;
  assign n18027 = ( n3847 & n17041 ) | ( n3847 & n18026 ) | ( n17041 & n18026 ) ;
  assign n18028 = n13570 ^ n2835 ^ n637 ;
  assign n18029 = ( n7290 & ~n17319 ) | ( n7290 & n18028 ) | ( ~n17319 & n18028 ) ;
  assign n18030 = n846 | n18029 ;
  assign n18031 = n18030 ^ n8314 ^ 1'b0 ;
  assign n18032 = n878 & ~n8200 ;
  assign n18033 = ( n10706 & n11478 ) | ( n10706 & n18032 ) | ( n11478 & n18032 ) ;
  assign n18034 = ( n721 & n4150 ) | ( n721 & n8697 ) | ( n4150 & n8697 ) ;
  assign n18035 = ( n5206 & n10620 ) | ( n5206 & n18034 ) | ( n10620 & n18034 ) ;
  assign n18036 = ( n620 & ~n2736 ) | ( n620 & n3111 ) | ( ~n2736 & n3111 ) ;
  assign n18037 = n15776 ^ n4318 ^ 1'b0 ;
  assign n18038 = n1905 | n10945 ;
  assign n18039 = n18037 | n18038 ;
  assign n18040 = ~n3151 & n17967 ;
  assign n18041 = n9262 & n18040 ;
  assign n18042 = n10738 ^ n5671 ^ 1'b0 ;
  assign n18043 = n15525 ^ x21 ^ 1'b0 ;
  assign n18044 = n15345 ^ n10918 ^ n1983 ;
  assign n18045 = n6447 | n15786 ;
  assign n18046 = n12968 | n15344 ;
  assign n18047 = n3392 & ~n7994 ;
  assign n18048 = n11227 ^ n887 ^ 1'b0 ;
  assign n18049 = n3708 | n18048 ;
  assign n18050 = n18049 ^ n6954 ^ n2957 ;
  assign n18051 = n17329 ^ n8281 ^ 1'b0 ;
  assign n18052 = n5228 & ~n10871 ;
  assign n18053 = n18052 ^ n7779 ^ 1'b0 ;
  assign n18054 = ( n5000 & n11108 ) | ( n5000 & n15278 ) | ( n11108 & n15278 ) ;
  assign n18055 = n18054 ^ n17221 ^ n1057 ;
  assign n18056 = n17670 ^ n4049 ^ n1193 ;
  assign n18057 = ( n5973 & n10687 ) | ( n5973 & ~n17623 ) | ( n10687 & ~n17623 ) ;
  assign n18058 = n8221 ^ n8126 ^ n7582 ;
  assign n18059 = n11211 ^ n2265 ^ 1'b0 ;
  assign n18060 = n3814 | n18059 ;
  assign n18061 = ( ~n5874 & n10981 ) | ( ~n5874 & n18060 ) | ( n10981 & n18060 ) ;
  assign n18062 = n6653 ^ n3897 ^ 1'b0 ;
  assign n18063 = ( n9316 & n16531 ) | ( n9316 & ~n18062 ) | ( n16531 & ~n18062 ) ;
  assign n18064 = ( ~n3496 & n6298 ) | ( ~n3496 & n18063 ) | ( n6298 & n18063 ) ;
  assign n18065 = ( n5327 & n9328 ) | ( n5327 & ~n11146 ) | ( n9328 & ~n11146 ) ;
  assign n18066 = n18065 ^ n17986 ^ n11378 ;
  assign n18067 = n9624 & ~n15455 ;
  assign n18068 = n15473 ^ n8380 ^ n2792 ;
  assign n18069 = n2740 & n2931 ;
  assign n18070 = n18069 ^ n6899 ^ 1'b0 ;
  assign n18071 = n18070 ^ n4014 ^ 1'b0 ;
  assign n18072 = n18068 | n18071 ;
  assign n18073 = n18072 ^ n11567 ^ n2377 ;
  assign n18074 = ( n3480 & ~n5209 ) | ( n3480 & n18073 ) | ( ~n5209 & n18073 ) ;
  assign n18075 = ( ~n1186 & n5616 ) | ( ~n1186 & n13512 ) | ( n5616 & n13512 ) ;
  assign n18076 = ( n6066 & n7809 ) | ( n6066 & ~n18075 ) | ( n7809 & ~n18075 ) ;
  assign n18077 = n8053 ^ n2211 ^ 1'b0 ;
  assign n18078 = ( n9958 & n18076 ) | ( n9958 & n18077 ) | ( n18076 & n18077 ) ;
  assign n18079 = n14239 ^ n2713 ^ n183 ;
  assign n18083 = ~n1642 & n16148 ;
  assign n18084 = ~n16658 & n18083 ;
  assign n18080 = ( ~x95 & n2916 ) | ( ~x95 & n3576 ) | ( n2916 & n3576 ) ;
  assign n18081 = n18080 ^ n12101 ^ n7209 ;
  assign n18082 = n5883 & n18081 ;
  assign n18085 = n18084 ^ n18082 ^ 1'b0 ;
  assign n18086 = n18085 ^ n17581 ^ n16694 ;
  assign n18087 = ( n2357 & ~n4467 ) | ( n2357 & n11369 ) | ( ~n4467 & n11369 ) ;
  assign n18088 = ( ~n3298 & n5697 ) | ( ~n3298 & n7192 ) | ( n5697 & n7192 ) ;
  assign n18089 = n13147 ^ n1895 ^ n235 ;
  assign n18090 = n5150 ^ n755 ^ 1'b0 ;
  assign n18091 = n18089 & ~n18090 ;
  assign n18092 = n18091 ^ n7968 ^ 1'b0 ;
  assign n18093 = ( ~n9448 & n18088 ) | ( ~n9448 & n18092 ) | ( n18088 & n18092 ) ;
  assign n18094 = n18093 ^ n11844 ^ n8565 ;
  assign n18095 = ( ~n8372 & n12455 ) | ( ~n8372 & n17947 ) | ( n12455 & n17947 ) ;
  assign n18096 = ( ~n7894 & n10966 ) | ( ~n7894 & n11897 ) | ( n10966 & n11897 ) ;
  assign n18097 = n15186 ^ n2849 ^ n2440 ;
  assign n18098 = ( n18095 & n18096 ) | ( n18095 & ~n18097 ) | ( n18096 & ~n18097 ) ;
  assign n18099 = ( n9277 & ~n15191 ) | ( n9277 & n17439 ) | ( ~n15191 & n17439 ) ;
  assign n18100 = n5711 & ~n13549 ;
  assign n18101 = n12588 & n12599 ;
  assign n18102 = ~n1125 & n5380 ;
  assign n18103 = n1486 | n4221 ;
  assign n18104 = n917 | n4444 ;
  assign n18105 = ( n6364 & n11338 ) | ( n6364 & n18104 ) | ( n11338 & n18104 ) ;
  assign n18106 = n7146 ^ n528 ^ 1'b0 ;
  assign n18107 = n11679 & ~n18106 ;
  assign n18108 = n14271 ^ n7202 ^ x90 ;
  assign n18109 = ( n16155 & ~n18107 ) | ( n16155 & n18108 ) | ( ~n18107 & n18108 ) ;
  assign n18110 = n2708 & n17986 ;
  assign n18111 = n18110 ^ n16155 ^ 1'b0 ;
  assign n18112 = n1560 & ~n18111 ;
  assign n18113 = n12387 ^ n11134 ^ n4740 ;
  assign n18114 = ( ~n4886 & n11498 ) | ( ~n4886 & n18113 ) | ( n11498 & n18113 ) ;
  assign n18115 = n10016 ^ n8810 ^ n2078 ;
  assign n18116 = ( n7100 & n10715 ) | ( n7100 & ~n12102 ) | ( n10715 & ~n12102 ) ;
  assign n18117 = n6049 & n14425 ;
  assign n18118 = n12380 ^ n11682 ^ n5586 ;
  assign n18134 = ( ~n1400 & n9555 ) | ( ~n1400 & n10237 ) | ( n9555 & n10237 ) ;
  assign n18133 = n13944 ^ n2173 ^ n1675 ;
  assign n18119 = n4470 ^ n385 ^ 1'b0 ;
  assign n18120 = n18119 ^ n12586 ^ 1'b0 ;
  assign n18121 = ~n5908 & n18120 ;
  assign n18122 = n571 | n7198 ;
  assign n18123 = n18122 ^ n3811 ^ 1'b0 ;
  assign n18124 = ( n196 & n4971 ) | ( n196 & n10988 ) | ( n4971 & n10988 ) ;
  assign n18125 = n18124 ^ n6364 ^ n596 ;
  assign n18126 = n11276 ^ n10670 ^ 1'b0 ;
  assign n18127 = n1142 & ~n18126 ;
  assign n18128 = n16687 ^ n9788 ^ n3277 ;
  assign n18129 = n270 & ~n1877 ;
  assign n18130 = ~n18128 & n18129 ;
  assign n18131 = ( ~n18125 & n18127 ) | ( ~n18125 & n18130 ) | ( n18127 & n18130 ) ;
  assign n18132 = ( n18121 & ~n18123 ) | ( n18121 & n18131 ) | ( ~n18123 & n18131 ) ;
  assign n18135 = n18134 ^ n18133 ^ n18132 ;
  assign n18136 = n7377 ^ n5358 ^ n710 ;
  assign n18137 = n18136 ^ n12063 ^ 1'b0 ;
  assign n18138 = ~n16466 & n18137 ;
  assign n18139 = ( n6172 & n12678 ) | ( n6172 & n18138 ) | ( n12678 & n18138 ) ;
  assign n18140 = n4396 | n6503 ;
  assign n18141 = n18140 ^ n12228 ^ n6234 ;
  assign n18142 = n4884 & ~n9519 ;
  assign n18143 = n3281 | n15278 ;
  assign n18144 = n18142 & ~n18143 ;
  assign n18145 = ( n1606 & ~n1800 ) | ( n1606 & n18144 ) | ( ~n1800 & n18144 ) ;
  assign n18146 = n6987 ^ n4079 ^ 1'b0 ;
  assign n18147 = n10070 & n18146 ;
  assign n18148 = n2664 & n4416 ;
  assign n18149 = n18148 ^ n13264 ^ 1'b0 ;
  assign n18150 = ( n5969 & n13218 ) | ( n5969 & n18149 ) | ( n13218 & n18149 ) ;
  assign n18151 = ( n8459 & n10085 ) | ( n8459 & ~n11373 ) | ( n10085 & ~n11373 ) ;
  assign n18152 = n18151 ^ n4954 ^ 1'b0 ;
  assign n18153 = n16973 ^ n9534 ^ n1998 ;
  assign n18155 = n4647 ^ n1847 ^ 1'b0 ;
  assign n18154 = n4085 & ~n13451 ;
  assign n18156 = n18155 ^ n18154 ^ 1'b0 ;
  assign n18157 = ~n18153 & n18156 ;
  assign n18158 = ( n6377 & ~n8654 ) | ( n6377 & n18157 ) | ( ~n8654 & n18157 ) ;
  assign n18159 = ( n1798 & ~n11931 ) | ( n1798 & n18158 ) | ( ~n11931 & n18158 ) ;
  assign n18160 = n18159 ^ n17043 ^ n15562 ;
  assign n18161 = ( n1613 & n4559 ) | ( n1613 & ~n11544 ) | ( n4559 & ~n11544 ) ;
  assign n18162 = n18161 ^ n11513 ^ 1'b0 ;
  assign n18163 = n15789 | n18162 ;
  assign n18164 = n1120 & n4030 ;
  assign n18165 = n1573 & n18164 ;
  assign n18166 = n10374 & ~n18165 ;
  assign n18167 = n18166 ^ n3910 ^ 1'b0 ;
  assign n18169 = n2887 ^ n1858 ^ 1'b0 ;
  assign n18170 = n2236 & ~n18169 ;
  assign n18168 = n3052 & n6605 ;
  assign n18171 = n18170 ^ n18168 ^ 1'b0 ;
  assign n18172 = ( ~n6749 & n16760 ) | ( ~n6749 & n18171 ) | ( n16760 & n18171 ) ;
  assign n18173 = ( n2117 & n6957 ) | ( n2117 & ~n16219 ) | ( n6957 & ~n16219 ) ;
  assign n18174 = ( n4141 & n11093 ) | ( n4141 & n18173 ) | ( n11093 & n18173 ) ;
  assign n18175 = n18174 ^ n9103 ^ 1'b0 ;
  assign n18176 = n14668 & n18175 ;
  assign n18177 = ( n7631 & ~n9493 ) | ( n7631 & n18176 ) | ( ~n9493 & n18176 ) ;
  assign n18185 = n16572 ^ n15563 ^ n12979 ;
  assign n18184 = n12540 ^ n3573 ^ 1'b0 ;
  assign n18180 = n1880 & n9224 ;
  assign n18181 = ~n1148 & n18180 ;
  assign n18178 = ( ~n966 & n5214 ) | ( ~n966 & n6688 ) | ( n5214 & n6688 ) ;
  assign n18179 = n18178 ^ n14588 ^ n1874 ;
  assign n18182 = n18181 ^ n18179 ^ 1'b0 ;
  assign n18183 = ( ~n7988 & n17407 ) | ( ~n7988 & n18182 ) | ( n17407 & n18182 ) ;
  assign n18186 = n18185 ^ n18184 ^ n18183 ;
  assign n18187 = n4899 & ~n7192 ;
  assign n18188 = n18187 ^ n16115 ^ n11963 ;
  assign n18189 = n7631 ^ n5648 ^ n1588 ;
  assign n18190 = ~n2115 & n4828 ;
  assign n18191 = n7002 & ~n9649 ;
  assign n18192 = n18191 ^ n12762 ^ 1'b0 ;
  assign n18193 = n14135 ^ n5822 ^ 1'b0 ;
  assign n18194 = n2071 & n18193 ;
  assign n18195 = n18194 ^ n12679 ^ 1'b0 ;
  assign n18196 = ( n14847 & n18192 ) | ( n14847 & n18195 ) | ( n18192 & n18195 ) ;
  assign n18197 = n1809 | n12085 ;
  assign n18198 = n11627 ^ n2949 ^ n1671 ;
  assign n18199 = ( n7775 & ~n18197 ) | ( n7775 & n18198 ) | ( ~n18197 & n18198 ) ;
  assign n18204 = n16784 ^ n14955 ^ n473 ;
  assign n18200 = n8280 ^ n4878 ^ n3469 ;
  assign n18201 = n8139 ^ n242 ^ 1'b0 ;
  assign n18202 = n17450 & ~n18201 ;
  assign n18203 = ( ~n463 & n18200 ) | ( ~n463 & n18202 ) | ( n18200 & n18202 ) ;
  assign n18205 = n18204 ^ n18203 ^ x71 ;
  assign n18206 = n2638 & n4056 ;
  assign n18207 = n1822 & n18206 ;
  assign n18208 = n18207 ^ n12904 ^ n2231 ;
  assign n18209 = n18208 ^ n11148 ^ n5942 ;
  assign n18210 = n11988 ^ n4209 ^ n1242 ;
  assign n18211 = n18210 ^ n10398 ^ n3531 ;
  assign n18212 = n4876 | n11208 ;
  assign n18213 = n3272 ^ n2590 ^ n1949 ;
  assign n18214 = n18213 ^ n14500 ^ n8584 ;
  assign n18215 = n5981 ^ n2585 ^ 1'b0 ;
  assign n18216 = n6992 & n18215 ;
  assign n18217 = n18216 ^ n2005 ^ 1'b0 ;
  assign n18218 = n18214 & ~n18217 ;
  assign n18219 = n17663 | n18218 ;
  assign n18220 = ( n3279 & n3792 ) | ( n3279 & ~n4031 ) | ( n3792 & ~n4031 ) ;
  assign n18221 = ( n977 & n15805 ) | ( n977 & ~n18220 ) | ( n15805 & ~n18220 ) ;
  assign n18222 = n18221 ^ n14844 ^ n5169 ;
  assign n18223 = ( n2235 & ~n7343 ) | ( n2235 & n18222 ) | ( ~n7343 & n18222 ) ;
  assign n18224 = ( ~n8402 & n11079 ) | ( ~n8402 & n18223 ) | ( n11079 & n18223 ) ;
  assign n18225 = n5525 ^ n2888 ^ n2164 ;
  assign n18226 = n2283 & n4970 ;
  assign n18227 = n18225 & n18226 ;
  assign n18228 = n13732 ^ n3267 ^ 1'b0 ;
  assign n18229 = n10899 ^ n5235 ^ 1'b0 ;
  assign n18232 = n14464 ^ n8781 ^ n7340 ;
  assign n18230 = ( ~n3672 & n5604 ) | ( ~n3672 & n8691 ) | ( n5604 & n8691 ) ;
  assign n18231 = ( ~n627 & n4565 ) | ( ~n627 & n18230 ) | ( n4565 & n18230 ) ;
  assign n18233 = n18232 ^ n18231 ^ 1'b0 ;
  assign n18234 = n13078 ^ x13 ^ 1'b0 ;
  assign n18235 = ~n16309 & n18234 ;
  assign n18236 = ~n5618 & n7785 ;
  assign n18237 = n1579 & n18236 ;
  assign n18238 = n5372 & ~n5568 ;
  assign n18239 = n12743 & n18238 ;
  assign n18240 = ( n5118 & n7118 ) | ( n5118 & ~n18239 ) | ( n7118 & ~n18239 ) ;
  assign n18241 = n7556 & n18240 ;
  assign n18242 = n18241 ^ n5689 ^ 1'b0 ;
  assign n18243 = ( n3603 & ~n18237 ) | ( n3603 & n18242 ) | ( ~n18237 & n18242 ) ;
  assign n18244 = n9574 & n11998 ;
  assign n18245 = n8769 & n18244 ;
  assign n18246 = n18245 ^ n4265 ^ 1'b0 ;
  assign n18247 = n18243 & ~n18246 ;
  assign n18248 = ( ~n18233 & n18235 ) | ( ~n18233 & n18247 ) | ( n18235 & n18247 ) ;
  assign n18249 = ( n852 & ~n1437 ) | ( n852 & n16819 ) | ( ~n1437 & n16819 ) ;
  assign n18250 = n18203 ^ n902 ^ 1'b0 ;
  assign n18251 = n5331 & n17801 ;
  assign n18252 = n18250 | n18251 ;
  assign n18253 = n14521 ^ n5999 ^ n2680 ;
  assign n18254 = n2069 & ~n8433 ;
  assign n18255 = n18254 ^ n3900 ^ 1'b0 ;
  assign n18256 = n18255 ^ n13967 ^ n3795 ;
  assign n18257 = ( n5335 & n18197 ) | ( n5335 & n18256 ) | ( n18197 & n18256 ) ;
  assign n18258 = ( n4623 & ~n7744 ) | ( n4623 & n17079 ) | ( ~n7744 & n17079 ) ;
  assign n18259 = ( ~n5324 & n5376 ) | ( ~n5324 & n9671 ) | ( n5376 & n9671 ) ;
  assign n18260 = ~n1634 & n18259 ;
  assign n18261 = ~x117 & n18260 ;
  assign n18262 = n18261 ^ n3052 ^ 1'b0 ;
  assign n18263 = n13825 ^ n11949 ^ n10246 ;
  assign n18264 = n18263 ^ n7923 ^ 1'b0 ;
  assign n18265 = n2231 & n18264 ;
  assign n18266 = ( n2573 & n6537 ) | ( n2573 & ~n11284 ) | ( n6537 & ~n11284 ) ;
  assign n18267 = ~n6310 & n18266 ;
  assign n18268 = n15274 & n18267 ;
  assign n18269 = n18268 ^ n17469 ^ n6479 ;
  assign n18270 = n12910 | n17327 ;
  assign n18271 = n3908 & ~n18270 ;
  assign n18272 = n18271 ^ n7463 ^ 1'b0 ;
  assign n18273 = n14553 ^ n9285 ^ n5361 ;
  assign n18274 = ~n1433 & n7533 ;
  assign n18275 = n18274 ^ n746 ^ 1'b0 ;
  assign n18276 = ( n13881 & ~n18273 ) | ( n13881 & n18275 ) | ( ~n18273 & n18275 ) ;
  assign n18277 = ( ~n576 & n2665 ) | ( ~n576 & n13276 ) | ( n2665 & n13276 ) ;
  assign n18278 = ( n3156 & n3698 ) | ( n3156 & n5242 ) | ( n3698 & n5242 ) ;
  assign n18279 = n18278 ^ n16190 ^ n10713 ;
  assign n18280 = ( n4176 & ~n4242 ) | ( n4176 & n8259 ) | ( ~n4242 & n8259 ) ;
  assign n18281 = ( n5214 & ~n7175 ) | ( n5214 & n18280 ) | ( ~n7175 & n18280 ) ;
  assign n18292 = n5692 ^ n2664 ^ n1703 ;
  assign n18282 = n16426 ^ n2032 ^ 1'b0 ;
  assign n18283 = ~n4341 & n18282 ;
  assign n18284 = n703 & ~n1359 ;
  assign n18285 = n2612 & n18284 ;
  assign n18286 = n18283 & ~n18285 ;
  assign n18287 = n18286 ^ n2322 ^ 1'b0 ;
  assign n18288 = n273 & n13839 ;
  assign n18289 = n18288 ^ n6444 ^ 1'b0 ;
  assign n18290 = n18289 ^ n6729 ^ 1'b0 ;
  assign n18291 = n18287 & ~n18290 ;
  assign n18293 = n18292 ^ n18291 ^ n6631 ;
  assign n18294 = n16263 ^ n3531 ^ 1'b0 ;
  assign n18295 = n4147 & n18294 ;
  assign n18296 = n2498 ^ n2368 ^ 1'b0 ;
  assign n18297 = ( n9524 & ~n16548 ) | ( n9524 & n18296 ) | ( ~n16548 & n18296 ) ;
  assign n18298 = n18297 ^ n11205 ^ n6444 ;
  assign n18299 = ( n4567 & n6063 ) | ( n4567 & ~n18298 ) | ( n6063 & ~n18298 ) ;
  assign n18300 = n4097 ^ n2998 ^ n2943 ;
  assign n18301 = n5172 ^ n3357 ^ n2805 ;
  assign n18302 = n5443 ^ n645 ^ 1'b0 ;
  assign n18303 = ~n1334 & n18302 ;
  assign n18304 = n18303 ^ n11948 ^ n8166 ;
  assign n18306 = n13609 ^ n823 ^ 1'b0 ;
  assign n18307 = ( n139 & ~n2149 ) | ( n139 & n18306 ) | ( ~n2149 & n18306 ) ;
  assign n18305 = n6900 & ~n10257 ;
  assign n18308 = n18307 ^ n18305 ^ n2054 ;
  assign n18309 = n4796 & n5843 ;
  assign n18310 = ~n4567 & n18309 ;
  assign n18311 = n18310 ^ n13952 ^ n13303 ;
  assign n18312 = ( n4576 & ~n11763 ) | ( n4576 & n13445 ) | ( ~n11763 & n13445 ) ;
  assign n18313 = n18312 ^ n10299 ^ 1'b0 ;
  assign n18314 = n18313 ^ n12852 ^ 1'b0 ;
  assign n18315 = n18314 ^ n8968 ^ 1'b0 ;
  assign n18316 = ~n6145 & n18315 ;
  assign n18317 = n11767 ^ n7556 ^ n1318 ;
  assign n18318 = n10752 ^ n5648 ^ n336 ;
  assign n18319 = n18318 ^ n17992 ^ n564 ;
  assign n18320 = ~n8319 & n18319 ;
  assign n18321 = n18317 & n18320 ;
  assign n18322 = n6203 ^ n2724 ^ 1'b0 ;
  assign n18323 = ~n11540 & n18322 ;
  assign n18324 = ( n7674 & n9682 ) | ( n7674 & ~n11577 ) | ( n9682 & ~n11577 ) ;
  assign n18325 = n3753 & n18324 ;
  assign n18326 = x49 & ~n18325 ;
  assign n18327 = n9553 & n18326 ;
  assign n18329 = n8849 ^ n8576 ^ n542 ;
  assign n18330 = n18329 ^ x111 ^ 1'b0 ;
  assign n18331 = ( ~n1771 & n9643 ) | ( ~n1771 & n18330 ) | ( n9643 & n18330 ) ;
  assign n18328 = n5005 & ~n12366 ;
  assign n18332 = n18331 ^ n18328 ^ n9811 ;
  assign n18333 = n9685 | n17370 ;
  assign n18334 = n18333 ^ n6850 ^ 1'b0 ;
  assign n18335 = ( n8045 & n12392 ) | ( n8045 & ~n18334 ) | ( n12392 & ~n18334 ) ;
  assign n18336 = n14224 ^ n10732 ^ n5421 ;
  assign n18337 = n3714 ^ n1627 ^ n440 ;
  assign n18338 = ( n9430 & ~n18336 ) | ( n9430 & n18337 ) | ( ~n18336 & n18337 ) ;
  assign n18339 = ~n3506 & n13999 ;
  assign n18340 = n18338 & n18339 ;
  assign n18341 = n5866 ^ n359 ^ 1'b0 ;
  assign n18342 = n13518 & n18341 ;
  assign n18343 = ~n600 & n18342 ;
  assign n18344 = ~n17728 & n18343 ;
  assign n18345 = n18344 ^ n14459 ^ 1'b0 ;
  assign n18346 = n18345 ^ n7358 ^ 1'b0 ;
  assign n18347 = ( n4197 & ~n4486 ) | ( n4197 & n4528 ) | ( ~n4486 & n4528 ) ;
  assign n18348 = ( x62 & n6314 ) | ( x62 & ~n18347 ) | ( n6314 & ~n18347 ) ;
  assign n18349 = ( ~n4310 & n4495 ) | ( ~n4310 & n18303 ) | ( n4495 & n18303 ) ;
  assign n18350 = n7081 & n18349 ;
  assign n18351 = n18350 ^ n4579 ^ 1'b0 ;
  assign n18352 = n6105 ^ n5324 ^ n725 ;
  assign n18353 = n4989 & n18352 ;
  assign n18354 = n18353 ^ n3599 ^ 1'b0 ;
  assign n18355 = n5307 ^ n2631 ^ x69 ;
  assign n18356 = n18355 ^ n13531 ^ n2610 ;
  assign n18357 = n4539 & n9865 ;
  assign n18358 = n1433 & n18357 ;
  assign n18359 = n1098 & ~n3388 ;
  assign n18360 = n18359 ^ n1559 ^ 1'b0 ;
  assign n18361 = n18360 ^ n1107 ^ 1'b0 ;
  assign n18362 = n5664 & n18361 ;
  assign n18363 = n18358 | n18362 ;
  assign n18364 = n2437 & n6758 ;
  assign n18365 = n18363 & n18364 ;
  assign n18368 = ( n3094 & n3373 ) | ( n3094 & ~n4490 ) | ( n3373 & ~n4490 ) ;
  assign n18366 = n4589 ^ n1871 ^ x46 ;
  assign n18367 = ~n1287 & n18366 ;
  assign n18369 = n18368 ^ n18367 ^ 1'b0 ;
  assign n18370 = n10458 ^ n9776 ^ 1'b0 ;
  assign n18371 = n12824 | n18370 ;
  assign n18372 = n10503 & n17771 ;
  assign n18373 = n18372 ^ n13942 ^ n4292 ;
  assign n18374 = ~n3413 & n6462 ;
  assign n18375 = n18374 ^ n9434 ^ 1'b0 ;
  assign n18376 = n18375 ^ n8519 ^ n5969 ;
  assign n18377 = n15701 ^ n11344 ^ 1'b0 ;
  assign n18378 = ( n1377 & n2580 ) | ( n1377 & ~n4624 ) | ( n2580 & ~n4624 ) ;
  assign n18379 = n18378 ^ n6766 ^ n1901 ;
  assign n18380 = n18091 ^ n4418 ^ 1'b0 ;
  assign n18381 = n10561 ^ n4453 ^ 1'b0 ;
  assign n18382 = n16652 & n18381 ;
  assign n18387 = n14750 ^ n12227 ^ n4353 ;
  assign n18383 = n708 | n7481 ;
  assign n18384 = n1484 & ~n18383 ;
  assign n18385 = n340 | n4792 ;
  assign n18386 = n18384 & ~n18385 ;
  assign n18388 = n18387 ^ n18386 ^ n4069 ;
  assign n18389 = n18382 & n18388 ;
  assign n18393 = n8848 ^ n8055 ^ n867 ;
  assign n18394 = n18393 ^ n9532 ^ n385 ;
  assign n18391 = n13967 ^ n5214 ^ x5 ;
  assign n18390 = n7837 | n10436 ;
  assign n18392 = n18391 ^ n18390 ^ n3642 ;
  assign n18395 = n18394 ^ n18392 ^ 1'b0 ;
  assign n18396 = n843 & ~n18395 ;
  assign n18397 = ~n3309 & n4170 ;
  assign n18398 = n16527 & n18397 ;
  assign n18399 = ( n407 & n5318 ) | ( n407 & ~n18398 ) | ( n5318 & ~n18398 ) ;
  assign n18400 = n10767 ^ n3998 ^ 1'b0 ;
  assign n18402 = n4796 & ~n6071 ;
  assign n18403 = ~n7806 & n18402 ;
  assign n18401 = ( ~n3600 & n4053 ) | ( ~n3600 & n8257 ) | ( n4053 & n8257 ) ;
  assign n18404 = n18403 ^ n18401 ^ n15300 ;
  assign n18405 = n18400 | n18404 ;
  assign n18409 = ( n3888 & n4984 ) | ( n3888 & n8854 ) | ( n4984 & n8854 ) ;
  assign n18408 = n11210 ^ n9788 ^ n6700 ;
  assign n18410 = n18409 ^ n18408 ^ n12478 ;
  assign n18407 = ( ~n1426 & n2749 ) | ( ~n1426 & n17376 ) | ( n2749 & n17376 ) ;
  assign n18406 = ~n8810 & n13920 ;
  assign n18411 = n18410 ^ n18407 ^ n18406 ;
  assign n18412 = n2115 | n6557 ;
  assign n18413 = ~n505 & n5349 ;
  assign n18414 = n394 & n18413 ;
  assign n18415 = ( n2193 & ~n6044 ) | ( n2193 & n14101 ) | ( ~n6044 & n14101 ) ;
  assign n18416 = ( n10242 & n18414 ) | ( n10242 & ~n18415 ) | ( n18414 & ~n18415 ) ;
  assign n18417 = ( n3640 & n18412 ) | ( n3640 & n18416 ) | ( n18412 & n18416 ) ;
  assign n18418 = ( n6261 & ~n7934 ) | ( n6261 & n18307 ) | ( ~n7934 & n18307 ) ;
  assign n18419 = ~n10555 & n18418 ;
  assign n18420 = n14238 & n14533 ;
  assign n18421 = n5942 & n18420 ;
  assign n18423 = ( n5719 & ~n8028 ) | ( n5719 & n14484 ) | ( ~n8028 & n14484 ) ;
  assign n18424 = n14359 ^ n9644 ^ 1'b0 ;
  assign n18425 = n18423 & ~n18424 ;
  assign n18422 = ~n3917 & n6273 ;
  assign n18426 = n18425 ^ n18422 ^ 1'b0 ;
  assign n18427 = n1212 & ~n6549 ;
  assign n18428 = n17509 ^ n15537 ^ 1'b0 ;
  assign n18429 = n18427 & n18428 ;
  assign n18430 = n11568 & ~n18429 ;
  assign n18434 = n1215 & ~n13646 ;
  assign n18431 = n8895 ^ n2689 ^ 1'b0 ;
  assign n18432 = n15486 ^ n3310 ^ 1'b0 ;
  assign n18433 = ( n12425 & n18431 ) | ( n12425 & ~n18432 ) | ( n18431 & ~n18432 ) ;
  assign n18435 = n18434 ^ n18433 ^ n16573 ;
  assign n18436 = n4871 ^ n1159 ^ 1'b0 ;
  assign n18437 = n3192 | n18436 ;
  assign n18438 = n4230 & n18437 ;
  assign n18439 = ~n9917 & n12366 ;
  assign n18440 = ( n1754 & n5381 ) | ( n1754 & ~n6724 ) | ( n5381 & ~n6724 ) ;
  assign n18441 = n18440 ^ n12208 ^ 1'b0 ;
  assign n18442 = n5409 & n18441 ;
  assign n18443 = n1487 | n3716 ;
  assign n18444 = n1519 & n18443 ;
  assign n18445 = ~n12855 & n18444 ;
  assign n18446 = ( ~n131 & n18442 ) | ( ~n131 & n18445 ) | ( n18442 & n18445 ) ;
  assign n18447 = n10730 & n10847 ;
  assign n18448 = n13089 & n18447 ;
  assign n18449 = n7546 ^ n5800 ^ 1'b0 ;
  assign n18450 = n11419 & ~n18449 ;
  assign n18452 = n11160 ^ n4991 ^ n3095 ;
  assign n18453 = n18452 ^ n16555 ^ n5070 ;
  assign n18454 = n18453 ^ n7306 ^ 1'b0 ;
  assign n18455 = n8888 & n18454 ;
  assign n18451 = n14264 ^ n2912 ^ n282 ;
  assign n18456 = n18455 ^ n18451 ^ 1'b0 ;
  assign n18457 = n18456 ^ n643 ^ x103 ;
  assign n18458 = n1384 | n9787 ;
  assign n18459 = n2176 & ~n18458 ;
  assign n18460 = n18459 ^ n12465 ^ n3021 ;
  assign n18461 = n17000 ^ n16358 ^ n3540 ;
  assign n18462 = ( n4000 & n11862 ) | ( n4000 & n18461 ) | ( n11862 & n18461 ) ;
  assign n18463 = n571 | n6808 ;
  assign n18464 = ( n6099 & ~n12913 ) | ( n6099 & n14464 ) | ( ~n12913 & n14464 ) ;
  assign n18465 = n10796 ^ n7373 ^ n2159 ;
  assign n18466 = ( n153 & n5302 ) | ( n153 & n5407 ) | ( n5302 & n5407 ) ;
  assign n18467 = ~n12910 & n18466 ;
  assign n18468 = ( n10926 & n17544 ) | ( n10926 & ~n18467 ) | ( n17544 & ~n18467 ) ;
  assign n18469 = n6419 ^ n3885 ^ 1'b0 ;
  assign n18470 = ( ~n10959 & n11779 ) | ( ~n10959 & n18469 ) | ( n11779 & n18469 ) ;
  assign n18471 = n16783 ^ n2073 ^ 1'b0 ;
  assign n18472 = ~n6348 & n18471 ;
  assign n18473 = ( n7435 & n15087 ) | ( n7435 & n18472 ) | ( n15087 & n18472 ) ;
  assign n18475 = n2654 ^ n1809 ^ n144 ;
  assign n18474 = n14051 ^ n5725 ^ n4480 ;
  assign n18476 = n18475 ^ n18474 ^ n10701 ;
  assign n18478 = ~n9796 & n14405 ;
  assign n18479 = n18478 ^ n14181 ^ 1'b0 ;
  assign n18477 = ~n1775 & n12261 ;
  assign n18480 = n18479 ^ n18477 ^ 1'b0 ;
  assign n18481 = ( x104 & n11453 ) | ( x104 & n14115 ) | ( n11453 & n14115 ) ;
  assign n18482 = ( n4652 & ~n8291 ) | ( n4652 & n15770 ) | ( ~n8291 & n15770 ) ;
  assign n18483 = n9652 ^ n8295 ^ 1'b0 ;
  assign n18484 = ~n6033 & n18483 ;
  assign n18485 = n11861 ^ n6443 ^ n1867 ;
  assign n18486 = ( ~n6547 & n11530 ) | ( ~n6547 & n18485 ) | ( n11530 & n18485 ) ;
  assign n18487 = ( ~n9649 & n18484 ) | ( ~n9649 & n18486 ) | ( n18484 & n18486 ) ;
  assign n18488 = ( n11508 & ~n11719 ) | ( n11508 & n12896 ) | ( ~n11719 & n12896 ) ;
  assign n18492 = n9780 ^ n4634 ^ n3239 ;
  assign n18493 = n18492 ^ n10651 ^ n4997 ;
  assign n18494 = n18493 ^ n2103 ^ n451 ;
  assign n18489 = ( n1480 & n2389 ) | ( n1480 & ~n2637 ) | ( n2389 & ~n2637 ) ;
  assign n18490 = n18489 ^ n3934 ^ 1'b0 ;
  assign n18491 = n2464 | n18490 ;
  assign n18495 = n18494 ^ n18491 ^ n17796 ;
  assign n18496 = n18495 ^ n10421 ^ n773 ;
  assign n18497 = ( n3891 & n15341 ) | ( n3891 & ~n16934 ) | ( n15341 & ~n16934 ) ;
  assign n18498 = ( n851 & n1688 ) | ( n851 & n4265 ) | ( n1688 & n4265 ) ;
  assign n18499 = n18498 ^ n17333 ^ 1'b0 ;
  assign n18501 = ~n7375 & n13989 ;
  assign n18502 = n18501 ^ n8921 ^ 1'b0 ;
  assign n18503 = ( n12396 & n17680 ) | ( n12396 & ~n18502 ) | ( n17680 & ~n18502 ) ;
  assign n18500 = ( n10718 & n14053 ) | ( n10718 & ~n14351 ) | ( n14053 & ~n14351 ) ;
  assign n18504 = n18503 ^ n18500 ^ n3049 ;
  assign n18505 = n7625 & ~n10533 ;
  assign n18506 = n11080 ^ n10152 ^ 1'b0 ;
  assign n18507 = ( n8211 & ~n16874 ) | ( n8211 & n18506 ) | ( ~n16874 & n18506 ) ;
  assign n18508 = ( ~n13215 & n18505 ) | ( ~n13215 & n18507 ) | ( n18505 & n18507 ) ;
  assign n18509 = x36 & ~n5070 ;
  assign n18510 = ~n5797 & n18509 ;
  assign n18511 = n12332 | n18510 ;
  assign n18512 = ( ~n2820 & n17822 ) | ( ~n2820 & n18511 ) | ( n17822 & n18511 ) ;
  assign n18513 = n16709 ^ n10290 ^ n3854 ;
  assign n18514 = n154 & n2446 ;
  assign n18515 = n2943 & ~n18514 ;
  assign n18516 = n12674 & n18515 ;
  assign n18517 = n15140 & ~n18516 ;
  assign n18518 = ~n2988 & n18517 ;
  assign n18522 = ( n4008 & n11487 ) | ( n4008 & ~n17063 ) | ( n11487 & ~n17063 ) ;
  assign n18523 = n18522 ^ n16747 ^ 1'b0 ;
  assign n18519 = n7657 | n10948 ;
  assign n18520 = n7849 | n18519 ;
  assign n18521 = n18520 ^ n17509 ^ n11687 ;
  assign n18524 = n18523 ^ n18521 ^ n2246 ;
  assign n18525 = ( n914 & n6018 ) | ( n914 & n18242 ) | ( n6018 & n18242 ) ;
  assign n18526 = n4250 & ~n7448 ;
  assign n18527 = n18526 ^ n12284 ^ n1242 ;
  assign n18528 = n17394 ^ n10448 ^ 1'b0 ;
  assign n18529 = n4342 | n18528 ;
  assign n18530 = ( ~n2296 & n10623 ) | ( ~n2296 & n18529 ) | ( n10623 & n18529 ) ;
  assign n18531 = n10048 & ~n18530 ;
  assign n18532 = n3482 | n18531 ;
  assign n18533 = n9581 | n10162 ;
  assign n18534 = n11041 ^ n10938 ^ n2759 ;
  assign n18535 = n18534 ^ n13455 ^ n6489 ;
  assign n18536 = n3380 & ~n18535 ;
  assign n18537 = n18536 ^ n6464 ^ n847 ;
  assign n18538 = n11747 ^ n6719 ^ n2128 ;
  assign n18542 = ( ~n5435 & n5956 ) | ( ~n5435 & n8704 ) | ( n5956 & n8704 ) ;
  assign n18543 = ( ~n3318 & n12990 ) | ( ~n3318 & n18542 ) | ( n12990 & n18542 ) ;
  assign n18539 = n933 | n7321 ;
  assign n18540 = n11855 | n18539 ;
  assign n18541 = n7669 & n18540 ;
  assign n18544 = n18543 ^ n18541 ^ 1'b0 ;
  assign n18545 = ~n18538 & n18544 ;
  assign n18546 = n18255 ^ n17227 ^ n15963 ;
  assign n18547 = n10234 ^ n4306 ^ 1'b0 ;
  assign n18548 = ~n18546 & n18547 ;
  assign n18549 = n13174 ^ n1518 ^ 1'b0 ;
  assign n18550 = ( ~n9123 & n11620 ) | ( ~n9123 & n18549 ) | ( n11620 & n18549 ) ;
  assign n18551 = n8614 & ~n10528 ;
  assign n18552 = n8029 ^ n7777 ^ 1'b0 ;
  assign n18553 = n5234 & ~n18552 ;
  assign n18554 = n13502 & n18553 ;
  assign n18555 = ( n3861 & ~n12807 ) | ( n3861 & n16599 ) | ( ~n12807 & n16599 ) ;
  assign n18556 = n8186 ^ n3375 ^ 1'b0 ;
  assign n18557 = n3857 | n18556 ;
  assign n18558 = n18557 ^ n2036 ^ 1'b0 ;
  assign n18559 = n14039 ^ n11326 ^ n6721 ;
  assign n18560 = ( n1428 & n1971 ) | ( n1428 & ~n8159 ) | ( n1971 & ~n8159 ) ;
  assign n18561 = n12456 ^ n3087 ^ 1'b0 ;
  assign n18562 = ( n1107 & n4894 ) | ( n1107 & n7533 ) | ( n4894 & n7533 ) ;
  assign n18563 = n3316 & n18562 ;
  assign n18564 = ~n18561 & n18563 ;
  assign n18565 = n5014 ^ n4168 ^ 1'b0 ;
  assign n18566 = n17079 ^ n2785 ^ 1'b0 ;
  assign n18567 = n18565 & ~n18566 ;
  assign n18568 = n18567 ^ n7890 ^ 1'b0 ;
  assign n18569 = n18568 ^ n544 ^ 1'b0 ;
  assign n18570 = n18569 ^ n9880 ^ n1099 ;
  assign n18571 = ( n5129 & n5774 ) | ( n5129 & n7091 ) | ( n5774 & n7091 ) ;
  assign n18572 = n1483 & n2410 ;
  assign n18573 = ( ~n11695 & n18571 ) | ( ~n11695 & n18572 ) | ( n18571 & n18572 ) ;
  assign n18574 = n5155 | n5763 ;
  assign n18575 = n13076 | n18574 ;
  assign n18576 = n15423 ^ n15159 ^ 1'b0 ;
  assign n18577 = n10465 & n18576 ;
  assign n18578 = n2192 ^ n1542 ^ 1'b0 ;
  assign n18579 = n11871 & n18578 ;
  assign n18580 = n1546 & ~n15901 ;
  assign n18581 = n18580 ^ n3083 ^ 1'b0 ;
  assign n18582 = n18251 & n18581 ;
  assign n18583 = n3681 | n7814 ;
  assign n18584 = ( ~n488 & n14634 ) | ( ~n488 & n18583 ) | ( n14634 & n18583 ) ;
  assign n18585 = ( ~n4305 & n5875 ) | ( ~n4305 & n6416 ) | ( n5875 & n6416 ) ;
  assign n18586 = n5434 ^ n3133 ^ n901 ;
  assign n18587 = n9341 ^ n8403 ^ 1'b0 ;
  assign n18588 = ~n9149 & n18587 ;
  assign n18589 = ( ~n13905 & n18586 ) | ( ~n13905 & n18588 ) | ( n18586 & n18588 ) ;
  assign n18590 = ( n5601 & ~n18585 ) | ( n5601 & n18589 ) | ( ~n18585 & n18589 ) ;
  assign n18591 = n12174 ^ n1645 ^ n709 ;
  assign n18592 = ( n1834 & n8704 ) | ( n1834 & n17340 ) | ( n8704 & n17340 ) ;
  assign n18593 = ( n7229 & ~n18591 ) | ( n7229 & n18592 ) | ( ~n18591 & n18592 ) ;
  assign n18594 = ( n6838 & ~n10562 ) | ( n6838 & n18200 ) | ( ~n10562 & n18200 ) ;
  assign n18595 = n18594 ^ n9119 ^ 1'b0 ;
  assign n18596 = ( n14418 & ~n15947 ) | ( n14418 & n18595 ) | ( ~n15947 & n18595 ) ;
  assign n18597 = n1557 | n10974 ;
  assign n18598 = ~n10665 & n18597 ;
  assign n18599 = n18598 ^ n2734 ^ 1'b0 ;
  assign n18600 = n230 | n7059 ;
  assign n18601 = n18599 | n18600 ;
  assign n18602 = n3353 ^ n487 ^ 1'b0 ;
  assign n18603 = n18602 ^ n9217 ^ n8826 ;
  assign n18604 = n18603 ^ n17036 ^ n4074 ;
  assign n18605 = ~n18601 & n18604 ;
  assign n18606 = n17745 ^ n9413 ^ n8585 ;
  assign n18607 = ( n6125 & n8775 ) | ( n6125 & n13190 ) | ( n8775 & n13190 ) ;
  assign n18608 = n14411 ^ n2423 ^ 1'b0 ;
  assign n18609 = n16686 & n18608 ;
  assign n18610 = ( n1690 & n2931 ) | ( n1690 & n14556 ) | ( n2931 & n14556 ) ;
  assign n18611 = n348 & n5754 ;
  assign n18612 = ( n14063 & n16687 ) | ( n14063 & n18611 ) | ( n16687 & n18611 ) ;
  assign n18613 = n794 & n9821 ;
  assign n18614 = n18613 ^ n4340 ^ 1'b0 ;
  assign n18615 = n10391 & ~n18614 ;
  assign n18616 = ( n16865 & ~n18612 ) | ( n16865 & n18615 ) | ( ~n18612 & n18615 ) ;
  assign n18617 = n9929 ^ n2923 ^ n1088 ;
  assign n18618 = n13929 ^ n13824 ^ n2775 ;
  assign n18619 = n18618 ^ n4996 ^ n3613 ;
  assign n18620 = n11679 ^ n8589 ^ 1'b0 ;
  assign n18621 = n17636 ^ n16438 ^ n1143 ;
  assign n18622 = n3661 & n7584 ;
  assign n18623 = ~n14867 & n18622 ;
  assign n18624 = n15539 & ~n18623 ;
  assign n18625 = ( ~n1525 & n7726 ) | ( ~n1525 & n11833 ) | ( n7726 & n11833 ) ;
  assign n18626 = n4980 | n18625 ;
  assign n18627 = ( n3666 & n13093 ) | ( n3666 & n16063 ) | ( n13093 & n16063 ) ;
  assign n18628 = n5635 & ~n11131 ;
  assign n18629 = n18628 ^ n18322 ^ 1'b0 ;
  assign n18630 = n2896 & ~n2917 ;
  assign n18631 = ~n18629 & n18630 ;
  assign n18632 = n12944 ^ n4953 ^ 1'b0 ;
  assign n18633 = ( n7100 & ~n14663 ) | ( n7100 & n18632 ) | ( ~n14663 & n18632 ) ;
  assign n18634 = n17929 ^ n4142 ^ n1100 ;
  assign n18635 = n10029 ^ n7399 ^ 1'b0 ;
  assign n18636 = n18635 ^ n12004 ^ n202 ;
  assign n18637 = n8498 ^ n7752 ^ 1'b0 ;
  assign n18638 = ( ~n1309 & n6382 ) | ( ~n1309 & n17178 ) | ( n6382 & n17178 ) ;
  assign n18639 = n5508 | n18638 ;
  assign n18640 = n7085 | n18639 ;
  assign n18641 = n18640 ^ n12598 ^ n3433 ;
  assign n18642 = ( n17137 & n18637 ) | ( n17137 & ~n18641 ) | ( n18637 & ~n18641 ) ;
  assign n18643 = ( n2469 & ~n4020 ) | ( n2469 & n18642 ) | ( ~n4020 & n18642 ) ;
  assign n18644 = ( ~n3053 & n12729 ) | ( ~n3053 & n13744 ) | ( n12729 & n13744 ) ;
  assign n18646 = n17825 ^ n6565 ^ 1'b0 ;
  assign n18645 = n8691 ^ n4708 ^ 1'b0 ;
  assign n18647 = n18646 ^ n18645 ^ n11736 ;
  assign n18648 = ( n5277 & n6034 ) | ( n5277 & ~n15665 ) | ( n6034 & ~n15665 ) ;
  assign n18649 = n18648 ^ n1609 ^ n837 ;
  assign n18650 = n8527 & n17503 ;
  assign n18651 = n18650 ^ n2389 ^ 1'b0 ;
  assign n18652 = n966 | n13662 ;
  assign n18653 = ~n14100 & n18652 ;
  assign n18654 = n18653 ^ n11587 ^ 1'b0 ;
  assign n18655 = n10618 & ~n11623 ;
  assign n18656 = ~n15907 & n18655 ;
  assign n18657 = n1822 | n2185 ;
  assign n18658 = n18657 ^ n14230 ^ 1'b0 ;
  assign n18659 = x88 & n1230 ;
  assign n18660 = n9128 & n18659 ;
  assign n18661 = n18660 ^ n4339 ^ 1'b0 ;
  assign n18662 = ( ~n1029 & n2640 ) | ( ~n1029 & n7852 ) | ( n2640 & n7852 ) ;
  assign n18663 = n18662 ^ n15895 ^ 1'b0 ;
  assign n18664 = ( ~n4868 & n8482 ) | ( ~n4868 & n9386 ) | ( n8482 & n9386 ) ;
  assign n18665 = n2988 | n18664 ;
  assign n18666 = n17325 ^ n10876 ^ n6529 ;
  assign n18667 = n7806 & n18666 ;
  assign n18668 = n18667 ^ n4681 ^ 1'b0 ;
  assign n18669 = n15135 ^ n13507 ^ n5967 ;
  assign n18670 = n15147 ^ n7875 ^ 1'b0 ;
  assign n18671 = n1522 & n17610 ;
  assign n18672 = ~n1366 & n18671 ;
  assign n18673 = n831 & n2568 ;
  assign n18674 = n18673 ^ n4970 ^ 1'b0 ;
  assign n18675 = n18674 ^ n12993 ^ n7098 ;
  assign n18676 = ( n12809 & n13881 ) | ( n12809 & n16509 ) | ( n13881 & n16509 ) ;
  assign n18677 = n6861 ^ n5609 ^ 1'b0 ;
  assign n18678 = n2185 ^ n641 ^ 1'b0 ;
  assign n18679 = ~n18677 & n18678 ;
  assign n18680 = ~n2579 & n18679 ;
  assign n18681 = n2398 & ~n5306 ;
  assign n18682 = ( n1651 & n9560 ) | ( n1651 & n18681 ) | ( n9560 & n18681 ) ;
  assign n18683 = n5578 | n14576 ;
  assign n18684 = n16838 & ~n18683 ;
  assign n18685 = n1659 & n18684 ;
  assign n18686 = n7725 ^ n386 ^ 1'b0 ;
  assign n18687 = n8488 | n18686 ;
  assign n18688 = n15352 | n18687 ;
  assign n18689 = ( ~x51 & n591 ) | ( ~x51 & n3148 ) | ( n591 & n3148 ) ;
  assign n18690 = n18689 ^ n15051 ^ n8425 ;
  assign n18694 = n4117 & n14193 ;
  assign n18691 = n14180 ^ n9112 ^ 1'b0 ;
  assign n18692 = n3644 & n18691 ;
  assign n18693 = n17770 & n18692 ;
  assign n18695 = n18694 ^ n18693 ^ n16808 ;
  assign n18696 = ( n748 & n2989 ) | ( n748 & ~n11975 ) | ( n2989 & ~n11975 ) ;
  assign n18697 = n16817 ^ n11541 ^ n8002 ;
  assign n18698 = ~n1350 & n12653 ;
  assign n18699 = ( n4561 & ~n11941 ) | ( n4561 & n18698 ) | ( ~n11941 & n18698 ) ;
  assign n18700 = ( ~n12324 & n18697 ) | ( ~n12324 & n18699 ) | ( n18697 & n18699 ) ;
  assign n18701 = n17151 ^ n4708 ^ 1'b0 ;
  assign n18702 = n235 & n18701 ;
  assign n18703 = n11927 & n15903 ;
  assign n18704 = ( n10830 & n18702 ) | ( n10830 & n18703 ) | ( n18702 & n18703 ) ;
  assign n18705 = ~n1085 & n1669 ;
  assign n18706 = n18705 ^ n14566 ^ 1'b0 ;
  assign n18707 = n13298 & n18706 ;
  assign n18708 = n4543 | n18707 ;
  assign n18709 = ( n1346 & ~n2941 ) | ( n1346 & n17586 ) | ( ~n2941 & n17586 ) ;
  assign n18710 = ~n11148 & n18709 ;
  assign n18711 = ( n451 & n2948 ) | ( n451 & n3295 ) | ( n2948 & n3295 ) ;
  assign n18712 = n4891 ^ n3131 ^ 1'b0 ;
  assign n18713 = n15206 & ~n18712 ;
  assign n18714 = ( n7855 & n8198 ) | ( n7855 & ~n12058 ) | ( n8198 & ~n12058 ) ;
  assign n18715 = ( n18711 & ~n18713 ) | ( n18711 & n18714 ) | ( ~n18713 & n18714 ) ;
  assign n18716 = ( n3975 & n10205 ) | ( n3975 & n18715 ) | ( n10205 & n18715 ) ;
  assign n18717 = ( ~n571 & n9354 ) | ( ~n571 & n16252 ) | ( n9354 & n16252 ) ;
  assign n18719 = n6639 ^ n277 ^ 1'b0 ;
  assign n18720 = n2763 | n18719 ;
  assign n18721 = ( n8482 & n18449 ) | ( n8482 & n18720 ) | ( n18449 & n18720 ) ;
  assign n18718 = n11283 & ~n14481 ;
  assign n18722 = n18721 ^ n18718 ^ 1'b0 ;
  assign n18723 = n17426 ^ n4972 ^ 1'b0 ;
  assign n18724 = n3362 | n18723 ;
  assign n18725 = n1800 & ~n18724 ;
  assign n18726 = n15585 & n18725 ;
  assign n18727 = ( ~x46 & n6990 ) | ( ~x46 & n13263 ) | ( n6990 & n13263 ) ;
  assign n18728 = n8309 ^ n4791 ^ n1120 ;
  assign n18729 = n18727 & ~n18728 ;
  assign n18730 = n18729 ^ n10333 ^ 1'b0 ;
  assign n18731 = n16462 | n17976 ;
  assign n18732 = n18730 & ~n18731 ;
  assign n18733 = ( n1085 & n7882 ) | ( n1085 & ~n12314 ) | ( n7882 & ~n12314 ) ;
  assign n18734 = n1798 | n10058 ;
  assign n18735 = n1663 | n18734 ;
  assign n18736 = ( n15110 & n18733 ) | ( n15110 & ~n18735 ) | ( n18733 & ~n18735 ) ;
  assign n18737 = n14307 | n18736 ;
  assign n18738 = ( n4800 & n14049 ) | ( n4800 & n14810 ) | ( n14049 & n14810 ) ;
  assign n18739 = ( n7940 & ~n9717 ) | ( n7940 & n11779 ) | ( ~n9717 & n11779 ) ;
  assign n18741 = n8279 ^ n6289 ^ n1708 ;
  assign n18740 = n7015 ^ n3130 ^ n2070 ;
  assign n18742 = n18741 ^ n18740 ^ 1'b0 ;
  assign n18743 = ( n5544 & ~n9292 ) | ( n5544 & n14770 ) | ( ~n9292 & n14770 ) ;
  assign n18744 = n9524 ^ n4702 ^ n280 ;
  assign n18745 = n18744 ^ n6810 ^ n2366 ;
  assign n18746 = ~n3089 & n18745 ;
  assign n18747 = n17979 ^ n6172 ^ 1'b0 ;
  assign n18748 = ( n11118 & n14301 ) | ( n11118 & ~n14872 ) | ( n14301 & ~n14872 ) ;
  assign n18749 = n15931 & ~n18748 ;
  assign n18750 = ~n9175 & n18749 ;
  assign n18751 = ~n7563 & n8904 ;
  assign n18752 = ~x126 & n18751 ;
  assign n18753 = n233 & n4540 ;
  assign n18754 = n9418 | n18753 ;
  assign n18755 = n18754 ^ n7843 ^ 1'b0 ;
  assign n18756 = ( n4556 & n18752 ) | ( n4556 & ~n18755 ) | ( n18752 & ~n18755 ) ;
  assign n18757 = n18756 ^ n16549 ^ n16288 ;
  assign n18758 = n5655 ^ n2965 ^ 1'b0 ;
  assign n18759 = n11763 | n18758 ;
  assign n18760 = ( n3140 & ~n11129 ) | ( n3140 & n18759 ) | ( ~n11129 & n18759 ) ;
  assign n18761 = n9792 ^ n5052 ^ 1'b0 ;
  assign n18762 = ( n6446 & n10174 ) | ( n6446 & ~n18761 ) | ( n10174 & ~n18761 ) ;
  assign n18763 = ( n1228 & ~n1291 ) | ( n1228 & n3395 ) | ( ~n1291 & n3395 ) ;
  assign n18764 = n18763 ^ n5808 ^ n3927 ;
  assign n18765 = n7292 ^ n3864 ^ n2491 ;
  assign n18766 = ( n13054 & n17305 ) | ( n13054 & ~n18765 ) | ( n17305 & ~n18765 ) ;
  assign n18767 = ~n5309 & n12377 ;
  assign n18768 = ~n2461 & n18767 ;
  assign n18769 = n4143 & n18768 ;
  assign n18770 = n17535 ^ n17466 ^ 1'b0 ;
  assign n18771 = n11225 | n16431 ;
  assign n18772 = n15338 ^ n13479 ^ n5559 ;
  assign n18773 = ( n9023 & n11144 ) | ( n9023 & ~n17315 ) | ( n11144 & ~n17315 ) ;
  assign n18774 = ~n11577 & n14688 ;
  assign n18775 = ( n6327 & n9369 ) | ( n6327 & ~n18774 ) | ( n9369 & ~n18774 ) ;
  assign n18776 = n5050 ^ n870 ^ n213 ;
  assign n18777 = n5929 | n18776 ;
  assign n18780 = ( n402 & n3056 ) | ( n402 & n3765 ) | ( n3056 & n3765 ) ;
  assign n18778 = n6325 & ~n15759 ;
  assign n18779 = n16437 & n18778 ;
  assign n18781 = n18780 ^ n18779 ^ 1'b0 ;
  assign n18782 = n10845 | n16978 ;
  assign n18783 = n18782 ^ n1067 ^ 1'b0 ;
  assign n18784 = ( n2954 & ~n6581 ) | ( n2954 & n18783 ) | ( ~n6581 & n18783 ) ;
  assign n18785 = ( x106 & n6134 ) | ( x106 & n10906 ) | ( n6134 & n10906 ) ;
  assign n18786 = ( ~n15502 & n18015 ) | ( ~n15502 & n18785 ) | ( n18015 & n18785 ) ;
  assign n18787 = n930 | n10568 ;
  assign n18788 = n18787 ^ n13072 ^ 1'b0 ;
  assign n18789 = ( n2279 & n2439 ) | ( n2279 & ~n3358 ) | ( n2439 & ~n3358 ) ;
  assign n18790 = n18789 ^ n17881 ^ n2952 ;
  assign n18791 = n12904 ^ n2907 ^ 1'b0 ;
  assign n18792 = n5358 & ~n18791 ;
  assign n18793 = n17530 ^ n3636 ^ n1024 ;
  assign n18794 = ( n589 & ~n5179 ) | ( n589 & n8058 ) | ( ~n5179 & n8058 ) ;
  assign n18795 = ~n14330 & n18794 ;
  assign n18796 = n18795 ^ n13458 ^ 1'b0 ;
  assign n18797 = n13036 ^ n8255 ^ n4459 ;
  assign n18798 = ( n6008 & n16748 ) | ( n6008 & ~n18797 ) | ( n16748 & ~n18797 ) ;
  assign n18799 = n9419 ^ n9336 ^ n5685 ;
  assign n18800 = n5697 & n6090 ;
  assign n18801 = n18800 ^ n3518 ^ 1'b0 ;
  assign n18802 = ( ~n3982 & n4015 ) | ( ~n3982 & n18801 ) | ( n4015 & n18801 ) ;
  assign n18803 = n4290 & n5279 ;
  assign n18804 = n18803 ^ n4029 ^ 1'b0 ;
  assign n18805 = n5313 | n18804 ;
  assign n18806 = ~n889 & n18805 ;
  assign n18807 = n6132 & n18806 ;
  assign n18808 = ( n5071 & ~n6816 ) | ( n5071 & n18807 ) | ( ~n6816 & n18807 ) ;
  assign n18809 = n14899 ^ n13912 ^ n8839 ;
  assign n18810 = n12053 ^ n8156 ^ n461 ;
  assign n18811 = n8509 ^ n4408 ^ 1'b0 ;
  assign n18812 = ~n18810 & n18811 ;
  assign n18813 = n8892 ^ n2216 ^ n611 ;
  assign n18814 = n18813 ^ n13297 ^ n6024 ;
  assign n18815 = n3573 & n18814 ;
  assign n18816 = n18815 ^ n4489 ^ 1'b0 ;
  assign n18817 = ( ~n11788 & n15225 ) | ( ~n11788 & n15859 ) | ( n15225 & n15859 ) ;
  assign n18818 = n5515 ^ n1938 ^ 1'b0 ;
  assign n18819 = n6538 ^ n4169 ^ 1'b0 ;
  assign n18820 = ~n17244 & n18819 ;
  assign n18821 = n18820 ^ n6851 ^ n2111 ;
  assign n18822 = ( ~n11465 & n11496 ) | ( ~n11465 & n11796 ) | ( n11496 & n11796 ) ;
  assign n18823 = n7426 ^ n2826 ^ 1'b0 ;
  assign n18824 = n17884 ^ n7419 ^ n4375 ;
  assign n18825 = ~n10435 & n16128 ;
  assign n18826 = n18825 ^ n17835 ^ 1'b0 ;
  assign n18827 = n17771 ^ n6031 ^ 1'b0 ;
  assign n18828 = n3906 | n18827 ;
  assign n18829 = n3626 ^ n320 ^ 1'b0 ;
  assign n18830 = ( n1174 & n1343 ) | ( n1174 & ~n18829 ) | ( n1343 & ~n18829 ) ;
  assign n18831 = ~n3646 & n17442 ;
  assign n18832 = n18830 & n18831 ;
  assign n18833 = n18832 ^ n11229 ^ n8359 ;
  assign n18834 = n2951 | n9293 ;
  assign n18835 = n18834 ^ n11829 ^ n6591 ;
  assign n18836 = n5377 | n12319 ;
  assign n18837 = n9352 & ~n18836 ;
  assign n18838 = ( n12817 & ~n17728 ) | ( n12817 & n18837 ) | ( ~n17728 & n18837 ) ;
  assign n18839 = ( n7058 & ~n17552 ) | ( n7058 & n18838 ) | ( ~n17552 & n18838 ) ;
  assign n18840 = n12497 ^ n5248 ^ n3324 ;
  assign n18841 = n18243 & n18840 ;
  assign n18842 = n16309 ^ n11903 ^ n4302 ;
  assign n18845 = n13845 ^ n9146 ^ 1'b0 ;
  assign n18846 = ~n11486 & n18845 ;
  assign n18843 = ( n1686 & n5882 ) | ( n1686 & ~n7735 ) | ( n5882 & ~n7735 ) ;
  assign n18844 = n7348 & n18843 ;
  assign n18847 = n18846 ^ n18844 ^ 1'b0 ;
  assign n18848 = n18847 ^ n13982 ^ n13773 ;
  assign n18851 = n3008 & n12771 ;
  assign n18852 = n18851 ^ n18000 ^ 1'b0 ;
  assign n18849 = n16587 ^ n5783 ^ 1'b0 ;
  assign n18850 = n4634 | n18849 ;
  assign n18853 = n18852 ^ n18850 ^ n4663 ;
  assign n18855 = n9617 ^ n1201 ^ 1'b0 ;
  assign n18854 = n14564 ^ n6580 ^ n6321 ;
  assign n18856 = n18855 ^ n18854 ^ n3518 ;
  assign n18857 = ( ~n6820 & n7734 ) | ( ~n6820 & n8251 ) | ( n7734 & n8251 ) ;
  assign n18858 = ( n3076 & n10029 ) | ( n3076 & ~n18857 ) | ( n10029 & ~n18857 ) ;
  assign n18859 = n11061 ^ n6685 ^ n2619 ;
  assign n18860 = ( n4231 & n10039 ) | ( n4231 & ~n18859 ) | ( n10039 & ~n18859 ) ;
  assign n18861 = n3935 & ~n15507 ;
  assign n18862 = ~n11916 & n18861 ;
  assign n18863 = n6106 ^ n2008 ^ n1625 ;
  assign n18864 = n13664 ^ n8211 ^ n2994 ;
  assign n18865 = ( n6977 & n18863 ) | ( n6977 & n18864 ) | ( n18863 & n18864 ) ;
  assign n18866 = ( n12763 & ~n18862 ) | ( n12763 & n18865 ) | ( ~n18862 & n18865 ) ;
  assign n18867 = n9198 ^ n5790 ^ n5178 ;
  assign n18868 = ~n8615 & n18867 ;
  assign n18869 = n18868 ^ n18697 ^ n10623 ;
  assign n18870 = n6195 ^ n1020 ^ 1'b0 ;
  assign n18871 = ~n11631 & n18870 ;
  assign n18872 = n10269 & n18871 ;
  assign n18873 = n15375 & n18872 ;
  assign n18874 = n11068 ^ n2149 ^ 1'b0 ;
  assign n18881 = n10120 ^ n8503 ^ n3900 ;
  assign n18880 = n6432 ^ n3370 ^ n1954 ;
  assign n18875 = n2566 | n9685 ;
  assign n18876 = n4823 & ~n18875 ;
  assign n18877 = n8684 & ~n18876 ;
  assign n18878 = n18877 ^ n15181 ^ 1'b0 ;
  assign n18879 = n8302 & ~n18878 ;
  assign n18882 = n18881 ^ n18880 ^ n18879 ;
  assign n18883 = n1994 | n3889 ;
  assign n18884 = n18883 ^ n6029 ^ n2162 ;
  assign n18885 = ( n4805 & n15142 ) | ( n4805 & ~n18884 ) | ( n15142 & ~n18884 ) ;
  assign n18886 = n18885 ^ n18679 ^ 1'b0 ;
  assign n18887 = n18882 & ~n18886 ;
  assign n18894 = n1331 & n8475 ;
  assign n18895 = n18894 ^ n13328 ^ n8210 ;
  assign n18889 = n331 & ~n9386 ;
  assign n18890 = n1283 & n18889 ;
  assign n18891 = n18890 ^ n3270 ^ n3241 ;
  assign n18888 = n8321 | n11942 ;
  assign n18892 = n18891 ^ n18888 ^ 1'b0 ;
  assign n18893 = n15736 & ~n18892 ;
  assign n18896 = n18895 ^ n18893 ^ 1'b0 ;
  assign n18897 = n9997 ^ n3458 ^ n1259 ;
  assign n18905 = n18382 ^ n9988 ^ n1229 ;
  assign n18903 = n18797 ^ n9743 ^ n3981 ;
  assign n18904 = ( n6918 & n13497 ) | ( n6918 & n18903 ) | ( n13497 & n18903 ) ;
  assign n18898 = n10869 ^ n810 ^ 1'b0 ;
  assign n18899 = ~n9777 & n18898 ;
  assign n18900 = n18899 ^ n18073 ^ n16041 ;
  assign n18901 = n18138 & ~n18900 ;
  assign n18902 = n5656 & n18901 ;
  assign n18906 = n18905 ^ n18904 ^ n18902 ;
  assign n18907 = ~n4236 & n4607 ;
  assign n18908 = n16900 ^ n13700 ^ n3081 ;
  assign n18909 = ( n7121 & n9458 ) | ( n7121 & n17906 ) | ( n9458 & n17906 ) ;
  assign n18910 = n1017 & ~n15677 ;
  assign n18911 = n14969 & n18910 ;
  assign n18912 = n11521 ^ n7437 ^ n2337 ;
  assign n18913 = n8841 & n18912 ;
  assign n18914 = n18913 ^ n16946 ^ 1'b0 ;
  assign n18915 = ~n1940 & n18914 ;
  assign n18918 = n148 & n967 ;
  assign n18919 = n3059 & n18918 ;
  assign n18920 = n18919 ^ n5885 ^ 1'b0 ;
  assign n18921 = ~n1074 & n18920 ;
  assign n18916 = n417 & ~n4510 ;
  assign n18917 = n18916 ^ n6899 ^ 1'b0 ;
  assign n18922 = n18921 ^ n18917 ^ n1878 ;
  assign n18923 = n18922 ^ n11587 ^ n7086 ;
  assign n18924 = n18923 ^ n7957 ^ 1'b0 ;
  assign n18925 = n17265 ^ n11862 ^ x38 ;
  assign n18930 = ( n5389 & n11691 ) | ( n5389 & n18070 ) | ( n11691 & n18070 ) ;
  assign n18926 = ( n4844 & ~n13246 ) | ( n4844 & n16286 ) | ( ~n13246 & n16286 ) ;
  assign n18927 = n2894 | n18926 ;
  assign n18928 = n18927 ^ n2404 ^ 1'b0 ;
  assign n18929 = n18928 ^ n13521 ^ n851 ;
  assign n18931 = n18930 ^ n18929 ^ n5896 ;
  assign n18932 = n6715 ^ n267 ^ 1'b0 ;
  assign n18933 = ( n1648 & ~n9757 ) | ( n1648 & n13848 ) | ( ~n9757 & n13848 ) ;
  assign n18934 = ( ~n453 & n13818 ) | ( ~n453 & n15399 ) | ( n13818 & n15399 ) ;
  assign n18935 = n6237 & n18934 ;
  assign n18936 = n18933 | n18935 ;
  assign n18937 = n18932 & ~n18936 ;
  assign n18938 = ( n1015 & ~n2363 ) | ( n1015 & n6961 ) | ( ~n2363 & n6961 ) ;
  assign n18939 = n18938 ^ n2767 ^ n1314 ;
  assign n18940 = n13955 ^ n13243 ^ n6111 ;
  assign n18941 = ( n3599 & n4304 ) | ( n3599 & ~n11660 ) | ( n4304 & ~n11660 ) ;
  assign n18942 = n2179 | n18941 ;
  assign n18943 = n14839 | n18942 ;
  assign n18944 = ( n1486 & n4927 ) | ( n1486 & ~n11536 ) | ( n4927 & ~n11536 ) ;
  assign n18945 = ( n4919 & n8699 ) | ( n4919 & n18944 ) | ( n8699 & n18944 ) ;
  assign n18946 = ( n15314 & n16321 ) | ( n15314 & n18945 ) | ( n16321 & n18945 ) ;
  assign n18947 = n18946 ^ n11181 ^ n7296 ;
  assign n18948 = n18586 ^ n4191 ^ n2862 ;
  assign n18949 = n18948 ^ n17665 ^ 1'b0 ;
  assign n18951 = n11236 ^ n8681 ^ 1'b0 ;
  assign n18952 = n5027 & n18951 ;
  assign n18953 = ( n1565 & n11821 ) | ( n1565 & n18952 ) | ( n11821 & n18952 ) ;
  assign n18950 = n18303 ^ n14727 ^ 1'b0 ;
  assign n18954 = n18953 ^ n18950 ^ n2765 ;
  assign n18955 = ( n6656 & n10720 ) | ( n6656 & n11864 ) | ( n10720 & n11864 ) ;
  assign n18956 = ( n4467 & n6748 ) | ( n4467 & n8513 ) | ( n6748 & n8513 ) ;
  assign n18957 = n15144 | n18956 ;
  assign n18958 = ( n12732 & n13659 ) | ( n12732 & n18957 ) | ( n13659 & n18957 ) ;
  assign n18959 = ( n7216 & n7962 ) | ( n7216 & n18958 ) | ( n7962 & n18958 ) ;
  assign n18962 = n13331 ^ n10526 ^ n6692 ;
  assign n18960 = n11315 & ~n16189 ;
  assign n18961 = ~n14823 & n18960 ;
  assign n18963 = n18962 ^ n18961 ^ n5442 ;
  assign n18964 = n12399 ^ n9441 ^ 1'b0 ;
  assign n18965 = n18964 ^ n8318 ^ n7269 ;
  assign n18966 = ( n5643 & ~n15578 ) | ( n5643 & n17542 ) | ( ~n15578 & n17542 ) ;
  assign n18967 = ~n6538 & n17017 ;
  assign n18968 = ~n18966 & n18967 ;
  assign n18969 = n2016 | n17280 ;
  assign n18970 = n2716 | n18969 ;
  assign n18971 = ~n959 & n2596 ;
  assign n18972 = n18971 ^ n495 ^ 1'b0 ;
  assign n18973 = ( n2792 & n12504 ) | ( n2792 & n18972 ) | ( n12504 & n18972 ) ;
  assign n18974 = n18343 ^ n17400 ^ n16572 ;
  assign n18976 = n10937 ^ n7977 ^ n4329 ;
  assign n18977 = ( n5678 & ~n18541 ) | ( n5678 & n18976 ) | ( ~n18541 & n18976 ) ;
  assign n18975 = n6477 & ~n16387 ;
  assign n18978 = n18977 ^ n18975 ^ 1'b0 ;
  assign n18979 = n15151 ^ n4470 ^ 1'b0 ;
  assign n18980 = n3795 & ~n18979 ;
  assign n18981 = ( ~n1795 & n4804 ) | ( ~n1795 & n18980 ) | ( n4804 & n18980 ) ;
  assign n18982 = ( n8084 & n8412 ) | ( n8084 & n10730 ) | ( n8412 & n10730 ) ;
  assign n18983 = ( n954 & ~n18981 ) | ( n954 & n18982 ) | ( ~n18981 & n18982 ) ;
  assign n18984 = n17611 & ~n18983 ;
  assign n18985 = n18984 ^ n2812 ^ 1'b0 ;
  assign n18986 = n11211 ^ n7577 ^ n1028 ;
  assign n18987 = n8624 ^ n716 ^ 1'b0 ;
  assign n18992 = n9834 ^ n5374 ^ n3318 ;
  assign n18993 = n9404 & n18992 ;
  assign n18994 = n15993 & n18993 ;
  assign n18990 = ( n6640 & ~n8552 ) | ( n6640 & n8839 ) | ( ~n8552 & n8839 ) ;
  assign n18991 = n15798 & ~n18990 ;
  assign n18995 = n18994 ^ n18991 ^ 1'b0 ;
  assign n18988 = ~n5523 & n11622 ;
  assign n18989 = ~n9892 & n18988 ;
  assign n18996 = n18995 ^ n18989 ^ n1940 ;
  assign n18997 = n6521 ^ n2747 ^ 1'b0 ;
  assign n18999 = n4154 ^ n827 ^ 1'b0 ;
  assign n19000 = n3723 & n18999 ;
  assign n18998 = n11503 ^ n6956 ^ n6697 ;
  assign n19001 = n19000 ^ n18998 ^ n12983 ;
  assign n19002 = n19001 ^ n17531 ^ x34 ;
  assign n19003 = ( n4150 & ~n5429 ) | ( n4150 & n19002 ) | ( ~n5429 & n19002 ) ;
  assign n19004 = ~n13969 & n16273 ;
  assign n19005 = ~n3329 & n14006 ;
  assign n19006 = n19005 ^ n3666 ^ n709 ;
  assign n19007 = n19006 ^ n13034 ^ n4469 ;
  assign n19008 = n19007 ^ n3866 ^ n1773 ;
  assign n19009 = n19008 ^ n9010 ^ n7892 ;
  assign n19010 = n3208 | n6990 ;
  assign n19011 = n19010 ^ n7868 ^ n4926 ;
  assign n19012 = n9105 ^ n5655 ^ 1'b0 ;
  assign n19015 = ~n13276 & n18992 ;
  assign n19013 = ( ~n4905 & n5449 ) | ( ~n4905 & n9549 ) | ( n5449 & n9549 ) ;
  assign n19014 = ~n16688 & n19013 ;
  assign n19016 = n19015 ^ n19014 ^ 1'b0 ;
  assign n19017 = n3926 & n4503 ;
  assign n19018 = n10942 ^ n10034 ^ 1'b0 ;
  assign n19019 = n19017 | n19018 ;
  assign n19020 = ( n2646 & n3670 ) | ( n2646 & ~n17376 ) | ( n3670 & ~n17376 ) ;
  assign n19021 = n14988 ^ n1763 ^ 1'b0 ;
  assign n19022 = n19021 ^ n9897 ^ n9227 ;
  assign n19023 = ( n2670 & n14240 ) | ( n2670 & ~n19022 ) | ( n14240 & ~n19022 ) ;
  assign n19024 = ( n5876 & ~n16066 ) | ( n5876 & n19023 ) | ( ~n16066 & n19023 ) ;
  assign n19025 = n6062 & ~n18393 ;
  assign n19027 = n12139 ^ n6024 ^ n2754 ;
  assign n19028 = ( n4115 & n17394 ) | ( n4115 & ~n19027 ) | ( n17394 & ~n19027 ) ;
  assign n19026 = ( ~n2592 & n4905 ) | ( ~n2592 & n13804 ) | ( n4905 & n13804 ) ;
  assign n19029 = n19028 ^ n19026 ^ n1467 ;
  assign n19030 = n12454 ^ n6907 ^ n2039 ;
  assign n19032 = n13437 ^ n9632 ^ n2665 ;
  assign n19031 = n8314 ^ n6910 ^ 1'b0 ;
  assign n19033 = n19032 ^ n19031 ^ n986 ;
  assign n19034 = n8919 | n15902 ;
  assign n19035 = n19034 ^ n12266 ^ n10618 ;
  assign n19036 = ( x67 & n568 ) | ( x67 & n6713 ) | ( n568 & n6713 ) ;
  assign n19037 = n8695 & n19036 ;
  assign n19038 = n7277 & n19037 ;
  assign n19039 = n14974 ^ n10438 ^ n9898 ;
  assign n19040 = ( n2810 & n7928 ) | ( n2810 & n19039 ) | ( n7928 & n19039 ) ;
  assign n19046 = ~n7947 & n17382 ;
  assign n19047 = n19046 ^ n12945 ^ n3014 ;
  assign n19043 = ( n3085 & ~n9059 ) | ( n3085 & n10641 ) | ( ~n9059 & n10641 ) ;
  assign n19042 = x9 & n6440 ;
  assign n19044 = n19043 ^ n19042 ^ n6487 ;
  assign n19041 = ( ~n2036 & n7114 ) | ( ~n2036 & n9643 ) | ( n7114 & n9643 ) ;
  assign n19045 = n19044 ^ n19041 ^ 1'b0 ;
  assign n19048 = n19047 ^ n19045 ^ n14401 ;
  assign n19049 = ( n5812 & ~n19040 ) | ( n5812 & n19048 ) | ( ~n19040 & n19048 ) ;
  assign n19050 = n19049 ^ n11755 ^ 1'b0 ;
  assign n19051 = ~n2404 & n19050 ;
  assign n19052 = n14389 ^ n6568 ^ n3061 ;
  assign n19053 = n3268 & ~n18469 ;
  assign n19054 = n19053 ^ n8136 ^ 1'b0 ;
  assign n19055 = n19054 ^ n12075 ^ 1'b0 ;
  assign n19056 = ~n10405 & n19055 ;
  assign n19057 = ~n16371 & n19056 ;
  assign n19059 = n2917 | n4657 ;
  assign n19058 = ( ~n636 & n8888 ) | ( ~n636 & n18382 ) | ( n8888 & n18382 ) ;
  assign n19060 = n19059 ^ n19058 ^ n2531 ;
  assign n19061 = ( ~n1808 & n15090 ) | ( ~n1808 & n18401 ) | ( n15090 & n18401 ) ;
  assign n19062 = n18213 ^ n9133 ^ n1395 ;
  assign n19063 = n17145 ^ n2590 ^ 1'b0 ;
  assign n19064 = n1771 | n19063 ;
  assign n19065 = ( n7333 & n9653 ) | ( n7333 & n19064 ) | ( n9653 & n19064 ) ;
  assign n19066 = ( n2897 & n19062 ) | ( n2897 & ~n19065 ) | ( n19062 & ~n19065 ) ;
  assign n19067 = ( n3165 & ~n3529 ) | ( n3165 & n10659 ) | ( ~n3529 & n10659 ) ;
  assign n19068 = n17737 ^ n10460 ^ n1361 ;
  assign n19069 = ( n3227 & n13549 ) | ( n3227 & ~n19068 ) | ( n13549 & ~n19068 ) ;
  assign n19070 = n9344 | n19069 ;
  assign n19071 = n19067 & ~n19070 ;
  assign n19072 = n5999 ^ n3697 ^ x110 ;
  assign n19073 = ~n766 & n19072 ;
  assign n19074 = n17283 ^ n5707 ^ x89 ;
  assign n19075 = ( ~n7416 & n17020 ) | ( ~n7416 & n19074 ) | ( n17020 & n19074 ) ;
  assign n19077 = ( n3533 & n5802 ) | ( n3533 & ~n13335 ) | ( n5802 & ~n13335 ) ;
  assign n19078 = ( n184 & n2178 ) | ( n184 & ~n19077 ) | ( n2178 & ~n19077 ) ;
  assign n19076 = n3654 ^ n2685 ^ n2163 ;
  assign n19079 = n19078 ^ n19076 ^ n13270 ;
  assign n19080 = n10392 ^ n1418 ^ 1'b0 ;
  assign n19081 = n19080 ^ n1621 ^ n146 ;
  assign n19082 = ( n9443 & n10971 ) | ( n9443 & n17707 ) | ( n10971 & n17707 ) ;
  assign n19083 = n14151 ^ n5777 ^ n2823 ;
  assign n19084 = ( n3265 & ~n8396 ) | ( n3265 & n19083 ) | ( ~n8396 & n19083 ) ;
  assign n19085 = n514 & n11087 ;
  assign n19086 = n19085 ^ n11067 ^ n5935 ;
  assign n19087 = n19086 ^ n11199 ^ n6285 ;
  assign n19088 = ( n12076 & n17344 ) | ( n12076 & ~n19087 ) | ( n17344 & ~n19087 ) ;
  assign n19089 = ( n4346 & ~n19084 ) | ( n4346 & n19088 ) | ( ~n19084 & n19088 ) ;
  assign n19090 = ( n1822 & ~n3738 ) | ( n1822 & n15060 ) | ( ~n3738 & n15060 ) ;
  assign n19091 = n12414 ^ n5596 ^ n1755 ;
  assign n19092 = n19091 ^ n7013 ^ 1'b0 ;
  assign n19093 = ~n12455 & n19092 ;
  assign n19094 = ( n9443 & n19090 ) | ( n9443 & ~n19093 ) | ( n19090 & ~n19093 ) ;
  assign n19095 = n5379 & n19094 ;
  assign n19096 = ~n640 & n19095 ;
  assign n19097 = n8462 & n12648 ;
  assign n19098 = ~n2801 & n19097 ;
  assign n19099 = n3348 ^ n748 ^ 1'b0 ;
  assign n19100 = n19099 ^ n14947 ^ n6078 ;
  assign n19101 = ( ~n12509 & n13728 ) | ( ~n12509 & n19100 ) | ( n13728 & n19100 ) ;
  assign n19102 = ( n4067 & ~n19098 ) | ( n4067 & n19101 ) | ( ~n19098 & n19101 ) ;
  assign n19104 = ~n2501 & n10566 ;
  assign n19105 = ~n2972 & n19104 ;
  assign n19106 = n3330 | n19105 ;
  assign n19107 = n19106 ^ n6150 ^ 1'b0 ;
  assign n19103 = ( n3947 & n8082 ) | ( n3947 & n14146 ) | ( n8082 & n14146 ) ;
  assign n19108 = n19107 ^ n19103 ^ 1'b0 ;
  assign n19109 = n17606 ^ n10730 ^ n5554 ;
  assign n19110 = n18198 ^ n17401 ^ 1'b0 ;
  assign n19111 = n13833 ^ n6754 ^ n440 ;
  assign n19112 = n3252 & n16194 ;
  assign n19113 = ( n2790 & n19111 ) | ( n2790 & n19112 ) | ( n19111 & n19112 ) ;
  assign n19114 = n8794 & n18284 ;
  assign n19115 = ~n10746 & n10786 ;
  assign n19116 = n3748 & n19115 ;
  assign n19117 = n19116 ^ n18233 ^ n6897 ;
  assign n19118 = n1647 | n19117 ;
  assign n19119 = n19118 ^ n9586 ^ 1'b0 ;
  assign n19120 = n6966 ^ n6043 ^ 1'b0 ;
  assign n19121 = n11814 | n19120 ;
  assign n19122 = n6058 | n15412 ;
  assign n19123 = n19122 ^ n2234 ^ 1'b0 ;
  assign n19124 = n16833 ^ n10106 ^ 1'b0 ;
  assign n19125 = n721 & n954 ;
  assign n19126 = ( n7704 & n8010 ) | ( n7704 & ~n8862 ) | ( n8010 & ~n8862 ) ;
  assign n19127 = n8865 ^ n6661 ^ 1'b0 ;
  assign n19128 = n19126 | n19127 ;
  assign n19129 = ( n6510 & n11393 ) | ( n6510 & n19128 ) | ( n11393 & n19128 ) ;
  assign n19130 = ( n1366 & n5356 ) | ( n1366 & ~n19129 ) | ( n5356 & ~n19129 ) ;
  assign n19131 = n13304 ^ n4257 ^ 1'b0 ;
  assign n19133 = n17895 ^ n13695 ^ n1856 ;
  assign n19132 = n201 & n3381 ;
  assign n19134 = n19133 ^ n19132 ^ 1'b0 ;
  assign n19135 = n15264 ^ n11920 ^ n10708 ;
  assign n19136 = n382 & n19135 ;
  assign n19139 = n8629 & ~n13475 ;
  assign n19140 = n721 & n7713 ;
  assign n19141 = ~n19139 & n19140 ;
  assign n19137 = ( n2816 & ~n3705 ) | ( n2816 & n17106 ) | ( ~n3705 & n17106 ) ;
  assign n19138 = n1571 | n19137 ;
  assign n19142 = n19141 ^ n19138 ^ 1'b0 ;
  assign n19143 = ( n5132 & n19136 ) | ( n5132 & n19142 ) | ( n19136 & n19142 ) ;
  assign n19144 = n5658 ^ n2077 ^ 1'b0 ;
  assign n19145 = n18842 | n19144 ;
  assign n19146 = n19143 & ~n19145 ;
  assign n19147 = ( ~n9382 & n14669 ) | ( ~n9382 & n14950 ) | ( n14669 & n14950 ) ;
  assign n19148 = n8537 ^ n3959 ^ 1'b0 ;
  assign n19149 = ( n2360 & ~n3735 ) | ( n2360 & n10102 ) | ( ~n3735 & n10102 ) ;
  assign n19150 = ( ~n5381 & n10271 ) | ( ~n5381 & n15772 ) | ( n10271 & n15772 ) ;
  assign n19151 = ( n13938 & n18763 ) | ( n13938 & ~n19150 ) | ( n18763 & ~n19150 ) ;
  assign n19153 = n1882 & n5524 ;
  assign n19154 = ~n3537 & n19153 ;
  assign n19155 = n19154 ^ n9579 ^ n2491 ;
  assign n19152 = n4687 | n9541 ;
  assign n19156 = n19155 ^ n19152 ^ 1'b0 ;
  assign n19160 = n7429 | n14745 ;
  assign n19161 = n751 & ~n19160 ;
  assign n19157 = n13004 & n14877 ;
  assign n19158 = n1337 & n19157 ;
  assign n19159 = n19158 ^ n7844 ^ n131 ;
  assign n19162 = n19161 ^ n19159 ^ n6975 ;
  assign n19163 = ~n12427 & n19162 ;
  assign n19164 = ~n19156 & n19163 ;
  assign n19165 = n15648 ^ n14402 ^ n1540 ;
  assign n19166 = n4989 ^ n3779 ^ 1'b0 ;
  assign n19167 = n19165 & n19166 ;
  assign n19168 = ( ~n8520 & n12856 ) | ( ~n8520 & n14392 ) | ( n12856 & n14392 ) ;
  assign n19169 = n19168 ^ n11371 ^ 1'b0 ;
  assign n19170 = ~n5281 & n19169 ;
  assign n19171 = n11078 & ~n13109 ;
  assign n19172 = n19171 ^ x90 ^ 1'b0 ;
  assign n19173 = n6149 | n19172 ;
  assign n19174 = n19173 ^ n12352 ^ x27 ;
  assign n19175 = ~n2198 & n19174 ;
  assign n19176 = n19175 ^ n4830 ^ n434 ;
  assign n19177 = ( ~n2989 & n8475 ) | ( ~n2989 & n17059 ) | ( n8475 & n17059 ) ;
  assign n19178 = n4246 ^ n1033 ^ 1'b0 ;
  assign n19179 = ( n1708 & n16808 ) | ( n1708 & n19178 ) | ( n16808 & n19178 ) ;
  assign n19180 = ( n4078 & n13480 ) | ( n4078 & n19179 ) | ( n13480 & n19179 ) ;
  assign n19181 = n17127 ^ n3390 ^ n851 ;
  assign n19182 = n19181 ^ n16148 ^ n931 ;
  assign n19183 = n19182 ^ n4930 ^ n1414 ;
  assign n19184 = ( n4495 & n5525 ) | ( n4495 & ~n19183 ) | ( n5525 & ~n19183 ) ;
  assign n19185 = n6467 & n17450 ;
  assign n19186 = n19185 ^ n6363 ^ 1'b0 ;
  assign n19187 = n4674 & ~n15130 ;
  assign n19188 = ~n19186 & n19187 ;
  assign n19189 = n10718 | n14206 ;
  assign n19190 = ( n9887 & n15697 ) | ( n9887 & n19189 ) | ( n15697 & n19189 ) ;
  assign n19191 = n5024 ^ n3044 ^ n1207 ;
  assign n19192 = n7332 ^ n2234 ^ 1'b0 ;
  assign n19193 = n493 & ~n19192 ;
  assign n19194 = ( n1051 & ~n19191 ) | ( n1051 & n19193 ) | ( ~n19191 & n19193 ) ;
  assign n19195 = ( n4666 & ~n6403 ) | ( n4666 & n12650 ) | ( ~n6403 & n12650 ) ;
  assign n19196 = n8786 ^ n2907 ^ x100 ;
  assign n19197 = ( ~n6733 & n15065 ) | ( ~n6733 & n19196 ) | ( n15065 & n19196 ) ;
  assign n19198 = n16726 ^ n3853 ^ n430 ;
  assign n19199 = ( ~n11739 & n15246 ) | ( ~n11739 & n19198 ) | ( n15246 & n19198 ) ;
  assign n19200 = n17020 & ~n19199 ;
  assign n19202 = ( n3076 & n6530 ) | ( n3076 & ~n15825 ) | ( n6530 & ~n15825 ) ;
  assign n19201 = ( n11297 & n16491 ) | ( n11297 & ~n18891 ) | ( n16491 & ~n18891 ) ;
  assign n19203 = n19202 ^ n19201 ^ n15783 ;
  assign n19204 = ( n1889 & n12742 ) | ( n1889 & ~n18265 ) | ( n12742 & ~n18265 ) ;
  assign n19205 = ~n5364 & n8306 ;
  assign n19206 = n19204 & n19205 ;
  assign n19207 = n7154 | n18823 ;
  assign n19209 = n15460 ^ n14973 ^ 1'b0 ;
  assign n19208 = n3862 & ~n11819 ;
  assign n19210 = n19209 ^ n19208 ^ 1'b0 ;
  assign n19211 = n19210 ^ n12451 ^ 1'b0 ;
  assign n19212 = n19207 & n19211 ;
  assign n19213 = ~n1485 & n4437 ;
  assign n19214 = n16754 ^ n8852 ^ 1'b0 ;
  assign n19215 = n7853 & ~n19214 ;
  assign n19216 = n19215 ^ n3337 ^ 1'b0 ;
  assign n19217 = ( ~n3501 & n11760 ) | ( ~n3501 & n18185 ) | ( n11760 & n18185 ) ;
  assign n19218 = n15465 ^ n15444 ^ n348 ;
  assign n19219 = n18871 ^ n713 ^ 1'b0 ;
  assign n19220 = ~n9726 & n19219 ;
  assign n19221 = n19220 ^ n10384 ^ n6260 ;
  assign n19222 = n14741 ^ n7052 ^ n4963 ;
  assign n19223 = ( ~n864 & n2754 ) | ( ~n864 & n6274 ) | ( n2754 & n6274 ) ;
  assign n19224 = ( n4446 & n19222 ) | ( n4446 & n19223 ) | ( n19222 & n19223 ) ;
  assign n19225 = n2427 | n19224 ;
  assign n19226 = n19225 ^ n737 ^ 1'b0 ;
  assign n19227 = ( n5062 & n11792 ) | ( n5062 & ~n19226 ) | ( n11792 & ~n19226 ) ;
  assign n19228 = n11706 ^ n2930 ^ 1'b0 ;
  assign n19229 = n9802 & ~n19228 ;
  assign n19230 = n12072 ^ n10550 ^ 1'b0 ;
  assign n19231 = n19229 & ~n19230 ;
  assign n19232 = n7209 ^ n4524 ^ n3707 ;
  assign n19233 = ( ~n2721 & n6138 ) | ( ~n2721 & n9738 ) | ( n6138 & n9738 ) ;
  assign n19234 = n19233 ^ n18656 ^ 1'b0 ;
  assign n19235 = n19232 & ~n19234 ;
  assign n19236 = ( x65 & n1252 ) | ( x65 & ~n2425 ) | ( n1252 & ~n2425 ) ;
  assign n19237 = ( ~n2302 & n6173 ) | ( ~n2302 & n19236 ) | ( n6173 & n19236 ) ;
  assign n19238 = ( ~n3081 & n6274 ) | ( ~n3081 & n17254 ) | ( n6274 & n17254 ) ;
  assign n19239 = n18912 ^ n4225 ^ n3460 ;
  assign n19240 = ( n1525 & ~n4085 ) | ( n1525 & n9254 ) | ( ~n4085 & n9254 ) ;
  assign n19241 = ~n2212 & n19240 ;
  assign n19242 = n6971 & n19241 ;
  assign n19243 = ~n4717 & n19242 ;
  assign n19244 = n19243 ^ n2762 ^ n1161 ;
  assign n19245 = n2018 ^ n354 ^ 1'b0 ;
  assign n19246 = n9118 ^ n8992 ^ n1794 ;
  assign n19247 = ~n9330 & n19246 ;
  assign n19248 = ~n19245 & n19247 ;
  assign n19249 = n2126 ^ n1679 ^ 1'b0 ;
  assign n19250 = ~n5415 & n19249 ;
  assign n19251 = ( ~n2714 & n12144 ) | ( ~n2714 & n15213 ) | ( n12144 & n15213 ) ;
  assign n19252 = n9048 & n11984 ;
  assign n19253 = n19252 ^ n2316 ^ 1'b0 ;
  assign n19254 = ( n3395 & n6701 ) | ( n3395 & ~n8865 ) | ( n6701 & ~n8865 ) ;
  assign n19255 = ( n789 & n19253 ) | ( n789 & n19254 ) | ( n19253 & n19254 ) ;
  assign n19257 = ( n699 & n1780 ) | ( n699 & n5948 ) | ( n1780 & n5948 ) ;
  assign n19258 = n19257 ^ n5915 ^ 1'b0 ;
  assign n19259 = ( ~n1480 & n6465 ) | ( ~n1480 & n19258 ) | ( n6465 & n19258 ) ;
  assign n19256 = n14206 ^ n7902 ^ n3316 ;
  assign n19260 = n19259 ^ n19256 ^ n7948 ;
  assign n19263 = ( ~n1465 & n2541 ) | ( ~n1465 & n4667 ) | ( n2541 & n4667 ) ;
  assign n19264 = n1476 | n19263 ;
  assign n19265 = n19264 ^ n14956 ^ 1'b0 ;
  assign n19266 = n2801 & ~n19265 ;
  assign n19261 = n11819 | n14618 ;
  assign n19262 = n19261 ^ n12271 ^ 1'b0 ;
  assign n19267 = n19266 ^ n19262 ^ n10830 ;
  assign n19268 = n7757 ^ n5192 ^ n638 ;
  assign n19269 = n19268 ^ n19238 ^ 1'b0 ;
  assign n19270 = n8244 & ~n18432 ;
  assign n19271 = n10229 & n19270 ;
  assign n19272 = n14603 | n15049 ;
  assign n19273 = n19272 ^ n5093 ^ 1'b0 ;
  assign n19274 = n19271 | n19273 ;
  assign n19275 = ( ~n2813 & n7584 ) | ( ~n2813 & n14340 ) | ( n7584 & n14340 ) ;
  assign n19276 = n4227 ^ n3458 ^ n3083 ;
  assign n19277 = ( ~n1290 & n19275 ) | ( ~n1290 & n19276 ) | ( n19275 & n19276 ) ;
  assign n19278 = n19277 ^ n10858 ^ 1'b0 ;
  assign n19282 = n2619 ^ n1280 ^ n333 ;
  assign n19280 = n7568 | n10110 ;
  assign n19281 = ( n3365 & n11182 ) | ( n3365 & ~n19280 ) | ( n11182 & ~n19280 ) ;
  assign n19283 = n19282 ^ n19281 ^ n857 ;
  assign n19279 = n12666 ^ n4527 ^ 1'b0 ;
  assign n19284 = n19283 ^ n19279 ^ n10680 ;
  assign n19285 = n19284 ^ n4495 ^ 1'b0 ;
  assign n19286 = ( n4832 & n9222 ) | ( n4832 & ~n11241 ) | ( n9222 & ~n11241 ) ;
  assign n19287 = n14184 ^ n4606 ^ 1'b0 ;
  assign n19288 = n16327 & n19287 ;
  assign n19289 = n4363 | n8855 ;
  assign n19290 = n19289 ^ n2152 ^ 1'b0 ;
  assign n19291 = ~n13227 & n16395 ;
  assign n19292 = n19291 ^ n10944 ^ 1'b0 ;
  assign n19295 = ( x43 & n3510 ) | ( x43 & ~n3867 ) | ( n3510 & ~n3867 ) ;
  assign n19293 = ( ~n1617 & n1638 ) | ( ~n1617 & n7301 ) | ( n1638 & n7301 ) ;
  assign n19294 = n13628 & ~n19293 ;
  assign n19296 = n19295 ^ n19294 ^ n1753 ;
  assign n19297 = n17973 ^ n6087 ^ 1'b0 ;
  assign n19298 = n3534 & ~n19297 ;
  assign n19299 = ~n19296 & n19298 ;
  assign n19300 = ( ~n650 & n1969 ) | ( ~n650 & n14420 ) | ( n1969 & n14420 ) ;
  assign n19301 = n19300 ^ n11241 ^ 1'b0 ;
  assign n19302 = n19301 ^ n15949 ^ n8868 ;
  assign n19303 = ( ~n2097 & n7620 ) | ( ~n2097 & n11128 ) | ( n7620 & n11128 ) ;
  assign n19304 = n17531 ^ n12502 ^ n6873 ;
  assign n19305 = n19304 ^ n11748 ^ n3704 ;
  assign n19306 = n19058 ^ n6509 ^ n6385 ;
  assign n19307 = n436 | n14939 ;
  assign n19308 = n19307 ^ n8826 ^ 1'b0 ;
  assign n19309 = n4504 & n9584 ;
  assign n19310 = n11623 & n19309 ;
  assign n19311 = n16091 & ~n19310 ;
  assign n19312 = n19311 ^ n12703 ^ 1'b0 ;
  assign n19313 = n3081 | n16495 ;
  assign n19314 = ( n330 & n3058 ) | ( n330 & n5986 ) | ( n3058 & n5986 ) ;
  assign n19315 = ~n13430 & n19314 ;
  assign n19316 = n2606 & n19315 ;
  assign n19317 = n19316 ^ n11318 ^ 1'b0 ;
  assign n19318 = ~n7404 & n19317 ;
  assign n19319 = ( n17431 & n18745 ) | ( n17431 & ~n19318 ) | ( n18745 & ~n19318 ) ;
  assign n19320 = n5228 ^ n4116 ^ x34 ;
  assign n19321 = n18864 ^ n10261 ^ n3653 ;
  assign n19322 = n18514 ^ n2960 ^ n1667 ;
  assign n19323 = ( n306 & n8041 ) | ( n306 & ~n19322 ) | ( n8041 & ~n19322 ) ;
  assign n19324 = ( n459 & n6508 ) | ( n459 & ~n11834 ) | ( n6508 & ~n11834 ) ;
  assign n19325 = n7943 | n17325 ;
  assign n19326 = n19325 ^ n10075 ^ 1'b0 ;
  assign n19329 = n7688 ^ n4344 ^ n1047 ;
  assign n19330 = n1612 & ~n1738 ;
  assign n19331 = n19329 & n19330 ;
  assign n19332 = n19331 ^ n17284 ^ 1'b0 ;
  assign n19327 = n13866 ^ n3824 ^ n2906 ;
  assign n19328 = n378 & n19327 ;
  assign n19333 = n19332 ^ n19328 ^ 1'b0 ;
  assign n19334 = n2772 & ~n14975 ;
  assign n19335 = n4915 & n19334 ;
  assign n19336 = ~n2292 & n19335 ;
  assign n19337 = n19336 ^ n7161 ^ n6752 ;
  assign n19338 = ~n4240 & n8097 ;
  assign n19339 = n19338 ^ n7260 ^ 1'b0 ;
  assign n19340 = n4161 & n19339 ;
  assign n19341 = n9598 & ~n11100 ;
  assign n19342 = ~n4744 & n19341 ;
  assign n19343 = n19342 ^ n4430 ^ 1'b0 ;
  assign n19344 = ~n17025 & n19343 ;
  assign n19345 = n11236 | n13198 ;
  assign n19346 = n19344 | n19345 ;
  assign n19347 = ( n1840 & n19340 ) | ( n1840 & n19346 ) | ( n19340 & n19346 ) ;
  assign n19348 = n9727 ^ n5075 ^ n3306 ;
  assign n19349 = n19348 ^ n16751 ^ 1'b0 ;
  assign n19350 = ~n4656 & n8632 ;
  assign n19351 = n19350 ^ n1824 ^ 1'b0 ;
  assign n19352 = ( ~n3409 & n19198 ) | ( ~n3409 & n19351 ) | ( n19198 & n19351 ) ;
  assign n19353 = n5787 ^ n1434 ^ n1231 ;
  assign n19354 = ( n8520 & n15429 ) | ( n8520 & ~n16840 ) | ( n15429 & ~n16840 ) ;
  assign n19357 = ( n1773 & n3828 ) | ( n1773 & n8324 ) | ( n3828 & n8324 ) ;
  assign n19355 = n9352 ^ n4743 ^ 1'b0 ;
  assign n19356 = n827 & ~n19355 ;
  assign n19358 = n19357 ^ n19356 ^ n3927 ;
  assign n19359 = n19358 ^ n9702 ^ n2607 ;
  assign n19360 = n18821 ^ n733 ^ 1'b0 ;
  assign n19361 = n10756 & ~n19360 ;
  assign n19362 = n9677 ^ n6546 ^ n4332 ;
  assign n19363 = ( ~n3319 & n12570 ) | ( ~n3319 & n19362 ) | ( n12570 & n19362 ) ;
  assign n19364 = n19363 ^ n14177 ^ n713 ;
  assign n19365 = n5075 ^ n4947 ^ n3670 ;
  assign n19366 = ~n11676 & n19365 ;
  assign n19367 = n19366 ^ n17803 ^ n4105 ;
  assign n19368 = n3758 ^ n1027 ^ 1'b0 ;
  assign n19369 = ~n4851 & n19368 ;
  assign n19370 = n3556 & n19369 ;
  assign n19371 = n19370 ^ n11051 ^ n6034 ;
  assign n19372 = ( n4014 & ~n15710 ) | ( n4014 & n19371 ) | ( ~n15710 & n19371 ) ;
  assign n19373 = n762 & ~n2486 ;
  assign n19374 = n19373 ^ n8109 ^ 1'b0 ;
  assign n19375 = ( ~n8241 & n12842 ) | ( ~n8241 & n19374 ) | ( n12842 & n19374 ) ;
  assign n19376 = ( n4132 & n10094 ) | ( n4132 & n19375 ) | ( n10094 & n19375 ) ;
  assign n19377 = ~n10959 & n19376 ;
  assign n19378 = n19377 ^ n17405 ^ 1'b0 ;
  assign n19379 = ( x6 & n5236 ) | ( x6 & ~n19378 ) | ( n5236 & ~n19378 ) ;
  assign n19380 = ~n8937 & n14101 ;
  assign n19381 = n19380 ^ n18203 ^ 1'b0 ;
  assign n19382 = ( n1400 & n6792 ) | ( n1400 & n7880 ) | ( n6792 & n7880 ) ;
  assign n19383 = n17287 | n19382 ;
  assign n19387 = ( n1460 & n5319 ) | ( n1460 & ~n5721 ) | ( n5319 & ~n5721 ) ;
  assign n19384 = n13579 & n18992 ;
  assign n19385 = n4159 & n19384 ;
  assign n19386 = n19385 ^ n14329 ^ n3350 ;
  assign n19388 = n19387 ^ n19386 ^ 1'b0 ;
  assign n19389 = n19388 ^ n18455 ^ n11129 ;
  assign n19390 = n496 | n11456 ;
  assign n19391 = ( ~n4392 & n9987 ) | ( ~n4392 & n12221 ) | ( n9987 & n12221 ) ;
  assign n19392 = n19391 ^ n10992 ^ 1'b0 ;
  assign n19393 = ~n6790 & n19392 ;
  assign n19394 = n4061 ^ n1940 ^ 1'b0 ;
  assign n19395 = ( ~n8996 & n12118 ) | ( ~n8996 & n19394 ) | ( n12118 & n19394 ) ;
  assign n19396 = n12213 & ~n19395 ;
  assign n19397 = n5381 ^ n3600 ^ n2847 ;
  assign n19398 = n19397 ^ n5930 ^ 1'b0 ;
  assign n19402 = n18489 ^ n7017 ^ n2585 ;
  assign n19399 = n8630 ^ n7281 ^ n2848 ;
  assign n19400 = ~n1390 & n5469 ;
  assign n19401 = n19399 & n19400 ;
  assign n19403 = n19402 ^ n19401 ^ n15772 ;
  assign n19404 = ( n5719 & n10890 ) | ( n5719 & ~n11334 ) | ( n10890 & ~n11334 ) ;
  assign n19405 = n7725 & n19404 ;
  assign n19406 = ~n647 & n19405 ;
  assign n19407 = n4078 ^ n3237 ^ 1'b0 ;
  assign n19408 = n8649 & n19407 ;
  assign n19409 = ~n1223 & n6805 ;
  assign n19410 = ~n19408 & n19409 ;
  assign n19411 = ( n1914 & ~n2774 ) | ( n1914 & n5797 ) | ( ~n2774 & n5797 ) ;
  assign n19412 = ~n1075 & n19411 ;
  assign n19413 = ~n6369 & n19412 ;
  assign n19414 = ( ~n10829 & n13002 ) | ( ~n10829 & n17834 ) | ( n13002 & n17834 ) ;
  assign n19415 = n16336 ^ n13732 ^ n8584 ;
  assign n19416 = n19415 ^ n18068 ^ n15893 ;
  assign n19417 = ( n377 & n19414 ) | ( n377 & ~n19416 ) | ( n19414 & ~n19416 ) ;
  assign n19420 = ( n6858 & n10298 ) | ( n6858 & ~n12713 ) | ( n10298 & ~n12713 ) ;
  assign n19418 = ( n1921 & ~n3543 ) | ( n1921 & n7594 ) | ( ~n3543 & n7594 ) ;
  assign n19419 = n19418 ^ n15640 ^ n5126 ;
  assign n19421 = n19420 ^ n19419 ^ n17990 ;
  assign n19422 = ( ~n2760 & n5731 ) | ( ~n2760 & n19421 ) | ( n5731 & n19421 ) ;
  assign n19423 = n19422 ^ n10978 ^ n8421 ;
  assign n19424 = ( n4814 & ~n9386 ) | ( n4814 & n15390 ) | ( ~n9386 & n15390 ) ;
  assign n19425 = n12209 & n19424 ;
  assign n19426 = n19425 ^ n3799 ^ 1'b0 ;
  assign n19427 = n19426 ^ n8653 ^ n7453 ;
  assign n19428 = n9322 ^ n5972 ^ n4240 ;
  assign n19429 = n5005 | n18222 ;
  assign n19430 = n13053 & ~n13096 ;
  assign n19431 = ~n1378 & n19430 ;
  assign n19432 = ~n4055 & n10116 ;
  assign n19433 = n13780 & n19432 ;
  assign n19434 = ( n5558 & n5998 ) | ( n5558 & ~n9559 ) | ( n5998 & ~n9559 ) ;
  assign n19435 = ~n1234 & n19434 ;
  assign n19436 = n19435 ^ n14677 ^ 1'b0 ;
  assign n19437 = n19436 ^ n10940 ^ n3544 ;
  assign n19438 = ( n11536 & n19433 ) | ( n11536 & ~n19437 ) | ( n19433 & ~n19437 ) ;
  assign n19439 = n3156 & ~n6564 ;
  assign n19440 = ( n255 & ~n1613 ) | ( n255 & n17209 ) | ( ~n1613 & n17209 ) ;
  assign n19441 = n2562 & n10176 ;
  assign n19442 = n19441 ^ n4750 ^ 1'b0 ;
  assign n19443 = ( n19439 & ~n19440 ) | ( n19439 & n19442 ) | ( ~n19440 & n19442 ) ;
  assign n19444 = ( n1123 & ~n3317 ) | ( n1123 & n16587 ) | ( ~n3317 & n16587 ) ;
  assign n19445 = n19444 ^ n19023 ^ n13385 ;
  assign n19446 = n6661 ^ n4850 ^ n3757 ;
  assign n19448 = n4271 ^ n1120 ^ 1'b0 ;
  assign n19447 = ( n8302 & ~n9691 ) | ( n8302 & n11909 ) | ( ~n9691 & n11909 ) ;
  assign n19449 = n19448 ^ n19447 ^ n10503 ;
  assign n19450 = ( n1363 & n6004 ) | ( n1363 & ~n19449 ) | ( n6004 & ~n19449 ) ;
  assign n19451 = n16921 ^ n6770 ^ 1'b0 ;
  assign n19452 = ~n2022 & n4437 ;
  assign n19453 = ~n6325 & n19452 ;
  assign n19454 = n11342 & ~n19453 ;
  assign n19455 = n19454 ^ n15375 ^ 1'b0 ;
  assign n19457 = n9497 ^ n7853 ^ n5527 ;
  assign n19456 = ~n430 & n3875 ;
  assign n19458 = n19457 ^ n19456 ^ 1'b0 ;
  assign n19459 = ( n820 & n17338 ) | ( n820 & ~n19127 ) | ( n17338 & ~n19127 ) ;
  assign n19460 = n19459 ^ n5438 ^ n1826 ;
  assign n19465 = n18602 ^ n9423 ^ 1'b0 ;
  assign n19464 = n11446 ^ n9488 ^ n2884 ;
  assign n19462 = n7442 ^ n7426 ^ 1'b0 ;
  assign n19461 = ( n7218 & n8449 ) | ( n7218 & n8720 ) | ( n8449 & n8720 ) ;
  assign n19463 = n19462 ^ n19461 ^ n18922 ;
  assign n19466 = n19465 ^ n19464 ^ n19463 ;
  assign n19467 = n7685 & ~n10598 ;
  assign n19468 = n15607 & n19467 ;
  assign n19469 = n19468 ^ n19171 ^ n13076 ;
  assign n19470 = n14860 ^ n9979 ^ n7582 ;
  assign n19472 = n1927 | n3089 ;
  assign n19473 = n19472 ^ n809 ^ 1'b0 ;
  assign n19471 = ( n6153 & n8012 ) | ( n6153 & ~n15451 ) | ( n8012 & ~n15451 ) ;
  assign n19474 = n19473 ^ n19471 ^ n14485 ;
  assign n19475 = n693 | n7488 ;
  assign n19476 = n19475 ^ n12185 ^ 1'b0 ;
  assign n19477 = x102 & n19476 ;
  assign n19478 = n9021 ^ n8978 ^ n7805 ;
  assign n19479 = n19478 ^ n5756 ^ 1'b0 ;
  assign n19480 = n19477 & ~n19479 ;
  assign n19482 = ( n2732 & n3117 ) | ( n2732 & ~n8045 ) | ( n3117 & ~n8045 ) ;
  assign n19481 = n7264 | n10280 ;
  assign n19483 = n19482 ^ n19481 ^ 1'b0 ;
  assign n19484 = ~n4197 & n19483 ;
  assign n19485 = ( n2563 & n3544 ) | ( n2563 & n9464 ) | ( n3544 & n9464 ) ;
  assign n19486 = n9851 ^ n1361 ^ 1'b0 ;
  assign n19487 = n16277 ^ n8498 ^ 1'b0 ;
  assign n19488 = n12013 & ~n19487 ;
  assign n19489 = ( n441 & n3744 ) | ( n441 & ~n8045 ) | ( n3744 & ~n8045 ) ;
  assign n19490 = n1476 | n1552 ;
  assign n19491 = ( ~n8786 & n19489 ) | ( ~n8786 & n19490 ) | ( n19489 & n19490 ) ;
  assign n19492 = ( n10383 & ~n12532 ) | ( n10383 & n19491 ) | ( ~n12532 & n19491 ) ;
  assign n19493 = n6519 & ~n19492 ;
  assign n19494 = ~n7512 & n8475 ;
  assign n19495 = n19494 ^ n1877 ^ 1'b0 ;
  assign n19496 = ~n9004 & n19495 ;
  assign n19497 = n19496 ^ n5963 ^ 1'b0 ;
  assign n19498 = n13780 ^ n5586 ^ n2302 ;
  assign n19499 = n13811 ^ n2315 ^ n1606 ;
  assign n19500 = n19499 ^ n1336 ^ 1'b0 ;
  assign n19501 = n4690 ^ n1327 ^ 1'b0 ;
  assign n19502 = ( n9890 & n19348 ) | ( n9890 & n19501 ) | ( n19348 & n19501 ) ;
  assign n19503 = ( n1516 & n12635 ) | ( n1516 & n19502 ) | ( n12635 & n19502 ) ;
  assign n19504 = n19503 ^ n15978 ^ n13942 ;
  assign n19505 = n9647 & ~n19504 ;
  assign n19506 = ( n761 & ~n11442 ) | ( n761 & n17923 ) | ( ~n11442 & n17923 ) ;
  assign n19507 = n14035 ^ n5436 ^ 1'b0 ;
  assign n19508 = n19507 ^ n15241 ^ 1'b0 ;
  assign n19509 = n12010 ^ n2016 ^ n1301 ;
  assign n19510 = ( n2551 & n9856 ) | ( n2551 & n15606 ) | ( n9856 & n15606 ) ;
  assign n19511 = n8208 ^ n7843 ^ 1'b0 ;
  assign n19512 = n11829 & n19511 ;
  assign n19513 = n1731 | n3794 ;
  assign n19514 = n6084 | n19513 ;
  assign n19515 = n14734 ^ n3787 ^ n1474 ;
  assign n19516 = ( n8744 & n19514 ) | ( n8744 & ~n19515 ) | ( n19514 & ~n19515 ) ;
  assign n19517 = n11648 | n19516 ;
  assign n19518 = n19512 | n19517 ;
  assign n19519 = n9959 | n13365 ;
  assign n19520 = n19519 ^ n3434 ^ 1'b0 ;
  assign n19521 = ( n4961 & ~n10015 ) | ( n4961 & n15216 ) | ( ~n10015 & n15216 ) ;
  assign n19522 = n5710 ^ n966 ^ x7 ;
  assign n19523 = n19522 ^ n10537 ^ n10257 ;
  assign n19524 = ( ~n11508 & n16114 ) | ( ~n11508 & n19523 ) | ( n16114 & n19523 ) ;
  assign n19525 = n10931 ^ n1899 ^ 1'b0 ;
  assign n19526 = ( n16221 & ~n19524 ) | ( n16221 & n19525 ) | ( ~n19524 & n19525 ) ;
  assign n19527 = n1125 & ~n1864 ;
  assign n19528 = n5955 & n13074 ;
  assign n19529 = ( n1227 & n11506 ) | ( n1227 & n16126 ) | ( n11506 & n16126 ) ;
  assign n19530 = n1227 & ~n5531 ;
  assign n19531 = ~n19529 & n19530 ;
  assign n19532 = ( x60 & ~n988 ) | ( x60 & n1326 ) | ( ~n988 & n1326 ) ;
  assign n19533 = n12829 ^ n10872 ^ n3465 ;
  assign n19534 = n19533 ^ n7487 ^ 1'b0 ;
  assign n19535 = n15799 & ~n19534 ;
  assign n19536 = n19535 ^ n11179 ^ 1'b0 ;
  assign n19537 = ~n4477 & n19536 ;
  assign n19538 = n19532 & n19537 ;
  assign n19539 = ~n4976 & n7265 ;
  assign n19540 = n4000 & n19539 ;
  assign n19541 = n19540 ^ n4114 ^ n1122 ;
  assign n19542 = n18368 ^ n10614 ^ 1'b0 ;
  assign n19543 = n19541 & ~n19542 ;
  assign n19544 = n13753 ^ x82 ^ 1'b0 ;
  assign n19545 = n6756 & ~n19544 ;
  assign n19546 = n19545 ^ n393 ^ 1'b0 ;
  assign n19547 = n5140 ^ n3957 ^ 1'b0 ;
  assign n19548 = ~n9904 & n19547 ;
  assign n19549 = n5624 & n19548 ;
  assign n19550 = n11091 ^ n9617 ^ 1'b0 ;
  assign n19551 = n19549 | n19550 ;
  assign n19552 = ( ~n8081 & n19546 ) | ( ~n8081 & n19551 ) | ( n19546 & n19551 ) ;
  assign n19553 = ( n2896 & n9430 ) | ( n2896 & n9706 ) | ( n9430 & n9706 ) ;
  assign n19555 = ( n1854 & n9664 ) | ( n1854 & n12097 ) | ( n9664 & n12097 ) ;
  assign n19554 = ( n4675 & ~n5763 ) | ( n4675 & n9526 ) | ( ~n5763 & n9526 ) ;
  assign n19556 = n19555 ^ n19554 ^ n4913 ;
  assign n19557 = n15060 ^ n2357 ^ 1'b0 ;
  assign n19558 = ( ~n8915 & n18586 ) | ( ~n8915 & n19557 ) | ( n18586 & n19557 ) ;
  assign n19561 = n7337 ^ n1982 ^ n1273 ;
  assign n19559 = ( n5997 & n13423 ) | ( n5997 & ~n16532 ) | ( n13423 & ~n16532 ) ;
  assign n19560 = ( n11527 & n16125 ) | ( n11527 & ~n19559 ) | ( n16125 & ~n19559 ) ;
  assign n19562 = n19561 ^ n19560 ^ n2041 ;
  assign n19563 = n16004 ^ n13869 ^ n9850 ;
  assign n19564 = n4974 ^ n4788 ^ n3286 ;
  assign n19565 = n19564 ^ n1917 ^ 1'b0 ;
  assign n19566 = n15990 ^ n13125 ^ 1'b0 ;
  assign n19567 = n3211 & ~n8168 ;
  assign n19568 = ~n2713 & n3217 ;
  assign n19569 = n19568 ^ n14726 ^ 1'b0 ;
  assign n19570 = n19569 ^ n6666 ^ n2870 ;
  assign n19571 = ( n17482 & n19006 ) | ( n17482 & ~n19570 ) | ( n19006 & ~n19570 ) ;
  assign n19572 = n12798 ^ n6968 ^ 1'b0 ;
  assign n19579 = n7948 & n8545 ;
  assign n19580 = n13097 & n19579 ;
  assign n19573 = ~n2246 & n9651 ;
  assign n19574 = n19573 ^ n13325 ^ 1'b0 ;
  assign n19575 = ( n9231 & ~n16188 ) | ( n9231 & n16667 ) | ( ~n16188 & n16667 ) ;
  assign n19576 = ( n352 & n2316 ) | ( n352 & n12124 ) | ( n2316 & n12124 ) ;
  assign n19577 = ( ~n19094 & n19575 ) | ( ~n19094 & n19576 ) | ( n19575 & n19576 ) ;
  assign n19578 = ( n10968 & n19574 ) | ( n10968 & ~n19577 ) | ( n19574 & ~n19577 ) ;
  assign n19581 = n19580 ^ n19578 ^ n6881 ;
  assign n19582 = n14653 ^ n10941 ^ n5723 ;
  assign n19585 = n7125 ^ n3384 ^ 1'b0 ;
  assign n19583 = n13641 ^ n1216 ^ 1'b0 ;
  assign n19584 = n12928 | n19583 ;
  assign n19586 = n19585 ^ n19584 ^ n10214 ;
  assign n19587 = n10324 & n13722 ;
  assign n19588 = ( n3033 & n15554 ) | ( n3033 & n19387 ) | ( n15554 & n19387 ) ;
  assign n19589 = ~n1226 & n1679 ;
  assign n19590 = n19589 ^ n7427 ^ 1'b0 ;
  assign n19591 = n8026 ^ n719 ^ 1'b0 ;
  assign n19592 = n9404 & ~n19591 ;
  assign n19593 = n6802 & n14770 ;
  assign n19594 = ~n7744 & n19593 ;
  assign n19595 = ( n8057 & n11903 ) | ( n8057 & n16808 ) | ( n11903 & n16808 ) ;
  assign n19596 = n19595 ^ n8966 ^ 1'b0 ;
  assign n19597 = n3392 ^ n2464 ^ n292 ;
  assign n19598 = n4093 & ~n10906 ;
  assign n19599 = n19598 ^ n1261 ^ 1'b0 ;
  assign n19600 = n19597 & n19599 ;
  assign n19601 = ~n15110 & n19600 ;
  assign n19602 = n19601 ^ n15271 ^ n597 ;
  assign n19603 = ~n2524 & n15662 ;
  assign n19604 = ( n3327 & n11725 ) | ( n3327 & ~n13763 ) | ( n11725 & ~n13763 ) ;
  assign n19605 = ( n2063 & n13473 ) | ( n2063 & n18953 ) | ( n13473 & n18953 ) ;
  assign n19608 = ~n8638 & n18193 ;
  assign n19606 = ( n6032 & n9146 ) | ( n6032 & n11590 ) | ( n9146 & n11590 ) ;
  assign n19607 = ~n10375 & n19606 ;
  assign n19609 = n19608 ^ n19607 ^ 1'b0 ;
  assign n19610 = n1783 ^ n1619 ^ 1'b0 ;
  assign n19611 = n5657 & ~n19610 ;
  assign n19612 = n8187 ^ n3108 ^ 1'b0 ;
  assign n19613 = n9977 & ~n19612 ;
  assign n19614 = n19613 ^ n4177 ^ 1'b0 ;
  assign n19615 = n13960 ^ n11888 ^ 1'b0 ;
  assign n19616 = n1595 | n19615 ;
  assign n19617 = n11019 ^ n6543 ^ 1'b0 ;
  assign n19618 = n12172 ^ n7180 ^ n266 ;
  assign n19619 = n19618 ^ n5717 ^ 1'b0 ;
  assign n19620 = n9190 & n19619 ;
  assign n19621 = n19620 ^ n5050 ^ n1431 ;
  assign n19622 = n19621 ^ n18852 ^ n5968 ;
  assign n19623 = ( ~n19616 & n19617 ) | ( ~n19616 & n19622 ) | ( n19617 & n19622 ) ;
  assign n19624 = n3526 ^ n564 ^ 1'b0 ;
  assign n19625 = n14695 & n19624 ;
  assign n19626 = n3532 | n6606 ;
  assign n19627 = n8565 & ~n19626 ;
  assign n19628 = ( n4984 & n10193 ) | ( n4984 & ~n19627 ) | ( n10193 & ~n19627 ) ;
  assign n19629 = ( n10010 & n16138 ) | ( n10010 & ~n19628 ) | ( n16138 & ~n19628 ) ;
  assign n19630 = n3432 & n8614 ;
  assign n19631 = n5373 & ~n11684 ;
  assign n19632 = n17526 ^ n9651 ^ 1'b0 ;
  assign n19633 = n13897 | n19632 ;
  assign n19634 = n6644 & n19633 ;
  assign n19635 = n14186 & ~n17466 ;
  assign n19636 = n19635 ^ n6485 ^ 1'b0 ;
  assign n19637 = ( n4563 & n6885 ) | ( n4563 & n14772 ) | ( n6885 & n14772 ) ;
  assign n19638 = n19637 ^ n8625 ^ n3935 ;
  assign n19639 = n19638 ^ n4029 ^ 1'b0 ;
  assign n19648 = n5706 ^ n5344 ^ 1'b0 ;
  assign n19640 = ( n4646 & n5233 ) | ( n4646 & n6860 ) | ( n5233 & n6860 ) ;
  assign n19641 = n19640 ^ n8530 ^ n3919 ;
  assign n19642 = n15532 ^ n3052 ^ n151 ;
  assign n19643 = n19642 ^ n5797 ^ 1'b0 ;
  assign n19644 = n1522 & n19643 ;
  assign n19645 = n19644 ^ n10242 ^ 1'b0 ;
  assign n19646 = n19645 ^ n4585 ^ 1'b0 ;
  assign n19647 = ( n17258 & n19641 ) | ( n17258 & n19646 ) | ( n19641 & n19646 ) ;
  assign n19649 = n19648 ^ n19647 ^ n2884 ;
  assign n19650 = n19649 ^ n14226 ^ 1'b0 ;
  assign n19651 = n8339 ^ n1534 ^ 1'b0 ;
  assign n19652 = n5238 ^ n1060 ^ 1'b0 ;
  assign n19653 = n5980 & n19652 ;
  assign n19654 = n19653 ^ n5312 ^ n264 ;
  assign n19655 = n5379 ^ n3861 ^ 1'b0 ;
  assign n19656 = n8625 & ~n19655 ;
  assign n19657 = n19249 | n19656 ;
  assign n19658 = n6820 ^ n3551 ^ 1'b0 ;
  assign n19659 = ~n3317 & n19658 ;
  assign n19660 = n19659 ^ n13686 ^ 1'b0 ;
  assign n19661 = n16290 ^ n4924 ^ 1'b0 ;
  assign n19662 = n18660 ^ n13962 ^ n177 ;
  assign n19663 = n6551 | n16211 ;
  assign n19664 = n5169 | n6839 ;
  assign n19665 = n19664 ^ n14736 ^ 1'b0 ;
  assign n19667 = n1987 | n17922 ;
  assign n19668 = n19667 ^ n9209 ^ 1'b0 ;
  assign n19666 = n5332 | n11735 ;
  assign n19669 = n19668 ^ n19666 ^ 1'b0 ;
  assign n19670 = n5639 ^ n2014 ^ 1'b0 ;
  assign n19671 = ~n5624 & n19670 ;
  assign n19672 = n18953 ^ n2760 ^ n1805 ;
  assign n19673 = n19672 ^ n15327 ^ n8025 ;
  assign n19674 = n2676 & ~n19673 ;
  assign n19675 = ( n5782 & n19671 ) | ( n5782 & n19674 ) | ( n19671 & n19674 ) ;
  assign n19676 = ( n15937 & n17529 ) | ( n15937 & ~n17729 ) | ( n17529 & ~n17729 ) ;
  assign n19677 = n19374 ^ n9829 ^ n4630 ;
  assign n19678 = ~n1495 & n1509 ;
  assign n19679 = n19678 ^ n19284 ^ 1'b0 ;
  assign n19680 = n12980 ^ n3615 ^ 1'b0 ;
  assign n19681 = ~n5815 & n19680 ;
  assign n19682 = n5218 & ~n13163 ;
  assign n19683 = ~n19681 & n19682 ;
  assign n19684 = n5423 | n19683 ;
  assign n19685 = n19684 ^ n8619 ^ 1'b0 ;
  assign n19686 = n657 | n12707 ;
  assign n19687 = n19686 ^ n13035 ^ n2216 ;
  assign n19688 = ( n1060 & ~n10154 ) | ( n1060 & n19687 ) | ( ~n10154 & n19687 ) ;
  assign n19689 = ( n9993 & n14115 ) | ( n9993 & n16327 ) | ( n14115 & n16327 ) ;
  assign n19690 = n18505 ^ n4579 ^ 1'b0 ;
  assign n19691 = ( ~n2452 & n6901 ) | ( ~n2452 & n19690 ) | ( n6901 & n19690 ) ;
  assign n19698 = ( n5950 & n7014 ) | ( n5950 & ~n13686 ) | ( n7014 & ~n13686 ) ;
  assign n19699 = n19698 ^ n1553 ^ 1'b0 ;
  assign n19700 = ~n14778 & n19699 ;
  assign n19692 = ( n602 & ~n6995 ) | ( n602 & n15170 ) | ( ~n6995 & n15170 ) ;
  assign n19693 = n19692 ^ n14233 ^ n9584 ;
  assign n19694 = ( n378 & n1644 ) | ( n378 & ~n19693 ) | ( n1644 & ~n19693 ) ;
  assign n19695 = ( n1994 & n7252 ) | ( n1994 & ~n8029 ) | ( n7252 & ~n8029 ) ;
  assign n19696 = n9564 | n19695 ;
  assign n19697 = n19694 & ~n19696 ;
  assign n19701 = n19700 ^ n19697 ^ n12312 ;
  assign n19702 = ~n4223 & n11805 ;
  assign n19703 = n10766 | n19702 ;
  assign n19704 = n6610 ^ n6411 ^ n238 ;
  assign n19705 = ~n7511 & n10641 ;
  assign n19706 = n15859 | n19705 ;
  assign n19707 = n19704 | n19706 ;
  assign n19708 = n18130 ^ n17045 ^ n12906 ;
  assign n19709 = n19708 ^ n6198 ^ 1'b0 ;
  assign n19710 = n6416 ^ n1818 ^ 1'b0 ;
  assign n19711 = n13684 & n19710 ;
  assign n19712 = ( n2653 & ~n13894 ) | ( n2653 & n18776 ) | ( ~n13894 & n18776 ) ;
  assign n19713 = n17738 ^ n4610 ^ n4024 ;
  assign n19714 = ( n11024 & ~n17088 ) | ( n11024 & n19713 ) | ( ~n17088 & n19713 ) ;
  assign n19715 = ( n962 & ~n19076 ) | ( n962 & n19714 ) | ( ~n19076 & n19714 ) ;
  assign n19716 = ( n19263 & n19712 ) | ( n19263 & ~n19715 ) | ( n19712 & ~n19715 ) ;
  assign n19717 = ( n3900 & ~n11671 ) | ( n3900 & n18415 ) | ( ~n11671 & n18415 ) ;
  assign n19718 = n350 & ~n930 ;
  assign n19719 = ~n8981 & n19718 ;
  assign n19720 = ( n12593 & n14215 ) | ( n12593 & n19719 ) | ( n14215 & n19719 ) ;
  assign n19721 = n19720 ^ n4538 ^ n4478 ;
  assign n19722 = n4503 ^ n3596 ^ 1'b0 ;
  assign n19723 = ( ~n11398 & n16260 ) | ( ~n11398 & n19722 ) | ( n16260 & n19722 ) ;
  assign n19724 = ( n3739 & n11388 ) | ( n3739 & n11474 ) | ( n11388 & n11474 ) ;
  assign n19725 = n15690 ^ n8166 ^ n165 ;
  assign n19726 = ~n3469 & n19725 ;
  assign n19727 = n19724 & n19726 ;
  assign n19728 = ( n1295 & n14848 ) | ( n1295 & n15657 ) | ( n14848 & n15657 ) ;
  assign n19729 = n19728 ^ n15908 ^ n11232 ;
  assign n19730 = n17946 ^ n17796 ^ n130 ;
  assign n19731 = n19730 ^ n1078 ^ 1'b0 ;
  assign n19732 = n10830 ^ n4977 ^ n4915 ;
  assign n19733 = n12889 & n19732 ;
  assign n19734 = n11839 & n19733 ;
  assign n19735 = n12455 ^ n10083 ^ 1'b0 ;
  assign n19736 = n1076 | n19735 ;
  assign n19737 = n7901 | n19736 ;
  assign n19738 = n19737 ^ n6288 ^ 1'b0 ;
  assign n19739 = n17283 ^ n433 ^ 1'b0 ;
  assign n19740 = n3166 & n19739 ;
  assign n19741 = n16510 ^ n7098 ^ 1'b0 ;
  assign n19742 = n17098 ^ n1745 ^ x110 ;
  assign n19743 = ( n5694 & n14505 ) | ( n5694 & n19742 ) | ( n14505 & n19742 ) ;
  assign n19744 = n19743 ^ n19257 ^ n4633 ;
  assign n19745 = n2818 & ~n11272 ;
  assign n19746 = n19745 ^ n3324 ^ 1'b0 ;
  assign n19747 = n19746 ^ n15476 ^ n14226 ;
  assign n19749 = n10257 ^ n3179 ^ n3073 ;
  assign n19748 = n8292 & n9053 ;
  assign n19750 = n19749 ^ n19748 ^ n7935 ;
  assign n19751 = n10996 ^ n8295 ^ n2314 ;
  assign n19752 = n19751 ^ n4440 ^ 1'b0 ;
  assign n19753 = n11026 ^ n542 ^ 1'b0 ;
  assign n19754 = n19752 | n19753 ;
  assign n19755 = n15964 ^ n1352 ^ 1'b0 ;
  assign n19756 = n18187 & ~n19755 ;
  assign n19766 = ( n738 & n5292 ) | ( n738 & ~n9440 ) | ( n5292 & ~n9440 ) ;
  assign n19767 = n10110 ^ n7289 ^ n1982 ;
  assign n19768 = n19767 ^ n8084 ^ n6233 ;
  assign n19769 = n19766 | n19768 ;
  assign n19770 = n6180 & ~n19769 ;
  assign n19757 = n17106 & n19046 ;
  assign n19758 = ~n10788 & n19757 ;
  assign n19759 = n5345 & ~n18255 ;
  assign n19760 = n19759 ^ n3250 ^ 1'b0 ;
  assign n19762 = n5150 ^ n3495 ^ 1'b0 ;
  assign n19761 = n2631 ^ n1638 ^ n902 ;
  assign n19763 = n19762 ^ n19761 ^ n15324 ;
  assign n19764 = n19763 ^ n17867 ^ n14899 ;
  assign n19765 = ( n19758 & ~n19760 ) | ( n19758 & n19764 ) | ( ~n19760 & n19764 ) ;
  assign n19771 = n19770 ^ n19765 ^ n1913 ;
  assign n19772 = n15312 & ~n16123 ;
  assign n19773 = ( n2710 & n6518 ) | ( n2710 & ~n10954 ) | ( n6518 & ~n10954 ) ;
  assign n19774 = n12813 ^ n694 ^ 1'b0 ;
  assign n19775 = n19773 & n19774 ;
  assign n19776 = n12738 | n13852 ;
  assign n19777 = n15221 ^ n6016 ^ 1'b0 ;
  assign n19778 = n19776 & n19777 ;
  assign n19779 = x80 & n5696 ;
  assign n19780 = n19779 ^ n163 ^ 1'b0 ;
  assign n19781 = n16549 ^ n8268 ^ n5324 ;
  assign n19782 = n17069 ^ n4400 ^ n3893 ;
  assign n19783 = ( n12251 & n15830 ) | ( n12251 & n19782 ) | ( n15830 & n19782 ) ;
  assign n19784 = n15167 ^ n9324 ^ 1'b0 ;
  assign n19785 = ( n2085 & n2295 ) | ( n2085 & n3831 ) | ( n2295 & n3831 ) ;
  assign n19786 = n5003 ^ n4567 ^ 1'b0 ;
  assign n19787 = x82 & ~n19786 ;
  assign n19788 = n5469 & n19787 ;
  assign n19789 = ( ~n12256 & n19785 ) | ( ~n12256 & n19788 ) | ( n19785 & n19788 ) ;
  assign n19790 = n19789 ^ n9694 ^ n2597 ;
  assign n19791 = n711 & n1394 ;
  assign n19792 = n17695 & n19791 ;
  assign n19793 = n4259 ^ n1291 ^ n357 ;
  assign n19794 = n19793 ^ n12189 ^ 1'b0 ;
  assign n19795 = n4808 & ~n19794 ;
  assign n19796 = ~n2812 & n9109 ;
  assign n19797 = ~n19795 & n19796 ;
  assign n19798 = ( ~n5849 & n14979 ) | ( ~n5849 & n19797 ) | ( n14979 & n19797 ) ;
  assign n19799 = n19798 ^ n17656 ^ n3557 ;
  assign n19800 = ( n4871 & n11770 ) | ( n4871 & n13404 ) | ( n11770 & n13404 ) ;
  assign n19801 = n10580 ^ n8996 ^ 1'b0 ;
  assign n19802 = n4945 & n19801 ;
  assign n19803 = n19802 ^ n17323 ^ n8330 ;
  assign n19804 = n7294 ^ n7215 ^ 1'b0 ;
  assign n19805 = n1068 & ~n6351 ;
  assign n19806 = ( n196 & n4406 ) | ( n196 & n19805 ) | ( n4406 & n19805 ) ;
  assign n19807 = n5480 & n7164 ;
  assign n19809 = n9011 ^ n7771 ^ n6553 ;
  assign n19808 = n4818 | n6216 ;
  assign n19810 = n19809 ^ n19808 ^ 1'b0 ;
  assign n19811 = n9595 | n19810 ;
  assign n19812 = n5545 ^ n4225 ^ 1'b0 ;
  assign n19813 = n13517 & n19812 ;
  assign n19814 = n14231 ^ n14200 ^ 1'b0 ;
  assign n19816 = ( ~n1842 & n6704 ) | ( ~n1842 & n7759 ) | ( n6704 & n7759 ) ;
  assign n19815 = n6000 ^ n4299 ^ n1784 ;
  assign n19817 = n19816 ^ n19815 ^ n9538 ;
  assign n19818 = ( n592 & n5126 ) | ( n592 & n7399 ) | ( n5126 & n7399 ) ;
  assign n19819 = n19818 ^ n15509 ^ 1'b0 ;
  assign n19820 = n407 & n5678 ;
  assign n19821 = n11654 ^ n1301 ^ 1'b0 ;
  assign n19822 = n16012 | n19821 ;
  assign n19823 = ( n5218 & n11330 ) | ( n5218 & ~n13882 ) | ( n11330 & ~n13882 ) ;
  assign n19824 = ( n3139 & ~n15794 ) | ( n3139 & n15831 ) | ( ~n15794 & n15831 ) ;
  assign n19825 = n19824 ^ n12648 ^ n12027 ;
  assign n19826 = n13991 ^ n12545 ^ 1'b0 ;
  assign n19827 = n662 | n15250 ;
  assign n19828 = n5896 ^ n4684 ^ n2689 ;
  assign n19829 = n19828 ^ n4314 ^ 1'b0 ;
  assign n19830 = n19829 ^ n13028 ^ n6165 ;
  assign n19831 = n6363 | n19830 ;
  assign n19832 = ( ~n5344 & n7890 ) | ( ~n5344 & n16676 ) | ( n7890 & n16676 ) ;
  assign n19833 = n19832 ^ n11236 ^ n4608 ;
  assign n19834 = n8029 ^ n3767 ^ n2469 ;
  assign n19835 = n14401 ^ n5178 ^ x61 ;
  assign n19836 = ( n926 & n19834 ) | ( n926 & ~n19835 ) | ( n19834 & ~n19835 ) ;
  assign n19837 = ( n8444 & ~n12218 ) | ( n8444 & n14646 ) | ( ~n12218 & n14646 ) ;
  assign n19838 = n19837 ^ n14240 ^ n5576 ;
  assign n19839 = n2075 & n13414 ;
  assign n19840 = n19839 ^ n14998 ^ 1'b0 ;
  assign n19841 = n2917 ^ n2710 ^ 1'b0 ;
  assign n19842 = n19841 ^ n17340 ^ n1334 ;
  assign n19843 = ( n19838 & ~n19840 ) | ( n19838 & n19842 ) | ( ~n19840 & n19842 ) ;
  assign n19844 = n14246 | n17059 ;
  assign n19845 = n19844 ^ n16327 ^ 1'b0 ;
  assign n19846 = n1864 | n18278 ;
  assign n19847 = n19845 | n19846 ;
  assign n19848 = n2219 & n2615 ;
  assign n19849 = n5044 & n5771 ;
  assign n19850 = n19849 ^ n17021 ^ 1'b0 ;
  assign n19851 = ( ~n6819 & n8493 ) | ( ~n6819 & n9525 ) | ( n8493 & n9525 ) ;
  assign n19852 = n12654 ^ n5602 ^ 1'b0 ;
  assign n19853 = ( n3022 & n18864 ) | ( n3022 & n19852 ) | ( n18864 & n19852 ) ;
  assign n19854 = n7852 & n12604 ;
  assign n19855 = ( n8891 & n17014 ) | ( n8891 & ~n19854 ) | ( n17014 & ~n19854 ) ;
  assign n19856 = ( n4275 & ~n7205 ) | ( n4275 & n17043 ) | ( ~n7205 & n17043 ) ;
  assign n19857 = ( n1099 & ~n2825 ) | ( n1099 & n7489 ) | ( ~n2825 & n7489 ) ;
  assign n19858 = ~n9052 & n19857 ;
  assign n19859 = n10028 ^ n1972 ^ 1'b0 ;
  assign n19861 = ( n4041 & n4624 ) | ( n4041 & n12348 ) | ( n4624 & n12348 ) ;
  assign n19860 = ~n3477 & n10533 ;
  assign n19862 = n19861 ^ n19860 ^ 1'b0 ;
  assign n19863 = n19862 ^ n18714 ^ n12005 ;
  assign n19864 = n15635 & ~n18668 ;
  assign n19865 = n19864 ^ n6685 ^ 1'b0 ;
  assign n19866 = ~n1211 & n2667 ;
  assign n19867 = n19866 ^ n1573 ^ 1'b0 ;
  assign n19868 = n19867 ^ n10583 ^ n643 ;
  assign n19869 = n19868 ^ n2417 ^ 1'b0 ;
  assign n19870 = ( n3742 & n8152 ) | ( n3742 & ~n19869 ) | ( n8152 & ~n19869 ) ;
  assign n19875 = n1238 | n11819 ;
  assign n19876 = ( n640 & n14995 ) | ( n640 & n19875 ) | ( n14995 & n19875 ) ;
  assign n19871 = n13830 ^ n12356 ^ n2428 ;
  assign n19872 = n19871 ^ n3301 ^ 1'b0 ;
  assign n19873 = ~n3597 & n19872 ;
  assign n19874 = n19873 ^ n1187 ^ 1'b0 ;
  assign n19877 = n19876 ^ n19874 ^ n3026 ;
  assign n19878 = ( n5703 & n11061 ) | ( n5703 & ~n13783 ) | ( n11061 & ~n13783 ) ;
  assign n19882 = n7080 ^ n741 ^ 1'b0 ;
  assign n19883 = n10600 | n19882 ;
  assign n19879 = ~n2519 & n2732 ;
  assign n19880 = n19879 ^ n5777 ^ 1'b0 ;
  assign n19881 = ( n10157 & n12534 ) | ( n10157 & ~n19880 ) | ( n12534 & ~n19880 ) ;
  assign n19884 = n19883 ^ n19881 ^ n3025 ;
  assign n19885 = n13337 ^ n1546 ^ n148 ;
  assign n19886 = ( n19878 & n19884 ) | ( n19878 & ~n19885 ) | ( n19884 & ~n19885 ) ;
  assign n19887 = n7944 ^ n137 ^ 1'b0 ;
  assign n19888 = n442 | n6129 ;
  assign n19889 = n19888 ^ n8715 ^ 1'b0 ;
  assign n19890 = n19889 ^ n14232 ^ 1'b0 ;
  assign n19891 = n1340 & n19890 ;
  assign n19894 = ( n201 & n6544 ) | ( n201 & ~n7603 ) | ( n6544 & ~n7603 ) ;
  assign n19892 = n8781 ^ n196 ^ 1'b0 ;
  assign n19893 = ~n11741 & n19892 ;
  assign n19895 = n19894 ^ n19893 ^ n9585 ;
  assign n19896 = ( n1445 & ~n5713 ) | ( n1445 & n13908 ) | ( ~n5713 & n13908 ) ;
  assign n19897 = ( n5132 & n13037 ) | ( n5132 & ~n19896 ) | ( n13037 & ~n19896 ) ;
  assign n19898 = ( n2891 & n12844 ) | ( n2891 & n19897 ) | ( n12844 & n19897 ) ;
  assign n19899 = ~n1517 & n7809 ;
  assign n19900 = n19899 ^ n13456 ^ 1'b0 ;
  assign n19901 = n15993 ^ n5241 ^ n3827 ;
  assign n19902 = n1758 & ~n11058 ;
  assign n19903 = n19902 ^ n13099 ^ 1'b0 ;
  assign n19904 = n3500 & ~n18297 ;
  assign n19905 = n367 & ~n19904 ;
  assign n19906 = ~n7073 & n19905 ;
  assign n19907 = ( n7421 & n19903 ) | ( n7421 & ~n19906 ) | ( n19903 & ~n19906 ) ;
  assign n19908 = ( ~x57 & n5759 ) | ( ~x57 & n10238 ) | ( n5759 & n10238 ) ;
  assign n19909 = ( n15696 & ~n17745 ) | ( n15696 & n19908 ) | ( ~n17745 & n19908 ) ;
  assign n19910 = n16691 ^ n2575 ^ n386 ;
  assign n19911 = n19910 ^ n1369 ^ 1'b0 ;
  assign n19912 = n5514 & n19911 ;
  assign n19913 = n4746 & ~n10588 ;
  assign n19914 = ~n16696 & n19913 ;
  assign n19915 = ~n16354 & n19914 ;
  assign n19916 = ~n8448 & n19915 ;
  assign n19917 = ( n13803 & ~n17667 ) | ( n13803 & n18693 ) | ( ~n17667 & n18693 ) ;
  assign n19918 = n14198 ^ n4690 ^ n2083 ;
  assign n19919 = ( ~n8214 & n8695 ) | ( ~n8214 & n17059 ) | ( n8695 & n17059 ) ;
  assign n19920 = n14379 ^ n3076 ^ 1'b0 ;
  assign n19921 = n19919 & n19920 ;
  assign n19924 = n7154 ^ n4976 ^ n746 ;
  assign n19922 = n3145 & n3442 ;
  assign n19923 = ~n14190 & n19922 ;
  assign n19925 = n19924 ^ n19923 ^ n4830 ;
  assign n19926 = n12843 ^ n1542 ^ 1'b0 ;
  assign n19927 = ( n4551 & n9237 ) | ( n4551 & n19926 ) | ( n9237 & n19926 ) ;
  assign n19935 = ( ~n308 & n3053 ) | ( ~n308 & n4649 ) | ( n3053 & n4649 ) ;
  assign n19930 = n4066 ^ n428 ^ 1'b0 ;
  assign n19931 = n760 & ~n19930 ;
  assign n19932 = n19931 ^ n5868 ^ 1'b0 ;
  assign n19933 = n17674 & ~n19932 ;
  assign n19928 = n3340 | n17703 ;
  assign n19929 = n19928 ^ n4720 ^ 1'b0 ;
  assign n19934 = n19933 ^ n19929 ^ 1'b0 ;
  assign n19936 = n19935 ^ n19934 ^ 1'b0 ;
  assign n19939 = n4053 ^ n3597 ^ 1'b0 ;
  assign n19938 = ( n603 & n6484 ) | ( n603 & n7749 ) | ( n6484 & n7749 ) ;
  assign n19937 = ~n1067 & n10118 ;
  assign n19940 = n19939 ^ n19938 ^ n19937 ;
  assign n19941 = n329 & ~n6187 ;
  assign n19942 = n19941 ^ n2668 ^ 1'b0 ;
  assign n19943 = n19942 ^ n19427 ^ n8591 ;
  assign n19944 = n4487 ^ n4434 ^ n1739 ;
  assign n19945 = ( n8036 & n17098 ) | ( n8036 & n19944 ) | ( n17098 & n19944 ) ;
  assign n19946 = n19945 ^ n10855 ^ n6183 ;
  assign n19948 = n13899 ^ n5894 ^ n4727 ;
  assign n19949 = ( n4041 & ~n11093 ) | ( n4041 & n19948 ) | ( ~n11093 & n19948 ) ;
  assign n19950 = n1728 & ~n4097 ;
  assign n19951 = n19950 ^ n16419 ^ n13321 ;
  assign n19952 = n19949 & ~n19951 ;
  assign n19953 = ~n17727 & n19952 ;
  assign n19947 = n4313 & ~n12234 ;
  assign n19954 = n19953 ^ n19947 ^ 1'b0 ;
  assign n19955 = n19686 ^ n14425 ^ n10488 ;
  assign n19956 = n19955 ^ n16711 ^ 1'b0 ;
  assign n19957 = n14872 & n19956 ;
  assign n19958 = n8495 ^ n1980 ^ n852 ;
  assign n19959 = n9887 ^ n1113 ^ 1'b0 ;
  assign n19960 = ~n19958 & n19959 ;
  assign n19961 = n5818 ^ n4765 ^ n4667 ;
  assign n19962 = n19081 ^ n14290 ^ n2236 ;
  assign n19963 = ( n8216 & n9068 ) | ( n8216 & ~n9826 ) | ( n9068 & ~n9826 ) ;
  assign n19964 = ~n14209 & n19963 ;
  assign n19965 = ( ~n5056 & n12954 ) | ( ~n5056 & n19964 ) | ( n12954 & n19964 ) ;
  assign n19966 = n15593 ^ n5638 ^ n2118 ;
  assign n19967 = n19966 ^ n11698 ^ n11369 ;
  assign n19968 = ( ~n8433 & n17335 ) | ( ~n8433 & n19967 ) | ( n17335 & n19967 ) ;
  assign n19969 = n16747 ^ n10816 ^ n6644 ;
  assign n19970 = n19969 ^ n9710 ^ n2703 ;
  assign n19971 = ( n491 & ~n8335 ) | ( n491 & n13389 ) | ( ~n8335 & n13389 ) ;
  assign n19972 = ( n4646 & n13818 ) | ( n4646 & n19971 ) | ( n13818 & n19971 ) ;
  assign n19973 = ( ~n4304 & n19970 ) | ( ~n4304 & n19972 ) | ( n19970 & n19972 ) ;
  assign n19974 = n6892 ^ n4804 ^ 1'b0 ;
  assign n19976 = n10440 ^ n8426 ^ n8049 ;
  assign n19975 = n14456 ^ n8527 ^ x107 ;
  assign n19977 = n19976 ^ n19975 ^ n17516 ;
  assign n19979 = n16352 ^ n2376 ^ 1'b0 ;
  assign n19978 = n7460 ^ n2267 ^ 1'b0 ;
  assign n19980 = n19979 ^ n19978 ^ 1'b0 ;
  assign n19981 = n7435 ^ n7165 ^ 1'b0 ;
  assign n19982 = ~n916 & n2336 ;
  assign n19983 = ( n847 & n3657 ) | ( n847 & n3883 ) | ( n3657 & n3883 ) ;
  assign n19984 = n13103 & n19983 ;
  assign n19985 = n19984 ^ n14549 ^ 1'b0 ;
  assign n19986 = n5543 | n19985 ;
  assign n19987 = n4925 ^ n3788 ^ 1'b0 ;
  assign n19988 = n19987 ^ n11413 ^ n3651 ;
  assign n19989 = ( n9172 & n14678 ) | ( n9172 & n19988 ) | ( n14678 & n19988 ) ;
  assign n19993 = ( n12788 & n13333 ) | ( n12788 & n16086 ) | ( n13333 & n16086 ) ;
  assign n19994 = n9733 & ~n19993 ;
  assign n19995 = n19994 ^ n9624 ^ 1'b0 ;
  assign n19990 = n6813 ^ n6462 ^ 1'b0 ;
  assign n19991 = n6396 | n14656 ;
  assign n19992 = n19990 | n19991 ;
  assign n19996 = n19995 ^ n19992 ^ n9567 ;
  assign n19997 = n346 | n1418 ;
  assign n19998 = ( n1416 & n15382 ) | ( n1416 & ~n19997 ) | ( n15382 & ~n19997 ) ;
  assign n19999 = n4651 ^ n2391 ^ n1931 ;
  assign n20000 = n14420 ^ n13439 ^ n2984 ;
  assign n20001 = n18476 ^ n14653 ^ n11349 ;
  assign n20002 = ( n8827 & ~n10492 ) | ( n8827 & n15960 ) | ( ~n10492 & n15960 ) ;
  assign n20003 = ( n2645 & n5535 ) | ( n2645 & n7275 ) | ( n5535 & n7275 ) ;
  assign n20004 = n20003 ^ n2411 ^ n1481 ;
  assign n20005 = ~n8052 & n9327 ;
  assign n20006 = n20005 ^ n4588 ^ 1'b0 ;
  assign n20007 = n20006 ^ n6975 ^ n1441 ;
  assign n20008 = n455 & ~n20007 ;
  assign n20009 = n5527 ^ n4864 ^ 1'b0 ;
  assign n20010 = n10307 | n20009 ;
  assign n20011 = n4617 | n20010 ;
  assign n20012 = n20011 ^ n15525 ^ 1'b0 ;
  assign n20013 = n5336 & ~n11395 ;
  assign n20014 = n15550 & n20013 ;
  assign n20015 = ( ~n4697 & n11548 ) | ( ~n4697 & n13615 ) | ( n11548 & n13615 ) ;
  assign n20016 = n19039 & ~n20015 ;
  assign n20017 = n20014 & n20016 ;
  assign n20018 = ( ~n6024 & n8486 ) | ( ~n6024 & n13365 ) | ( n8486 & n13365 ) ;
  assign n20019 = n965 & ~n2803 ;
  assign n20020 = n17801 ^ n4562 ^ 1'b0 ;
  assign n20024 = n11222 ^ n4467 ^ 1'b0 ;
  assign n20021 = ( n1734 & n5480 ) | ( n1734 & ~n11933 ) | ( n5480 & ~n11933 ) ;
  assign n20022 = n20021 ^ n12374 ^ n11888 ;
  assign n20023 = n3486 | n20022 ;
  assign n20025 = n20024 ^ n20023 ^ 1'b0 ;
  assign n20026 = n7788 | n12798 ;
  assign n20027 = n20026 ^ n14033 ^ n3671 ;
  assign n20028 = n20027 ^ n11902 ^ n403 ;
  assign n20029 = n3901 & ~n14190 ;
  assign n20031 = ~n1852 & n4074 ;
  assign n20032 = n1953 & n20031 ;
  assign n20030 = n5742 ^ n313 ^ 1'b0 ;
  assign n20033 = n20032 ^ n20030 ^ n12024 ;
  assign n20034 = n378 & ~n9408 ;
  assign n20035 = ~n9613 & n20034 ;
  assign n20036 = n12144 & n15435 ;
  assign n20037 = n1376 & n20036 ;
  assign n20038 = ~n16925 & n20012 ;
  assign n20039 = n6703 & n20038 ;
  assign n20040 = n11318 ^ n10825 ^ n1613 ;
  assign n20041 = n20040 ^ n11005 ^ 1'b0 ;
  assign n20042 = n8570 & ~n13545 ;
  assign n20043 = n20042 ^ n9121 ^ 1'b0 ;
  assign n20044 = n3203 ^ n242 ^ 1'b0 ;
  assign n20045 = ~n20043 & n20044 ;
  assign n20046 = x31 & ~n3281 ;
  assign n20047 = n20046 ^ n19357 ^ 1'b0 ;
  assign n20048 = n12867 ^ n4378 ^ n4252 ;
  assign n20049 = n10162 ^ n9555 ^ n4200 ;
  assign n20050 = n11369 ^ n9665 ^ 1'b0 ;
  assign n20051 = ~n6020 & n20050 ;
  assign n20052 = n5121 ^ n4731 ^ n728 ;
  assign n20053 = ~n3069 & n4573 ;
  assign n20054 = n3758 & n20053 ;
  assign n20055 = ( n1258 & n1910 ) | ( n1258 & n14125 ) | ( n1910 & n14125 ) ;
  assign n20056 = n20055 ^ n3175 ^ 1'b0 ;
  assign n20057 = n15896 & n20056 ;
  assign n20058 = ( ~n14261 & n20054 ) | ( ~n14261 & n20057 ) | ( n20054 & n20057 ) ;
  assign n20059 = ( n18952 & ~n20052 ) | ( n18952 & n20058 ) | ( ~n20052 & n20058 ) ;
  assign n20060 = ( n16408 & n20051 ) | ( n16408 & ~n20059 ) | ( n20051 & ~n20059 ) ;
  assign n20061 = n16436 ^ n10270 ^ 1'b0 ;
  assign n20062 = ( n9237 & ~n18153 ) | ( n9237 & n20061 ) | ( ~n18153 & n20061 ) ;
  assign n20063 = ( ~n2092 & n14556 ) | ( ~n2092 & n20062 ) | ( n14556 & n20062 ) ;
  assign n20064 = n15731 ^ n5875 ^ n5041 ;
  assign n20065 = n14660 ^ n11486 ^ 1'b0 ;
  assign n20066 = n7801 & n19088 ;
  assign n20067 = n20066 ^ n3350 ^ 1'b0 ;
  assign n20069 = n15403 ^ n8211 ^ n1597 ;
  assign n20068 = n866 | n14364 ;
  assign n20070 = n20069 ^ n20068 ^ 1'b0 ;
  assign n20071 = ( n11856 & n12534 ) | ( n11856 & ~n13390 ) | ( n12534 & ~n13390 ) ;
  assign n20072 = ( n1882 & n2853 ) | ( n1882 & n5462 ) | ( n2853 & n5462 ) ;
  assign n20073 = ~n14986 & n16808 ;
  assign n20074 = n20073 ^ n15418 ^ 1'b0 ;
  assign n20075 = ( n16321 & n20072 ) | ( n16321 & n20074 ) | ( n20072 & n20074 ) ;
  assign n20076 = ( ~n940 & n2159 ) | ( ~n940 & n4794 ) | ( n2159 & n4794 ) ;
  assign n20077 = n818 & n11222 ;
  assign n20078 = n5004 ^ n1547 ^ 1'b0 ;
  assign n20079 = n20077 | n20078 ;
  assign n20080 = n6055 & ~n20079 ;
  assign n20081 = ( n15360 & n20076 ) | ( n15360 & n20080 ) | ( n20076 & n20080 ) ;
  assign n20082 = n19793 ^ n10626 ^ n4798 ;
  assign n20083 = n20082 ^ n8094 ^ n6106 ;
  assign n20084 = n16927 ^ n16111 ^ n15301 ;
  assign n20086 = ( n9215 & ~n11406 ) | ( n9215 & n16571 ) | ( ~n11406 & n16571 ) ;
  assign n20085 = n271 & ~n8376 ;
  assign n20087 = n20086 ^ n20085 ^ 1'b0 ;
  assign n20088 = n20087 ^ n9865 ^ n5415 ;
  assign n20089 = ( n10322 & n13261 ) | ( n10322 & n14927 ) | ( n13261 & n14927 ) ;
  assign n20090 = n20089 ^ n19690 ^ n4821 ;
  assign n20091 = n7677 ^ n1901 ^ 1'b0 ;
  assign n20092 = n11701 ^ n10892 ^ n2910 ;
  assign n20093 = ( n468 & n828 ) | ( n468 & n2045 ) | ( n828 & n2045 ) ;
  assign n20094 = n12557 & ~n20093 ;
  assign n20095 = ( n20091 & n20092 ) | ( n20091 & ~n20094 ) | ( n20092 & ~n20094 ) ;
  assign n20096 = n3528 & n6403 ;
  assign n20097 = n20096 ^ n11641 ^ 1'b0 ;
  assign n20103 = n7701 ^ n3919 ^ n1869 ;
  assign n20104 = ( ~n7767 & n14192 ) | ( ~n7767 & n20103 ) | ( n14192 & n20103 ) ;
  assign n20099 = ( n801 & n1258 ) | ( n801 & ~n2754 ) | ( n1258 & ~n2754 ) ;
  assign n20100 = n20099 ^ n7094 ^ n1842 ;
  assign n20101 = ( n1474 & n3119 ) | ( n1474 & ~n10878 ) | ( n3119 & ~n10878 ) ;
  assign n20102 = ( n3786 & ~n20100 ) | ( n3786 & n20101 ) | ( ~n20100 & n20101 ) ;
  assign n20105 = n20104 ^ n20102 ^ n1957 ;
  assign n20098 = n5570 & n5669 ;
  assign n20106 = n20105 ^ n20098 ^ 1'b0 ;
  assign n20107 = n7522 | n11027 ;
  assign n20108 = n329 | n20107 ;
  assign n20109 = n386 & ~n16359 ;
  assign n20110 = n1106 & n20109 ;
  assign n20111 = n20110 ^ n423 ^ 1'b0 ;
  assign n20112 = n1635 & ~n20111 ;
  assign n20113 = n4103 ^ n3250 ^ x99 ;
  assign n20114 = ( n2292 & ~n20112 ) | ( n2292 & n20113 ) | ( ~n20112 & n20113 ) ;
  assign n20115 = n20114 ^ n7035 ^ 1'b0 ;
  assign n20116 = n20108 & ~n20115 ;
  assign n20117 = n1273 & n6807 ;
  assign n20118 = n6558 | n20117 ;
  assign n20119 = n19834 ^ n14644 ^ n4589 ;
  assign n20120 = ( ~n1180 & n20118 ) | ( ~n1180 & n20119 ) | ( n20118 & n20119 ) ;
  assign n20121 = ( n6271 & n7836 ) | ( n6271 & ~n20120 ) | ( n7836 & ~n20120 ) ;
  assign n20122 = n5787 | n9030 ;
  assign n20123 = n347 & n10313 ;
  assign n20124 = ~n7601 & n20123 ;
  assign n20125 = n20124 ^ n11172 ^ n2749 ;
  assign n20126 = n20125 ^ n4157 ^ 1'b0 ;
  assign n20127 = n20126 ^ n13456 ^ n9860 ;
  assign n20128 = ( ~n8020 & n18427 ) | ( ~n8020 & n19068 ) | ( n18427 & n19068 ) ;
  assign n20129 = n17102 ^ n5775 ^ 1'b0 ;
  assign n20130 = n9301 | n20129 ;
  assign n20131 = n11889 ^ n11312 ^ n6462 ;
  assign n20132 = n1353 | n8216 ;
  assign n20133 = n12098 ^ n5478 ^ n1959 ;
  assign n20134 = n20133 ^ n18299 ^ 1'b0 ;
  assign n20135 = ( n4244 & n14590 ) | ( n4244 & ~n18702 ) | ( n14590 & ~n18702 ) ;
  assign n20136 = n3786 & n15005 ;
  assign n20137 = n20135 & n20136 ;
  assign n20138 = n17933 ^ n14051 ^ n1839 ;
  assign n20139 = n141 & n6974 ;
  assign n20140 = ( n160 & n5387 ) | ( n160 & ~n10922 ) | ( n5387 & ~n10922 ) ;
  assign n20141 = n10200 ^ n2701 ^ n734 ;
  assign n20142 = n4473 ^ n1543 ^ 1'b0 ;
  assign n20143 = n20141 & ~n20142 ;
  assign n20144 = n20143 ^ n15694 ^ n14967 ;
  assign n20145 = ( n4196 & n15607 ) | ( n4196 & n19951 ) | ( n15607 & n19951 ) ;
  assign n20146 = n2294 ^ n2025 ^ 1'b0 ;
  assign n20147 = n10583 & n20146 ;
  assign n20150 = ( ~n1769 & n8035 ) | ( ~n1769 & n19620 ) | ( n8035 & n19620 ) ;
  assign n20151 = ( n6004 & n13758 ) | ( n6004 & n20150 ) | ( n13758 & n20150 ) ;
  assign n20152 = n20151 ^ n13053 ^ n3816 ;
  assign n20148 = n19310 ^ n11679 ^ n10955 ;
  assign n20149 = n14269 & n20148 ;
  assign n20153 = n20152 ^ n20149 ^ n2075 ;
  assign n20154 = n10973 ^ n1217 ^ n705 ;
  assign n20155 = ( n8958 & ~n13478 ) | ( n8958 & n20154 ) | ( ~n13478 & n20154 ) ;
  assign n20156 = ( n13646 & n18059 ) | ( n13646 & ~n20155 ) | ( n18059 & ~n20155 ) ;
  assign n20157 = ( n5909 & n6409 ) | ( n5909 & n10682 ) | ( n6409 & n10682 ) ;
  assign n20158 = n8335 & n20157 ;
  assign n20159 = ~n12046 & n12074 ;
  assign n20160 = n11960 | n20159 ;
  assign n20161 = ~n15761 & n20160 ;
  assign n20162 = n20054 ^ n13056 ^ n563 ;
  assign n20163 = n4555 & ~n9199 ;
  assign n20164 = n7303 & ~n18224 ;
  assign n20165 = n20164 ^ n14803 ^ 1'b0 ;
  assign n20166 = ( n20162 & n20163 ) | ( n20162 & ~n20165 ) | ( n20163 & ~n20165 ) ;
  assign n20167 = n7169 & n9757 ;
  assign n20168 = n11236 & n20167 ;
  assign n20169 = n20168 ^ n11225 ^ 1'b0 ;
  assign n20170 = ( n8362 & n14932 ) | ( n8362 & n20169 ) | ( n14932 & n20169 ) ;
  assign n20171 = n20170 ^ n11213 ^ n4669 ;
  assign n20174 = ( n2402 & ~n2555 ) | ( n2402 & n7098 ) | ( ~n2555 & n7098 ) ;
  assign n20175 = ~n3464 & n11273 ;
  assign n20176 = ( n13541 & n20174 ) | ( n13541 & ~n20175 ) | ( n20174 & ~n20175 ) ;
  assign n20172 = n16687 ^ n10561 ^ n4006 ;
  assign n20173 = ( ~n4800 & n9245 ) | ( ~n4800 & n20172 ) | ( n9245 & n20172 ) ;
  assign n20177 = n20176 ^ n20173 ^ n6485 ;
  assign n20178 = n213 & n5524 ;
  assign n20179 = n20178 ^ n18328 ^ 1'b0 ;
  assign n20181 = ( n456 & ~n2822 ) | ( n456 & n2962 ) | ( ~n2822 & n2962 ) ;
  assign n20180 = ( n4451 & n14510 ) | ( n4451 & n16136 ) | ( n14510 & n16136 ) ;
  assign n20182 = n20181 ^ n20180 ^ n12935 ;
  assign n20183 = n10383 ^ n1391 ^ 1'b0 ;
  assign n20189 = n3188 | n4117 ;
  assign n20190 = n20189 ^ n5407 ^ 1'b0 ;
  assign n20191 = n20190 ^ n18523 ^ n13736 ;
  assign n20184 = ( n3899 & n5604 ) | ( n3899 & n5650 ) | ( n5604 & n5650 ) ;
  assign n20185 = n20184 ^ n15579 ^ n4988 ;
  assign n20186 = n20185 ^ n2339 ^ 1'b0 ;
  assign n20187 = n4281 & n20186 ;
  assign n20188 = n6633 & n20187 ;
  assign n20192 = n20191 ^ n20188 ^ 1'b0 ;
  assign n20193 = n12023 ^ n4475 ^ 1'b0 ;
  assign n20194 = n971 & ~n20193 ;
  assign n20195 = n20194 ^ n13852 ^ 1'b0 ;
  assign n20196 = n10402 & ~n14724 ;
  assign n20198 = ~n3284 & n3949 ;
  assign n20199 = n6116 & n20198 ;
  assign n20197 = n19758 ^ n16969 ^ n1130 ;
  assign n20200 = n20199 ^ n20197 ^ n17251 ;
  assign n20201 = ~n11995 & n12095 ;
  assign n20202 = n14025 ^ n9900 ^ n3870 ;
  assign n20203 = ( n13900 & ~n20201 ) | ( n13900 & n20202 ) | ( ~n20201 & n20202 ) ;
  assign n20204 = ( n2618 & n18876 ) | ( n2618 & ~n19477 ) | ( n18876 & ~n19477 ) ;
  assign n20205 = ( ~n17304 & n17969 ) | ( ~n17304 & n20204 ) | ( n17969 & n20204 ) ;
  assign n20206 = n3734 & n8282 ;
  assign n20207 = n15084 & n20206 ;
  assign n20208 = ( ~n3667 & n5046 ) | ( ~n3667 & n7230 ) | ( n5046 & n7230 ) ;
  assign n20209 = n8614 ^ n7605 ^ 1'b0 ;
  assign n20210 = n15352 & n20209 ;
  assign n20211 = n5489 ^ n3057 ^ n1638 ;
  assign n20212 = ( n4886 & n19564 ) | ( n4886 & n20211 ) | ( n19564 & n20211 ) ;
  assign n20213 = n20212 ^ n8055 ^ 1'b0 ;
  assign n20216 = n7902 ^ n4761 ^ n3153 ;
  assign n20214 = ( ~n7299 & n14900 ) | ( ~n7299 & n16753 ) | ( n14900 & n16753 ) ;
  assign n20215 = n8921 & n20214 ;
  assign n20217 = n20216 ^ n20215 ^ n994 ;
  assign n20218 = n7049 ^ n2089 ^ 1'b0 ;
  assign n20219 = n2032 | n20218 ;
  assign n20220 = n9367 | n20219 ;
  assign n20221 = n20220 ^ n6309 ^ 1'b0 ;
  assign n20222 = ( ~n2884 & n14063 ) | ( ~n2884 & n20221 ) | ( n14063 & n20221 ) ;
  assign n20223 = n20222 ^ n14483 ^ n10470 ;
  assign n20225 = ( n282 & n5103 ) | ( n282 & n17137 ) | ( n5103 & n17137 ) ;
  assign n20226 = ( ~n6248 & n16232 ) | ( ~n6248 & n20225 ) | ( n16232 & n20225 ) ;
  assign n20227 = n20226 ^ n9250 ^ n746 ;
  assign n20228 = n20227 ^ n17315 ^ n5898 ;
  assign n20224 = ~n15559 & n15785 ;
  assign n20229 = n20228 ^ n20224 ^ 1'b0 ;
  assign n20238 = n7377 & ~n14725 ;
  assign n20233 = ( n2396 & ~n3926 ) | ( n2396 & n9802 ) | ( ~n3926 & n9802 ) ;
  assign n20234 = ( n2239 & ~n4130 ) | ( n2239 & n7917 ) | ( ~n4130 & n7917 ) ;
  assign n20235 = n20234 ^ n143 ^ x51 ;
  assign n20236 = ( ~n17185 & n20233 ) | ( ~n17185 & n20235 ) | ( n20233 & n20235 ) ;
  assign n20231 = n5702 ^ n4152 ^ n4101 ;
  assign n20232 = ( n495 & n6967 ) | ( n495 & n20231 ) | ( n6967 & n20231 ) ;
  assign n20237 = n20236 ^ n20232 ^ n1033 ;
  assign n20230 = n942 & ~n9053 ;
  assign n20239 = n20238 ^ n20237 ^ n20230 ;
  assign n20240 = n14306 ^ n11042 ^ n7382 ;
  assign n20241 = n9812 | n20240 ;
  assign n20242 = n11929 ^ n10961 ^ 1'b0 ;
  assign n20243 = n900 | n14986 ;
  assign n20244 = n6720 | n20243 ;
  assign n20245 = n12464 & n20244 ;
  assign n20246 = ~n20242 & n20245 ;
  assign n20250 = n11706 ^ n3723 ^ n2608 ;
  assign n20251 = ( n11496 & n17370 ) | ( n11496 & n20250 ) | ( n17370 & n20250 ) ;
  assign n20247 = n1153 | n3393 ;
  assign n20248 = n5692 & ~n20247 ;
  assign n20249 = ( n3049 & ~n6786 ) | ( n3049 & n20248 ) | ( ~n6786 & n20248 ) ;
  assign n20252 = n20251 ^ n20249 ^ n1462 ;
  assign n20253 = n12707 ^ n3296 ^ 1'b0 ;
  assign n20254 = ( ~n17816 & n20252 ) | ( ~n17816 & n20253 ) | ( n20252 & n20253 ) ;
  assign n20255 = n15572 ^ n9602 ^ n7063 ;
  assign n20256 = ( n3737 & ~n15710 ) | ( n3737 & n20255 ) | ( ~n15710 & n20255 ) ;
  assign n20257 = n5738 & n18520 ;
  assign n20258 = n9556 & n20257 ;
  assign n20259 = n20258 ^ n18329 ^ 1'b0 ;
  assign n20260 = ~n1461 & n6927 ;
  assign n20261 = n8906 & n20260 ;
  assign n20262 = ( n19620 & n20259 ) | ( n19620 & n20261 ) | ( n20259 & n20261 ) ;
  assign n20263 = n12514 ^ n10629 ^ n6985 ;
  assign n20264 = ~n545 & n20263 ;
  assign n20265 = n19875 ^ n18883 ^ n9215 ;
  assign n20269 = n1183 & n13824 ;
  assign n20266 = ~n4468 & n12792 ;
  assign n20267 = n20266 ^ n4991 ^ 1'b0 ;
  assign n20268 = n1796 & n20267 ;
  assign n20270 = n20269 ^ n20268 ^ n17052 ;
  assign n20271 = n1865 & n18612 ;
  assign n20272 = n8489 ^ n7868 ^ 1'b0 ;
  assign n20273 = ~n20271 & n20272 ;
  assign n20274 = n9247 ^ n7272 ^ 1'b0 ;
  assign n20275 = n15100 ^ n6503 ^ 1'b0 ;
  assign n20276 = n20274 & ~n20275 ;
  assign n20277 = ( n2733 & n8473 ) | ( n2733 & ~n12662 ) | ( n8473 & ~n12662 ) ;
  assign n20278 = n14492 & ~n20277 ;
  assign n20279 = n20278 ^ n6785 ^ 1'b0 ;
  assign n20280 = ( ~n3305 & n9692 ) | ( ~n3305 & n17917 ) | ( n9692 & n17917 ) ;
  assign n20281 = n20280 ^ n9036 ^ n7705 ;
  assign n20283 = n14932 ^ n13414 ^ n10772 ;
  assign n20282 = n11182 ^ n1984 ^ n472 ;
  assign n20284 = n20283 ^ n20282 ^ n2996 ;
  assign n20285 = n9245 ^ n3689 ^ n1893 ;
  assign n20286 = ( n2542 & ~n10222 ) | ( n2542 & n20285 ) | ( ~n10222 & n20285 ) ;
  assign n20287 = n20286 ^ n11864 ^ n4012 ;
  assign n20288 = n4486 | n15656 ;
  assign n20289 = n20288 ^ n18296 ^ 1'b0 ;
  assign n20290 = n11806 ^ n3861 ^ 1'b0 ;
  assign n20291 = n18922 | n20290 ;
  assign n20292 = n4093 & ~n5969 ;
  assign n20293 = n20292 ^ n6350 ^ 1'b0 ;
  assign n20294 = n20293 ^ n3929 ^ n1880 ;
  assign n20295 = n20294 ^ n2114 ^ 1'b0 ;
  assign n20296 = n8833 & ~n20295 ;
  assign n20297 = n19985 ^ n18566 ^ n7673 ;
  assign n20299 = n657 & n1597 ;
  assign n20298 = ~n12428 & n15245 ;
  assign n20300 = n20299 ^ n20298 ^ 1'b0 ;
  assign n20301 = n15232 ^ n4614 ^ n3176 ;
  assign n20302 = ( n3530 & n16770 ) | ( n3530 & ~n20301 ) | ( n16770 & ~n20301 ) ;
  assign n20303 = n10080 ^ n5291 ^ n4481 ;
  assign n20304 = ( n3546 & ~n11267 ) | ( n3546 & n19782 ) | ( ~n11267 & n19782 ) ;
  assign n20306 = n12382 ^ n8815 ^ n7088 ;
  assign n20305 = n10333 ^ n6032 ^ 1'b0 ;
  assign n20307 = n20306 ^ n20305 ^ 1'b0 ;
  assign n20308 = ( n2221 & ~n9919 ) | ( n2221 & n10099 ) | ( ~n9919 & n10099 ) ;
  assign n20309 = n6165 & n15841 ;
  assign n20310 = n15930 ^ n1516 ^ 1'b0 ;
  assign n20311 = ~n1445 & n20310 ;
  assign n20313 = n5310 ^ n5193 ^ n411 ;
  assign n20312 = n7761 ^ n4228 ^ n1064 ;
  assign n20314 = n20313 ^ n20312 ^ n1238 ;
  assign n20315 = n20314 ^ n11897 ^ 1'b0 ;
  assign n20316 = n20315 ^ n8018 ^ n5023 ;
  assign n20317 = n6180 ^ n4721 ^ 1'b0 ;
  assign n20318 = ( n19408 & ~n20204 ) | ( n19408 & n20317 ) | ( ~n20204 & n20317 ) ;
  assign n20322 = n18174 ^ n10079 ^ n4836 ;
  assign n20320 = n14226 ^ n7638 ^ n897 ;
  assign n20319 = n12978 ^ n11512 ^ 1'b0 ;
  assign n20321 = n20320 ^ n20319 ^ n20022 ;
  assign n20323 = n20322 ^ n20321 ^ n10480 ;
  assign n20324 = n4980 | n10959 ;
  assign n20325 = n19993 & ~n20324 ;
  assign n20326 = n20325 ^ n10619 ^ n5325 ;
  assign n20327 = ( n4155 & n7752 ) | ( n4155 & ~n15300 ) | ( n7752 & ~n15300 ) ;
  assign n20328 = n5593 ^ n4641 ^ n165 ;
  assign n20329 = n7549 & ~n20328 ;
  assign n20330 = ( n16392 & n20327 ) | ( n16392 & ~n20329 ) | ( n20327 & ~n20329 ) ;
  assign n20331 = ~n3200 & n3967 ;
  assign n20332 = n13124 ^ n3122 ^ n1018 ;
  assign n20333 = ( ~n7956 & n11935 ) | ( ~n7956 & n20332 ) | ( n11935 & n20332 ) ;
  assign n20334 = n20333 ^ n7036 ^ 1'b0 ;
  assign n20335 = n17605 & n20334 ;
  assign n20336 = ( ~n12802 & n20331 ) | ( ~n12802 & n20335 ) | ( n20331 & n20335 ) ;
  assign n20337 = n16930 ^ n2406 ^ 1'b0 ;
  assign n20338 = n7909 | n20337 ;
  assign n20339 = n1833 & ~n14766 ;
  assign n20340 = n20339 ^ n2744 ^ 1'b0 ;
  assign n20341 = n20340 ^ n18874 ^ 1'b0 ;
  assign n20342 = n14547 & ~n20341 ;
  assign n20343 = n13508 ^ n3739 ^ 1'b0 ;
  assign n20344 = n11478 & ~n20343 ;
  assign n20345 = ( n7098 & ~n8947 ) | ( n7098 & n10392 ) | ( ~n8947 & n10392 ) ;
  assign n20346 = ~n14986 & n19295 ;
  assign n20347 = n8153 ^ n4778 ^ 1'b0 ;
  assign n20348 = ( ~n3501 & n9997 ) | ( ~n3501 & n12911 ) | ( n9997 & n12911 ) ;
  assign n20349 = n5836 ^ n3874 ^ 1'b0 ;
  assign n20350 = n20349 ^ n19725 ^ n11876 ;
  assign n20351 = n6884 ^ n2984 ^ 1'b0 ;
  assign n20352 = ( n11774 & n14812 ) | ( n11774 & ~n20351 ) | ( n14812 & ~n20351 ) ;
  assign n20353 = ( ~x19 & n9195 ) | ( ~x19 & n20352 ) | ( n9195 & n20352 ) ;
  assign n20354 = n15077 ^ n9907 ^ 1'b0 ;
  assign n20355 = n2452 & ~n20354 ;
  assign n20356 = n20355 ^ n2005 ^ 1'b0 ;
  assign n20357 = n11473 & ~n20356 ;
  assign n20358 = ( ~n4230 & n6133 ) | ( ~n4230 & n8888 ) | ( n6133 & n8888 ) ;
  assign n20359 = n20358 ^ n17208 ^ x52 ;
  assign n20360 = ( n5434 & n7194 ) | ( n5434 & ~n12201 ) | ( n7194 & ~n12201 ) ;
  assign n20361 = n20360 ^ n17377 ^ n4973 ;
  assign n20362 = n3188 | n20361 ;
  assign n20363 = n2224 | n20362 ;
  assign n20364 = ~n4229 & n20363 ;
  assign n20365 = ~n20359 & n20364 ;
  assign n20366 = n6252 | n17374 ;
  assign n20367 = n20366 ^ n8078 ^ 1'b0 ;
  assign n20368 = n13834 ^ n8794 ^ 1'b0 ;
  assign n20369 = ( n2009 & ~n9900 ) | ( n2009 & n20368 ) | ( ~n9900 & n20368 ) ;
  assign n20370 = ( n9941 & n10274 ) | ( n9941 & n16619 ) | ( n10274 & n16619 ) ;
  assign n20371 = n6343 ^ n1638 ^ n296 ;
  assign n20372 = ( n870 & ~n3643 ) | ( n870 & n20371 ) | ( ~n3643 & n20371 ) ;
  assign n20373 = ( n2781 & n20370 ) | ( n2781 & n20372 ) | ( n20370 & n20372 ) ;
  assign n20374 = n13643 ^ n6066 ^ 1'b0 ;
  assign n20375 = n6844 & ~n10055 ;
  assign n20376 = n16590 ^ n9999 ^ n3804 ;
  assign n20377 = ~n10009 & n20376 ;
  assign n20378 = ~n20375 & n20377 ;
  assign n20379 = n2061 & ~n17674 ;
  assign n20380 = n6208 & ~n13622 ;
  assign n20382 = n3581 & n7148 ;
  assign n20383 = ~n2693 & n20382 ;
  assign n20384 = n20383 ^ n1623 ^ n755 ;
  assign n20385 = n20384 ^ n9900 ^ n8719 ;
  assign n20381 = ( ~n4366 & n7130 ) | ( ~n4366 & n12094 ) | ( n7130 & n12094 ) ;
  assign n20386 = n20385 ^ n20381 ^ n12476 ;
  assign n20387 = ~n6364 & n20386 ;
  assign n20388 = ( n19628 & n20380 ) | ( n19628 & ~n20387 ) | ( n20380 & ~n20387 ) ;
  assign n20389 = n1337 & n14698 ;
  assign n20390 = ( ~n1234 & n3766 ) | ( ~n1234 & n6120 ) | ( n3766 & n6120 ) ;
  assign n20391 = n17896 | n20390 ;
  assign n20392 = n15262 & ~n20391 ;
  assign n20393 = ~n5318 & n8857 ;
  assign n20394 = n20393 ^ n542 ^ 1'b0 ;
  assign n20401 = ~n4188 & n12266 ;
  assign n20402 = n7686 & n20401 ;
  assign n20403 = ( n5332 & n7636 ) | ( n5332 & n20402 ) | ( n7636 & n20402 ) ;
  assign n20398 = ( n129 & ~n2408 ) | ( n129 & n3496 ) | ( ~n2408 & n3496 ) ;
  assign n20399 = ( n3136 & n4360 ) | ( n3136 & ~n20398 ) | ( n4360 & ~n20398 ) ;
  assign n20395 = n526 | n5509 ;
  assign n20396 = n11867 & ~n20395 ;
  assign n20397 = n17770 | n20396 ;
  assign n20400 = n20399 ^ n20397 ^ 1'b0 ;
  assign n20404 = n20403 ^ n20400 ^ n7050 ;
  assign n20405 = n14474 & n20006 ;
  assign n20406 = n20405 ^ n2898 ^ n2097 ;
  assign n20407 = n6039 ^ n4152 ^ n1187 ;
  assign n20408 = n20407 ^ n19183 ^ n4074 ;
  assign n20409 = n17443 ^ n11355 ^ 1'b0 ;
  assign n20410 = n2580 ^ n553 ^ 1'b0 ;
  assign n20411 = n11988 | n20410 ;
  assign n20412 = n14717 ^ n9117 ^ n6544 ;
  assign n20413 = n5724 & n7419 ;
  assign n20414 = n20413 ^ n866 ^ 1'b0 ;
  assign n20415 = ~n20412 & n20414 ;
  assign n20418 = ( n2145 & ~n6104 ) | ( n2145 & n6145 ) | ( ~n6104 & n6145 ) ;
  assign n20416 = n6275 ^ n1828 ^ 1'b0 ;
  assign n20417 = ~n7341 & n20416 ;
  assign n20419 = n20418 ^ n20417 ^ n8717 ;
  assign n20420 = n18317 ^ n12938 ^ 1'b0 ;
  assign n20421 = n20419 & n20420 ;
  assign n20422 = n20421 ^ n16543 ^ n5313 ;
  assign n20423 = n7304 & ~n9259 ;
  assign n20424 = n14424 ^ n5530 ^ n3464 ;
  assign n20425 = n20424 ^ n13372 ^ n7787 ;
  assign n20426 = n20425 ^ n13463 ^ n8691 ;
  assign n20427 = n20426 ^ n17063 ^ n14754 ;
  assign n20428 = n20399 ^ n15152 ^ n659 ;
  assign n20429 = n2857 | n9060 ;
  assign n20430 = ( n3573 & ~n7976 ) | ( n3573 & n20429 ) | ( ~n7976 & n20429 ) ;
  assign n20431 = n20430 ^ n2946 ^ 1'b0 ;
  assign n20432 = n2599 | n20431 ;
  assign n20433 = n3052 & n10407 ;
  assign n20434 = n10390 & n20433 ;
  assign n20435 = ( n11102 & ~n18885 ) | ( n11102 & n20434 ) | ( ~n18885 & n20434 ) ;
  assign n20436 = ( n2433 & n4734 ) | ( n2433 & ~n14484 ) | ( n4734 & ~n14484 ) ;
  assign n20437 = ( n7316 & ~n19691 ) | ( n7316 & n20436 ) | ( ~n19691 & n20436 ) ;
  assign n20449 = ( n495 & ~n15203 ) | ( n495 & n16322 ) | ( ~n15203 & n16322 ) ;
  assign n20446 = n2400 ^ n1697 ^ n1390 ;
  assign n20447 = n20446 ^ n8609 ^ 1'b0 ;
  assign n20448 = ( n1624 & ~n13440 ) | ( n1624 & n20447 ) | ( ~n13440 & n20447 ) ;
  assign n20438 = ( n1915 & n5827 ) | ( n1915 & ~n8461 ) | ( n5827 & ~n8461 ) ;
  assign n20439 = n20438 ^ n14206 ^ n8295 ;
  assign n20440 = n1286 & ~n5725 ;
  assign n20441 = n11089 & n20440 ;
  assign n20442 = ( ~n1571 & n8473 ) | ( ~n1571 & n8567 ) | ( n8473 & n8567 ) ;
  assign n20443 = n8739 & ~n20442 ;
  assign n20444 = n15162 & n20443 ;
  assign n20445 = ( n20439 & ~n20441 ) | ( n20439 & n20444 ) | ( ~n20441 & n20444 ) ;
  assign n20450 = n20449 ^ n20448 ^ n20445 ;
  assign n20451 = n18337 ^ n14443 ^ n13072 ;
  assign n20452 = ( n5945 & n7141 ) | ( n5945 & ~n20451 ) | ( n7141 & ~n20451 ) ;
  assign n20453 = n10136 ^ n8402 ^ n6960 ;
  assign n20454 = n20453 ^ n7827 ^ n3523 ;
  assign n20455 = n20454 ^ n17163 ^ n10489 ;
  assign n20456 = n16896 ^ n8780 ^ n1959 ;
  assign n20457 = ( n1027 & n7569 ) | ( n1027 & n20456 ) | ( n7569 & n20456 ) ;
  assign n20458 = n20457 ^ n12621 ^ n2827 ;
  assign n20459 = ( ~n1125 & n1126 ) | ( ~n1125 & n15006 ) | ( n1126 & n15006 ) ;
  assign n20460 = n6845 ^ n4228 ^ n3138 ;
  assign n20461 = ( ~n799 & n3129 ) | ( ~n799 & n11087 ) | ( n3129 & n11087 ) ;
  assign n20462 = n20461 ^ n8300 ^ n8252 ;
  assign n20463 = n8275 | n20462 ;
  assign n20464 = ( n1407 & ~n4014 ) | ( n1407 & n12643 ) | ( ~n4014 & n12643 ) ;
  assign n20465 = n7780 & n20464 ;
  assign n20466 = n16494 & n20465 ;
  assign n20470 = ( ~n468 & n4731 ) | ( ~n468 & n7031 ) | ( n4731 & n7031 ) ;
  assign n20468 = n17134 ^ n2205 ^ n1379 ;
  assign n20469 = n16310 & ~n20468 ;
  assign n20471 = n20470 ^ n20469 ^ 1'b0 ;
  assign n20467 = n4104 | n7269 ;
  assign n20472 = n20471 ^ n20467 ^ 1'b0 ;
  assign n20475 = ( ~n4292 & n5740 ) | ( ~n4292 & n10718 ) | ( n5740 & n10718 ) ;
  assign n20473 = n1416 | n10431 ;
  assign n20474 = n20473 ^ n10830 ^ 1'b0 ;
  assign n20476 = n20475 ^ n20474 ^ n6222 ;
  assign n20477 = n4333 ^ n2035 ^ n969 ;
  assign n20478 = n10176 ^ n5368 ^ n4077 ;
  assign n20479 = ( n13865 & ~n20477 ) | ( n13865 & n20478 ) | ( ~n20477 & n20478 ) ;
  assign n20480 = n20479 ^ n761 ^ 1'b0 ;
  assign n20481 = n13031 ^ n3967 ^ n359 ;
  assign n20482 = ~n9116 & n20481 ;
  assign n20483 = n20482 ^ n9835 ^ 1'b0 ;
  assign n20484 = n4756 | n10575 ;
  assign n20485 = n20484 ^ n9767 ^ 1'b0 ;
  assign n20486 = n20483 & n20485 ;
  assign n20487 = n20486 ^ n1134 ^ 1'b0 ;
  assign n20488 = n20418 ^ n6690 ^ 1'b0 ;
  assign n20489 = ~n14386 & n20488 ;
  assign n20490 = ( n5924 & ~n5968 ) | ( n5924 & n14187 ) | ( ~n5968 & n14187 ) ;
  assign n20491 = n20490 ^ n1197 ^ 1'b0 ;
  assign n20492 = n2457 & n5079 ;
  assign n20493 = n20492 ^ n4611 ^ 1'b0 ;
  assign n20494 = n13953 ^ n12081 ^ n11942 ;
  assign n20495 = n20494 ^ n6253 ^ 1'b0 ;
  assign n20496 = n20493 & n20495 ;
  assign n20497 = n1251 | n3466 ;
  assign n20498 = n2798 | n20497 ;
  assign n20499 = n20498 ^ n18261 ^ n10555 ;
  assign n20500 = n20499 ^ n15012 ^ 1'b0 ;
  assign n20501 = n15544 ^ n1313 ^ n994 ;
  assign n20502 = n5945 ^ n1785 ^ 1'b0 ;
  assign n20503 = n20502 ^ n11352 ^ n4520 ;
  assign n20504 = n18080 | n20503 ;
  assign n20505 = ( ~n10013 & n11078 ) | ( ~n10013 & n13953 ) | ( n11078 & n13953 ) ;
  assign n20506 = n12428 ^ n4564 ^ 1'b0 ;
  assign n20507 = n8886 & ~n20506 ;
  assign n20511 = n8354 & ~n13198 ;
  assign n20512 = ~n6485 & n20511 ;
  assign n20508 = ~n153 & n4236 ;
  assign n20509 = ( n5322 & n20436 ) | ( n5322 & ~n20508 ) | ( n20436 & ~n20508 ) ;
  assign n20510 = n20509 ^ n14206 ^ n213 ;
  assign n20513 = n20512 ^ n20510 ^ n19875 ;
  assign n20514 = ~n6099 & n20513 ;
  assign n20515 = n20514 ^ n10590 ^ 1'b0 ;
  assign n20516 = ( n1712 & n4181 ) | ( n1712 & n4734 ) | ( n4181 & n4734 ) ;
  assign n20517 = n20516 ^ n19522 ^ n8382 ;
  assign n20518 = n5389 ^ x98 ^ 1'b0 ;
  assign n20519 = n20517 | n20518 ;
  assign n20520 = n20519 ^ n11235 ^ 1'b0 ;
  assign n20521 = n13580 ^ n9147 ^ 1'b0 ;
  assign n20522 = ( n486 & ~n1372 ) | ( n486 & n5447 ) | ( ~n1372 & n5447 ) ;
  assign n20523 = n3697 ^ x91 ^ 1'b0 ;
  assign n20524 = n6923 & ~n20523 ;
  assign n20525 = ( n4610 & n20522 ) | ( n4610 & ~n20524 ) | ( n20522 & ~n20524 ) ;
  assign n20526 = n14500 ^ n14128 ^ n2844 ;
  assign n20527 = ~n2734 & n19235 ;
  assign n20528 = ~n13891 & n20527 ;
  assign n20532 = ~n5254 & n18952 ;
  assign n20533 = ~n139 & n20532 ;
  assign n20529 = n2041 | n3318 ;
  assign n20530 = n4135 | n20529 ;
  assign n20531 = ( n4580 & n7941 ) | ( n4580 & ~n20530 ) | ( n7941 & ~n20530 ) ;
  assign n20534 = n20533 ^ n20531 ^ n8819 ;
  assign n20535 = ( n2479 & ~n2541 ) | ( n2479 & n13741 ) | ( ~n2541 & n13741 ) ;
  assign n20536 = n20535 ^ n9845 ^ n1644 ;
  assign n20537 = ~n3637 & n8594 ;
  assign n20538 = n3877 | n8590 ;
  assign n20539 = n15919 ^ n7947 ^ 1'b0 ;
  assign n20540 = n20538 & ~n20539 ;
  assign n20541 = n20540 ^ n11393 ^ n6251 ;
  assign n20542 = n20537 & n20541 ;
  assign n20543 = n2789 | n7890 ;
  assign n20544 = n19871 ^ n4474 ^ n562 ;
  assign n20545 = ( ~n1066 & n4504 ) | ( ~n1066 & n20544 ) | ( n4504 & n20544 ) ;
  assign n20546 = ~n646 & n20228 ;
  assign n20547 = ( n20543 & n20545 ) | ( n20543 & n20546 ) | ( n20545 & n20546 ) ;
  assign n20550 = n5387 & ~n7612 ;
  assign n20551 = n2047 & n20550 ;
  assign n20548 = n8381 ^ n7414 ^ 1'b0 ;
  assign n20549 = n14266 & ~n20548 ;
  assign n20552 = n20551 ^ n20549 ^ n19612 ;
  assign n20553 = ( n3804 & n8164 ) | ( n3804 & ~n14354 ) | ( n8164 & ~n14354 ) ;
  assign n20555 = n1226 | n5973 ;
  assign n20554 = n10179 & n18378 ;
  assign n20556 = n20555 ^ n20554 ^ 1'b0 ;
  assign n20557 = n15676 | n19935 ;
  assign n20558 = n20557 ^ n13757 ^ n8242 ;
  assign n20559 = n9856 | n13192 ;
  assign n20560 = n5117 & n20559 ;
  assign n20561 = ~n20558 & n20560 ;
  assign n20562 = n20561 ^ n8337 ^ 1'b0 ;
  assign n20563 = n18150 | n20562 ;
  assign n20569 = ( n367 & n10139 ) | ( n367 & ~n14331 ) | ( n10139 & ~n14331 ) ;
  assign n20565 = n11312 & ~n17247 ;
  assign n20566 = n12271 & ~n18431 ;
  assign n20567 = ( n1941 & n20565 ) | ( n1941 & ~n20566 ) | ( n20565 & ~n20566 ) ;
  assign n20568 = n20567 ^ n16616 ^ n11342 ;
  assign n20564 = n6066 | n6918 ;
  assign n20570 = n20569 ^ n20568 ^ n20564 ;
  assign n20571 = n7522 ^ n3606 ^ n1407 ;
  assign n20572 = n20571 ^ n17538 ^ n10752 ;
  assign n20573 = ( ~n6083 & n6242 ) | ( ~n6083 & n20572 ) | ( n6242 & n20572 ) ;
  assign n20574 = ( n6199 & ~n13160 ) | ( n6199 & n20573 ) | ( ~n13160 & n20573 ) ;
  assign n20575 = n7845 ^ n1298 ^ n1069 ;
  assign n20576 = n12786 ^ n3570 ^ n2283 ;
  assign n20577 = n17665 & ~n20576 ;
  assign n20578 = ( n2668 & ~n11166 ) | ( n2668 & n20577 ) | ( ~n11166 & n20577 ) ;
  assign n20579 = n16656 ^ n223 ^ 1'b0 ;
  assign n20580 = ( ~n8878 & n16897 ) | ( ~n8878 & n20579 ) | ( n16897 & n20579 ) ;
  assign n20581 = ( n20575 & n20578 ) | ( n20575 & n20580 ) | ( n20578 & n20580 ) ;
  assign n20582 = n4804 & ~n6233 ;
  assign n20583 = n12316 & ~n14979 ;
  assign n20584 = n20583 ^ n17525 ^ n4273 ;
  assign n20585 = ( ~n5196 & n10868 ) | ( ~n5196 & n20584 ) | ( n10868 & n20584 ) ;
  assign n20586 = n8943 ^ n8527 ^ n5324 ;
  assign n20587 = n20586 ^ n2821 ^ 1'b0 ;
  assign n20588 = ~n12422 & n20587 ;
  assign n20590 = ( x31 & n4234 ) | ( x31 & n5308 ) | ( n4234 & n5308 ) ;
  assign n20589 = n1285 & ~n15735 ;
  assign n20591 = n20590 ^ n20589 ^ 1'b0 ;
  assign n20592 = n1565 | n20591 ;
  assign n20595 = ~n1670 & n10232 ;
  assign n20596 = n20595 ^ n14673 ^ 1'b0 ;
  assign n20593 = ( n1233 & n2366 ) | ( n1233 & ~n12016 ) | ( n2366 & ~n12016 ) ;
  assign n20594 = n5686 | n20593 ;
  assign n20597 = n20596 ^ n20594 ^ 1'b0 ;
  assign n20599 = n2370 ^ n2175 ^ 1'b0 ;
  assign n20600 = n2025 & n20599 ;
  assign n20598 = n1425 & n16476 ;
  assign n20601 = n20600 ^ n20598 ^ 1'b0 ;
  assign n20602 = n3134 & ~n5405 ;
  assign n20603 = ~n2338 & n20602 ;
  assign n20604 = ( n7437 & n20601 ) | ( n7437 & n20603 ) | ( n20601 & n20603 ) ;
  assign n20605 = n13843 ^ n9206 ^ n6172 ;
  assign n20606 = n14687 & ~n16934 ;
  assign n20607 = n2404 & n20606 ;
  assign n20614 = ( ~n2293 & n6984 ) | ( ~n2293 & n20396 ) | ( n6984 & n20396 ) ;
  assign n20615 = n11383 & ~n20614 ;
  assign n20616 = n20615 ^ n14906 ^ 1'b0 ;
  assign n20617 = ( ~n280 & n3571 ) | ( ~n280 & n20616 ) | ( n3571 & n20616 ) ;
  assign n20608 = n4663 & n8385 ;
  assign n20609 = ~n12171 & n20608 ;
  assign n20610 = n20609 ^ n4250 ^ 1'b0 ;
  assign n20611 = n20610 ^ n10563 ^ n5226 ;
  assign n20612 = n20611 ^ n2341 ^ 1'b0 ;
  assign n20613 = n3986 & ~n20612 ;
  assign n20618 = n20617 ^ n20613 ^ n13965 ;
  assign n20620 = n5365 | n5644 ;
  assign n20621 = n5997 & ~n20620 ;
  assign n20622 = n20621 ^ n822 ^ 1'b0 ;
  assign n20619 = ~n5661 & n20274 ;
  assign n20623 = n20622 ^ n20619 ^ 1'b0 ;
  assign n20624 = n20623 ^ n9338 ^ 1'b0 ;
  assign n20625 = ~n20618 & n20624 ;
  assign n20626 = n5854 ^ n5265 ^ n4881 ;
  assign n20627 = ~n10843 & n20626 ;
  assign n20628 = n7984 & n20627 ;
  assign n20629 = n10692 & ~n20628 ;
  assign n20630 = n3782 & n20629 ;
  assign n20631 = n9703 ^ n6942 ^ 1'b0 ;
  assign n20635 = ( n3794 & ~n4834 ) | ( n3794 & n10825 ) | ( ~n4834 & n10825 ) ;
  assign n20634 = n5426 & ~n7264 ;
  assign n20632 = ( n883 & n1373 ) | ( n883 & ~n6880 ) | ( n1373 & ~n6880 ) ;
  assign n20633 = ( ~n1468 & n8458 ) | ( ~n1468 & n20632 ) | ( n8458 & n20632 ) ;
  assign n20636 = n20635 ^ n20634 ^ n20633 ;
  assign n20637 = ( n1524 & ~n3518 ) | ( n1524 & n18733 ) | ( ~n3518 & n18733 ) ;
  assign n20638 = n15593 ^ n13679 ^ n11752 ;
  assign n20639 = ( n8266 & ~n8571 ) | ( n8266 & n15258 ) | ( ~n8571 & n15258 ) ;
  assign n20640 = ~n8888 & n20639 ;
  assign n20641 = ( n1306 & n7467 ) | ( n1306 & ~n16746 ) | ( n7467 & ~n16746 ) ;
  assign n20642 = n20641 ^ n11732 ^ 1'b0 ;
  assign n20643 = n2308 & ~n13136 ;
  assign n20644 = n20642 & n20643 ;
  assign n20645 = n6449 | n20644 ;
  assign n20646 = n20645 ^ n2332 ^ 1'b0 ;
  assign n20647 = n7874 ^ n6782 ^ 1'b0 ;
  assign n20648 = n13022 | n20647 ;
  assign n20649 = n487 | n11339 ;
  assign n20650 = n20649 ^ n267 ^ 1'b0 ;
  assign n20651 = ( n1277 & ~n4177 ) | ( n1277 & n20650 ) | ( ~n4177 & n20650 ) ;
  assign n20652 = ~n7381 & n20651 ;
  assign n20656 = ( x75 & n981 ) | ( x75 & ~n7927 ) | ( n981 & ~n7927 ) ;
  assign n20653 = ( n3005 & n3098 ) | ( n3005 & n9355 ) | ( n3098 & n9355 ) ;
  assign n20654 = ( n2636 & n3153 ) | ( n2636 & ~n3516 ) | ( n3153 & ~n3516 ) ;
  assign n20655 = ( n7270 & ~n20653 ) | ( n7270 & n20654 ) | ( ~n20653 & n20654 ) ;
  assign n20657 = n20656 ^ n20655 ^ n18783 ;
  assign n20658 = n6621 ^ n4738 ^ 1'b0 ;
  assign n20659 = n20658 ^ n9809 ^ 1'b0 ;
  assign n20660 = n4336 & n20659 ;
  assign n20661 = n20660 ^ n3322 ^ 1'b0 ;
  assign n20662 = n13800 & ~n20661 ;
  assign n20663 = n12209 | n20662 ;
  assign n20664 = ( ~n524 & n2362 ) | ( ~n524 & n4485 ) | ( n2362 & n4485 ) ;
  assign n20665 = n17325 ^ n10461 ^ n3147 ;
  assign n20666 = n20664 & ~n20665 ;
  assign n20667 = n20666 ^ n9729 ^ 1'b0 ;
  assign n20668 = n3272 ^ n1061 ^ 1'b0 ;
  assign n20669 = n5398 | n20668 ;
  assign n20670 = ( n6203 & n17763 ) | ( n6203 & n20669 ) | ( n17763 & n20669 ) ;
  assign n20671 = ( n13178 & n20611 ) | ( n13178 & n20670 ) | ( n20611 & n20670 ) ;
  assign n20672 = n16129 ^ n13733 ^ n1228 ;
  assign n20673 = n3352 & ~n4729 ;
  assign n20674 = n20673 ^ n1140 ^ 1'b0 ;
  assign n20675 = n4814 | n20674 ;
  assign n20676 = ( n1876 & ~n18863 ) | ( n1876 & n20675 ) | ( ~n18863 & n20675 ) ;
  assign n20677 = ~n7984 & n12992 ;
  assign n20678 = n19809 & n20677 ;
  assign n20679 = n20678 ^ n10110 ^ 1'b0 ;
  assign n20680 = n12246 & n20679 ;
  assign n20681 = n9797 ^ n2135 ^ 1'b0 ;
  assign n20682 = n6396 ^ n1712 ^ 1'b0 ;
  assign n20683 = n20681 & n20682 ;
  assign n20685 = n8843 | n11447 ;
  assign n20686 = n20685 ^ n17785 ^ 1'b0 ;
  assign n20684 = ~n8531 & n9174 ;
  assign n20687 = n20686 ^ n20684 ^ 1'b0 ;
  assign n20688 = n20687 ^ n14669 ^ 1'b0 ;
  assign n20689 = n7507 | n7795 ;
  assign n20691 = n8033 ^ n4342 ^ n1052 ;
  assign n20692 = n20691 ^ n3886 ^ 1'b0 ;
  assign n20690 = n666 & ~n4143 ;
  assign n20693 = n20692 ^ n20690 ^ 1'b0 ;
  assign n20694 = n9925 & ~n19654 ;
  assign n20695 = n14230 & n20694 ;
  assign n20696 = n12326 ^ n4683 ^ 1'b0 ;
  assign n20697 = n20696 ^ n17222 ^ n1920 ;
  assign n20698 = ( n7678 & n11431 ) | ( n7678 & n19502 ) | ( n11431 & n19502 ) ;
  assign n20699 = n16128 ^ n3872 ^ 1'b0 ;
  assign n20700 = n5741 ^ n3022 ^ 1'b0 ;
  assign n20701 = n20700 ^ n10520 ^ n6069 ;
  assign n20702 = n20701 ^ n4632 ^ 1'b0 ;
  assign n20703 = ( n6416 & n8764 ) | ( n6416 & n20702 ) | ( n8764 & n20702 ) ;
  assign n20704 = n20703 ^ n15568 ^ 1'b0 ;
  assign n20705 = n20699 | n20704 ;
  assign n20706 = ( n7117 & n16236 ) | ( n7117 & ~n18155 ) | ( n16236 & ~n18155 ) ;
  assign n20707 = n19981 ^ n11375 ^ 1'b0 ;
  assign n20708 = n20706 & ~n20707 ;
  assign n20709 = n5398 ^ n3947 ^ n1574 ;
  assign n20710 = n10635 | n13205 ;
  assign n20711 = n20710 ^ n632 ^ 1'b0 ;
  assign n20717 = n3726 ^ n3599 ^ 1'b0 ;
  assign n20718 = ~n4447 & n20717 ;
  assign n20712 = n13848 ^ n3032 ^ 1'b0 ;
  assign n20713 = n6148 & n18562 ;
  assign n20714 = n20713 ^ n13971 ^ 1'b0 ;
  assign n20715 = ( n3926 & n4279 ) | ( n3926 & ~n20714 ) | ( n4279 & ~n20714 ) ;
  assign n20716 = ( n10921 & n20712 ) | ( n10921 & ~n20715 ) | ( n20712 & ~n20715 ) ;
  assign n20719 = n20718 ^ n20716 ^ n18220 ;
  assign n20720 = n13665 ^ n11708 ^ 1'b0 ;
  assign n20721 = n1340 & ~n2077 ;
  assign n20722 = n20720 & n20721 ;
  assign n20723 = ( n2016 & n3164 ) | ( n2016 & ~n20722 ) | ( n3164 & ~n20722 ) ;
  assign n20724 = n1929 & ~n20723 ;
  assign n20725 = ~n5254 & n16237 ;
  assign n20726 = n20725 ^ n11739 ^ 1'b0 ;
  assign n20727 = ~n16165 & n20726 ;
  assign n20728 = n20727 ^ n18366 ^ n1669 ;
  assign n20729 = n15121 ^ n8496 ^ 1'b0 ;
  assign n20730 = n6067 | n6602 ;
  assign n20731 = n20730 ^ n1069 ^ x106 ;
  assign n20732 = ( n5354 & n12035 ) | ( n5354 & ~n20731 ) | ( n12035 & ~n20731 ) ;
  assign n20733 = n4816 | n16087 ;
  assign n20734 = n20733 ^ n4876 ^ 1'b0 ;
  assign n20735 = n10318 ^ n2946 ^ 1'b0 ;
  assign n20736 = n20735 ^ n18242 ^ n15020 ;
  assign n20737 = n20736 ^ n14505 ^ n10449 ;
  assign n20738 = ( ~n9355 & n10734 ) | ( ~n9355 & n18418 ) | ( n10734 & n18418 ) ;
  assign n20739 = ( n386 & n1340 ) | ( n386 & n5913 ) | ( n1340 & n5913 ) ;
  assign n20740 = ( n3640 & ~n13435 ) | ( n3640 & n20739 ) | ( ~n13435 & n20739 ) ;
  assign n20741 = n6995 ^ n5442 ^ n4268 ;
  assign n20742 = n14260 ^ n8674 ^ n4779 ;
  assign n20743 = ~n20741 & n20742 ;
  assign n20744 = n8330 & n20743 ;
  assign n20745 = ~n8416 & n18619 ;
  assign n20746 = n12148 & n20745 ;
  assign n20747 = ( n5858 & ~n11978 ) | ( n5858 & n16136 ) | ( ~n11978 & n16136 ) ;
  assign n20748 = n547 & n2375 ;
  assign n20749 = n10190 & n20748 ;
  assign n20750 = n20749 ^ n9467 ^ n564 ;
  assign n20751 = n20750 ^ n12928 ^ n1780 ;
  assign n20754 = n7706 ^ n1367 ^ n996 ;
  assign n20752 = n16823 ^ n600 ^ 1'b0 ;
  assign n20753 = n15435 & n20752 ;
  assign n20755 = n20754 ^ n20753 ^ n6794 ;
  assign n20758 = n18059 ^ n5270 ^ n5097 ;
  assign n20756 = ( ~n8911 & n13171 ) | ( ~n8911 & n19264 ) | ( n13171 & n19264 ) ;
  assign n20757 = ( n10975 & n17875 ) | ( n10975 & n20756 ) | ( n17875 & n20756 ) ;
  assign n20759 = n20758 ^ n20757 ^ 1'b0 ;
  assign n20760 = n9120 ^ n385 ^ 1'b0 ;
  assign n20761 = n20760 ^ n17296 ^ n7791 ;
  assign n20762 = ~n8200 & n11130 ;
  assign n20763 = n20762 ^ n6481 ^ 1'b0 ;
  assign n20764 = ( ~n2514 & n6092 ) | ( ~n2514 & n6897 ) | ( n6092 & n6897 ) ;
  assign n20765 = n20764 ^ n7561 ^ n7503 ;
  assign n20766 = ( n695 & n9452 ) | ( n695 & ~n9562 ) | ( n9452 & ~n9562 ) ;
  assign n20767 = ( n3627 & n16252 ) | ( n3627 & ~n20766 ) | ( n16252 & ~n20766 ) ;
  assign n20768 = n20765 | n20767 ;
  assign n20769 = ( n7849 & n8559 ) | ( n7849 & n12663 ) | ( n8559 & n12663 ) ;
  assign n20772 = n9937 ^ n6504 ^ n1750 ;
  assign n20770 = ( n6480 & n9682 ) | ( n6480 & n10892 ) | ( n9682 & n10892 ) ;
  assign n20771 = n8406 & ~n20770 ;
  assign n20773 = n20772 ^ n20771 ^ 1'b0 ;
  assign n20774 = n20773 ^ n9432 ^ n3950 ;
  assign n20775 = n4052 ^ n1433 ^ 1'b0 ;
  assign n20776 = ~n2386 & n20775 ;
  assign n20777 = ( n17478 & n18946 ) | ( n17478 & n20776 ) | ( n18946 & n20776 ) ;
  assign n20778 = ~n2049 & n16969 ;
  assign n20779 = ( n7823 & n16870 ) | ( n7823 & ~n20778 ) | ( n16870 & ~n20778 ) ;
  assign n20780 = n7392 ^ n3805 ^ n1191 ;
  assign n20781 = ( ~n593 & n16193 ) | ( ~n593 & n20780 ) | ( n16193 & n20780 ) ;
  assign n20782 = n5063 | n11444 ;
  assign n20783 = n11468 & ~n20782 ;
  assign n20784 = n8060 ^ n5121 ^ 1'b0 ;
  assign n20785 = ~n2578 & n20784 ;
  assign n20786 = n20259 ^ n9031 ^ 1'b0 ;
  assign n20787 = n7920 | n20786 ;
  assign n20788 = n6562 ^ n4570 ^ 1'b0 ;
  assign n20789 = ( ~n3543 & n12053 ) | ( ~n3543 & n14957 ) | ( n12053 & n14957 ) ;
  assign n20790 = n18394 & ~n20789 ;
  assign n20791 = n20790 ^ n19558 ^ n14246 ;
  assign n20792 = n19111 ^ n8010 ^ n7437 ;
  assign n20793 = n20792 ^ n19032 ^ n435 ;
  assign n20794 = n17968 ^ n7357 ^ 1'b0 ;
  assign n20795 = n11594 | n20794 ;
  assign n20796 = ( ~n10920 & n11894 ) | ( ~n10920 & n13406 ) | ( n11894 & n13406 ) ;
  assign n20797 = n7033 | n14277 ;
  assign n20798 = n20797 ^ n20170 ^ 1'b0 ;
  assign n20799 = n20798 ^ n11406 ^ n3183 ;
  assign n20800 = ( n10682 & n20796 ) | ( n10682 & ~n20799 ) | ( n20796 & ~n20799 ) ;
  assign n20801 = n19993 ^ n7673 ^ 1'b0 ;
  assign n20802 = ( n1027 & n5812 ) | ( n1027 & ~n20801 ) | ( n5812 & ~n20801 ) ;
  assign n20813 = ( n7807 & ~n8785 ) | ( n7807 & n9229 ) | ( ~n8785 & n9229 ) ;
  assign n20808 = n1738 & ~n4170 ;
  assign n20809 = n440 & ~n2257 ;
  assign n20810 = ~n774 & n20809 ;
  assign n20811 = ( n13575 & n20808 ) | ( n13575 & ~n20810 ) | ( n20808 & ~n20810 ) ;
  assign n20812 = n20811 ^ n5318 ^ n3757 ;
  assign n20804 = ( n410 & n13126 ) | ( n410 & n16800 ) | ( n13126 & n16800 ) ;
  assign n20803 = ( n11334 & n11825 ) | ( n11334 & n18591 ) | ( n11825 & n18591 ) ;
  assign n20805 = n20804 ^ n20803 ^ n4361 ;
  assign n20806 = n20805 ^ n20074 ^ n7155 ;
  assign n20807 = ( n13458 & ~n17207 ) | ( n13458 & n20806 ) | ( ~n17207 & n20806 ) ;
  assign n20814 = n20813 ^ n20812 ^ n20807 ;
  assign n20815 = n19949 & ~n20730 ;
  assign n20816 = ~n4217 & n20815 ;
  assign n20818 = ( n6612 & n10523 ) | ( n6612 & ~n12055 ) | ( n10523 & ~n12055 ) ;
  assign n20819 = n10309 ^ n1800 ^ 1'b0 ;
  assign n20820 = n7098 | n20819 ;
  assign n20821 = ( ~n1646 & n20818 ) | ( ~n1646 & n20820 ) | ( n20818 & n20820 ) ;
  assign n20817 = n760 & ~n13986 ;
  assign n20822 = n20821 ^ n20817 ^ 1'b0 ;
  assign n20823 = n20078 ^ n5820 ^ 1'b0 ;
  assign n20825 = n4271 ^ n2593 ^ n1142 ;
  assign n20824 = ( n3834 & n7739 ) | ( n3834 & n10512 ) | ( n7739 & n10512 ) ;
  assign n20826 = n20825 ^ n20824 ^ n2707 ;
  assign n20828 = n13809 ^ n1951 ^ n1485 ;
  assign n20829 = n20828 ^ n17264 ^ n1365 ;
  assign n20830 = ( n7134 & n9765 ) | ( n7134 & n20829 ) | ( n9765 & n20829 ) ;
  assign n20827 = n18200 ^ n9471 ^ n2149 ;
  assign n20831 = n20830 ^ n20827 ^ n18753 ;
  assign n20832 = n13349 | n20124 ;
  assign n20833 = n20832 ^ n19414 ^ 1'b0 ;
  assign n20834 = n4636 ^ n4135 ^ n2320 ;
  assign n20835 = ( n477 & ~n9729 ) | ( n477 & n16114 ) | ( ~n9729 & n16114 ) ;
  assign n20836 = n9729 ^ n4732 ^ n3660 ;
  assign n20837 = ~n4679 & n11776 ;
  assign n20838 = n15768 & n20837 ;
  assign n20839 = n20838 ^ n18832 ^ n15396 ;
  assign n20840 = n5644 ^ n4754 ^ 1'b0 ;
  assign n20841 = n17727 ^ n8433 ^ 1'b0 ;
  assign n20842 = n4882 & ~n14326 ;
  assign n20843 = n20842 ^ n10116 ^ 1'b0 ;
  assign n20844 = n9030 | n20843 ;
  assign n20845 = n4790 | n20844 ;
  assign n20846 = n4848 & ~n20845 ;
  assign n20847 = n3090 ^ n1402 ^ n1125 ;
  assign n20848 = n1533 & n6733 ;
  assign n20849 = n20847 & n20848 ;
  assign n20850 = ( ~n3569 & n3796 ) | ( ~n3569 & n5851 ) | ( n3796 & n5851 ) ;
  assign n20851 = ( ~n13857 & n17688 ) | ( ~n13857 & n20850 ) | ( n17688 & n20850 ) ;
  assign n20852 = n20851 ^ n19549 ^ 1'b0 ;
  assign n20853 = n7771 ^ n5209 ^ 1'b0 ;
  assign n20854 = n4895 & n7323 ;
  assign n20855 = n20854 ^ n8038 ^ n892 ;
  assign n20856 = n12737 ^ n10684 ^ 1'b0 ;
  assign n20857 = n20855 & ~n20856 ;
  assign n20858 = n7466 ^ n6001 ^ n2551 ;
  assign n20859 = n20858 ^ n14687 ^ 1'b0 ;
  assign n20860 = n9369 & ~n20859 ;
  assign n20861 = n9615 & ~n20860 ;
  assign n20862 = n4380 ^ x47 ^ 1'b0 ;
  assign n20863 = n20862 ^ n16477 ^ n3399 ;
  assign n20864 = ( n5133 & ~n11222 ) | ( n5133 & n12173 ) | ( ~n11222 & n12173 ) ;
  assign n20865 = n20864 ^ n13278 ^ n8411 ;
  assign n20866 = n4141 | n20865 ;
  assign n20867 = n20866 ^ n16481 ^ 1'b0 ;
  assign n20868 = ( ~x60 & n1955 ) | ( ~x60 & n4956 ) | ( n1955 & n4956 ) ;
  assign n20869 = n20868 ^ n2338 ^ n1003 ;
  assign n20870 = n20869 ^ n3427 ^ 1'b0 ;
  assign n20871 = n365 & ~n3752 ;
  assign n20872 = n20871 ^ n3991 ^ 1'b0 ;
  assign n20873 = ~n20870 & n20872 ;
  assign n20874 = n20867 & n20873 ;
  assign n20875 = ~n20863 & n20874 ;
  assign n20876 = ( n4646 & n13077 ) | ( n4646 & n15593 ) | ( n13077 & n15593 ) ;
  assign n20877 = n3430 & n7018 ;
  assign n20878 = n20877 ^ n12372 ^ 1'b0 ;
  assign n20879 = n20878 ^ n17650 ^ n12347 ;
  assign n20880 = n20879 ^ n12835 ^ 1'b0 ;
  assign n20881 = n15272 ^ n4108 ^ 1'b0 ;
  assign n20882 = ( ~n3286 & n5012 ) | ( ~n3286 & n20881 ) | ( n5012 & n20881 ) ;
  assign n20883 = n9986 ^ n7416 ^ 1'b0 ;
  assign n20884 = ~n11494 & n20883 ;
  assign n20885 = n20882 & n20884 ;
  assign n20886 = ~n14065 & n20885 ;
  assign n20887 = n17120 ^ n10823 ^ n6357 ;
  assign n20892 = n7175 ^ n2531 ^ 1'b0 ;
  assign n20890 = ~n3822 & n18157 ;
  assign n20891 = n8533 & n20890 ;
  assign n20888 = x84 & n761 ;
  assign n20889 = n20888 ^ n15271 ^ n6528 ;
  assign n20893 = n20892 ^ n20891 ^ n20889 ;
  assign n20894 = ~n20887 & n20893 ;
  assign n20895 = ( n132 & n4126 ) | ( n132 & ~n12075 ) | ( n4126 & ~n12075 ) ;
  assign n20896 = n20895 ^ n18745 ^ 1'b0 ;
  assign n20897 = ~n285 & n10580 ;
  assign n20898 = n20897 ^ n1179 ^ 1'b0 ;
  assign n20899 = ~n11460 & n20898 ;
  assign n20900 = n2597 & n5375 ;
  assign n20901 = ( n8153 & n15501 ) | ( n8153 & n20641 ) | ( n15501 & n20641 ) ;
  assign n20902 = n18717 ^ n8231 ^ n6187 ;
  assign n20903 = n9258 | n12636 ;
  assign n20904 = n20903 ^ n1723 ^ 1'b0 ;
  assign n20905 = n10583 ^ n6572 ^ 1'b0 ;
  assign n20906 = n19798 ^ n11741 ^ n5436 ;
  assign n20914 = ( n3427 & n4765 ) | ( n3427 & n10071 ) | ( n4765 & n10071 ) ;
  assign n20907 = n3472 | n7825 ;
  assign n20908 = n7585 ^ n5405 ^ n3658 ;
  assign n20909 = ( n2343 & n2535 ) | ( n2343 & ~n6099 ) | ( n2535 & ~n6099 ) ;
  assign n20910 = n20909 ^ n7033 ^ n1938 ;
  assign n20911 = n20910 ^ n6126 ^ 1'b0 ;
  assign n20912 = n20908 & n20911 ;
  assign n20913 = ( n18575 & n20907 ) | ( n18575 & ~n20912 ) | ( n20907 & ~n20912 ) ;
  assign n20915 = n20914 ^ n20913 ^ n18195 ;
  assign n20916 = n7034 ^ n1032 ^ x59 ;
  assign n20917 = n1113 & n5086 ;
  assign n20918 = n20917 ^ n2198 ^ 1'b0 ;
  assign n20919 = n6540 & ~n20918 ;
  assign n20920 = n20919 ^ n18378 ^ n14921 ;
  assign n20921 = ( n15410 & ~n19159 ) | ( n15410 & n20804 ) | ( ~n19159 & n20804 ) ;
  assign n20922 = ( n4528 & n5926 ) | ( n4528 & ~n6347 ) | ( n5926 & ~n6347 ) ;
  assign n20923 = ~n15062 & n20922 ;
  assign n20924 = ~n19564 & n20923 ;
  assign n20929 = n16091 ^ n13799 ^ n2880 ;
  assign n20925 = n433 & ~n3408 ;
  assign n20926 = n20925 ^ n737 ^ 1'b0 ;
  assign n20927 = n14438 & n20926 ;
  assign n20928 = ( n10774 & n11530 ) | ( n10774 & ~n20927 ) | ( n11530 & ~n20927 ) ;
  assign n20930 = n20929 ^ n20928 ^ n8220 ;
  assign n20931 = n7224 ^ n1207 ^ 1'b0 ;
  assign n20932 = n20930 & n20931 ;
  assign n20933 = ~n4014 & n15771 ;
  assign n20934 = n20933 ^ n9938 ^ n8594 ;
  assign n20935 = n6596 ^ n4265 ^ n813 ;
  assign n20936 = n20935 ^ n6665 ^ n1074 ;
  assign n20937 = ( n11966 & n15050 ) | ( n11966 & n16193 ) | ( n15050 & n16193 ) ;
  assign n20938 = n20937 ^ n9841 ^ n2061 ;
  assign n20939 = n7031 ^ n3948 ^ 1'b0 ;
  assign n20940 = ( n225 & ~n566 ) | ( n225 & n2765 ) | ( ~n566 & n2765 ) ;
  assign n20941 = ( n1939 & n5177 ) | ( n1939 & ~n8754 ) | ( n5177 & ~n8754 ) ;
  assign n20942 = n20941 ^ n11929 ^ 1'b0 ;
  assign n20943 = ( n20939 & ~n20940 ) | ( n20939 & n20942 ) | ( ~n20940 & n20942 ) ;
  assign n20944 = n8954 & n20943 ;
  assign n20945 = n20944 ^ n3894 ^ 1'b0 ;
  assign n20946 = n10030 & n14855 ;
  assign n20947 = n15873 ^ n1058 ^ 1'b0 ;
  assign n20948 = ~n20946 & n20947 ;
  assign n20949 = n14084 ^ n12981 ^ 1'b0 ;
  assign n20950 = n7626 & n20949 ;
  assign n20951 = ( ~n3103 & n4189 ) | ( ~n3103 & n8745 ) | ( n4189 & n8745 ) ;
  assign n20952 = ( ~n1795 & n2032 ) | ( ~n1795 & n20951 ) | ( n2032 & n20951 ) ;
  assign n20953 = n20950 & n20952 ;
  assign n20954 = n5464 & n15550 ;
  assign n20960 = n379 | n826 ;
  assign n20957 = ( n1633 & n14101 ) | ( n1633 & n15879 ) | ( n14101 & n15879 ) ;
  assign n20955 = n8895 ^ n6886 ^ n3750 ;
  assign n20956 = n20955 ^ n4738 ^ 1'b0 ;
  assign n20958 = n20957 ^ n20956 ^ n810 ;
  assign n20959 = ( n298 & ~n988 ) | ( n298 & n20958 ) | ( ~n988 & n20958 ) ;
  assign n20961 = n20960 ^ n20959 ^ n20263 ;
  assign n20962 = n9379 & ~n9674 ;
  assign n20963 = n3014 ^ n976 ^ 1'b0 ;
  assign n20964 = n15843 & ~n20963 ;
  assign n20965 = n20964 ^ n5285 ^ n4092 ;
  assign n20966 = ( ~n2235 & n3666 ) | ( ~n2235 & n9247 ) | ( n3666 & n9247 ) ;
  assign n20967 = n20966 ^ n13337 ^ n8579 ;
  assign n20968 = n11326 | n20967 ;
  assign n20969 = n20968 ^ n5263 ^ 1'b0 ;
  assign n20970 = n1482 & n12372 ;
  assign n20976 = n5945 ^ n3000 ^ 1'b0 ;
  assign n20977 = n4941 & ~n20976 ;
  assign n20978 = n7661 ^ n4210 ^ n3758 ;
  assign n20979 = ( n16555 & ~n20977 ) | ( n16555 & n20978 ) | ( ~n20977 & n20978 ) ;
  assign n20971 = ( ~n1763 & n2964 ) | ( ~n1763 & n9988 ) | ( n2964 & n9988 ) ;
  assign n20972 = ( x31 & n9297 ) | ( x31 & ~n20971 ) | ( n9297 & ~n20971 ) ;
  assign n20973 = n20972 ^ n17541 ^ n565 ;
  assign n20974 = n20973 ^ n20252 ^ n676 ;
  assign n20975 = ( n9120 & n10425 ) | ( n9120 & ~n20974 ) | ( n10425 & ~n20974 ) ;
  assign n20980 = n20979 ^ n20975 ^ n13762 ;
  assign n20981 = n1395 & n3058 ;
  assign n20982 = n20981 ^ n1256 ^ 1'b0 ;
  assign n20983 = n20982 ^ n14490 ^ 1'b0 ;
  assign n20984 = ( ~n3019 & n6275 ) | ( ~n3019 & n6498 ) | ( n6275 & n6498 ) ;
  assign n20985 = ( n507 & n2685 ) | ( n507 & n7511 ) | ( n2685 & n7511 ) ;
  assign n20986 = n20985 ^ n16426 ^ n3464 ;
  assign n20987 = ( n6580 & n20984 ) | ( n6580 & n20986 ) | ( n20984 & n20986 ) ;
  assign n20988 = ( ~n2707 & n6766 ) | ( ~n2707 & n20987 ) | ( n6766 & n20987 ) ;
  assign n20992 = ( n1039 & ~n2039 ) | ( n1039 & n2893 ) | ( ~n2039 & n2893 ) ;
  assign n20989 = n6018 ^ n5714 ^ 1'b0 ;
  assign n20990 = n20989 ^ n13465 ^ n10291 ;
  assign n20991 = ~n9302 & n20990 ;
  assign n20993 = n20992 ^ n20991 ^ n11059 ;
  assign n20994 = n5380 & n20993 ;
  assign n20995 = ~n8199 & n20994 ;
  assign n20996 = n20995 ^ n20650 ^ n6586 ;
  assign n20997 = ( ~x36 & n6504 ) | ( ~x36 & n16136 ) | ( n6504 & n16136 ) ;
  assign n20998 = n18733 & ~n20997 ;
  assign n21002 = n4044 & ~n4946 ;
  assign n21003 = n21002 ^ n6355 ^ 1'b0 ;
  assign n20999 = ~n825 & n1055 ;
  assign n21000 = n20999 ^ n10269 ^ 1'b0 ;
  assign n21001 = n1418 & n21000 ;
  assign n21004 = n21003 ^ n21001 ^ 1'b0 ;
  assign n21005 = n6912 ^ n5602 ^ n1580 ;
  assign n21006 = ~n1550 & n21005 ;
  assign n21007 = ( ~n5985 & n8983 ) | ( ~n5985 & n12040 ) | ( n8983 & n12040 ) ;
  assign n21008 = n19694 & ~n21007 ;
  assign n21009 = n21008 ^ n9490 ^ n9116 ;
  assign n21010 = ( n199 & ~n7563 ) | ( n199 & n21009 ) | ( ~n7563 & n21009 ) ;
  assign n21011 = n19459 ^ n11823 ^ n2366 ;
  assign n21012 = n19627 ^ n15838 ^ n1381 ;
  assign n21013 = n21012 ^ n11161 ^ 1'b0 ;
  assign n21014 = ~n9761 & n21013 ;
  assign n21017 = n10618 ^ n1561 ^ 1'b0 ;
  assign n21018 = ( ~n816 & n5490 ) | ( ~n816 & n21017 ) | ( n5490 & n21017 ) ;
  assign n21015 = n11010 ^ n5041 ^ 1'b0 ;
  assign n21016 = n21015 ^ n9335 ^ 1'b0 ;
  assign n21019 = n21018 ^ n21016 ^ n4593 ;
  assign n21023 = n1240 | n1836 ;
  assign n21024 = ~n17636 & n21023 ;
  assign n21020 = ( ~n220 & n2882 ) | ( ~n220 & n11597 ) | ( n2882 & n11597 ) ;
  assign n21021 = n21020 ^ n7175 ^ n3798 ;
  assign n21022 = n21021 ^ n18479 ^ n851 ;
  assign n21025 = n21024 ^ n21022 ^ n6385 ;
  assign n21026 = n5443 | n19441 ;
  assign n21027 = n21026 ^ n11568 ^ n4529 ;
  assign n21030 = n11844 ^ n8855 ^ n5180 ;
  assign n21028 = ~n3130 & n12933 ;
  assign n21029 = n9339 & ~n21028 ;
  assign n21031 = n21030 ^ n21029 ^ 1'b0 ;
  assign n21032 = n13253 ^ n6572 ^ 1'b0 ;
  assign n21033 = x39 & n21032 ;
  assign n21034 = n10404 ^ n10329 ^ 1'b0 ;
  assign n21039 = n20811 ^ n18829 ^ n13562 ;
  assign n21038 = n16318 ^ n7301 ^ n2061 ;
  assign n21036 = ( n2264 & ~n4744 ) | ( n2264 & n5526 ) | ( ~n4744 & n5526 ) ;
  assign n21035 = x43 | n12348 ;
  assign n21037 = n21036 ^ n21035 ^ n15065 ;
  assign n21040 = n21039 ^ n21038 ^ n21037 ;
  assign n21041 = n8336 ^ n6495 ^ n3925 ;
  assign n21042 = ( ~n1630 & n19453 ) | ( ~n1630 & n21041 ) | ( n19453 & n21041 ) ;
  assign n21047 = ( ~n6931 & n8090 ) | ( ~n6931 & n13977 ) | ( n8090 & n13977 ) ;
  assign n21048 = n21047 ^ n7052 ^ n2653 ;
  assign n21043 = x74 & n9043 ;
  assign n21044 = n857 | n2162 ;
  assign n21045 = n21043 & ~n21044 ;
  assign n21046 = n21045 ^ n1875 ^ n383 ;
  assign n21049 = n21048 ^ n21046 ^ n18368 ;
  assign n21053 = ~n1670 & n8785 ;
  assign n21054 = n15512 | n21053 ;
  assign n21050 = ( n8038 & n9652 ) | ( n8038 & n11185 ) | ( n9652 & n11185 ) ;
  assign n21051 = ~n551 & n13866 ;
  assign n21052 = n21050 | n21051 ;
  assign n21055 = n21054 ^ n21052 ^ n13831 ;
  assign n21056 = n8865 ^ n1851 ^ n1298 ;
  assign n21057 = n11889 ^ n5267 ^ n487 ;
  assign n21058 = ( n4991 & n21056 ) | ( n4991 & ~n21057 ) | ( n21056 & ~n21057 ) ;
  assign n21059 = ( ~n12280 & n13778 ) | ( ~n12280 & n21058 ) | ( n13778 & n21058 ) ;
  assign n21060 = n975 ^ x115 ^ 1'b0 ;
  assign n21061 = n6953 & n13234 ;
  assign n21062 = n19760 & ~n21061 ;
  assign n21063 = ~n6078 & n21062 ;
  assign n21064 = ( n301 & ~n20665 ) | ( n301 & n21063 ) | ( ~n20665 & n21063 ) ;
  assign n21067 = n14273 ^ n10873 ^ n3281 ;
  assign n21065 = n169 & ~n4191 ;
  assign n21066 = n1102 | n21065 ;
  assign n21068 = n21067 ^ n21066 ^ n584 ;
  assign n21069 = n8697 ^ n3449 ^ 1'b0 ;
  assign n21070 = ( n2771 & ~n8411 ) | ( n2771 & n10257 ) | ( ~n8411 & n10257 ) ;
  assign n21071 = ( ~n4170 & n5216 ) | ( ~n4170 & n21070 ) | ( n5216 & n21070 ) ;
  assign n21072 = n3376 & ~n5725 ;
  assign n21073 = n21072 ^ n10669 ^ 1'b0 ;
  assign n21074 = ( ~n2503 & n6228 ) | ( ~n2503 & n21073 ) | ( n6228 & n21073 ) ;
  assign n21075 = ( ~n9708 & n10934 ) | ( ~n9708 & n13045 ) | ( n10934 & n13045 ) ;
  assign n21076 = ~n3221 & n21075 ;
  assign n21077 = ( n1290 & n7148 ) | ( n1290 & ~n21076 ) | ( n7148 & ~n21076 ) ;
  assign n21078 = ( n1991 & n7631 ) | ( n1991 & n18879 ) | ( n7631 & n18879 ) ;
  assign n21079 = n13891 ^ n12534 ^ n1999 ;
  assign n21080 = n7158 & ~n8027 ;
  assign n21081 = ~n21079 & n21080 ;
  assign n21082 = n15274 ^ n11763 ^ 1'b0 ;
  assign n21083 = ~n5360 & n21082 ;
  assign n21084 = n21083 ^ n1265 ^ 1'b0 ;
  assign n21085 = n21081 | n21084 ;
  assign n21086 = ( ~n1822 & n8973 ) | ( ~n1822 & n21085 ) | ( n8973 & n21085 ) ;
  assign n21087 = n17609 ^ n15742 ^ n8290 ;
  assign n21088 = ( n791 & n15274 ) | ( n791 & ~n21087 ) | ( n15274 & ~n21087 ) ;
  assign n21089 = n2752 & n20641 ;
  assign n21090 = n21089 ^ n7013 ^ 1'b0 ;
  assign n21091 = n13198 ^ n1653 ^ 1'b0 ;
  assign n21092 = n9584 & n21091 ;
  assign n21093 = ~n16956 & n21092 ;
  assign n21094 = n10575 | n11935 ;
  assign n21095 = n21094 ^ n10993 ^ 1'b0 ;
  assign n21096 = n21095 ^ n8346 ^ 1'b0 ;
  assign n21097 = n161 | n1484 ;
  assign n21098 = n4839 & n21097 ;
  assign n21099 = n17853 ^ n1404 ^ 1'b0 ;
  assign n21100 = ( n8313 & n9490 ) | ( n8313 & ~n13152 ) | ( n9490 & ~n13152 ) ;
  assign n21101 = n15379 ^ n14357 ^ n6128 ;
  assign n21102 = n5558 | n21101 ;
  assign n21103 = n11862 & ~n21102 ;
  assign n21104 = ( n12708 & n17235 ) | ( n12708 & ~n21103 ) | ( n17235 & ~n21103 ) ;
  assign n21106 = ( n1459 & n9999 ) | ( n1459 & ~n17464 ) | ( n9999 & ~n17464 ) ;
  assign n21105 = n2542 & n4536 ;
  assign n21107 = n21106 ^ n21105 ^ 1'b0 ;
  assign n21108 = n576 & ~n3906 ;
  assign n21109 = n12660 ^ n11273 ^ n8302 ;
  assign n21110 = n21109 ^ n6711 ^ 1'b0 ;
  assign n21111 = ( ~n1582 & n16309 ) | ( ~n1582 & n18005 ) | ( n16309 & n18005 ) ;
  assign n21112 = ~n12451 & n13223 ;
  assign n21113 = n21112 ^ n5016 ^ 1'b0 ;
  assign n21114 = n8534 ^ n5334 ^ n2965 ;
  assign n21115 = ~n18776 & n19380 ;
  assign n21116 = n21018 ^ n7747 ^ 1'b0 ;
  assign n21117 = n21116 ^ n15635 ^ 1'b0 ;
  assign n21118 = n21115 & ~n21117 ;
  assign n21119 = n21118 ^ n14030 ^ 1'b0 ;
  assign n21120 = n21114 & n21119 ;
  assign n21121 = ( ~n4415 & n7862 ) | ( ~n4415 & n14287 ) | ( n7862 & n14287 ) ;
  assign n21122 = ( n4580 & ~n5862 ) | ( n4580 & n6011 ) | ( ~n5862 & n6011 ) ;
  assign n21123 = n21122 ^ n10716 ^ 1'b0 ;
  assign n21124 = n21121 & n21123 ;
  assign n21125 = n21124 ^ n13468 ^ n12590 ;
  assign n21126 = n6051 ^ n4525 ^ 1'b0 ;
  assign n21127 = n1311 | n21126 ;
  assign n21128 = n21127 ^ n11032 ^ n10334 ;
  assign n21129 = ( n1854 & n5726 ) | ( n1854 & n19297 ) | ( n5726 & n19297 ) ;
  assign n21133 = n13889 ^ n11419 ^ n5583 ;
  assign n21132 = ( ~n482 & n5798 ) | ( ~n482 & n18765 ) | ( n5798 & n18765 ) ;
  assign n21134 = n21133 ^ n21132 ^ 1'b0 ;
  assign n21135 = n11774 & ~n21134 ;
  assign n21130 = n8978 & ~n13051 ;
  assign n21131 = n17389 & ~n21130 ;
  assign n21136 = n21135 ^ n21131 ^ 1'b0 ;
  assign n21137 = ( ~n6071 & n12630 ) | ( ~n6071 & n18852 ) | ( n12630 & n18852 ) ;
  assign n21138 = n9715 ^ n6045 ^ n2581 ;
  assign n21139 = ( n1191 & ~n10355 ) | ( n1191 & n21138 ) | ( ~n10355 & n21138 ) ;
  assign n21140 = n10903 ^ n5478 ^ n1444 ;
  assign n21141 = n18425 & n18588 ;
  assign n21142 = n21141 ^ n14380 ^ 1'b0 ;
  assign n21143 = ~n21140 & n21142 ;
  assign n21152 = n15086 ^ n12227 ^ n10916 ;
  assign n21153 = n21152 ^ n10282 ^ n9411 ;
  assign n21144 = n20436 ^ n13746 ^ n10988 ;
  assign n21145 = n3064 ^ n716 ^ 1'b0 ;
  assign n21146 = n2346 & n21145 ;
  assign n21147 = ( n6135 & ~n7849 ) | ( n6135 & n21146 ) | ( ~n7849 & n21146 ) ;
  assign n21148 = ~n11623 & n21147 ;
  assign n21149 = n21144 & n21148 ;
  assign n21150 = n1289 | n21149 ;
  assign n21151 = n21150 ^ n18892 ^ 1'b0 ;
  assign n21154 = n21153 ^ n21151 ^ n18352 ;
  assign n21155 = ~n218 & n14910 ;
  assign n21156 = ( n3558 & n17433 ) | ( n3558 & n21155 ) | ( n17433 & n21155 ) ;
  assign n21157 = n21156 ^ n18256 ^ 1'b0 ;
  assign n21158 = ( ~n4474 & n14368 ) | ( ~n4474 & n14815 ) | ( n14368 & n14815 ) ;
  assign n21159 = n21158 ^ n20475 ^ n3240 ;
  assign n21160 = ( n6556 & ~n10451 ) | ( n6556 & n21159 ) | ( ~n10451 & n21159 ) ;
  assign n21161 = n13821 & ~n21160 ;
  assign n21162 = n21161 ^ n3096 ^ 1'b0 ;
  assign n21163 = n10110 ^ n4115 ^ 1'b0 ;
  assign n21164 = n16017 ^ n9281 ^ n3599 ;
  assign n21165 = ( n2421 & n7367 ) | ( n2421 & n8005 ) | ( n7367 & n8005 ) ;
  assign n21166 = ( n3786 & n20742 ) | ( n3786 & ~n21165 ) | ( n20742 & ~n21165 ) ;
  assign n21167 = ( n3335 & n11276 ) | ( n3335 & n17733 ) | ( n11276 & n17733 ) ;
  assign n21168 = n15995 ^ n5820 ^ 1'b0 ;
  assign n21169 = n21168 ^ n16227 ^ n4302 ;
  assign n21170 = ( ~n1306 & n5615 ) | ( ~n1306 & n13214 ) | ( n5615 & n13214 ) ;
  assign n21171 = n21170 ^ n18505 ^ n9505 ;
  assign n21172 = n4834 & n12627 ;
  assign n21173 = n7264 ^ n1607 ^ n1069 ;
  assign n21174 = n11536 ^ n2516 ^ 1'b0 ;
  assign n21175 = ~n17266 & n21174 ;
  assign n21176 = ( ~n21172 & n21173 ) | ( ~n21172 & n21175 ) | ( n21173 & n21175 ) ;
  assign n21177 = n1589 & ~n21176 ;
  assign n21178 = ( n12359 & n13715 ) | ( n12359 & n16747 ) | ( n13715 & n16747 ) ;
  assign n21180 = n4810 ^ n2809 ^ n2738 ;
  assign n21179 = n13338 ^ n10311 ^ n1785 ;
  assign n21181 = n21180 ^ n21179 ^ 1'b0 ;
  assign n21182 = ~n14421 & n21181 ;
  assign n21183 = ~n21178 & n21182 ;
  assign n21184 = ~n8200 & n18026 ;
  assign n21185 = ~n9719 & n21184 ;
  assign n21186 = n12449 ^ n10379 ^ 1'b0 ;
  assign n21187 = n6056 & n17830 ;
  assign n21188 = ~n17291 & n21187 ;
  assign n21193 = n2733 | n16654 ;
  assign n21189 = n8632 ^ n2364 ^ 1'b0 ;
  assign n21190 = n19434 ^ n2958 ^ 1'b0 ;
  assign n21191 = n21189 & ~n21190 ;
  assign n21192 = n16338 & n21191 ;
  assign n21194 = n21193 ^ n21192 ^ 1'b0 ;
  assign n21195 = n17431 | n19058 ;
  assign n21196 = n21195 ^ n12788 ^ 1'b0 ;
  assign n21197 = n12490 ^ n9482 ^ n1102 ;
  assign n21198 = n5051 & ~n5870 ;
  assign n21199 = n1676 | n12191 ;
  assign n21201 = n1980 | n14936 ;
  assign n21202 = n8590 | n21201 ;
  assign n21200 = n5261 | n19995 ;
  assign n21203 = n21202 ^ n21200 ^ 1'b0 ;
  assign n21206 = n14729 ^ n161 ^ 1'b0 ;
  assign n21207 = n19374 & ~n21206 ;
  assign n21208 = ( n2779 & n12023 ) | ( n2779 & ~n21207 ) | ( n12023 & ~n21207 ) ;
  assign n21204 = ( n4245 & n6148 ) | ( n4245 & n16023 ) | ( n6148 & n16023 ) ;
  assign n21205 = ~n1101 & n21204 ;
  assign n21209 = n21208 ^ n21205 ^ 1'b0 ;
  assign n21210 = n1139 & ~n9943 ;
  assign n21211 = n9184 ^ n5424 ^ n1465 ;
  assign n21212 = n21211 ^ n17688 ^ n1686 ;
  assign n21213 = ( n3365 & n8072 ) | ( n3365 & ~n21212 ) | ( n8072 & ~n21212 ) ;
  assign n21214 = ~n8865 & n15772 ;
  assign n21215 = n4339 & n11476 ;
  assign n21216 = n21215 ^ n10445 ^ 1'b0 ;
  assign n21217 = ( n13414 & n14312 ) | ( n13414 & ~n21216 ) | ( n14312 & ~n21216 ) ;
  assign n21219 = ( ~n1159 & n1534 ) | ( ~n1159 & n8102 ) | ( n1534 & n8102 ) ;
  assign n21218 = n17745 ^ n14456 ^ n11260 ;
  assign n21220 = n21219 ^ n21218 ^ n17866 ;
  assign n21221 = n21220 ^ n17020 ^ n11083 ;
  assign n21222 = n7262 ^ n164 ^ x121 ;
  assign n21223 = n16374 ^ n4249 ^ n1170 ;
  assign n21224 = n21223 ^ n9384 ^ 1'b0 ;
  assign n21225 = n8560 & n21224 ;
  assign n21226 = n7218 ^ n1399 ^ 1'b0 ;
  assign n21227 = ~n13358 & n21226 ;
  assign n21228 = ~n14232 & n21227 ;
  assign n21231 = n740 | n2610 ;
  assign n21232 = n21231 ^ n645 ^ 1'b0 ;
  assign n21233 = ( n4056 & n12627 ) | ( n4056 & n21232 ) | ( n12627 & n21232 ) ;
  assign n21229 = n12827 ^ n7824 ^ n7644 ;
  assign n21230 = n21229 ^ n18514 ^ n14810 ;
  assign n21234 = n21233 ^ n21230 ^ n5883 ;
  assign n21235 = n9248 ^ n3895 ^ 1'b0 ;
  assign n21236 = n21235 ^ n15441 ^ 1'b0 ;
  assign n21237 = n17515 ^ n5622 ^ n5361 ;
  assign n21238 = ( n9790 & ~n16298 ) | ( n9790 & n16914 ) | ( ~n16298 & n16914 ) ;
  assign n21239 = n8599 & n18025 ;
  assign n21240 = n21239 ^ n6578 ^ 1'b0 ;
  assign n21241 = ( n8615 & n11884 ) | ( n8615 & ~n12856 ) | ( n11884 & ~n12856 ) ;
  assign n21242 = n12752 & n21241 ;
  assign n21243 = ( n3725 & ~n4298 ) | ( n3725 & n4502 ) | ( ~n4298 & n4502 ) ;
  assign n21244 = n4924 | n21243 ;
  assign n21245 = ( n300 & n930 ) | ( n300 & n6640 ) | ( n930 & n6640 ) ;
  assign n21246 = n21245 ^ n19653 ^ n2258 ;
  assign n21247 = n21244 & ~n21246 ;
  assign n21248 = n21247 ^ n16155 ^ 1'b0 ;
  assign n21249 = ( n9701 & ~n10458 ) | ( n9701 & n19951 ) | ( ~n10458 & n19951 ) ;
  assign n21250 = ( n9644 & n21248 ) | ( n9644 & ~n21249 ) | ( n21248 & ~n21249 ) ;
  assign n21251 = ~n4659 & n20654 ;
  assign n21252 = n4330 & n8583 ;
  assign n21253 = ( ~n9443 & n11600 ) | ( ~n9443 & n12382 ) | ( n11600 & n12382 ) ;
  assign n21254 = ( ~n3606 & n15669 ) | ( ~n3606 & n16134 ) | ( n15669 & n16134 ) ;
  assign n21255 = ~n6584 & n8468 ;
  assign n21256 = n3814 & n21255 ;
  assign n21257 = ( n3580 & n8042 ) | ( n3580 & ~n21256 ) | ( n8042 & ~n21256 ) ;
  assign n21258 = n2830 ^ n1949 ^ 1'b0 ;
  assign n21259 = ~n21257 & n21258 ;
  assign n21260 = ( n2013 & n9976 ) | ( n2013 & n21259 ) | ( n9976 & n21259 ) ;
  assign n21261 = n8653 | n17275 ;
  assign n21262 = n21261 ^ n10343 ^ 1'b0 ;
  assign n21263 = n3840 | n9565 ;
  assign n21264 = n2167 | n21263 ;
  assign n21265 = n10099 & n21264 ;
  assign n21266 = ~n9247 & n21265 ;
  assign n21267 = ( n8203 & n16629 ) | ( n8203 & n20475 ) | ( n16629 & n20475 ) ;
  assign n21268 = n21267 ^ n16746 ^ n565 ;
  assign n21269 = n21268 ^ n18797 ^ 1'b0 ;
  assign n21271 = n6008 ^ n3439 ^ 1'b0 ;
  assign n21272 = ( ~n5756 & n17244 ) | ( ~n5756 & n21271 ) | ( n17244 & n21271 ) ;
  assign n21270 = n17506 ^ n16174 ^ n12719 ;
  assign n21273 = n21272 ^ n21270 ^ n14782 ;
  assign n21275 = n15930 ^ n9215 ^ n706 ;
  assign n21274 = n13981 ^ n9895 ^ n7531 ;
  assign n21276 = n21275 ^ n21274 ^ n4431 ;
  assign n21277 = n21276 ^ n20508 ^ n12976 ;
  assign n21278 = ( ~n2493 & n3195 ) | ( ~n2493 & n5313 ) | ( n3195 & n5313 ) ;
  assign n21279 = ~n5496 & n7297 ;
  assign n21280 = ~n1963 & n15435 ;
  assign n21281 = n21280 ^ n16557 ^ n15850 ;
  assign n21282 = ( n4077 & n4853 ) | ( n4077 & ~n14931 ) | ( n4853 & ~n14931 ) ;
  assign n21283 = n9481 ^ n6938 ^ 1'b0 ;
  assign n21284 = n21282 | n21283 ;
  assign n21285 = n12517 ^ n11297 ^ n3318 ;
  assign n21286 = n459 & n21285 ;
  assign n21287 = n21286 ^ n18522 ^ 1'b0 ;
  assign n21288 = n2388 | n7878 ;
  assign n21289 = n21288 ^ n7303 ^ 1'b0 ;
  assign n21290 = n1989 ^ n360 ^ 1'b0 ;
  assign n21291 = n14588 & ~n21290 ;
  assign n21292 = n21291 ^ n503 ^ 1'b0 ;
  assign n21293 = n13802 | n21292 ;
  assign n21294 = n18693 | n21293 ;
  assign n21295 = n17374 ^ n14486 ^ n1441 ;
  assign n21296 = n1834 | n16438 ;
  assign n21298 = n854 | n5429 ;
  assign n21299 = x2 | n21298 ;
  assign n21300 = n21299 ^ n4984 ^ n4511 ;
  assign n21297 = n476 & ~n8231 ;
  assign n21301 = n21300 ^ n21297 ^ 1'b0 ;
  assign n21302 = n14149 | n14196 ;
  assign n21303 = ~n21301 & n21302 ;
  assign n21304 = n21303 ^ n9947 ^ 1'b0 ;
  assign n21305 = n18442 & n19910 ;
  assign n21306 = n1391 & ~n3174 ;
  assign n21307 = ( n2922 & n21305 ) | ( n2922 & ~n21306 ) | ( n21305 & ~n21306 ) ;
  assign n21308 = n14239 & ~n21307 ;
  assign n21309 = n21308 ^ n1829 ^ 1'b0 ;
  assign n21310 = ( n1032 & n1869 ) | ( n1032 & n18864 ) | ( n1869 & n18864 ) ;
  assign n21311 = n16152 | n21310 ;
  assign n21312 = n4721 ^ n4575 ^ n3941 ;
  assign n21313 = n21312 ^ n8828 ^ n5701 ;
  assign n21314 = n21313 ^ n9076 ^ n5438 ;
  assign n21315 = n6973 & n15827 ;
  assign n21316 = ~n11638 & n21315 ;
  assign n21317 = n8914 ^ n8653 ^ n8085 ;
  assign n21318 = n14408 & ~n21317 ;
  assign n21319 = ( n7127 & n21316 ) | ( n7127 & n21318 ) | ( n21316 & n21318 ) ;
  assign n21320 = ( n13660 & ~n16059 ) | ( n13660 & n17221 ) | ( ~n16059 & n17221 ) ;
  assign n21321 = ( ~n4652 & n6762 ) | ( ~n4652 & n21320 ) | ( n6762 & n21320 ) ;
  assign n21322 = n14474 ^ n6441 ^ n310 ;
  assign n21323 = n2239 ^ n1868 ^ 1'b0 ;
  assign n21324 = n7377 & n21323 ;
  assign n21325 = n2068 & n21324 ;
  assign n21326 = n8935 | n19585 ;
  assign n21327 = ( n4488 & ~n17979 ) | ( n4488 & n21326 ) | ( ~n17979 & n21326 ) ;
  assign n21331 = n3887 ^ n3444 ^ 1'b0 ;
  assign n21330 = ( n7621 & ~n8081 ) | ( n7621 & n11705 ) | ( ~n8081 & n11705 ) ;
  assign n21328 = n12912 ^ n10722 ^ 1'b0 ;
  assign n21329 = n3442 & ~n21328 ;
  assign n21332 = n21331 ^ n21330 ^ n21329 ;
  assign n21333 = n20155 ^ n7763 ^ 1'b0 ;
  assign n21334 = n4447 ^ n3679 ^ n365 ;
  assign n21335 = n1544 ^ n584 ^ 1'b0 ;
  assign n21336 = ~n1141 & n21335 ;
  assign n21337 = ( n11915 & ~n21334 ) | ( n11915 & n21336 ) | ( ~n21334 & n21336 ) ;
  assign n21338 = n14379 ^ n9905 ^ n639 ;
  assign n21339 = n13594 & ~n21338 ;
  assign n21340 = n21339 ^ n19715 ^ 1'b0 ;
  assign n21341 = n6561 ^ n2043 ^ 1'b0 ;
  assign n21342 = n13544 & ~n21341 ;
  assign n21343 = ~n12553 & n21342 ;
  assign n21344 = n6630 & ~n6935 ;
  assign n21345 = n9561 & n21344 ;
  assign n21346 = n13942 ^ n607 ^ 1'b0 ;
  assign n21347 = n4979 | n21346 ;
  assign n21348 = n9685 | n12082 ;
  assign n21349 = n8401 | n21348 ;
  assign n21350 = ~n9291 & n19492 ;
  assign n21351 = ( n6576 & ~n21349 ) | ( n6576 & n21350 ) | ( ~n21349 & n21350 ) ;
  assign n21357 = n5900 & ~n13830 ;
  assign n21353 = n8362 ^ n2587 ^ n880 ;
  assign n21354 = n21353 ^ n5833 ^ 1'b0 ;
  assign n21355 = n6601 | n21354 ;
  assign n21352 = n6987 | n21274 ;
  assign n21356 = n21355 ^ n21352 ^ 1'b0 ;
  assign n21358 = n21357 ^ n21356 ^ n315 ;
  assign n21363 = n15204 & ~n19903 ;
  assign n21359 = n8399 ^ n6552 ^ n3725 ;
  assign n21360 = n21359 ^ n21229 ^ n9723 ;
  assign n21361 = ~n2837 & n21360 ;
  assign n21362 = ~n3910 & n21361 ;
  assign n21364 = n21363 ^ n21362 ^ 1'b0 ;
  assign n21365 = ( n1430 & n16262 ) | ( n1430 & n21191 ) | ( n16262 & n21191 ) ;
  assign n21366 = n9752 | n13148 ;
  assign n21367 = n21366 ^ n20117 ^ 1'b0 ;
  assign n21368 = n10438 | n21367 ;
  assign n21369 = n21368 ^ n15133 ^ 1'b0 ;
  assign n21370 = n13692 ^ n1258 ^ n766 ;
  assign n21371 = n187 & ~n21370 ;
  assign n21372 = ( n4771 & n5667 ) | ( n4771 & ~n21371 ) | ( n5667 & ~n21371 ) ;
  assign n21373 = n19747 ^ n5133 ^ n2915 ;
  assign n21374 = n21229 ^ n10557 ^ n8620 ;
  assign n21375 = ( n17686 & ~n20426 ) | ( n17686 & n21374 ) | ( ~n20426 & n21374 ) ;
  assign n21376 = n19068 ^ n6194 ^ 1'b0 ;
  assign n21377 = ( n7641 & n13365 ) | ( n7641 & ~n21376 ) | ( n13365 & ~n21376 ) ;
  assign n21378 = n13447 ^ n11778 ^ 1'b0 ;
  assign n21379 = ~n16565 & n21378 ;
  assign n21380 = n7049 & n8396 ;
  assign n21381 = n21380 ^ n2414 ^ 1'b0 ;
  assign n21382 = n9177 ^ n4007 ^ n2145 ;
  assign n21383 = ( n1413 & ~n15159 ) | ( n1413 & n21382 ) | ( ~n15159 & n21382 ) ;
  assign n21384 = n18972 & n21383 ;
  assign n21385 = n21384 ^ n2957 ^ 1'b0 ;
  assign n21386 = ~n8903 & n15811 ;
  assign n21387 = ( n10624 & n20327 ) | ( n10624 & ~n21386 ) | ( n20327 & ~n21386 ) ;
  assign n21388 = n16944 ^ n12352 ^ n761 ;
  assign n21389 = n21388 ^ n7584 ^ 1'b0 ;
  assign n21390 = n4899 ^ n1119 ^ 1'b0 ;
  assign n21391 = ~n1527 & n21390 ;
  assign n21392 = n21391 ^ n6809 ^ n1409 ;
  assign n21393 = n1517 | n7607 ;
  assign n21394 = ( n494 & n4886 ) | ( n494 & ~n17605 ) | ( n4886 & ~n17605 ) ;
  assign n21395 = ( n5452 & n21393 ) | ( n5452 & ~n21394 ) | ( n21393 & ~n21394 ) ;
  assign n21396 = ~n448 & n18157 ;
  assign n21397 = n21396 ^ n954 ^ 1'b0 ;
  assign n21398 = n3062 & n10131 ;
  assign n21399 = n10411 ^ n4306 ^ 1'b0 ;
  assign n21400 = n21398 & n21399 ;
  assign n21401 = ( x27 & n3096 ) | ( x27 & n7523 ) | ( n3096 & n7523 ) ;
  assign n21402 = ( ~n5074 & n13293 ) | ( ~n5074 & n14815 ) | ( n13293 & n14815 ) ;
  assign n21403 = ( ~n6975 & n18829 ) | ( ~n6975 & n21402 ) | ( n18829 & n21402 ) ;
  assign n21404 = ~n9554 & n19448 ;
  assign n21405 = n14601 ^ n11204 ^ n4990 ;
  assign n21406 = ( n3347 & ~n21404 ) | ( n3347 & n21405 ) | ( ~n21404 & n21405 ) ;
  assign n21407 = ( ~n3271 & n7473 ) | ( ~n3271 & n14798 ) | ( n7473 & n14798 ) ;
  assign n21408 = ( n741 & n8953 ) | ( n741 & n21407 ) | ( n8953 & n21407 ) ;
  assign n21409 = n5632 & n21408 ;
  assign n21410 = n13457 & n21409 ;
  assign n21411 = n2118 & ~n6893 ;
  assign n21412 = n1165 & n6023 ;
  assign n21413 = n21412 ^ n1893 ^ 1'b0 ;
  assign n21414 = n8900 | n21127 ;
  assign n21415 = n11985 & ~n15806 ;
  assign n21416 = ( n4191 & ~n9906 ) | ( n4191 & n21415 ) | ( ~n9906 & n21415 ) ;
  assign n21417 = n6081 | n11701 ;
  assign n21418 = n11304 | n21417 ;
  assign n21419 = ( n5421 & n6479 ) | ( n5421 & n21418 ) | ( n6479 & n21418 ) ;
  assign n21420 = ( n1362 & n3286 ) | ( n1362 & n3822 ) | ( n3286 & n3822 ) ;
  assign n21421 = ( ~n2050 & n6020 ) | ( ~n2050 & n11089 ) | ( n6020 & n11089 ) ;
  assign n21422 = n21085 ^ n13462 ^ n10221 ;
  assign n21423 = ( n21420 & n21421 ) | ( n21420 & ~n21422 ) | ( n21421 & ~n21422 ) ;
  assign n21424 = ( n5543 & n7912 ) | ( n5543 & n20478 ) | ( n7912 & n20478 ) ;
  assign n21430 = n9323 ^ n9070 ^ 1'b0 ;
  assign n21428 = ( ~n3087 & n4839 ) | ( ~n3087 & n5557 ) | ( n4839 & n5557 ) ;
  assign n21427 = n3348 | n16711 ;
  assign n21429 = n21428 ^ n21427 ^ x78 ;
  assign n21425 = ( ~n1203 & n4265 ) | ( ~n1203 & n11947 ) | ( n4265 & n11947 ) ;
  assign n21426 = n21425 ^ n5658 ^ n5071 ;
  assign n21431 = n21430 ^ n21429 ^ n21426 ;
  assign n21432 = n709 & ~n1741 ;
  assign n21433 = n21431 & n21432 ;
  assign n21434 = n4724 | n10381 ;
  assign n21435 = n12287 ^ n1591 ^ 1'b0 ;
  assign n21436 = ~n10845 & n21435 ;
  assign n21437 = n10916 ^ n9006 ^ n789 ;
  assign n21438 = n21436 & n21437 ;
  assign n21439 = n21438 ^ n12242 ^ 1'b0 ;
  assign n21440 = ( n1633 & n10459 ) | ( n1633 & n21026 ) | ( n10459 & n21026 ) ;
  assign n21441 = n4565 ^ n3234 ^ n3166 ;
  assign n21442 = n12243 ^ n1563 ^ n372 ;
  assign n21443 = n21442 ^ n7632 ^ n2434 ;
  assign n21444 = ( ~n2216 & n9909 ) | ( ~n2216 & n13425 ) | ( n9909 & n13425 ) ;
  assign n21445 = ( n21441 & ~n21443 ) | ( n21441 & n21444 ) | ( ~n21443 & n21444 ) ;
  assign n21446 = ( n1561 & ~n3568 ) | ( n1561 & n21445 ) | ( ~n3568 & n21445 ) ;
  assign n21448 = n8943 ^ n1021 ^ n901 ;
  assign n21447 = n3929 & ~n4358 ;
  assign n21449 = n21448 ^ n21447 ^ 1'b0 ;
  assign n21450 = ( ~n510 & n4120 ) | ( ~n510 & n13134 ) | ( n4120 & n13134 ) ;
  assign n21451 = ( n1194 & n7229 ) | ( n1194 & n14927 ) | ( n7229 & n14927 ) ;
  assign n21455 = ( n2820 & n5864 ) | ( n2820 & n10303 ) | ( n5864 & n10303 ) ;
  assign n21454 = ~n5477 & n15133 ;
  assign n21452 = ( n1186 & n4641 ) | ( n1186 & ~n9850 ) | ( n4641 & ~n9850 ) ;
  assign n21453 = n21452 ^ n12595 ^ n421 ;
  assign n21456 = n21455 ^ n21454 ^ n21453 ;
  assign n21457 = n14887 | n21456 ;
  assign n21458 = n17662 ^ n6764 ^ 1'b0 ;
  assign n21459 = ~n4810 & n21458 ;
  assign n21460 = n8679 ^ n5527 ^ n609 ;
  assign n21461 = n13419 ^ n5826 ^ n4179 ;
  assign n21462 = ( n15349 & n21460 ) | ( n15349 & ~n21461 ) | ( n21460 & ~n21461 ) ;
  assign n21463 = n3762 ^ n572 ^ 1'b0 ;
  assign n21464 = n586 & ~n21463 ;
  assign n21465 = n21464 ^ n16567 ^ 1'b0 ;
  assign n21466 = n8537 | n20280 ;
  assign n21467 = n21465 | n21466 ;
  assign n21468 = n21467 ^ n20583 ^ n9480 ;
  assign n21469 = n1637 | n14184 ;
  assign n21470 = ( n3526 & n6734 ) | ( n3526 & n8531 ) | ( n6734 & n8531 ) ;
  assign n21471 = n15063 | n21470 ;
  assign n21472 = n11525 | n21471 ;
  assign n21477 = n21170 ^ n13630 ^ 1'b0 ;
  assign n21473 = n11810 & n12032 ;
  assign n21474 = n4532 & n21473 ;
  assign n21475 = ( n6371 & n10272 ) | ( n6371 & ~n21474 ) | ( n10272 & ~n21474 ) ;
  assign n21476 = n21475 ^ n17917 ^ 1'b0 ;
  assign n21478 = n21477 ^ n21476 ^ 1'b0 ;
  assign n21479 = ( n4296 & n9163 ) | ( n4296 & n21478 ) | ( n9163 & n21478 ) ;
  assign n21480 = ( n12008 & n21472 ) | ( n12008 & n21479 ) | ( n21472 & n21479 ) ;
  assign n21481 = n14304 ^ n8021 ^ 1'b0 ;
  assign n21482 = ~n20991 & n21481 ;
  assign n21483 = ( n1184 & n2080 ) | ( n1184 & n9688 ) | ( n2080 & n9688 ) ;
  assign n21484 = n2159 & n9549 ;
  assign n21485 = ~n8641 & n21484 ;
  assign n21486 = ( n2364 & n3117 ) | ( n2364 & n4777 ) | ( n3117 & n4777 ) ;
  assign n21487 = n6828 ^ n3821 ^ n2375 ;
  assign n21488 = ~n10195 & n11829 ;
  assign n21489 = n21488 ^ n308 ^ 1'b0 ;
  assign n21490 = n21489 ^ n6253 ^ n2313 ;
  assign n21491 = ( n21486 & n21487 ) | ( n21486 & n21490 ) | ( n21487 & n21490 ) ;
  assign n21492 = ( n2490 & n8992 ) | ( n2490 & n16277 ) | ( n8992 & n16277 ) ;
  assign n21493 = ( n7760 & n9355 ) | ( n7760 & n10792 ) | ( n9355 & n10792 ) ;
  assign n21494 = n15225 ^ n9302 ^ 1'b0 ;
  assign n21495 = n12226 & n21494 ;
  assign n21496 = n19368 ^ n16720 ^ 1'b0 ;
  assign n21497 = n10469 ^ n10381 ^ n2957 ;
  assign n21498 = n21497 ^ n10422 ^ n8619 ;
  assign n21499 = n4302 & ~n5927 ;
  assign n21500 = ( ~n4179 & n5312 ) | ( ~n4179 & n21499 ) | ( n5312 & n21499 ) ;
  assign n21501 = n21500 ^ n5321 ^ n4739 ;
  assign n21502 = n12860 ^ n8393 ^ n3214 ;
  assign n21503 = n21501 | n21502 ;
  assign n21504 = n21503 ^ n11982 ^ 1'b0 ;
  assign n21505 = ( n5265 & ~n11867 ) | ( n5265 & n14408 ) | ( ~n11867 & n14408 ) ;
  assign n21506 = n21504 & n21505 ;
  assign n21507 = n11974 & n13269 ;
  assign n21508 = n21507 ^ n14910 ^ 1'b0 ;
  assign n21509 = n21508 ^ n19260 ^ n7106 ;
  assign n21510 = n2664 | n21155 ;
  assign n21511 = n21036 ^ n2524 ^ 1'b0 ;
  assign n21512 = n10619 ^ n9255 ^ 1'b0 ;
  assign n21513 = n21511 & n21512 ;
  assign n21514 = ~n17780 & n21513 ;
  assign n21515 = ~n3410 & n21514 ;
  assign n21516 = n13809 ^ n11635 ^ n6854 ;
  assign n21517 = n1162 & ~n18881 ;
  assign n21518 = ( n3460 & n14716 ) | ( n3460 & ~n21517 ) | ( n14716 & ~n21517 ) ;
  assign n21519 = ( ~x76 & n12328 ) | ( ~x76 & n21028 ) | ( n12328 & n21028 ) ;
  assign n21520 = ( n1152 & ~n21518 ) | ( n1152 & n21519 ) | ( ~n21518 & n21519 ) ;
  assign n21521 = n18938 ^ n5240 ^ n4490 ;
  assign n21522 = n21521 ^ n9473 ^ n6497 ;
  assign n21523 = n3769 ^ n3699 ^ 1'b0 ;
  assign n21524 = ( n6809 & n9894 ) | ( n6809 & ~n21523 ) | ( n9894 & ~n21523 ) ;
  assign n21525 = n5405 & n20169 ;
  assign n21526 = n15825 & n21525 ;
  assign n21527 = n1620 & ~n11957 ;
  assign n21528 = n21527 ^ n3747 ^ 1'b0 ;
  assign n21529 = n648 & n12539 ;
  assign n21530 = n21529 ^ n17088 ^ 1'b0 ;
  assign n21531 = n21530 ^ n19375 ^ n15754 ;
  assign n21532 = ( n7217 & n9608 ) | ( n7217 & n15049 ) | ( n9608 & n15049 ) ;
  assign n21533 = n4964 ^ n1059 ^ 1'b0 ;
  assign n21534 = n21532 | n21533 ;
  assign n21535 = n21534 ^ n16865 ^ n5805 ;
  assign n21536 = n21535 ^ n12501 ^ n7193 ;
  assign n21537 = n2517 & ~n3868 ;
  assign n21538 = n21537 ^ n12622 ^ 1'b0 ;
  assign n21539 = n7735 ^ n3495 ^ n3337 ;
  assign n21540 = n21539 ^ n8973 ^ n2482 ;
  assign n21541 = ~n9209 & n21540 ;
  assign n21542 = n4676 & n21541 ;
  assign n21543 = n16673 ^ n7816 ^ n6599 ;
  assign n21544 = n21543 ^ n14620 ^ n8448 ;
  assign n21545 = n21544 ^ n19259 ^ n1920 ;
  assign n21547 = n3212 | n11739 ;
  assign n21548 = n12105 | n21547 ;
  assign n21546 = n20340 ^ n15628 ^ n2145 ;
  assign n21549 = n21548 ^ n21546 ^ n10161 ;
  assign n21550 = ~n6358 & n9678 ;
  assign n21551 = n21550 ^ n11902 ^ n1685 ;
  assign n21552 = n16914 & n21551 ;
  assign n21553 = n4202 | n5551 ;
  assign n21554 = n21553 ^ n5061 ^ 1'b0 ;
  assign n21555 = ( n3630 & n6116 ) | ( n3630 & ~n21554 ) | ( n6116 & ~n21554 ) ;
  assign n21557 = ~n2760 & n11827 ;
  assign n21558 = n21557 ^ n2937 ^ 1'b0 ;
  assign n21556 = n21499 ^ n10993 ^ 1'b0 ;
  assign n21559 = n21558 ^ n21556 ^ n319 ;
  assign n21560 = n1051 | n1608 ;
  assign n21561 = ( n1354 & n19705 ) | ( n1354 & ~n21560 ) | ( n19705 & ~n21560 ) ;
  assign n21562 = n13752 & ~n17588 ;
  assign n21563 = ( n17098 & ~n21320 ) | ( n17098 & n21562 ) | ( ~n21320 & n21562 ) ;
  assign n21564 = ( n2602 & n5321 ) | ( n2602 & n20955 ) | ( n5321 & n20955 ) ;
  assign n21565 = n9442 & ~n17404 ;
  assign n21566 = n21565 ^ n4597 ^ 1'b0 ;
  assign n21567 = ( n2024 & n17616 ) | ( n2024 & n19465 ) | ( n17616 & n19465 ) ;
  assign n21568 = n17231 & n21567 ;
  assign n21569 = n6867 & n21568 ;
  assign n21573 = n19374 ^ n9176 ^ 1'b0 ;
  assign n21570 = n10094 ^ n8024 ^ 1'b0 ;
  assign n21571 = ~n10402 & n21570 ;
  assign n21572 = n21571 ^ n16596 ^ 1'b0 ;
  assign n21574 = n21573 ^ n21572 ^ 1'b0 ;
  assign n21575 = n16125 ^ n10001 ^ 1'b0 ;
  assign n21576 = n6135 & ~n21575 ;
  assign n21577 = ~n9907 & n21576 ;
  assign n21578 = n2035 & n21577 ;
  assign n21579 = n21578 ^ n18594 ^ n856 ;
  assign n21580 = ( ~n222 & n1634 ) | ( ~n222 & n4730 ) | ( n1634 & n4730 ) ;
  assign n21581 = n11623 ^ n2317 ^ 1'b0 ;
  assign n21582 = ( n1216 & n6420 ) | ( n1216 & n15848 ) | ( n6420 & n15848 ) ;
  assign n21583 = ( ~n5195 & n9659 ) | ( ~n5195 & n20810 ) | ( n9659 & n20810 ) ;
  assign n21584 = n6397 | n21583 ;
  assign n21585 = n21582 & ~n21584 ;
  assign n21586 = n15363 & ~n18907 ;
  assign n21587 = ~n5071 & n21586 ;
  assign n21588 = n8413 | n14606 ;
  assign n21589 = n2801 | n21588 ;
  assign n21593 = n3039 & ~n8082 ;
  assign n21592 = n15099 ^ n10534 ^ 1'b0 ;
  assign n21594 = n21593 ^ n21592 ^ n15969 ;
  assign n21595 = n7106 | n21594 ;
  assign n21590 = n21207 ^ n18018 ^ n5328 ;
  assign n21591 = n5703 & n21590 ;
  assign n21596 = n21595 ^ n21591 ^ 1'b0 ;
  assign n21597 = n699 & n3840 ;
  assign n21598 = n1361 | n2671 ;
  assign n21599 = n21598 ^ n4857 ^ 1'b0 ;
  assign n21600 = n21597 | n21599 ;
  assign n21601 = ( n2267 & ~n5307 ) | ( n2267 & n21600 ) | ( ~n5307 & n21600 ) ;
  assign n21602 = ~n6344 & n8763 ;
  assign n21603 = n12500 & n21602 ;
  assign n21604 = n21603 ^ n13040 ^ x29 ;
  assign n21605 = n5618 ^ n5525 ^ n4555 ;
  assign n21607 = ( n3871 & n4193 ) | ( n3871 & ~n12412 ) | ( n4193 & ~n12412 ) ;
  assign n21608 = n1268 | n21607 ;
  assign n21606 = n3689 | n4476 ;
  assign n21609 = n21608 ^ n21606 ^ 1'b0 ;
  assign n21611 = n533 | n6550 ;
  assign n21612 = n21611 ^ n3049 ^ 1'b0 ;
  assign n21613 = ( n1735 & ~n6213 ) | ( n1735 & n21612 ) | ( ~n6213 & n21612 ) ;
  assign n21610 = n4864 | n16198 ;
  assign n21614 = n21613 ^ n21610 ^ n5849 ;
  assign n21617 = n1062 | n6816 ;
  assign n21618 = n6927 & ~n21617 ;
  assign n21619 = n21618 ^ n6263 ^ 1'b0 ;
  assign n21615 = x74 & ~n5449 ;
  assign n21616 = n21615 ^ n9812 ^ 1'b0 ;
  assign n21620 = n21619 ^ n21616 ^ n5731 ;
  assign n21621 = n2780 ^ n1780 ^ n928 ;
  assign n21622 = n21621 ^ n798 ^ 1'b0 ;
  assign n21623 = n7088 | n21622 ;
  assign n21624 = n21620 & ~n21623 ;
  assign n21625 = n21624 ^ n8500 ^ 1'b0 ;
  assign n21626 = ( n1259 & n1668 ) | ( n1259 & n5915 ) | ( n1668 & n5915 ) ;
  assign n21627 = ( n13952 & n17397 ) | ( n13952 & n21626 ) | ( n17397 & n21626 ) ;
  assign n21628 = n16257 | n21627 ;
  assign n21629 = n11136 & ~n13952 ;
  assign n21630 = n21629 ^ n8045 ^ 1'b0 ;
  assign n21631 = n5180 ^ n2771 ^ n218 ;
  assign n21632 = n20108 & ~n21631 ;
  assign n21633 = n21632 ^ n21359 ^ 1'b0 ;
  assign n21634 = n12918 & n21633 ;
  assign n21635 = ( n2238 & n7209 ) | ( n2238 & ~n9462 ) | ( n7209 & ~n9462 ) ;
  assign n21636 = ( ~n1529 & n16895 ) | ( ~n1529 & n21635 ) | ( n16895 & n21635 ) ;
  assign n21637 = ( n2356 & n5453 ) | ( n2356 & n11929 ) | ( n5453 & n11929 ) ;
  assign n21638 = ( n16150 & ~n20985 ) | ( n16150 & n21026 ) | ( ~n20985 & n21026 ) ;
  assign n21639 = ( n1046 & n10176 ) | ( n1046 & n19232 ) | ( n10176 & n19232 ) ;
  assign n21640 = n2852 & n19155 ;
  assign n21641 = ~n21639 & n21640 ;
  assign n21642 = n12742 | n21641 ;
  assign n21643 = ( n917 & n21638 ) | ( n917 & n21642 ) | ( n21638 & n21642 ) ;
  assign n21644 = ( ~n2283 & n12825 ) | ( ~n2283 & n21643 ) | ( n12825 & n21643 ) ;
  assign n21645 = ( n1973 & ~n16429 ) | ( n1973 & n19088 ) | ( ~n16429 & n19088 ) ;
  assign n21646 = n17336 ^ n13518 ^ 1'b0 ;
  assign n21647 = n13176 & ~n21646 ;
  assign n21648 = ( n8313 & n8585 ) | ( n8313 & ~n9898 ) | ( n8585 & ~n9898 ) ;
  assign n21649 = n17391 ^ n4756 ^ 1'b0 ;
  assign n21650 = n21648 & n21649 ;
  assign n21651 = ( n1476 & n1618 ) | ( n1476 & n15520 ) | ( n1618 & n15520 ) ;
  assign n21652 = ( n15166 & ~n19924 ) | ( n15166 & n21651 ) | ( ~n19924 & n21651 ) ;
  assign n21653 = ( n3805 & n12226 ) | ( n3805 & n18214 ) | ( n12226 & n18214 ) ;
  assign n21654 = n21653 ^ n9432 ^ n5245 ;
  assign n21655 = ( n135 & n21652 ) | ( n135 & n21654 ) | ( n21652 & n21654 ) ;
  assign n21658 = ( ~n1001 & n5360 ) | ( ~n1001 & n11328 ) | ( n5360 & n11328 ) ;
  assign n21656 = n4681 ^ n3603 ^ 1'b0 ;
  assign n21657 = n21656 ^ n16654 ^ n9541 ;
  assign n21659 = n21658 ^ n21657 ^ n21560 ;
  assign n21660 = n13352 ^ n11834 ^ n7953 ;
  assign n21663 = ( n1518 & n5136 ) | ( n1518 & ~n6310 ) | ( n5136 & ~n6310 ) ;
  assign n21664 = n1459 & n21663 ;
  assign n21665 = ~n1186 & n21664 ;
  assign n21661 = n389 & n2665 ;
  assign n21662 = ~n14388 & n21661 ;
  assign n21666 = n21665 ^ n21662 ^ n15272 ;
  assign n21667 = n5864 ^ n3901 ^ n3330 ;
  assign n21668 = n21667 ^ n12851 ^ n11883 ;
  assign n21669 = ( n6086 & n15166 ) | ( n6086 & ~n19036 ) | ( n15166 & ~n19036 ) ;
  assign n21670 = n15949 & n21669 ;
  assign n21671 = n21670 ^ n20080 ^ 1'b0 ;
  assign n21672 = x50 & ~n14769 ;
  assign n21673 = n3742 & n21672 ;
  assign n21674 = n13896 ^ n665 ^ 1'b0 ;
  assign n21675 = ~n21673 & n21674 ;
  assign n21676 = n4504 ^ n4164 ^ n1779 ;
  assign n21677 = n21676 ^ n20091 ^ n8500 ;
  assign n21678 = ( n6457 & ~n11134 ) | ( n6457 & n11392 ) | ( ~n11134 & n11392 ) ;
  assign n21679 = n21678 ^ n16800 ^ 1'b0 ;
  assign n21680 = n7951 | n21679 ;
  assign n21681 = ( n3598 & ~n21677 ) | ( n3598 & n21680 ) | ( ~n21677 & n21680 ) ;
  assign n21682 = n18652 ^ n16543 ^ n4798 ;
  assign n21683 = ( ~n1955 & n10616 ) | ( ~n1955 & n12613 ) | ( n10616 & n12613 ) ;
  assign n21684 = ( n2439 & n6543 ) | ( n2439 & n21683 ) | ( n6543 & n21683 ) ;
  assign n21686 = n5784 | n7758 ;
  assign n21687 = n5525 & ~n21686 ;
  assign n21685 = ~n5437 & n9153 ;
  assign n21688 = n21687 ^ n21685 ^ 1'b0 ;
  assign n21689 = n4357 & ~n5438 ;
  assign n21690 = n21689 ^ n4593 ^ 1'b0 ;
  assign n21691 = ( n6997 & n21688 ) | ( n6997 & n21690 ) | ( n21688 & n21690 ) ;
  assign n21692 = n1885 & n8914 ;
  assign n21693 = n3052 & n21692 ;
  assign n21694 = n1779 & n19101 ;
  assign n21695 = ~n398 & n21694 ;
  assign n21696 = ( ~n204 & n2214 ) | ( ~n204 & n21695 ) | ( n2214 & n21695 ) ;
  assign n21697 = ( n6645 & n15504 ) | ( n6645 & n20669 ) | ( n15504 & n20669 ) ;
  assign n21698 = n20827 ^ n926 ^ 1'b0 ;
  assign n21699 = ~n5509 & n21698 ;
  assign n21700 = n21018 ^ n7814 ^ n1702 ;
  assign n21701 = n7560 & n21700 ;
  assign n21702 = n17174 | n21701 ;
  assign n21703 = n6505 | n21702 ;
  assign n21704 = n15603 ^ n13876 ^ n2188 ;
  assign n21705 = ( n5783 & n21703 ) | ( n5783 & n21704 ) | ( n21703 & n21704 ) ;
  assign n21706 = n12105 ^ n4640 ^ n4344 ;
  assign n21707 = n21706 ^ n18063 ^ n9190 ;
  assign n21708 = ( n7092 & n16339 ) | ( n7092 & n20299 ) | ( n16339 & n20299 ) ;
  assign n21709 = n2670 & n21708 ;
  assign n21711 = ( n573 & n4353 ) | ( n573 & ~n9301 ) | ( n4353 & ~n9301 ) ;
  assign n21710 = n15824 ^ n4442 ^ 1'b0 ;
  assign n21712 = n21711 ^ n21710 ^ n14113 ;
  assign n21713 = n2151 ^ n1924 ^ n1302 ;
  assign n21714 = n1531 & n21713 ;
  assign n21715 = ~n1291 & n21714 ;
  assign n21717 = n2439 ^ n409 ^ 1'b0 ;
  assign n21718 = n4088 | n21717 ;
  assign n21719 = n21718 ^ n18511 ^ n4562 ;
  assign n21716 = n5931 & n9509 ;
  assign n21720 = n21719 ^ n21716 ^ 1'b0 ;
  assign n21721 = ( n5613 & n6971 ) | ( n5613 & ~n21720 ) | ( n6971 & ~n21720 ) ;
  assign n21722 = ( n21712 & n21715 ) | ( n21712 & ~n21721 ) | ( n21715 & ~n21721 ) ;
  assign n21723 = n7867 & ~n21722 ;
  assign n21724 = n14044 ^ n4517 ^ 1'b0 ;
  assign n21725 = ( ~n5646 & n14582 ) | ( ~n5646 & n21724 ) | ( n14582 & n21724 ) ;
  assign n21726 = n17513 | n18726 ;
  assign n21727 = n9713 & ~n21726 ;
  assign n21728 = n10413 ^ n3093 ^ n1238 ;
  assign n21729 = ~n18503 & n21728 ;
  assign n21730 = n6977 ^ n3384 ^ n2614 ;
  assign n21731 = n19253 ^ n13358 ^ n3140 ;
  assign n21732 = n16503 ^ n818 ^ 1'b0 ;
  assign n21733 = ~n21731 & n21732 ;
  assign n21734 = n16561 | n21733 ;
  assign n21735 = ( n12284 & n17825 ) | ( n12284 & n21734 ) | ( n17825 & n21734 ) ;
  assign n21738 = n17961 ^ n15691 ^ n15578 ;
  assign n21736 = n3395 ^ n3205 ^ 1'b0 ;
  assign n21737 = n21736 ^ n3169 ^ 1'b0 ;
  assign n21739 = n21738 ^ n21737 ^ n3049 ;
  assign n21740 = ( n11797 & ~n13184 ) | ( n11797 & n13256 ) | ( ~n13184 & n13256 ) ;
  assign n21741 = ( n6675 & n11414 ) | ( n6675 & ~n11454 ) | ( n11414 & ~n11454 ) ;
  assign n21742 = n21741 ^ n9077 ^ n7198 ;
  assign n21743 = n21742 ^ n9354 ^ n4943 ;
  assign n21744 = n10412 ^ n280 ^ 1'b0 ;
  assign n21745 = n6142 & ~n21744 ;
  assign n21746 = ~n12185 & n21745 ;
  assign n21747 = n21743 & n21746 ;
  assign n21748 = ~n4614 & n11129 ;
  assign n21749 = n21748 ^ n12700 ^ 1'b0 ;
  assign n21750 = n9180 & ~n19768 ;
  assign n21751 = n14912 ^ n8781 ^ n6032 ;
  assign n21752 = ( n8324 & ~n21750 ) | ( n8324 & n21751 ) | ( ~n21750 & n21751 ) ;
  assign n21756 = n8864 ^ n2943 ^ n1871 ;
  assign n21757 = ( n8485 & n8546 ) | ( n8485 & n21756 ) | ( n8546 & n21756 ) ;
  assign n21753 = n3853 | n5020 ;
  assign n21754 = n13622 ^ n2220 ^ 1'b0 ;
  assign n21755 = n21753 & n21754 ;
  assign n21758 = n21757 ^ n21755 ^ n4221 ;
  assign n21759 = n5915 ^ n2503 ^ 1'b0 ;
  assign n21760 = n16676 ^ n7148 ^ 1'b0 ;
  assign n21762 = ~n3417 & n7400 ;
  assign n21763 = n21762 ^ n15626 ^ 1'b0 ;
  assign n21761 = n17431 ^ n16214 ^ 1'b0 ;
  assign n21764 = n21763 ^ n21761 ^ n10140 ;
  assign n21765 = n12427 ^ n3011 ^ n2989 ;
  assign n21766 = n2678 | n5103 ;
  assign n21767 = n21766 ^ n329 ^ 1'b0 ;
  assign n21768 = ( n9607 & n21765 ) | ( n9607 & n21767 ) | ( n21765 & n21767 ) ;
  assign n21769 = ( n5857 & n15568 ) | ( n5857 & n21768 ) | ( n15568 & n21768 ) ;
  assign n21770 = n10626 ^ n5917 ^ n5233 ;
  assign n21773 = ~n5910 & n6034 ;
  assign n21774 = n9382 & n21773 ;
  assign n21775 = n21774 ^ n1228 ^ 1'b0 ;
  assign n21776 = ~n2578 & n21775 ;
  assign n21771 = n20234 ^ n14287 ^ n5235 ;
  assign n21772 = n3284 | n21771 ;
  assign n21777 = n21776 ^ n21772 ^ n2896 ;
  assign n21778 = n21770 & n21777 ;
  assign n21779 = n16165 | n21778 ;
  assign n21780 = ( n4581 & n13700 ) | ( n4581 & ~n17323 ) | ( n13700 & ~n17323 ) ;
  assign n21781 = n1621 & ~n21780 ;
  assign n21782 = n21781 ^ n7507 ^ 1'b0 ;
  assign n21792 = n2981 ^ n2452 ^ 1'b0 ;
  assign n21790 = ( n3049 & n10421 ) | ( n3049 & n16932 ) | ( n10421 & n16932 ) ;
  assign n21791 = n15167 & ~n21790 ;
  assign n21793 = n21792 ^ n21791 ^ 1'b0 ;
  assign n21783 = n7552 ^ n7352 ^ n2338 ;
  assign n21784 = n21783 ^ n436 ^ 1'b0 ;
  assign n21785 = n2914 & ~n21784 ;
  assign n21786 = ( ~n4991 & n10855 ) | ( ~n4991 & n21785 ) | ( n10855 & n21785 ) ;
  assign n21787 = n10212 | n20730 ;
  assign n21788 = n19692 & ~n21787 ;
  assign n21789 = ( n4100 & n21786 ) | ( n4100 & n21788 ) | ( n21786 & n21788 ) ;
  assign n21794 = n21793 ^ n21789 ^ n14200 ;
  assign n21795 = n10440 ^ n8597 ^ n3123 ;
  assign n21796 = n21795 ^ n8227 ^ n4019 ;
  assign n21798 = ( ~n796 & n4743 ) | ( ~n796 & n5349 ) | ( n4743 & n5349 ) ;
  assign n21797 = n2621 & n4043 ;
  assign n21799 = n21798 ^ n21797 ^ n11655 ;
  assign n21800 = n1278 & ~n8829 ;
  assign n21801 = n1645 & n21800 ;
  assign n21802 = n21801 ^ n3478 ^ 1'b0 ;
  assign n21803 = n21802 ^ n16979 ^ n2729 ;
  assign n21804 = n21803 ^ n2663 ^ n565 ;
  assign n21805 = n7912 ^ n7259 ^ n2810 ;
  assign n21806 = n16516 ^ n13554 ^ 1'b0 ;
  assign n21807 = n21805 | n21806 ;
  assign n21808 = n21807 ^ n11661 ^ 1'b0 ;
  assign n21809 = n12185 | n21808 ;
  assign n21810 = n14317 ^ n9312 ^ 1'b0 ;
  assign n21811 = n15327 | n21810 ;
  assign n21812 = n10947 & ~n21811 ;
  assign n21813 = n21812 ^ n12585 ^ 1'b0 ;
  assign n21814 = ~n9941 & n19028 ;
  assign n21815 = n10251 ^ n10006 ^ n2560 ;
  assign n21816 = n21815 ^ n15856 ^ n2429 ;
  assign n21817 = n21816 ^ n6593 ^ n5219 ;
  assign n21818 = n19854 ^ n18876 ^ n8140 ;
  assign n21819 = n7463 & ~n14707 ;
  assign n21820 = n21794 | n21819 ;
  assign n21821 = n11207 ^ n3437 ^ 1'b0 ;
  assign n21822 = ( ~n3944 & n14396 ) | ( ~n3944 & n21821 ) | ( n14396 & n21821 ) ;
  assign n21823 = n1638 | n7377 ;
  assign n21824 = n21823 ^ n20157 ^ n17597 ;
  assign n21825 = n19732 ^ n3776 ^ 1'b0 ;
  assign n21826 = n9200 ^ n1043 ^ 1'b0 ;
  assign n21827 = x43 & n10640 ;
  assign n21829 = n13686 ^ n3122 ^ n2518 ;
  assign n21828 = ~n4804 & n11473 ;
  assign n21830 = n21829 ^ n21828 ^ n4256 ;
  assign n21831 = n2990 & n14125 ;
  assign n21832 = n12200 & n21831 ;
  assign n21835 = ( n8155 & n8527 ) | ( n8155 & ~n18263 ) | ( n8527 & ~n18263 ) ;
  assign n21833 = n17384 ^ n4218 ^ 1'b0 ;
  assign n21834 = n9547 & n21833 ;
  assign n21836 = n21835 ^ n21834 ^ n11641 ;
  assign n21837 = n7223 ^ n4751 ^ n3604 ;
  assign n21838 = n605 & n12181 ;
  assign n21839 = n21838 ^ n4696 ^ 1'b0 ;
  assign n21840 = n16514 ^ n1574 ^ n496 ;
  assign n21841 = ( n21837 & ~n21839 ) | ( n21837 & n21840 ) | ( ~n21839 & n21840 ) ;
  assign n21842 = n434 | n1340 ;
  assign n21843 = n4570 & ~n21842 ;
  assign n21844 = ( n2887 & ~n14778 ) | ( n2887 & n19336 ) | ( ~n14778 & n19336 ) ;
  assign n21845 = n21844 ^ n1306 ^ 1'b0 ;
  assign n21846 = n10818 & n21845 ;
  assign n21847 = n8921 ^ n8493 ^ n1877 ;
  assign n21848 = ( n3510 & n20172 ) | ( n3510 & n21847 ) | ( n20172 & n21847 ) ;
  assign n21849 = ( n12213 & ~n13006 ) | ( n12213 & n21848 ) | ( ~n13006 & n21848 ) ;
  assign n21850 = n21849 ^ n1606 ^ 1'b0 ;
  assign n21851 = n12872 & n21850 ;
  assign n21852 = n15701 ^ n14464 ^ n13915 ;
  assign n21853 = n9326 ^ n8910 ^ 1'b0 ;
  assign n21854 = ~n5113 & n21853 ;
  assign n21855 = n11062 & n21854 ;
  assign n21856 = n9388 ^ n8226 ^ 1'b0 ;
  assign n21857 = n8845 & n21856 ;
  assign n21858 = n19368 ^ n13006 ^ n5599 ;
  assign n21859 = n7599 & n21858 ;
  assign n21860 = ~n1849 & n21859 ;
  assign n21861 = n18672 ^ n11280 ^ 1'b0 ;
  assign n21862 = n20234 & n21861 ;
  assign n21863 = n696 & ~n5502 ;
  assign n21864 = n21863 ^ n15754 ^ 1'b0 ;
  assign n21865 = ( n811 & ~n5777 ) | ( n811 & n10647 ) | ( ~n5777 & n10647 ) ;
  assign n21866 = n3377 | n3443 ;
  assign n21867 = n21866 ^ n3456 ^ 1'b0 ;
  assign n21868 = n7857 ^ n3657 ^ 1'b0 ;
  assign n21869 = n2285 & n21868 ;
  assign n21870 = ( n1204 & ~n13919 ) | ( n1204 & n21869 ) | ( ~n13919 & n21869 ) ;
  assign n21871 = ( n448 & ~n21867 ) | ( n448 & n21870 ) | ( ~n21867 & n21870 ) ;
  assign n21872 = n9162 ^ n4751 ^ n3035 ;
  assign n21873 = n18049 ^ n1789 ^ 1'b0 ;
  assign n21874 = ( n13700 & n14704 ) | ( n13700 & ~n21873 ) | ( n14704 & ~n21873 ) ;
  assign n21875 = n21874 ^ n10391 ^ 1'b0 ;
  assign n21876 = n21872 & ~n21875 ;
  assign n21877 = ( n16527 & ~n16702 ) | ( n16527 & n21876 ) | ( ~n16702 & n21876 ) ;
  assign n21879 = n5232 ^ n4205 ^ n242 ;
  assign n21880 = n4374 & n21879 ;
  assign n21881 = n21880 ^ n5547 ^ 1'b0 ;
  assign n21878 = n12973 ^ n10096 ^ n2402 ;
  assign n21882 = n21881 ^ n21878 ^ n2459 ;
  assign n21883 = n10328 ^ n9597 ^ n5533 ;
  assign n21884 = ( n7461 & ~n16568 ) | ( n7461 & n21883 ) | ( ~n16568 & n21883 ) ;
  assign n21885 = ( n10872 & n11546 ) | ( n10872 & ~n12361 ) | ( n11546 & ~n12361 ) ;
  assign n21886 = n14671 ^ n4126 ^ 1'b0 ;
  assign n21887 = n21885 & n21886 ;
  assign n21888 = ( n1311 & n3353 ) | ( n1311 & ~n7725 ) | ( n3353 & ~n7725 ) ;
  assign n21889 = n21330 ^ n12756 ^ n2978 ;
  assign n21890 = n10875 ^ n8520 ^ n2501 ;
  assign n21891 = n21890 ^ n14340 ^ n4994 ;
  assign n21893 = x98 | n4644 ;
  assign n21892 = n8299 ^ n7977 ^ 1'b0 ;
  assign n21894 = n21893 ^ n21892 ^ n12834 ;
  assign n21895 = ( n1867 & n19100 ) | ( n1867 & n21894 ) | ( n19100 & n21894 ) ;
  assign n21896 = n16123 ^ n15888 ^ n8507 ;
  assign n21897 = n21896 ^ n21099 ^ 1'b0 ;
  assign n21898 = n725 & ~n5918 ;
  assign n21899 = n21898 ^ n10696 ^ 1'b0 ;
  assign n21900 = n16106 ^ n13990 ^ n4256 ;
  assign n21901 = n11380 ^ n10379 ^ n561 ;
  assign n21902 = ( n2417 & ~n6821 ) | ( n2417 & n21901 ) | ( ~n6821 & n21901 ) ;
  assign n21903 = n21902 ^ n14702 ^ 1'b0 ;
  assign n21904 = n21900 & ~n21903 ;
  assign n21905 = n11002 ^ n630 ^ 1'b0 ;
  assign n21906 = n21778 & ~n21905 ;
  assign n21907 = n7198 & ~n12656 ;
  assign n21908 = n21907 ^ n4860 ^ 1'b0 ;
  assign n21909 = ( n1900 & n5496 ) | ( n1900 & ~n9765 ) | ( n5496 & ~n9765 ) ;
  assign n21910 = n21909 ^ n14932 ^ n8585 ;
  assign n21911 = ( n5114 & ~n6709 ) | ( n5114 & n8788 ) | ( ~n6709 & n8788 ) ;
  assign n21912 = n21911 ^ n6766 ^ n5045 ;
  assign n21913 = ( n3296 & n6599 ) | ( n3296 & n9723 ) | ( n6599 & n9723 ) ;
  assign n21914 = ( n3785 & n20501 ) | ( n3785 & n21913 ) | ( n20501 & n21913 ) ;
  assign n21916 = ( n2749 & n4846 ) | ( n2749 & ~n8069 ) | ( n4846 & ~n8069 ) ;
  assign n21915 = ( n6974 & ~n7481 ) | ( n6974 & n8007 ) | ( ~n7481 & n8007 ) ;
  assign n21917 = n21916 ^ n21915 ^ n11870 ;
  assign n21919 = ( ~n6499 & n11620 ) | ( ~n6499 & n15008 ) | ( n11620 & n15008 ) ;
  assign n21918 = n10634 ^ n346 ^ n300 ;
  assign n21920 = n21919 ^ n21918 ^ n19198 ;
  assign n21921 = n21920 ^ n8704 ^ 1'b0 ;
  assign n21922 = n13527 ^ n7098 ^ n5493 ;
  assign n21923 = ( n13419 & n16648 ) | ( n13419 & n21922 ) | ( n16648 & n21922 ) ;
  assign n21924 = n3041 & n14641 ;
  assign n21925 = n9682 | n13272 ;
  assign n21926 = n13399 & ~n21925 ;
  assign n21927 = ( ~n3380 & n21924 ) | ( ~n3380 & n21926 ) | ( n21924 & n21926 ) ;
  assign n21928 = ( n8045 & n8303 ) | ( n8045 & ~n20027 ) | ( n8303 & ~n20027 ) ;
  assign n21929 = n6510 | n10586 ;
  assign n21930 = n11359 ^ n6430 ^ n5156 ;
  assign n21931 = n13876 ^ n13419 ^ n3078 ;
  assign n21932 = ( n6646 & ~n13301 ) | ( n6646 & n13627 ) | ( ~n13301 & n13627 ) ;
  assign n21933 = ( n21930 & n21931 ) | ( n21930 & ~n21932 ) | ( n21931 & ~n21932 ) ;
  assign n21934 = n20535 ^ n13695 ^ n7905 ;
  assign n21935 = ( ~n648 & n2971 ) | ( ~n648 & n7638 ) | ( n2971 & n7638 ) ;
  assign n21936 = ~n6524 & n6887 ;
  assign n21937 = ( n10050 & ~n21301 ) | ( n10050 & n21936 ) | ( ~n21301 & n21936 ) ;
  assign n21938 = n21937 ^ n4087 ^ 1'b0 ;
  assign n21939 = n18862 | n21938 ;
  assign n21940 = ( n13723 & n21935 ) | ( n13723 & n21939 ) | ( n21935 & n21939 ) ;
  assign n21941 = n2837 & n21121 ;
  assign n21942 = ( n1533 & n3670 ) | ( n1533 & n9237 ) | ( n3670 & n9237 ) ;
  assign n21943 = ( n2912 & n4588 ) | ( n2912 & ~n21942 ) | ( n4588 & ~n21942 ) ;
  assign n21944 = n16128 & ~n21943 ;
  assign n21945 = ~n638 & n5412 ;
  assign n21946 = n21945 ^ n9126 ^ 1'b0 ;
  assign n21947 = n18461 ^ n17661 ^ n8889 ;
  assign n21948 = n21947 ^ n4757 ^ 1'b0 ;
  assign n21949 = n21946 & n21948 ;
  assign n21950 = n19358 ^ n14503 ^ n332 ;
  assign n21951 = n3126 & n12458 ;
  assign n21952 = n540 & n21951 ;
  assign n21953 = ( n7744 & ~n12574 ) | ( n7744 & n21952 ) | ( ~n12574 & n21952 ) ;
  assign n21954 = ( n11920 & ~n15390 ) | ( n11920 & n17891 ) | ( ~n15390 & n17891 ) ;
  assign n21955 = ( n7277 & n11350 ) | ( n7277 & ~n14649 ) | ( n11350 & ~n14649 ) ;
  assign n21956 = n21955 ^ n8272 ^ 1'b0 ;
  assign n21957 = ~n877 & n2520 ;
  assign n21958 = n6311 & n21957 ;
  assign n21959 = n7036 ^ n3714 ^ 1'b0 ;
  assign n21960 = n14053 ^ n9965 ^ 1'b0 ;
  assign n21961 = n13767 ^ n3072 ^ 1'b0 ;
  assign n21962 = n2827 | n19758 ;
  assign n21963 = n1712 | n21713 ;
  assign n21964 = n1037 & ~n21963 ;
  assign n21965 = n10603 | n11322 ;
  assign n21966 = n11058 & ~n21965 ;
  assign n21967 = n15433 ^ n2547 ^ 1'b0 ;
  assign n21968 = n1219 & ~n21967 ;
  assign n21969 = ~n10647 & n21968 ;
  assign n21970 = n8705 & n16812 ;
  assign n21971 = n14290 & n21970 ;
  assign n21972 = n1396 | n9043 ;
  assign n21973 = n21972 ^ n2545 ^ 1'b0 ;
  assign n21974 = n21973 ^ n12821 ^ n9050 ;
  assign n21975 = n7368 ^ n5876 ^ n3432 ;
  assign n21976 = n14578 ^ n5727 ^ 1'b0 ;
  assign n21977 = n5943 | n21976 ;
  assign n21978 = n21486 ^ n13249 ^ n8609 ;
  assign n21979 = n3390 & ~n20522 ;
  assign n21980 = ( ~n16844 & n18531 ) | ( ~n16844 & n21979 ) | ( n18531 & n21979 ) ;
  assign n21989 = n17579 ^ n12821 ^ n5979 ;
  assign n21988 = n20059 ^ n4823 ^ n2437 ;
  assign n21981 = n13254 ^ n8868 ^ n2568 ;
  assign n21984 = ~n3556 & n4622 ;
  assign n21985 = n21984 ^ n9572 ^ n8957 ;
  assign n21982 = ( n1012 & ~n9672 ) | ( n1012 & n10127 ) | ( ~n9672 & n10127 ) ;
  assign n21983 = ~n1005 & n21982 ;
  assign n21986 = n21985 ^ n21983 ^ 1'b0 ;
  assign n21987 = n21981 | n21986 ;
  assign n21990 = n21989 ^ n21988 ^ n21987 ;
  assign n21991 = n294 & n14734 ;
  assign n21992 = n6054 & n21991 ;
  assign n21993 = n21992 ^ n9988 ^ 1'b0 ;
  assign n21994 = ( n6408 & ~n17870 ) | ( n6408 & n21993 ) | ( ~n17870 & n21993 ) ;
  assign n21995 = n10455 ^ n7751 ^ 1'b0 ;
  assign n21996 = n6759 & ~n21995 ;
  assign n21997 = n15539 ^ n10725 ^ n4227 ;
  assign n21998 = ( n308 & n5877 ) | ( n308 & ~n6939 ) | ( n5877 & ~n6939 ) ;
  assign n21999 = ( n1085 & n5759 ) | ( n1085 & n11825 ) | ( n5759 & n11825 ) ;
  assign n22000 = ( ~n12793 & n19736 ) | ( ~n12793 & n21999 ) | ( n19736 & n21999 ) ;
  assign n22001 = n1625 & ~n7700 ;
  assign n22002 = n1280 & n1534 ;
  assign n22003 = ~n19240 & n22002 ;
  assign n22004 = ( n1759 & ~n14930 ) | ( n1759 & n22003 ) | ( ~n14930 & n22003 ) ;
  assign n22005 = n7947 & n9588 ;
  assign n22006 = n605 & n18553 ;
  assign n22007 = n20960 & n22006 ;
  assign n22008 = ( ~n4521 & n22005 ) | ( ~n4521 & n22007 ) | ( n22005 & n22007 ) ;
  assign n22009 = n8602 ^ n5648 ^ 1'b0 ;
  assign n22010 = ~n5580 & n22009 ;
  assign n22011 = ~n3266 & n15785 ;
  assign n22012 = ~n2281 & n22011 ;
  assign n22013 = ( n13125 & n16491 ) | ( n13125 & n20101 ) | ( n16491 & n20101 ) ;
  assign n22014 = n7821 & ~n17771 ;
  assign n22015 = n6603 & ~n8328 ;
  assign n22016 = n22015 ^ n8950 ^ 1'b0 ;
  assign n22017 = ( n10640 & n19939 ) | ( n10640 & n22016 ) | ( n19939 & n22016 ) ;
  assign n22018 = ( n4799 & n5053 ) | ( n4799 & n7777 ) | ( n5053 & n7777 ) ;
  assign n22019 = n20535 ^ n14182 ^ n9797 ;
  assign n22020 = n17628 ^ n13114 ^ n13077 ;
  assign n22021 = n2844 & n9580 ;
  assign n22022 = n22021 ^ n2375 ^ 1'b0 ;
  assign n22023 = n17819 | n22022 ;
  assign n22024 = n22023 ^ n2406 ^ 1'b0 ;
  assign n22025 = ~n1666 & n17025 ;
  assign n22026 = ( x51 & n1898 ) | ( x51 & ~n10818 ) | ( n1898 & ~n10818 ) ;
  assign n22027 = n22026 ^ n1413 ^ 1'b0 ;
  assign n22028 = ~n22025 & n22027 ;
  assign n22029 = n531 & n4051 ;
  assign n22030 = ~n3732 & n14190 ;
  assign n22031 = n22030 ^ n8749 ^ 1'b0 ;
  assign n22032 = ( n2660 & ~n22029 ) | ( n2660 & n22031 ) | ( ~n22029 & n22031 ) ;
  assign n22033 = ( ~x18 & n2895 ) | ( ~x18 & n10605 ) | ( n2895 & n10605 ) ;
  assign n22034 = n7944 ^ n5286 ^ 1'b0 ;
  assign n22035 = n10241 | n22034 ;
  assign n22036 = ( n157 & n4012 ) | ( n157 & ~n22035 ) | ( n4012 & ~n22035 ) ;
  assign n22037 = ( n7013 & ~n7938 ) | ( n7013 & n14453 ) | ( ~n7938 & n14453 ) ;
  assign n22038 = ( n2197 & ~n10010 ) | ( n2197 & n22037 ) | ( ~n10010 & n22037 ) ;
  assign n22039 = ( n1677 & n6487 ) | ( n1677 & ~n17085 ) | ( n6487 & ~n17085 ) ;
  assign n22040 = n11613 ^ n10513 ^ 1'b0 ;
  assign n22041 = n22040 ^ n11546 ^ 1'b0 ;
  assign n22042 = n22039 | n22041 ;
  assign n22043 = n6322 ^ n378 ^ 1'b0 ;
  assign n22044 = ~n20320 & n22043 ;
  assign n22045 = n20575 ^ n3657 ^ 1'b0 ;
  assign n22046 = ~n11978 & n22045 ;
  assign n22047 = ( n4440 & n5407 ) | ( n4440 & ~n6064 ) | ( n5407 & ~n6064 ) ;
  assign n22048 = n22047 ^ n21180 ^ n11834 ;
  assign n22049 = n15825 ^ n14306 ^ n1040 ;
  assign n22050 = ( n328 & n1550 ) | ( n328 & n12465 ) | ( n1550 & n12465 ) ;
  assign n22051 = n22050 ^ n19066 ^ n5801 ;
  assign n22052 = ~n3205 & n8652 ;
  assign n22053 = ( ~n8223 & n11691 ) | ( ~n8223 & n22052 ) | ( n11691 & n22052 ) ;
  assign n22054 = n14206 ^ n3563 ^ 1'b0 ;
  assign n22055 = n5690 | n22054 ;
  assign n22056 = n11211 & ~n22055 ;
  assign n22057 = n21944 | n22056 ;
  assign n22058 = n22057 ^ n14864 ^ 1'b0 ;
  assign n22059 = n3322 | n6390 ;
  assign n22060 = ~n840 & n13450 ;
  assign n22061 = n22060 ^ n3976 ^ 1'b0 ;
  assign n22062 = ( n4187 & n21543 ) | ( n4187 & n22061 ) | ( n21543 & n22061 ) ;
  assign n22063 = n18451 ^ n2943 ^ 1'b0 ;
  assign n22064 = n22063 ^ n10689 ^ n9788 ;
  assign n22065 = n2274 ^ n231 ^ 1'b0 ;
  assign n22066 = n22065 ^ n8454 ^ n4899 ;
  assign n22067 = ( ~n1092 & n11589 ) | ( ~n1092 & n22066 ) | ( n11589 & n22066 ) ;
  assign n22068 = n19107 ^ n12717 ^ n3000 ;
  assign n22069 = n22068 ^ n5820 ^ n5808 ;
  assign n22070 = n3934 & ~n16888 ;
  assign n22071 = n22070 ^ n2733 ^ 1'b0 ;
  assign n22072 = n22071 ^ n12489 ^ n1394 ;
  assign n22073 = ( n1047 & n16473 ) | ( n1047 & n22072 ) | ( n16473 & n22072 ) ;
  assign n22074 = n8620 ^ n4776 ^ n675 ;
  assign n22075 = ( x54 & n4931 ) | ( x54 & ~n8903 ) | ( n4931 & ~n8903 ) ;
  assign n22076 = n7317 ^ n605 ^ 1'b0 ;
  assign n22077 = n6406 | n22076 ;
  assign n22078 = n11409 ^ n7951 ^ n3770 ;
  assign n22079 = n12818 | n22078 ;
  assign n22080 = n6252 | n22079 ;
  assign n22081 = n22080 ^ n17268 ^ 1'b0 ;
  assign n22082 = n16200 ^ n3311 ^ 1'b0 ;
  assign n22083 = n16166 & n22082 ;
  assign n22084 = n8462 ^ n8128 ^ 1'b0 ;
  assign n22085 = n7600 & ~n22084 ;
  assign n22086 = n22085 ^ n18183 ^ 1'b0 ;
  assign n22087 = ( n7439 & n13301 ) | ( n7439 & n17657 ) | ( n13301 & n17657 ) ;
  assign n22088 = ( n9578 & n11988 ) | ( n9578 & ~n22087 ) | ( n11988 & ~n22087 ) ;
  assign n22089 = n4551 & ~n8073 ;
  assign n22090 = ( n1286 & ~n7319 ) | ( n1286 & n22089 ) | ( ~n7319 & n22089 ) ;
  assign n22091 = ( n1613 & ~n3879 ) | ( n1613 & n10201 ) | ( ~n3879 & n10201 ) ;
  assign n22092 = n12253 ^ n1217 ^ 1'b0 ;
  assign n22093 = n22091 | n22092 ;
  assign n22094 = n5872 | n22093 ;
  assign n22095 = n9544 & ~n22094 ;
  assign n22096 = ( n12649 & n21867 ) | ( n12649 & n22095 ) | ( n21867 & n22095 ) ;
  assign n22097 = n20094 ^ n18009 ^ n6732 ;
  assign n22098 = ( ~n4933 & n6120 ) | ( ~n4933 & n6307 ) | ( n6120 & n6307 ) ;
  assign n22099 = ( n8744 & n15037 ) | ( n8744 & ~n22098 ) | ( n15037 & ~n22098 ) ;
  assign n22100 = n13400 ^ n13222 ^ 1'b0 ;
  assign n22101 = n364 | n1301 ;
  assign n22102 = n6028 | n22101 ;
  assign n22103 = ~n690 & n5413 ;
  assign n22104 = n22103 ^ n9687 ^ 1'b0 ;
  assign n22105 = n22104 ^ n9422 ^ 1'b0 ;
  assign n22106 = n334 & ~n22105 ;
  assign n22107 = ( n1750 & ~n5444 ) | ( n1750 & n22106 ) | ( ~n5444 & n22106 ) ;
  assign n22108 = n12177 ^ n10651 ^ n10178 ;
  assign n22109 = ( n13451 & n13517 ) | ( n13451 & n22108 ) | ( n13517 & n22108 ) ;
  assign n22110 = ( n1573 & n8412 ) | ( n1573 & ~n10280 ) | ( n8412 & ~n10280 ) ;
  assign n22111 = n22110 ^ n3747 ^ 1'b0 ;
  assign n22113 = n19835 ^ n10891 ^ n6031 ;
  assign n22114 = n22113 ^ n7682 ^ 1'b0 ;
  assign n22112 = n14984 ^ n10416 ^ n7245 ;
  assign n22115 = n22114 ^ n22112 ^ n19263 ;
  assign n22116 = ( n4843 & n11991 ) | ( n4843 & n12196 ) | ( n11991 & n12196 ) ;
  assign n22117 = ( n529 & n5395 ) | ( n529 & n7454 ) | ( n5395 & n7454 ) ;
  assign n22118 = n17344 & n17856 ;
  assign n22119 = ~n4164 & n22118 ;
  assign n22120 = n22117 & ~n22119 ;
  assign n22121 = ( ~n1852 & n2569 ) | ( ~n1852 & n9388 ) | ( n2569 & n9388 ) ;
  assign n22122 = ( ~n17063 & n22120 ) | ( ~n17063 & n22121 ) | ( n22120 & n22121 ) ;
  assign n22123 = n18500 ^ n6511 ^ 1'b0 ;
  assign n22124 = n2903 | n4143 ;
  assign n22125 = n22124 ^ n1677 ^ 1'b0 ;
  assign n22126 = n22125 ^ n18136 ^ n535 ;
  assign n22127 = ~n6591 & n22126 ;
  assign n22128 = n9896 ^ n3726 ^ n1110 ;
  assign n22129 = n17394 ^ n12331 ^ 1'b0 ;
  assign n22130 = n22128 & ~n22129 ;
  assign n22131 = n22130 ^ n699 ^ n445 ;
  assign n22132 = n22131 ^ n8832 ^ 1'b0 ;
  assign n22133 = ( n7903 & n17690 ) | ( n7903 & ~n22132 ) | ( n17690 & ~n22132 ) ;
  assign n22135 = n12013 ^ n10120 ^ n2750 ;
  assign n22134 = ~n11811 & n11969 ;
  assign n22136 = n22135 ^ n22134 ^ 1'b0 ;
  assign n22137 = n21790 ^ n4939 ^ 1'b0 ;
  assign n22138 = n22136 | n22137 ;
  assign n22139 = ~n2398 & n6023 ;
  assign n22141 = n21047 ^ n11157 ^ n4953 ;
  assign n22140 = n1910 & ~n8211 ;
  assign n22142 = n22141 ^ n22140 ^ n12218 ;
  assign n22143 = n4457 ^ n588 ^ 1'b0 ;
  assign n22144 = ~n3830 & n21667 ;
  assign n22145 = n18756 ^ n13690 ^ 1'b0 ;
  assign n22146 = ( n4400 & n5347 ) | ( n4400 & ~n21815 ) | ( n5347 & ~n21815 ) ;
  assign n22147 = ( n7990 & n16872 ) | ( n7990 & ~n22146 ) | ( n16872 & ~n22146 ) ;
  assign n22148 = ( n12959 & ~n18992 ) | ( n12959 & n22147 ) | ( ~n18992 & n22147 ) ;
  assign n22149 = n11381 ^ n5612 ^ n4296 ;
  assign n22150 = n4164 ^ x62 ^ 1'b0 ;
  assign n22151 = n3508 | n22150 ;
  assign n22152 = ( n10582 & ~n22149 ) | ( n10582 & n22151 ) | ( ~n22149 & n22151 ) ;
  assign n22153 = n1242 & n12074 ;
  assign n22154 = n22153 ^ n13665 ^ 1'b0 ;
  assign n22155 = n20360 ^ n15485 ^ n4035 ;
  assign n22156 = n22155 ^ n13210 ^ 1'b0 ;
  assign n22157 = ~n4544 & n22156 ;
  assign n22158 = n22157 ^ n12737 ^ 1'b0 ;
  assign n22159 = n5100 & ~n5723 ;
  assign n22160 = ~n19618 & n22159 ;
  assign n22161 = n8403 ^ n7323 ^ n2912 ;
  assign n22163 = n12056 ^ n8358 ^ n1963 ;
  assign n22162 = n8954 ^ n5684 ^ n3069 ;
  assign n22164 = n22163 ^ n22162 ^ n14697 ;
  assign n22165 = ( n11041 & ~n19708 ) | ( n11041 & n22164 ) | ( ~n19708 & n22164 ) ;
  assign n22166 = n22161 | n22165 ;
  assign n22167 = n22160 & ~n22166 ;
  assign n22170 = n6183 ^ n2214 ^ n2154 ;
  assign n22171 = n22170 ^ n8938 ^ n2283 ;
  assign n22172 = n6537 | n22171 ;
  assign n22168 = ~n8636 & n20731 ;
  assign n22169 = n22168 ^ n4511 ^ 1'b0 ;
  assign n22173 = n22172 ^ n22169 ^ n8507 ;
  assign n22174 = n13333 ^ n7425 ^ 1'b0 ;
  assign n22175 = ( n10691 & n18755 ) | ( n10691 & ~n22174 ) | ( n18755 & ~n22174 ) ;
  assign n22176 = n22175 ^ n17139 ^ 1'b0 ;
  assign n22177 = n20912 ^ n19840 ^ n6481 ;
  assign n22179 = n1537 | n3045 ;
  assign n22180 = n22179 ^ n7567 ^ 1'b0 ;
  assign n22181 = n346 | n22180 ;
  assign n22178 = n473 & n3319 ;
  assign n22182 = n22181 ^ n22178 ^ n21919 ;
  assign n22183 = n12896 ^ n153 ^ 1'b0 ;
  assign n22184 = ~n18213 & n22183 ;
  assign n22185 = n22184 ^ n9788 ^ n4377 ;
  assign n22186 = ( n9995 & ~n13056 ) | ( n9995 & n22185 ) | ( ~n13056 & n22185 ) ;
  assign n22188 = n15901 ^ n13697 ^ 1'b0 ;
  assign n22187 = n5210 & ~n8966 ;
  assign n22189 = n22188 ^ n22187 ^ 1'b0 ;
  assign n22190 = n4888 & n12476 ;
  assign n22191 = ~n17654 & n22190 ;
  assign n22192 = n22191 ^ n1007 ^ 1'b0 ;
  assign n22193 = ( n4628 & n7347 ) | ( n4628 & n14233 ) | ( n7347 & n14233 ) ;
  assign n22194 = n6729 & n22193 ;
  assign n22195 = ( n1285 & ~n4083 ) | ( n1285 & n22194 ) | ( ~n4083 & n22194 ) ;
  assign n22196 = n17853 ^ n8320 ^ n3093 ;
  assign n22197 = ( n3452 & n10384 ) | ( n3452 & ~n14598 ) | ( n10384 & ~n14598 ) ;
  assign n22198 = n4681 & n4697 ;
  assign n22199 = n22198 ^ n6621 ^ 1'b0 ;
  assign n22200 = n22199 ^ n1908 ^ 1'b0 ;
  assign n22201 = n7073 ^ n6239 ^ 1'b0 ;
  assign n22202 = n22200 | n22201 ;
  assign n22203 = n10919 ^ n6728 ^ 1'b0 ;
  assign n22204 = n2506 & ~n22203 ;
  assign n22205 = n22204 ^ n10138 ^ 1'b0 ;
  assign n22206 = n22205 ^ n2265 ^ 1'b0 ;
  assign n22207 = n21778 & n22206 ;
  assign n22208 = ~n7201 & n22207 ;
  assign n22209 = ( ~n2029 & n4629 ) | ( ~n2029 & n10450 ) | ( n4629 & n10450 ) ;
  assign n22210 = n4598 & ~n22209 ;
  assign n22211 = ( n561 & n4874 ) | ( n561 & n12719 ) | ( n4874 & n12719 ) ;
  assign n22212 = ~n4715 & n22211 ;
  assign n22213 = n7947 & n22212 ;
  assign n22214 = ( n3998 & n8502 ) | ( n3998 & n14859 ) | ( n8502 & n14859 ) ;
  assign n22215 = n16821 ^ n12189 ^ 1'b0 ;
  assign n22216 = ( n938 & n2022 ) | ( n938 & ~n5604 ) | ( n2022 & ~n5604 ) ;
  assign n22217 = n22216 ^ n2638 ^ 1'b0 ;
  assign n22218 = n10878 ^ n10336 ^ n4102 ;
  assign n22219 = ~n8094 & n12263 ;
  assign n22220 = n5408 & ~n9280 ;
  assign n22221 = n1578 & n22220 ;
  assign n22222 = ( n571 & n2752 ) | ( n571 & ~n22221 ) | ( n2752 & ~n22221 ) ;
  assign n22223 = n10106 ^ n4087 ^ n3318 ;
  assign n22224 = n16086 ^ n865 ^ 1'b0 ;
  assign n22225 = x14 & n22224 ;
  assign n22226 = n22225 ^ n6407 ^ n1173 ;
  assign n22227 = ( n12725 & n22223 ) | ( n12725 & n22226 ) | ( n22223 & n22226 ) ;
  assign n22228 = n22227 ^ n6580 ^ 1'b0 ;
  assign n22229 = n22222 & n22228 ;
  assign n22230 = n12246 ^ n6399 ^ n1517 ;
  assign n22231 = n21589 ^ n7970 ^ 1'b0 ;
  assign n22232 = n22230 | n22231 ;
  assign n22234 = n1721 ^ n1573 ^ n698 ;
  assign n22233 = n855 | n3681 ;
  assign n22235 = n22234 ^ n22233 ^ 1'b0 ;
  assign n22236 = n22235 ^ n12143 ^ x25 ;
  assign n22237 = n22236 ^ n18510 ^ 1'b0 ;
  assign n22238 = n11706 | n22237 ;
  assign n22239 = n19022 ^ n14389 ^ n4064 ;
  assign n22240 = ( n9865 & n22238 ) | ( n9865 & ~n22239 ) | ( n22238 & ~n22239 ) ;
  assign n22241 = n4711 & ~n11270 ;
  assign n22242 = n22241 ^ n258 ^ 1'b0 ;
  assign n22243 = n22242 ^ n1034 ^ 1'b0 ;
  assign n22244 = ( ~n4755 & n7840 ) | ( ~n4755 & n12098 ) | ( n7840 & n12098 ) ;
  assign n22245 = n9816 & n13575 ;
  assign n22246 = ( n2803 & n3434 ) | ( n2803 & ~n18433 ) | ( n3434 & ~n18433 ) ;
  assign n22247 = n10503 & n22246 ;
  assign n22248 = n22247 ^ n7806 ^ 1'b0 ;
  assign n22249 = ~n8167 & n13628 ;
  assign n22250 = ( n3266 & n9779 ) | ( n3266 & ~n22199 ) | ( n9779 & ~n22199 ) ;
  assign n22251 = ( n400 & n918 ) | ( n400 & ~n9176 ) | ( n918 & ~n9176 ) ;
  assign n22252 = ( ~n15986 & n22250 ) | ( ~n15986 & n22251 ) | ( n22250 & n22251 ) ;
  assign n22253 = ( n488 & ~n3385 ) | ( n488 & n12372 ) | ( ~n3385 & n12372 ) ;
  assign n22254 = n20847 ^ n8018 ^ n7872 ;
  assign n22255 = n7724 ^ n3517 ^ n2790 ;
  assign n22256 = n6379 & ~n22255 ;
  assign n22257 = n3267 | n22256 ;
  assign n22258 = n11863 ^ n1987 ^ 1'b0 ;
  assign n22259 = n22258 ^ n20522 ^ n5551 ;
  assign n22260 = ( n1875 & n4600 ) | ( n1875 & n15646 ) | ( n4600 & n15646 ) ;
  assign n22261 = ( n22257 & ~n22259 ) | ( n22257 & n22260 ) | ( ~n22259 & n22260 ) ;
  assign n22262 = ( n5156 & n5651 ) | ( n5156 & n20306 ) | ( n5651 & n20306 ) ;
  assign n22263 = n22262 ^ n17090 ^ n4598 ;
  assign n22264 = n18440 ^ n13938 ^ n7004 ;
  assign n22265 = ( ~n7974 & n12635 ) | ( ~n7974 & n22264 ) | ( n12635 & n22264 ) ;
  assign n22266 = ( ~n6179 & n7294 ) | ( ~n6179 & n13870 ) | ( n7294 & n13870 ) ;
  assign n22270 = n12662 ^ n5400 ^ n4566 ;
  assign n22267 = n8931 ^ n4310 ^ n2009 ;
  assign n22268 = n15587 ^ n7004 ^ 1'b0 ;
  assign n22269 = n22267 & ~n22268 ;
  assign n22271 = n22270 ^ n22269 ^ n21597 ;
  assign n22272 = n11355 ^ n10448 ^ n1578 ;
  assign n22273 = n5450 & n16230 ;
  assign n22274 = ~n22272 & n22273 ;
  assign n22275 = n22274 ^ n9358 ^ n4269 ;
  assign n22276 = n17108 ^ n12004 ^ n3188 ;
  assign n22277 = ( ~n2765 & n7922 ) | ( ~n2765 & n22276 ) | ( n7922 & n22276 ) ;
  assign n22278 = ( n2425 & ~n3294 ) | ( n2425 & n12270 ) | ( ~n3294 & n12270 ) ;
  assign n22279 = n22278 ^ n3869 ^ 1'b0 ;
  assign n22280 = ( n2109 & ~n5544 ) | ( n2109 & n16250 ) | ( ~n5544 & n16250 ) ;
  assign n22281 = ~n14045 & n15492 ;
  assign n22282 = n22281 ^ n5448 ^ 1'b0 ;
  assign n22284 = x108 & ~n7627 ;
  assign n22285 = ( ~n168 & n14668 ) | ( ~n168 & n22284 ) | ( n14668 & n22284 ) ;
  assign n22283 = n3805 | n9134 ;
  assign n22286 = n22285 ^ n22283 ^ 1'b0 ;
  assign n22287 = n22286 ^ n21454 ^ n20977 ;
  assign n22288 = ~n9559 & n22287 ;
  assign n22289 = n22282 & n22288 ;
  assign n22290 = n8610 ^ x0 ^ 1'b0 ;
  assign n22291 = ~n977 & n22290 ;
  assign n22295 = n9254 ^ n5452 ^ n4392 ;
  assign n22292 = ( n7482 & ~n9162 ) | ( n7482 & n12935 ) | ( ~n9162 & n12935 ) ;
  assign n22293 = n22292 ^ n9458 ^ 1'b0 ;
  assign n22294 = ~n4356 & n22293 ;
  assign n22296 = n22295 ^ n22294 ^ n13997 ;
  assign n22297 = n9905 | n22296 ;
  assign n22298 = n22291 | n22297 ;
  assign n22304 = ( n1151 & ~n1613 ) | ( n1151 & n15684 ) | ( ~n1613 & n15684 ) ;
  assign n22305 = n2927 | n6811 ;
  assign n22306 = n22304 & ~n22305 ;
  assign n22299 = n266 & n11856 ;
  assign n22300 = n22299 ^ n13244 ^ 1'b0 ;
  assign n22301 = ( x75 & n5950 ) | ( x75 & ~n22300 ) | ( n5950 & ~n22300 ) ;
  assign n22302 = n22301 ^ n3022 ^ 1'b0 ;
  assign n22303 = n11453 & n22302 ;
  assign n22307 = n22306 ^ n22303 ^ n6912 ;
  assign n22308 = n365 & ~n5767 ;
  assign n22309 = ( ~n6957 & n19702 ) | ( ~n6957 & n22308 ) | ( n19702 & n22308 ) ;
  assign n22310 = ( n18011 & n21592 ) | ( n18011 & n22309 ) | ( n21592 & n22309 ) ;
  assign n22311 = ~n3893 & n4137 ;
  assign n22312 = n12151 | n13218 ;
  assign n22313 = n5122 & ~n13088 ;
  assign n22314 = n22312 & n22313 ;
  assign n22316 = n11795 ^ n293 ^ 1'b0 ;
  assign n22317 = n22316 ^ n2523 ^ n1522 ;
  assign n22315 = n12347 ^ n1907 ^ 1'b0 ;
  assign n22318 = n22317 ^ n22315 ^ n18170 ;
  assign n22319 = ( n2017 & n4175 ) | ( n2017 & ~n8164 ) | ( n4175 & ~n8164 ) ;
  assign n22320 = n3062 & ~n22319 ;
  assign n22321 = n22320 ^ n6090 ^ 1'b0 ;
  assign n22322 = ( n280 & ~n4513 ) | ( n280 & n22321 ) | ( ~n4513 & n22321 ) ;
  assign n22323 = n11086 ^ n5710 ^ n2700 ;
  assign n22324 = n22323 ^ n3786 ^ n3219 ;
  assign n22325 = n19985 & ~n22324 ;
  assign n22326 = n597 & n4850 ;
  assign n22327 = n22326 ^ n464 ^ 1'b0 ;
  assign n22328 = ( n3401 & n3977 ) | ( n3401 & n22327 ) | ( n3977 & n22327 ) ;
  assign n22329 = n22328 ^ n7553 ^ n4513 ;
  assign n22330 = ( n5209 & ~n6939 ) | ( n5209 & n15151 ) | ( ~n6939 & n15151 ) ;
  assign n22331 = n9612 ^ n1718 ^ 1'b0 ;
  assign n22332 = n20453 ^ n10535 ^ n971 ;
  assign n22333 = ~n728 & n1108 ;
  assign n22334 = n11299 & n22333 ;
  assign n22335 = ~n22332 & n22334 ;
  assign n22336 = n22335 ^ n20499 ^ n10736 ;
  assign n22337 = n22336 ^ n15029 ^ 1'b0 ;
  assign n22338 = n21935 ^ n3716 ^ n2909 ;
  assign n22339 = n1369 & n12512 ;
  assign n22340 = ( ~n6607 & n12821 ) | ( ~n6607 & n22339 ) | ( n12821 & n22339 ) ;
  assign n22341 = n17186 ^ n2846 ^ 1'b0 ;
  assign n22342 = ~n11380 & n22341 ;
  assign n22343 = n725 & n15932 ;
  assign n22344 = n22343 ^ n11432 ^ 1'b0 ;
  assign n22345 = ( n8952 & ~n22342 ) | ( n8952 & n22344 ) | ( ~n22342 & n22344 ) ;
  assign n22346 = ( n1597 & n5244 ) | ( n1597 & ~n8208 ) | ( n5244 & ~n8208 ) ;
  assign n22347 = n22346 ^ n5333 ^ n4381 ;
  assign n22348 = ( n18331 & ~n22345 ) | ( n18331 & n22347 ) | ( ~n22345 & n22347 ) ;
  assign n22349 = n8103 & n10092 ;
  assign n22350 = n22349 ^ n6238 ^ 1'b0 ;
  assign n22351 = n18857 ^ n14483 ^ 1'b0 ;
  assign n22352 = n19878 & ~n22351 ;
  assign n22353 = n18084 ^ n7266 ^ 1'b0 ;
  assign n22354 = ( n19787 & n20805 ) | ( n19787 & n21947 ) | ( n20805 & n21947 ) ;
  assign n22355 = n19236 ^ n6430 ^ 1'b0 ;
  assign n22356 = n11722 & ~n11844 ;
  assign n22357 = ~n11527 & n22356 ;
  assign n22358 = n18123 & ~n22357 ;
  assign n22359 = ( n3141 & ~n15686 ) | ( n3141 & n20399 ) | ( ~n15686 & n20399 ) ;
  assign n22360 = n22359 ^ n12659 ^ n3723 ;
  assign n22361 = n17346 ^ n11341 ^ n7724 ;
  assign n22362 = n5766 & n9717 ;
  assign n22363 = n21663 ^ n13529 ^ n4844 ;
  assign n22364 = n3462 ^ n329 ^ x86 ;
  assign n22366 = n10437 ^ n7333 ^ n602 ;
  assign n22365 = n12707 ^ n6077 ^ n5735 ;
  assign n22367 = n22366 ^ n22365 ^ 1'b0 ;
  assign n22368 = ( n3610 & ~n4592 ) | ( n3610 & n13674 ) | ( ~n4592 & n13674 ) ;
  assign n22371 = n22163 ^ n3935 ^ 1'b0 ;
  assign n22369 = ~n236 & n10451 ;
  assign n22370 = ~n2286 & n22369 ;
  assign n22372 = n22371 ^ n22370 ^ n15742 ;
  assign n22373 = n22372 ^ n19087 ^ 1'b0 ;
  assign n22374 = ( n7202 & n22368 ) | ( n7202 & n22373 ) | ( n22368 & n22373 ) ;
  assign n22375 = n22374 ^ n20143 ^ n1042 ;
  assign n22376 = n6783 & ~n21828 ;
  assign n22377 = n22376 ^ n3139 ^ 1'b0 ;
  assign n22378 = n6722 & ~n17933 ;
  assign n22379 = n4299 & n22378 ;
  assign n22380 = n8965 | n18495 ;
  assign n22381 = n1797 & n8480 ;
  assign n22382 = n22380 & n22381 ;
  assign n22383 = n17327 ^ n11564 ^ n4410 ;
  assign n22384 = n22383 ^ n14673 ^ n1745 ;
  assign n22385 = n7936 & ~n19708 ;
  assign n22386 = ~n18854 & n22385 ;
  assign n22387 = ( n2686 & ~n4515 ) | ( n2686 & n22386 ) | ( ~n4515 & n22386 ) ;
  assign n22388 = n17875 ^ n4818 ^ n846 ;
  assign n22389 = n12607 & ~n15970 ;
  assign n22390 = ~n22388 & n22389 ;
  assign n22391 = n5828 ^ n4290 ^ n3603 ;
  assign n22392 = ( n2276 & n13825 ) | ( n2276 & ~n22391 ) | ( n13825 & ~n22391 ) ;
  assign n22393 = n22390 & n22392 ;
  assign n22394 = n6187 ^ n5474 ^ n4231 ;
  assign n22406 = ( ~n975 & n2013 ) | ( ~n975 & n7582 ) | ( n2013 & n7582 ) ;
  assign n22404 = n3241 ^ n2260 ^ n317 ;
  assign n22405 = n22404 ^ n4993 ^ n1740 ;
  assign n22407 = n22406 ^ n22405 ^ n15815 ;
  assign n22402 = n14753 ^ n11579 ^ n4997 ;
  assign n22403 = n22402 ^ n10176 ^ n6734 ;
  assign n22395 = n11739 ^ n9419 ^ n2961 ;
  assign n22396 = n22395 ^ n18400 ^ n13490 ;
  assign n22397 = n13344 ^ n8116 ^ n6158 ;
  assign n22398 = ( n7800 & n9280 ) | ( n7800 & n22397 ) | ( n9280 & n22397 ) ;
  assign n22399 = ( n7669 & ~n15993 ) | ( n7669 & n22398 ) | ( ~n15993 & n22398 ) ;
  assign n22400 = ( n1676 & n13056 ) | ( n1676 & ~n22399 ) | ( n13056 & ~n22399 ) ;
  assign n22401 = ( ~n6675 & n22396 ) | ( ~n6675 & n22400 ) | ( n22396 & n22400 ) ;
  assign n22408 = n22407 ^ n22403 ^ n22401 ;
  assign n22409 = ( n1874 & ~n1920 ) | ( n1874 & n8588 ) | ( ~n1920 & n8588 ) ;
  assign n22410 = n20244 ^ n3662 ^ 1'b0 ;
  assign n22411 = n22409 & ~n22410 ;
  assign n22412 = ( n9199 & ~n15876 ) | ( n9199 & n18892 ) | ( ~n15876 & n18892 ) ;
  assign n22414 = n1891 & n6897 ;
  assign n22413 = ( n306 & n9267 ) | ( n306 & n15770 ) | ( n9267 & n15770 ) ;
  assign n22415 = n22414 ^ n22413 ^ n1260 ;
  assign n22416 = ( n4543 & n22412 ) | ( n4543 & n22415 ) | ( n22412 & n22415 ) ;
  assign n22417 = ( ~n1350 & n5199 ) | ( ~n1350 & n20102 ) | ( n5199 & n20102 ) ;
  assign n22418 = n15819 ^ n11840 ^ n4412 ;
  assign n22419 = n7517 | n8042 ;
  assign n22420 = ( n694 & n3259 ) | ( n694 & n18938 ) | ( n3259 & n18938 ) ;
  assign n22421 = n22420 ^ n14060 ^ 1'b0 ;
  assign n22422 = n22421 ^ n11235 ^ 1'b0 ;
  assign n22425 = ( n270 & n463 ) | ( n270 & ~n3014 ) | ( n463 & ~n3014 ) ;
  assign n22423 = ( n1567 & n1788 ) | ( n1567 & n6909 ) | ( n1788 & n6909 ) ;
  assign n22424 = n22423 ^ n5851 ^ n5563 ;
  assign n22426 = n22425 ^ n22424 ^ n7895 ;
  assign n22427 = n22032 ^ n2887 ^ 1'b0 ;
  assign n22428 = ~n22426 & n22427 ;
  assign n22429 = ~n6570 & n10941 ;
  assign n22430 = n7912 & n22429 ;
  assign n22431 = n16846 ^ n4052 ^ n2958 ;
  assign n22432 = n16761 ^ n2672 ^ 1'b0 ;
  assign n22433 = ( ~n3430 & n10037 ) | ( ~n3430 & n14289 ) | ( n10037 & n14289 ) ;
  assign n22434 = n3439 ^ n1318 ^ 1'b0 ;
  assign n22435 = ( ~n5249 & n15538 ) | ( ~n5249 & n22434 ) | ( n15538 & n22434 ) ;
  assign n22436 = n21109 ^ n13782 ^ n7603 ;
  assign n22437 = n7948 ^ n2058 ^ n1141 ;
  assign n22438 = n22437 ^ n10309 ^ n3038 ;
  assign n22439 = n13237 ^ n4731 ^ n1276 ;
  assign n22440 = n3719 ^ n1647 ^ 1'b0 ;
  assign n22441 = n22440 ^ n11889 ^ 1'b0 ;
  assign n22442 = n1931 & n6201 ;
  assign n22443 = ( n738 & ~n3387 ) | ( n738 & n15498 ) | ( ~n3387 & n15498 ) ;
  assign n22444 = ( n20324 & n22442 ) | ( n20324 & ~n22443 ) | ( n22442 & ~n22443 ) ;
  assign n22445 = n22120 ^ n11172 ^ n3518 ;
  assign n22446 = ( n418 & ~n22444 ) | ( n418 & n22445 ) | ( ~n22444 & n22445 ) ;
  assign n22449 = ( ~n8050 & n14772 ) | ( ~n8050 & n16800 ) | ( n14772 & n16800 ) ;
  assign n22447 = n10462 & n17777 ;
  assign n22448 = n2202 & n22447 ;
  assign n22450 = n22449 ^ n22448 ^ n14437 ;
  assign n22451 = ~n4778 & n8389 ;
  assign n22452 = n22451 ^ n19637 ^ 1'b0 ;
  assign n22453 = ( n1054 & ~n5021 ) | ( n1054 & n22452 ) | ( ~n5021 & n22452 ) ;
  assign n22454 = n7823 & ~n14633 ;
  assign n22455 = n22454 ^ n12750 ^ 1'b0 ;
  assign n22456 = n22455 ^ n19119 ^ 1'b0 ;
  assign n22457 = ~n8608 & n22456 ;
  assign n22458 = ( n2624 & n4625 ) | ( n2624 & n14192 ) | ( n4625 & n14192 ) ;
  assign n22459 = ~n13232 & n14939 ;
  assign n22460 = n11370 ^ n10209 ^ n2915 ;
  assign n22466 = n15360 ^ n12472 ^ n5360 ;
  assign n22467 = n22466 ^ n14669 ^ n8020 ;
  assign n22461 = n16477 ^ n12526 ^ 1'b0 ;
  assign n22462 = n18484 & ~n22461 ;
  assign n22463 = n22462 ^ n13928 ^ n1694 ;
  assign n22464 = n4827 & ~n22463 ;
  assign n22465 = n22464 ^ n791 ^ 1'b0 ;
  assign n22468 = n22467 ^ n22465 ^ n6287 ;
  assign n22469 = n4507 & ~n21554 ;
  assign n22470 = n22469 ^ n3804 ^ 1'b0 ;
  assign n22471 = ( n6347 & n15200 ) | ( n6347 & ~n22470 ) | ( n15200 & ~n22470 ) ;
  assign n22472 = ( n4894 & ~n9023 ) | ( n4894 & n19434 ) | ( ~n9023 & n19434 ) ;
  assign n22473 = n1642 | n9293 ;
  assign n22474 = n1086 | n22473 ;
  assign n22475 = n22474 ^ n17298 ^ 1'b0 ;
  assign n22476 = ( ~n10013 & n16646 ) | ( ~n10013 & n22475 ) | ( n16646 & n22475 ) ;
  assign n22477 = ( n4710 & n22472 ) | ( n4710 & ~n22476 ) | ( n22472 & ~n22476 ) ;
  assign n22478 = ~n3764 & n15969 ;
  assign n22479 = n22478 ^ n21533 ^ 1'b0 ;
  assign n22480 = n807 & ~n22479 ;
  assign n22481 = ~n19574 & n22480 ;
  assign n22482 = n14237 ^ n8587 ^ 1'b0 ;
  assign n22483 = n20474 & ~n22482 ;
  assign n22484 = n6226 ^ n2469 ^ 1'b0 ;
  assign n22485 = ~n6204 & n22484 ;
  assign n22486 = n22485 ^ n16913 ^ x49 ;
  assign n22487 = n4873 & n19174 ;
  assign n22488 = ( n3655 & ~n9890 ) | ( n3655 & n22487 ) | ( ~n9890 & n22487 ) ;
  assign n22489 = n3335 & n22488 ;
  assign n22490 = n22489 ^ n3739 ^ 1'b0 ;
  assign n22491 = n22490 ^ n15276 ^ 1'b0 ;
  assign n22492 = ( n1847 & n22486 ) | ( n1847 & n22491 ) | ( n22486 & n22491 ) ;
  assign n22493 = n6207 ^ n1570 ^ n1340 ;
  assign n22494 = n22493 ^ n3522 ^ 1'b0 ;
  assign n22495 = ~n16059 & n22494 ;
  assign n22496 = ( n2617 & n14769 ) | ( n2617 & n22495 ) | ( n14769 & n22495 ) ;
  assign n22497 = ( n6527 & n6927 ) | ( n6527 & ~n11338 ) | ( n6927 & ~n11338 ) ;
  assign n22498 = ( n383 & n13243 ) | ( n383 & n14897 ) | ( n13243 & n14897 ) ;
  assign n22499 = n6890 | n22498 ;
  assign n22500 = ( n4810 & n17727 ) | ( n4810 & n22227 ) | ( n17727 & n22227 ) ;
  assign n22501 = n18337 ^ n16565 ^ 1'b0 ;
  assign n22502 = ~n10007 & n22501 ;
  assign n22503 = n22502 ^ n4141 ^ 1'b0 ;
  assign n22504 = ( n2141 & n10955 ) | ( n2141 & n22503 ) | ( n10955 & n22503 ) ;
  assign n22505 = ( ~n8236 & n11490 ) | ( ~n8236 & n14470 ) | ( n11490 & n14470 ) ;
  assign n22506 = n11953 & n12605 ;
  assign n22507 = n22506 ^ n5562 ^ 1'b0 ;
  assign n22508 = n9897 & n22507 ;
  assign n22510 = n14450 ^ n10238 ^ 1'b0 ;
  assign n22509 = n9931 ^ n3061 ^ 1'b0 ;
  assign n22511 = n22510 ^ n22509 ^ n17991 ;
  assign n22517 = n8811 ^ n8786 ^ n5569 ;
  assign n22518 = ( ~n6982 & n14497 ) | ( ~n6982 & n22517 ) | ( n14497 & n22517 ) ;
  assign n22519 = n22518 ^ n15576 ^ n13299 ;
  assign n22513 = n11341 ^ n4549 ^ n3057 ;
  assign n22512 = ( ~n7571 & n8024 ) | ( ~n7571 & n16344 ) | ( n8024 & n16344 ) ;
  assign n22514 = n22513 ^ n22512 ^ n5302 ;
  assign n22515 = n22514 ^ n10872 ^ n1984 ;
  assign n22516 = ( n16665 & ~n18306 ) | ( n16665 & n22515 ) | ( ~n18306 & n22515 ) ;
  assign n22520 = n22519 ^ n22516 ^ n3083 ;
  assign n22521 = n9316 & n20805 ;
  assign n22522 = n22521 ^ n250 ^ 1'b0 ;
  assign n22524 = ( n1581 & n2464 ) | ( n1581 & ~n7845 ) | ( n2464 & ~n7845 ) ;
  assign n22523 = ( n2016 & ~n3327 ) | ( n2016 & n6789 ) | ( ~n3327 & n6789 ) ;
  assign n22525 = n22524 ^ n22523 ^ 1'b0 ;
  assign n22526 = n4630 & n14605 ;
  assign n22527 = ( n277 & n14368 ) | ( n277 & ~n19873 ) | ( n14368 & ~n19873 ) ;
  assign n22528 = ( ~n3197 & n5719 ) | ( ~n3197 & n22527 ) | ( n5719 & n22527 ) ;
  assign n22529 = n6642 ^ n3942 ^ n1213 ;
  assign n22530 = n387 | n12821 ;
  assign n22531 = n22530 ^ n2634 ^ n1308 ;
  assign n22532 = n11458 ^ n10703 ^ n343 ;
  assign n22533 = n8990 ^ n6959 ^ 1'b0 ;
  assign n22534 = ~n5291 & n22533 ;
  assign n22535 = n813 & n9550 ;
  assign n22536 = n12682 & n22535 ;
  assign n22537 = ( n2087 & n21338 ) | ( n2087 & n22536 ) | ( n21338 & n22536 ) ;
  assign n22538 = ~n16217 & n17276 ;
  assign n22539 = ( n3302 & ~n19107 ) | ( n3302 & n22538 ) | ( ~n19107 & n22538 ) ;
  assign n22540 = x63 & n7360 ;
  assign n22541 = n2503 | n22540 ;
  assign n22542 = n22541 ^ n16173 ^ n13603 ;
  assign n22543 = n5163 ^ n3166 ^ n1493 ;
  assign n22544 = ~n16315 & n22543 ;
  assign n22545 = ( n7644 & n8187 ) | ( n7644 & n18144 ) | ( n8187 & n18144 ) ;
  assign n22546 = n6886 ^ n1377 ^ 1'b0 ;
  assign n22547 = n405 | n22546 ;
  assign n22548 = ( ~n7787 & n12327 ) | ( ~n7787 & n22547 ) | ( n12327 & n22547 ) ;
  assign n22549 = ( n8371 & n14429 ) | ( n8371 & n18905 ) | ( n14429 & n18905 ) ;
  assign n22550 = n22549 ^ n17769 ^ n8425 ;
  assign n22551 = n1152 | n9936 ;
  assign n22552 = n22551 ^ n7408 ^ 1'b0 ;
  assign n22553 = ~n12380 & n22552 ;
  assign n22554 = n22553 ^ n20580 ^ n13665 ;
  assign n22555 = n16218 ^ n3533 ^ 1'b0 ;
  assign n22556 = ~n4544 & n22555 ;
  assign n22557 = n22556 ^ n1695 ^ 1'b0 ;
  assign n22558 = n21254 ^ n18476 ^ n1235 ;
  assign n22559 = ( n347 & n1382 ) | ( n347 & n15277 ) | ( n1382 & n15277 ) ;
  assign n22564 = n3311 & n5778 ;
  assign n22561 = n1413 | n11669 ;
  assign n22562 = n8473 & ~n22561 ;
  assign n22563 = ( n9436 & n14260 ) | ( n9436 & ~n22562 ) | ( n14260 & ~n22562 ) ;
  assign n22560 = ( n2257 & n2566 ) | ( n2257 & n10498 ) | ( n2566 & n10498 ) ;
  assign n22565 = n22564 ^ n22563 ^ n22560 ;
  assign n22566 = ( n17881 & n22559 ) | ( n17881 & ~n22565 ) | ( n22559 & ~n22565 ) ;
  assign n22567 = n5671 ^ n1127 ^ 1'b0 ;
  assign n22568 = n414 | n22567 ;
  assign n22569 = n9757 & n21913 ;
  assign n22570 = ~n22568 & n22569 ;
  assign n22571 = n8082 ^ n6898 ^ n6639 ;
  assign n22572 = n2946 | n3025 ;
  assign n22573 = n6380 & ~n22572 ;
  assign n22574 = ( n2950 & ~n11640 ) | ( n2950 & n22573 ) | ( ~n11640 & n22573 ) ;
  assign n22575 = n22574 ^ n15903 ^ n7106 ;
  assign n22577 = ~n2898 & n8383 ;
  assign n22578 = n1207 & n22577 ;
  assign n22576 = n14854 ^ n11723 ^ n10128 ;
  assign n22579 = n22578 ^ n22576 ^ n1042 ;
  assign n22580 = n15391 ^ n15322 ^ n2160 ;
  assign n22581 = n455 & n5687 ;
  assign n22582 = n22581 ^ n3203 ^ 1'b0 ;
  assign n22585 = n18255 ^ n1252 ^ n473 ;
  assign n22586 = ( n4592 & n15975 ) | ( n4592 & ~n20736 ) | ( n15975 & ~n20736 ) ;
  assign n22587 = n22585 & ~n22586 ;
  assign n22583 = ( n3947 & ~n17127 ) | ( n3947 & n18803 ) | ( ~n17127 & n18803 ) ;
  assign n22584 = n784 | n22583 ;
  assign n22588 = n22587 ^ n22584 ^ 1'b0 ;
  assign n22589 = n2761 | n3747 ;
  assign n22590 = n22589 ^ n18507 ^ 1'b0 ;
  assign n22591 = n7928 & ~n12958 ;
  assign n22592 = n14637 ^ n5583 ^ n4190 ;
  assign n22593 = ( ~n4008 & n18648 ) | ( ~n4008 & n22592 ) | ( n18648 & n22592 ) ;
  assign n22594 = n22593 ^ n16291 ^ 1'b0 ;
  assign n22595 = n16045 ^ n10746 ^ 1'b0 ;
  assign n22596 = n479 & n22595 ;
  assign n22597 = ~n4202 & n10650 ;
  assign n22598 = n22597 ^ n8866 ^ 1'b0 ;
  assign n22599 = n16899 ^ n10397 ^ 1'b0 ;
  assign n22600 = n18623 | n22599 ;
  assign n22601 = n14135 & ~n22600 ;
  assign n22602 = n1519 & n22601 ;
  assign n22603 = n1902 & ~n22602 ;
  assign n22604 = ( n22596 & ~n22598 ) | ( n22596 & n22603 ) | ( ~n22598 & n22603 ) ;
  assign n22605 = n17992 ^ n9251 ^ n8992 ;
  assign n22606 = n22605 ^ n11163 ^ n2159 ;
  assign n22607 = n22606 ^ n17991 ^ n7905 ;
  assign n22608 = n9178 & ~n12566 ;
  assign n22609 = n2902 & ~n17995 ;
  assign n22610 = n8218 & n22609 ;
  assign n22614 = n20989 ^ n3629 ^ n2331 ;
  assign n22611 = n11345 ^ n561 ^ 1'b0 ;
  assign n22612 = n2130 | n22611 ;
  assign n22613 = n711 & ~n22612 ;
  assign n22615 = n22614 ^ n22613 ^ 1'b0 ;
  assign n22616 = n22615 ^ n16050 ^ 1'b0 ;
  assign n22617 = n1309 & n5245 ;
  assign n22618 = n5181 & n22617 ;
  assign n22619 = ( n2568 & ~n15147 ) | ( n2568 & n22618 ) | ( ~n15147 & n22618 ) ;
  assign n22627 = ( n4072 & n4338 ) | ( n4072 & n4465 ) | ( n4338 & n4465 ) ;
  assign n22628 = ( n14464 & n22225 ) | ( n14464 & ~n22627 ) | ( n22225 & ~n22627 ) ;
  assign n22622 = n1440 & n12512 ;
  assign n22623 = ~n18603 & n22622 ;
  assign n22624 = ( n9362 & n13301 ) | ( n9362 & n22623 ) | ( n13301 & n22623 ) ;
  assign n22625 = n19402 ^ n4736 ^ 1'b0 ;
  assign n22626 = n22624 & n22625 ;
  assign n22620 = n5818 ^ n3997 ^ n3072 ;
  assign n22621 = ~n18810 & n22620 ;
  assign n22629 = n22628 ^ n22626 ^ n22621 ;
  assign n22630 = ~n6172 & n17593 ;
  assign n22631 = n8530 & n13575 ;
  assign n22632 = n6041 & n22631 ;
  assign n22633 = n22632 ^ n16670 ^ n5605 ;
  assign n22636 = n14788 ^ n11153 ^ n1719 ;
  assign n22637 = n280 & ~n22636 ;
  assign n22634 = n7806 ^ n2870 ^ 1'b0 ;
  assign n22635 = n322 & n22634 ;
  assign n22638 = n22637 ^ n22635 ^ n8098 ;
  assign n22639 = n2853 ^ n1185 ^ 1'b0 ;
  assign n22640 = ( ~n10306 & n14510 ) | ( ~n10306 & n19293 ) | ( n14510 & n19293 ) ;
  assign n22641 = n14125 & n22640 ;
  assign n22642 = n13811 ^ n8916 ^ 1'b0 ;
  assign n22643 = n17154 | n22642 ;
  assign n22644 = n6982 ^ n6200 ^ n947 ;
  assign n22645 = ~n167 & n16803 ;
  assign n22646 = ~n22644 & n22645 ;
  assign n22647 = ( n22641 & n22643 ) | ( n22641 & ~n22646 ) | ( n22643 & ~n22646 ) ;
  assign n22648 = n3736 & n7371 ;
  assign n22649 = ( ~n7984 & n8947 ) | ( ~n7984 & n9608 ) | ( n8947 & n9608 ) ;
  assign n22650 = ( n8927 & n12427 ) | ( n8927 & n22649 ) | ( n12427 & n22649 ) ;
  assign n22651 = ~n3227 & n9579 ;
  assign n22652 = n6728 ^ n5039 ^ 1'b0 ;
  assign n22653 = ( ~n4167 & n22651 ) | ( ~n4167 & n22652 ) | ( n22651 & n22652 ) ;
  assign n22654 = ( n1017 & n7757 ) | ( n1017 & n8785 ) | ( n7757 & n8785 ) ;
  assign n22655 = ( n9513 & ~n15736 ) | ( n9513 & n16953 ) | ( ~n15736 & n16953 ) ;
  assign n22656 = n3175 & ~n7582 ;
  assign n22657 = ( n7149 & ~n18641 ) | ( n7149 & n22656 ) | ( ~n18641 & n22656 ) ;
  assign n22658 = ~n737 & n7462 ;
  assign n22659 = n15422 ^ n4889 ^ 1'b0 ;
  assign n22660 = n22658 | n22659 ;
  assign n22661 = n17211 ^ n4687 ^ 1'b0 ;
  assign n22662 = n2404 | n22661 ;
  assign n22663 = ( n986 & n14246 ) | ( n986 & ~n16272 ) | ( n14246 & ~n16272 ) ;
  assign n22664 = ( n18002 & n22662 ) | ( n18002 & n22663 ) | ( n22662 & n22663 ) ;
  assign n22665 = n10725 ^ n6264 ^ n3431 ;
  assign n22666 = n3062 & ~n6031 ;
  assign n22667 = ( n14533 & n22665 ) | ( n14533 & n22666 ) | ( n22665 & n22666 ) ;
  assign n22668 = n16724 | n22667 ;
  assign n22669 = n19785 ^ n7898 ^ 1'b0 ;
  assign n22670 = n8473 | n22669 ;
  assign n22671 = ~n21508 & n22670 ;
  assign n22672 = n8315 ^ n5721 ^ 1'b0 ;
  assign n22673 = ( n1871 & n3526 ) | ( n1871 & ~n22672 ) | ( n3526 & ~n22672 ) ;
  assign n22674 = n22225 ^ n5113 ^ n3036 ;
  assign n22675 = ( n2643 & n6999 ) | ( n2643 & ~n22674 ) | ( n6999 & ~n22674 ) ;
  assign n22676 = ( ~n7194 & n22673 ) | ( ~n7194 & n22675 ) | ( n22673 & n22675 ) ;
  assign n22682 = n8779 & ~n10950 ;
  assign n22680 = n1441 & n5620 ;
  assign n22681 = ~n14556 & n22680 ;
  assign n22678 = n2798 ^ n2600 ^ n2103 ;
  assign n22677 = n10674 & n18921 ;
  assign n22679 = n22678 ^ n22677 ^ 1'b0 ;
  assign n22683 = n22682 ^ n22681 ^ n22679 ;
  assign n22684 = n22683 ^ n2445 ^ 1'b0 ;
  assign n22685 = ( n370 & ~n1449 ) | ( n370 & n4377 ) | ( ~n1449 & n4377 ) ;
  assign n22686 = n1089 & ~n4343 ;
  assign n22687 = ( n10732 & n17767 ) | ( n10732 & ~n22686 ) | ( n17767 & ~n22686 ) ;
  assign n22688 = ( n4116 & n22685 ) | ( n4116 & ~n22687 ) | ( n22685 & ~n22687 ) ;
  assign n22689 = n22688 ^ n14460 ^ n5544 ;
  assign n22690 = n19078 ^ n2866 ^ 1'b0 ;
  assign n22691 = n15830 & ~n22690 ;
  assign n22692 = ( n11009 & n13106 ) | ( n11009 & n22691 ) | ( n13106 & n22691 ) ;
  assign n22693 = n13433 ^ n13014 ^ 1'b0 ;
  assign n22694 = ~n602 & n4164 ;
  assign n22695 = n22693 & n22694 ;
  assign n22696 = n8833 & ~n22695 ;
  assign n22697 = ~n22692 & n22696 ;
  assign n22698 = n3037 & n6024 ;
  assign n22699 = n6987 & n22698 ;
  assign n22700 = n16321 ^ n14025 ^ n1133 ;
  assign n22701 = n22700 ^ n4799 ^ 1'b0 ;
  assign n22702 = n12032 & n22701 ;
  assign n22703 = x93 & n6560 ;
  assign n22704 = n22703 ^ n10177 ^ 1'b0 ;
  assign n22705 = ( n1201 & n8359 ) | ( n1201 & ~n22704 ) | ( n8359 & ~n22704 ) ;
  assign n22706 = n1747 & ~n8914 ;
  assign n22707 = ( ~n9777 & n11492 ) | ( ~n9777 & n22706 ) | ( n11492 & n22706 ) ;
  assign n22708 = n22707 ^ n15549 ^ n4639 ;
  assign n22709 = ( ~n19254 & n19329 ) | ( ~n19254 & n22708 ) | ( n19329 & n22708 ) ;
  assign n22710 = n2922 ^ n907 ^ 1'b0 ;
  assign n22711 = n4999 & n22710 ;
  assign n22712 = ( n13560 & n14036 ) | ( n13560 & n22711 ) | ( n14036 & n22711 ) ;
  assign n22713 = ( n17121 & n22709 ) | ( n17121 & ~n22712 ) | ( n22709 & ~n22712 ) ;
  assign n22714 = n12872 ^ n3824 ^ n531 ;
  assign n22715 = ( ~n471 & n11222 ) | ( ~n471 & n22714 ) | ( n11222 & n22714 ) ;
  assign n22716 = n22715 ^ n12999 ^ 1'b0 ;
  assign n22717 = n22716 ^ n9546 ^ n719 ;
  assign n22718 = ( ~n3589 & n10698 ) | ( ~n3589 & n15744 ) | ( n10698 & n15744 ) ;
  assign n22719 = ( n6146 & n8056 ) | ( n6146 & n9028 ) | ( n8056 & n9028 ) ;
  assign n22720 = ( n1482 & n10561 ) | ( n1482 & ~n10806 ) | ( n10561 & ~n10806 ) ;
  assign n22721 = n22720 ^ n9462 ^ n2772 ;
  assign n22722 = ( ~n8815 & n18060 ) | ( ~n8815 & n22721 ) | ( n18060 & n22721 ) ;
  assign n22723 = n1755 ^ n627 ^ 1'b0 ;
  assign n22724 = n22723 ^ n21885 ^ n159 ;
  assign n22725 = n13263 | n22724 ;
  assign n22726 = n19669 ^ n16986 ^ 1'b0 ;
  assign n22727 = n22725 & n22726 ;
  assign n22728 = n8717 ^ n5191 ^ 1'b0 ;
  assign n22729 = n17305 & n22728 ;
  assign n22730 = n6244 & n22729 ;
  assign n22731 = n22730 ^ n8372 ^ 1'b0 ;
  assign n22732 = n16672 & n17604 ;
  assign n22733 = n22732 ^ n7108 ^ 1'b0 ;
  assign n22734 = ( ~n3604 & n19162 ) | ( ~n3604 & n22733 ) | ( n19162 & n22733 ) ;
  assign n22735 = n2473 ^ n425 ^ 1'b0 ;
  assign n22736 = ( n1233 & n3388 ) | ( n1233 & ~n18964 ) | ( n3388 & ~n18964 ) ;
  assign n22737 = ( n8843 & n22735 ) | ( n8843 & n22736 ) | ( n22735 & n22736 ) ;
  assign n22738 = ( n981 & ~n4274 ) | ( n981 & n19224 ) | ( ~n4274 & n19224 ) ;
  assign n22739 = n16387 ^ n4917 ^ 1'b0 ;
  assign n22740 = ~n22738 & n22739 ;
  assign n22741 = n2523 & ~n7841 ;
  assign n22742 = n22741 ^ n2705 ^ 1'b0 ;
  assign n22743 = n22742 ^ n20316 ^ 1'b0 ;
  assign n22744 = n16746 & n22743 ;
  assign n22745 = n6949 ^ n1955 ^ 1'b0 ;
  assign n22746 = n15318 & ~n22745 ;
  assign n22747 = ~n9716 & n11500 ;
  assign n22748 = n14741 & n22747 ;
  assign n22749 = n22748 ^ n18540 ^ n18390 ;
  assign n22750 = n971 & n11622 ;
  assign n22751 = n22750 ^ n11284 ^ n11199 ;
  assign n22752 = n15926 ^ n10672 ^ n5038 ;
  assign n22753 = n22752 ^ n9727 ^ n6384 ;
  assign n22754 = n14988 ^ n8259 ^ 1'b0 ;
  assign n22755 = n22754 ^ n15660 ^ n7952 ;
  assign n22756 = n1024 & n3097 ;
  assign n22757 = n22756 ^ n2219 ^ 1'b0 ;
  assign n22758 = ( n11019 & n12412 ) | ( n11019 & n22757 ) | ( n12412 & n22757 ) ;
  assign n22759 = n2460 & ~n3261 ;
  assign n22760 = ~n3521 & n22759 ;
  assign n22761 = n22760 ^ n16139 ^ n763 ;
  assign n22762 = n11525 & ~n22761 ;
  assign n22763 = ( n5303 & n8266 ) | ( n5303 & n22762 ) | ( n8266 & n22762 ) ;
  assign n22764 = n22763 ^ n13774 ^ 1'b0 ;
  assign n22765 = n3449 | n15050 ;
  assign n22766 = n2900 | n2976 ;
  assign n22767 = n7608 & ~n22766 ;
  assign n22768 = ( n6728 & ~n8996 ) | ( n6728 & n22767 ) | ( ~n8996 & n22767 ) ;
  assign n22769 = n14745 ^ n6111 ^ 1'b0 ;
  assign n22770 = n22768 | n22769 ;
  assign n22775 = ~n11948 & n21202 ;
  assign n22771 = n18313 ^ n9856 ^ n4316 ;
  assign n22772 = n22771 ^ n3172 ^ n2802 ;
  assign n22773 = n22772 ^ n272 ^ 1'b0 ;
  assign n22774 = n12084 & ~n22773 ;
  assign n22776 = n22775 ^ n22774 ^ n9664 ;
  assign n22782 = n5032 & ~n6285 ;
  assign n22777 = ( n624 & n8038 ) | ( n624 & n18698 ) | ( n8038 & n18698 ) ;
  assign n22778 = n22777 ^ n14726 ^ n9984 ;
  assign n22779 = n1882 & n17160 ;
  assign n22780 = ~n22778 & n22779 ;
  assign n22781 = ( n1981 & ~n16966 ) | ( n1981 & n22780 ) | ( ~n16966 & n22780 ) ;
  assign n22783 = n22782 ^ n22781 ^ n7683 ;
  assign n22784 = n14732 ^ n13035 ^ n3991 ;
  assign n22785 = n9801 ^ n7760 ^ 1'b0 ;
  assign n22789 = n5751 ^ n2550 ^ 1'b0 ;
  assign n22787 = n2332 ^ n2039 ^ 1'b0 ;
  assign n22786 = n9338 ^ n8603 ^ 1'b0 ;
  assign n22788 = n22787 ^ n22786 ^ n20974 ;
  assign n22790 = n22789 ^ n22788 ^ n1116 ;
  assign n22791 = n13362 ^ n3666 ^ 1'b0 ;
  assign n22792 = ( n891 & n1494 ) | ( n891 & ~n22791 ) | ( n1494 & ~n22791 ) ;
  assign n22793 = ( n18261 & n19802 ) | ( n18261 & n22792 ) | ( n19802 & n22792 ) ;
  assign n22794 = n9665 ^ n1858 ^ n476 ;
  assign n22795 = ( n11714 & n11764 ) | ( n11714 & ~n22794 ) | ( n11764 & ~n22794 ) ;
  assign n22796 = n19069 ^ n891 ^ 1'b0 ;
  assign n22797 = ~n22795 & n22796 ;
  assign n22798 = n22797 ^ n20072 ^ n10721 ;
  assign n22802 = n5782 & ~n22540 ;
  assign n22800 = n5897 ^ x29 ^ 1'b0 ;
  assign n22799 = n17893 ^ n2324 ^ n1437 ;
  assign n22801 = n22800 ^ n22799 ^ n359 ;
  assign n22803 = n22802 ^ n22801 ^ 1'b0 ;
  assign n22804 = ( n3434 & n5384 ) | ( n3434 & ~n10267 ) | ( n5384 & ~n10267 ) ;
  assign n22805 = n22804 ^ n9235 ^ 1'b0 ;
  assign n22806 = n17488 | n22805 ;
  assign n22807 = n8193 & ~n20516 ;
  assign n22808 = n19210 ^ n17014 ^ 1'b0 ;
  assign n22809 = ( n12505 & ~n13410 ) | ( n12505 & n20987 ) | ( ~n13410 & n20987 ) ;
  assign n22810 = n21095 ^ n2519 ^ n1067 ;
  assign n22811 = ( n3422 & n22809 ) | ( n3422 & ~n22810 ) | ( n22809 & ~n22810 ) ;
  assign n22812 = n135 | n10768 ;
  assign n22813 = n22812 ^ n13780 ^ n12843 ;
  assign n22814 = n13275 ^ n1566 ^ 1'b0 ;
  assign n22817 = n789 | n4735 ;
  assign n22818 = ~n5398 & n22817 ;
  assign n22819 = ~n761 & n22818 ;
  assign n22816 = n12075 ^ n6777 ^ n1790 ;
  assign n22815 = ( x66 & n10244 ) | ( x66 & ~n14536 ) | ( n10244 & ~n14536 ) ;
  assign n22820 = n22819 ^ n22816 ^ n22815 ;
  assign n22821 = n16330 & ~n22164 ;
  assign n22822 = ~n22820 & n22821 ;
  assign n22823 = ( n1818 & n22814 ) | ( n1818 & n22822 ) | ( n22814 & n22822 ) ;
  assign n22824 = ( n13667 & n13815 ) | ( n13667 & n14682 ) | ( n13815 & n14682 ) ;
  assign n22825 = n8925 | n22824 ;
  assign n22826 = n2703 | n22825 ;
  assign n22827 = n2527 ^ n1517 ^ 1'b0 ;
  assign n22828 = ~n11614 & n22827 ;
  assign n22829 = ~n1280 & n22828 ;
  assign n22830 = n666 & ~n669 ;
  assign n22831 = n2769 & n22830 ;
  assign n22832 = n3318 ^ n488 ^ 1'b0 ;
  assign n22833 = n16015 ^ n11540 ^ n2316 ;
  assign n22834 = ( ~n13352 & n14735 ) | ( ~n13352 & n22833 ) | ( n14735 & n22833 ) ;
  assign n22835 = ( n22831 & n22832 ) | ( n22831 & n22834 ) | ( n22832 & n22834 ) ;
  assign n22836 = n20821 ^ n17248 ^ n2539 ;
  assign n22837 = n1176 | n20235 ;
  assign n22838 = ( ~n14233 & n19564 ) | ( ~n14233 & n22837 ) | ( n19564 & n22837 ) ;
  assign n22839 = n12973 ^ n2484 ^ 1'b0 ;
  assign n22840 = n3571 | n22839 ;
  assign n22841 = ( n1372 & n17418 ) | ( n1372 & n22840 ) | ( n17418 & n22840 ) ;
  assign n22842 = ( n7381 & n13790 ) | ( n7381 & n19316 ) | ( n13790 & n19316 ) ;
  assign n22843 = n20958 | n21334 ;
  assign n22844 = n1648 | n2322 ;
  assign n22845 = n2909 | n22844 ;
  assign n22846 = n22845 ^ n21180 ^ n16131 ;
  assign n22847 = n22540 ^ n2356 ^ n1025 ;
  assign n22848 = ( n7848 & n22846 ) | ( n7848 & n22847 ) | ( n22846 & n22847 ) ;
  assign n22849 = n20670 ^ n12354 ^ n1125 ;
  assign n22850 = n8278 ^ n2916 ^ 1'b0 ;
  assign n22851 = n22850 ^ n21115 ^ n10673 ;
  assign n22852 = n17174 ^ n16440 ^ n6020 ;
  assign n22853 = n8280 ^ n7845 ^ n5176 ;
  assign n22854 = n4891 & n10971 ;
  assign n22855 = n1023 | n22854 ;
  assign n22856 = n22853 & ~n22855 ;
  assign n22857 = n1519 & ~n16877 ;
  assign n22862 = ( ~n8646 & n10945 ) | ( ~n8646 & n11174 ) | ( n10945 & n11174 ) ;
  assign n22858 = n13358 ^ x82 ^ 1'b0 ;
  assign n22859 = n10329 ^ n9925 ^ n8298 ;
  assign n22860 = ( ~n19266 & n22858 ) | ( ~n19266 & n22859 ) | ( n22858 & n22859 ) ;
  assign n22861 = n22860 ^ n18343 ^ 1'b0 ;
  assign n22863 = n22862 ^ n22861 ^ n18425 ;
  assign n22864 = n20818 ^ n17875 ^ 1'b0 ;
  assign n22865 = n22863 | n22864 ;
  assign n22870 = ( ~n2213 & n5252 ) | ( ~n2213 & n8793 ) | ( n5252 & n8793 ) ;
  assign n22869 = ~n8358 & n15332 ;
  assign n22866 = n3712 ^ n1916 ^ 1'b0 ;
  assign n22867 = n17041 & ~n22866 ;
  assign n22868 = ( ~n10655 & n22285 ) | ( ~n10655 & n22867 ) | ( n22285 & n22867 ) ;
  assign n22871 = n22870 ^ n22869 ^ n22868 ;
  assign n22872 = ( n3340 & n22865 ) | ( n3340 & n22871 ) | ( n22865 & n22871 ) ;
  assign n22873 = ( ~n140 & n7396 ) | ( ~n140 & n9129 ) | ( n7396 & n9129 ) ;
  assign n22874 = n22873 ^ n4812 ^ n4556 ;
  assign n22875 = n7825 ^ n6548 ^ n2551 ;
  assign n22876 = ( n1009 & n4543 ) | ( n1009 & n5166 ) | ( n4543 & n5166 ) ;
  assign n22877 = n15105 & ~n17780 ;
  assign n22878 = n22876 & n22877 ;
  assign n22879 = n5041 ^ n4545 ^ 1'b0 ;
  assign n22880 = ( n1447 & n1947 ) | ( n1447 & ~n4343 ) | ( n1947 & ~n4343 ) ;
  assign n22881 = ( n14606 & n17181 ) | ( n14606 & n22880 ) | ( n17181 & n22880 ) ;
  assign n22882 = ( n2098 & n13721 ) | ( n2098 & ~n22881 ) | ( n13721 & ~n22881 ) ;
  assign n22883 = n13458 ^ n5402 ^ 1'b0 ;
  assign n22884 = ( n4920 & ~n5195 ) | ( n4920 & n6664 ) | ( ~n5195 & n6664 ) ;
  assign n22885 = n7502 & ~n9198 ;
  assign n22886 = ~n9363 & n22885 ;
  assign n22887 = ( n6042 & ~n22884 ) | ( n6042 & n22886 ) | ( ~n22884 & n22886 ) ;
  assign n22888 = n6473 ^ n3689 ^ n1425 ;
  assign n22889 = x12 & ~n22888 ;
  assign n22890 = ~n22887 & n22889 ;
  assign n22891 = n5927 | n22890 ;
  assign n22892 = n8152 | n22891 ;
  assign n22893 = ( n3963 & ~n9090 ) | ( n3963 & n14289 ) | ( ~n9090 & n14289 ) ;
  assign n22894 = n22893 ^ n4053 ^ n1205 ;
  assign n22895 = n15248 ^ n7299 ^ n1732 ;
  assign n22896 = ( ~n1920 & n5170 ) | ( ~n1920 & n15424 ) | ( n5170 & n15424 ) ;
  assign n22897 = n22896 ^ n11943 ^ n4353 ;
  assign n22898 = n6580 ^ n6388 ^ n643 ;
  assign n22899 = n22898 ^ n19258 ^ 1'b0 ;
  assign n22900 = n7791 | n22899 ;
  assign n22901 = ( n14423 & ~n15634 ) | ( n14423 & n22900 ) | ( ~n15634 & n22900 ) ;
  assign n22903 = n16165 ^ n7624 ^ n6908 ;
  assign n22902 = n12576 ^ n5563 ^ 1'b0 ;
  assign n22904 = n22903 ^ n22902 ^ n1996 ;
  assign n22905 = n15504 ^ n4143 ^ 1'b0 ;
  assign n22906 = ( x115 & ~n386 ) | ( x115 & n9379 ) | ( ~n386 & n9379 ) ;
  assign n22908 = n5157 ^ n3573 ^ 1'b0 ;
  assign n22907 = ~n5268 & n14012 ;
  assign n22909 = n22908 ^ n22907 ^ n2600 ;
  assign n22910 = ( n1541 & ~n14125 ) | ( n1541 & n19426 ) | ( ~n14125 & n19426 ) ;
  assign n22911 = n22909 | n22910 ;
  assign n22912 = ( x35 & ~n12432 ) | ( x35 & n14732 ) | ( ~n12432 & n14732 ) ;
  assign n22913 = ( n8248 & n22911 ) | ( n8248 & n22912 ) | ( n22911 & n22912 ) ;
  assign n22914 = n10402 ^ n4625 ^ 1'b0 ;
  assign n22915 = n1946 & n22914 ;
  assign n22916 = ~n12451 & n22915 ;
  assign n22917 = n17637 ^ n12032 ^ n2239 ;
  assign n22918 = n7548 | n22917 ;
  assign n22919 = n21398 ^ n9662 ^ n7348 ;
  assign n22920 = n10157 | n22919 ;
  assign n22921 = n22920 ^ n15559 ^ 1'b0 ;
  assign n22922 = ( n1958 & ~n16533 ) | ( n1958 & n22685 ) | ( ~n16533 & n22685 ) ;
  assign n22923 = n17084 ^ n10413 ^ n4624 ;
  assign n22924 = ( n1318 & n18310 ) | ( n1318 & ~n22923 ) | ( n18310 & ~n22923 ) ;
  assign n22925 = n2381 & ~n19175 ;
  assign n22926 = n2774 & n4564 ;
  assign n22927 = n22926 ^ n19010 ^ n9060 ;
  assign n22928 = n10721 ^ n8650 ^ 1'b0 ;
  assign n22929 = ~n1121 & n22928 ;
  assign n22930 = n22929 ^ n5246 ^ 1'b0 ;
  assign n22931 = n17111 & n22930 ;
  assign n22932 = n3415 & n22931 ;
  assign n22933 = ~n16521 & n22932 ;
  assign n22934 = n1242 & n12583 ;
  assign n22935 = n14844 & n22934 ;
  assign n22936 = n14414 ^ n12980 ^ 1'b0 ;
  assign n22937 = ( n21097 & n22935 ) | ( n21097 & ~n22936 ) | ( n22935 & ~n22936 ) ;
  assign n22938 = n22937 ^ n15006 ^ 1'b0 ;
  assign n22939 = n9481 | n22938 ;
  assign n22941 = n13463 ^ n1769 ^ x112 ;
  assign n22940 = n360 & ~n6041 ;
  assign n22942 = n22941 ^ n22940 ^ n14515 ;
  assign n22943 = n1713 ^ n609 ^ 1'b0 ;
  assign n22944 = n15691 ^ n10381 ^ n6430 ;
  assign n22945 = n22944 ^ n19489 ^ n9856 ;
  assign n22946 = ( ~n13727 & n22943 ) | ( ~n13727 & n22945 ) | ( n22943 & n22945 ) ;
  assign n22947 = n5630 ^ n4081 ^ 1'b0 ;
  assign n22948 = n22947 ^ n10486 ^ 1'b0 ;
  assign n22949 = ( n4877 & n7409 ) | ( n4877 & n14489 ) | ( n7409 & n14489 ) ;
  assign n22950 = n12284 ^ n6480 ^ n2941 ;
  assign n22951 = ( n20133 & n22949 ) | ( n20133 & ~n22950 ) | ( n22949 & ~n22950 ) ;
  assign n22952 = n14775 ^ n11682 ^ 1'b0 ;
  assign n22953 = n22951 | n22952 ;
  assign n22954 = n4181 | n4911 ;
  assign n22955 = n22954 ^ n12676 ^ 1'b0 ;
  assign n22956 = ~n12676 & n22955 ;
  assign n22957 = ~n2255 & n5603 ;
  assign n22958 = n13194 ^ n9829 ^ 1'b0 ;
  assign n22959 = n12391 ^ n9199 ^ n5891 ;
  assign n22960 = ( n6850 & n14208 ) | ( n6850 & ~n15641 ) | ( n14208 & ~n15641 ) ;
  assign n22961 = n22960 ^ n21745 ^ n6161 ;
  assign n22962 = ( ~n2391 & n9532 ) | ( ~n2391 & n19411 ) | ( n9532 & n19411 ) ;
  assign n22963 = n6666 | n22962 ;
  assign n22964 = n22963 ^ n703 ^ 1'b0 ;
  assign n22965 = n22964 ^ n16198 ^ n13235 ;
  assign n22966 = ( n3546 & n19849 ) | ( n3546 & ~n22965 ) | ( n19849 & ~n22965 ) ;
  assign n22967 = n17041 ^ n7847 ^ n356 ;
  assign n22970 = n13603 ^ n8425 ^ n4518 ;
  assign n22971 = n8793 ^ n7384 ^ 1'b0 ;
  assign n22972 = ~n22970 & n22971 ;
  assign n22968 = n20413 ^ n11208 ^ 1'b0 ;
  assign n22969 = ~n5863 & n22968 ;
  assign n22973 = n22972 ^ n22969 ^ 1'b0 ;
  assign n22974 = ( ~n3017 & n5672 ) | ( ~n3017 & n17434 ) | ( n5672 & n17434 ) ;
  assign n22975 = n20327 ^ n20249 ^ n14150 ;
  assign n22976 = n21772 ^ n1061 ^ 1'b0 ;
  assign n22977 = n14102 ^ n13763 ^ n633 ;
  assign n22978 = ( n2128 & ~n18263 ) | ( n2128 & n22977 ) | ( ~n18263 & n22977 ) ;
  assign n22979 = n22978 ^ n1468 ^ 1'b0 ;
  assign n22980 = n8380 & ~n19993 ;
  assign n22981 = n22980 ^ n7738 ^ 1'b0 ;
  assign n22982 = n9581 ^ n4290 ^ n2798 ;
  assign n22983 = n22982 ^ n19041 ^ n7757 ;
  assign n22984 = n16319 ^ n2638 ^ 1'b0 ;
  assign n22985 = n13351 ^ n9551 ^ 1'b0 ;
  assign n22986 = n22985 ^ n18195 ^ n6212 ;
  assign n22987 = ( ~n3257 & n5095 ) | ( ~n3257 & n7063 ) | ( n5095 & n7063 ) ;
  assign n22988 = n22987 ^ n8629 ^ n8618 ;
  assign n22989 = n22988 ^ n11065 ^ 1'b0 ;
  assign n22990 = n14660 & ~n15958 ;
  assign n22991 = n3507 ^ n3049 ^ 1'b0 ;
  assign n22992 = n13351 & ~n22991 ;
  assign n22993 = ~n9909 & n22992 ;
  assign n22994 = n16500 ^ n8469 ^ n3075 ;
  assign n22995 = n12284 & n22994 ;
  assign n22996 = n22995 ^ n753 ^ 1'b0 ;
  assign n22997 = n3991 & n15784 ;
  assign n22998 = n22997 ^ n10011 ^ x41 ;
  assign n22999 = n22998 ^ n18753 ^ 1'b0 ;
  assign n23000 = ( n9309 & ~n20157 ) | ( n9309 & n22999 ) | ( ~n20157 & n22999 ) ;
  assign n23008 = ( n1588 & n5706 ) | ( n1588 & ~n6879 ) | ( n5706 & ~n6879 ) ;
  assign n23009 = ( ~n4196 & n13651 ) | ( ~n4196 & n23008 ) | ( n13651 & n23008 ) ;
  assign n23006 = ( n4767 & n5193 ) | ( n4767 & n12586 ) | ( n5193 & n12586 ) ;
  assign n23007 = ( n7217 & ~n14695 ) | ( n7217 & n23006 ) | ( ~n14695 & n23006 ) ;
  assign n23001 = ( n1451 & n9717 ) | ( n1451 & n14660 ) | ( n9717 & n14660 ) ;
  assign n23002 = n7560 & ~n19979 ;
  assign n23003 = n2693 & n22199 ;
  assign n23004 = n8652 & n23003 ;
  assign n23005 = ( n23001 & n23002 ) | ( n23001 & ~n23004 ) | ( n23002 & ~n23004 ) ;
  assign n23010 = n23009 ^ n23007 ^ n23005 ;
  assign n23011 = n4306 ^ n942 ^ 1'b0 ;
  assign n23012 = n23011 ^ n16681 ^ n4289 ;
  assign n23013 = n17701 ^ n11598 ^ 1'b0 ;
  assign n23014 = n7825 & n23013 ;
  assign n23015 = ( ~n3593 & n6230 ) | ( ~n3593 & n7083 ) | ( n6230 & n7083 ) ;
  assign n23016 = ( n18151 & ~n23014 ) | ( n18151 & n23015 ) | ( ~n23014 & n23015 ) ;
  assign n23017 = n15473 | n22767 ;
  assign n23018 = n23017 ^ n17556 ^ 1'b0 ;
  assign n23019 = n23018 ^ n9408 ^ x38 ;
  assign n23020 = n11276 ^ n6858 ^ n3096 ;
  assign n23021 = n7234 ^ n300 ^ 1'b0 ;
  assign n23022 = n22165 | n23021 ;
  assign n23024 = n7944 & ~n12778 ;
  assign n23023 = ( n6179 & n16091 ) | ( n6179 & n20430 ) | ( n16091 & n20430 ) ;
  assign n23025 = n23024 ^ n23023 ^ n6027 ;
  assign n23026 = n8916 & n23025 ;
  assign n23027 = ~n6527 & n23026 ;
  assign n23028 = n2934 & n14388 ;
  assign n23029 = n21598 ^ n17928 ^ n17084 ;
  assign n23030 = n19541 ^ n9957 ^ n840 ;
  assign n23031 = n22194 ^ n11543 ^ 1'b0 ;
  assign n23032 = ( ~n23029 & n23030 ) | ( ~n23029 & n23031 ) | ( n23030 & n23031 ) ;
  assign n23033 = n7824 ^ n2192 ^ n148 ;
  assign n23034 = n9907 ^ n1507 ^ n822 ;
  assign n23035 = n23033 | n23034 ;
  assign n23036 = n18958 ^ n6364 ^ n896 ;
  assign n23037 = n23036 ^ n22256 ^ n15356 ;
  assign n23039 = n13373 ^ n12654 ^ n6209 ;
  assign n23038 = n305 & ~n14392 ;
  assign n23040 = n23039 ^ n23038 ^ 1'b0 ;
  assign n23041 = ( n5039 & n12843 ) | ( n5039 & ~n23040 ) | ( n12843 & ~n23040 ) ;
  assign n23042 = ~n5337 & n10948 ;
  assign n23043 = ( ~n510 & n6730 ) | ( ~n510 & n11134 ) | ( n6730 & n11134 ) ;
  assign n23050 = n3265 | n5374 ;
  assign n23051 = n23050 ^ n2440 ^ 1'b0 ;
  assign n23047 = ~n3782 & n6291 ;
  assign n23048 = n23047 ^ n1776 ^ 1'b0 ;
  assign n23049 = ( n1163 & n4988 ) | ( n1163 & ~n23048 ) | ( n4988 & ~n23048 ) ;
  assign n23044 = n1637 & n11852 ;
  assign n23045 = n23044 ^ n5987 ^ 1'b0 ;
  assign n23046 = ( n4398 & n21020 ) | ( n4398 & ~n23045 ) | ( n21020 & ~n23045 ) ;
  assign n23052 = n23051 ^ n23049 ^ n23046 ;
  assign n23053 = ( n6103 & n9644 ) | ( n6103 & n22652 ) | ( n9644 & n22652 ) ;
  assign n23054 = ( n20452 & n23052 ) | ( n20452 & n23053 ) | ( n23052 & n23053 ) ;
  assign n23055 = n19939 ^ n6888 ^ 1'b0 ;
  assign n23056 = n23054 | n23055 ;
  assign n23057 = ( n5337 & n6766 ) | ( n5337 & n14998 ) | ( n6766 & n14998 ) ;
  assign n23058 = ~n10805 & n23057 ;
  assign n23059 = n16144 & n23058 ;
  assign n23060 = ~n8072 & n11938 ;
  assign n23061 = ( n7872 & ~n9722 ) | ( n7872 & n23060 ) | ( ~n9722 & n23060 ) ;
  assign n23062 = n2205 | n23061 ;
  assign n23063 = n23062 ^ n6917 ^ 1'b0 ;
  assign n23064 = n343 & n5372 ;
  assign n23065 = n23064 ^ n7046 ^ 1'b0 ;
  assign n23066 = n14409 ^ n3610 ^ n1542 ;
  assign n23067 = n21427 ^ n12544 ^ n4015 ;
  assign n23069 = ( n1788 & ~n13298 ) | ( n1788 & n20349 ) | ( ~n13298 & n20349 ) ;
  assign n23068 = n365 & n20610 ;
  assign n23070 = n23069 ^ n23068 ^ n18121 ;
  assign n23071 = ( n2306 & ~n4754 ) | ( n2306 & n14060 ) | ( ~n4754 & n14060 ) ;
  assign n23072 = n11476 ^ n6125 ^ 1'b0 ;
  assign n23073 = n5394 & ~n23072 ;
  assign n23074 = ~n21249 & n23073 ;
  assign n23075 = n8834 | n23074 ;
  assign n23076 = n3018 & ~n23075 ;
  assign n23077 = n3522 & n11299 ;
  assign n23078 = n23077 ^ n2543 ^ 1'b0 ;
  assign n23079 = n18170 ^ n4843 ^ 1'b0 ;
  assign n23080 = n23078 & ~n23079 ;
  assign n23081 = ( ~n4610 & n6521 ) | ( ~n4610 & n13783 ) | ( n6521 & n13783 ) ;
  assign n23082 = n23081 ^ n11653 ^ n4247 ;
  assign n23083 = n2578 & n5038 ;
  assign n23084 = ( n15623 & ~n17930 ) | ( n15623 & n23083 ) | ( ~n17930 & n23083 ) ;
  assign n23085 = n4373 ^ n813 ^ n252 ;
  assign n23086 = ( x34 & n9590 ) | ( x34 & ~n23085 ) | ( n9590 & ~n23085 ) ;
  assign n23087 = ( n10048 & ~n12105 ) | ( n10048 & n23086 ) | ( ~n12105 & n23086 ) ;
  assign n23088 = n23087 ^ n18110 ^ n1642 ;
  assign n23089 = n23088 ^ n11345 ^ 1'b0 ;
  assign n23090 = ( ~n18866 & n19403 ) | ( ~n18866 & n23089 ) | ( n19403 & n23089 ) ;
  assign n23091 = n17158 ^ n3776 ^ n3011 ;
  assign n23092 = n5384 & n5947 ;
  assign n23093 = n23092 ^ n5168 ^ 1'b0 ;
  assign n23094 = n23093 ^ n7252 ^ 1'b0 ;
  assign n23095 = ~n13525 & n23094 ;
  assign n23096 = n23095 ^ n12793 ^ n729 ;
  assign n23097 = n23096 ^ n18850 ^ n17012 ;
  assign n23098 = n18266 & n22746 ;
  assign n23099 = n23098 ^ n6000 ^ 1'b0 ;
  assign n23100 = n8183 ^ n3079 ^ 1'b0 ;
  assign n23101 = ~n669 & n14961 ;
  assign n23102 = n23101 ^ n3834 ^ 1'b0 ;
  assign n23103 = n5095 & n14660 ;
  assign n23104 = n4048 & n23103 ;
  assign n23105 = ( n12762 & n23102 ) | ( n12762 & ~n23104 ) | ( n23102 & ~n23104 ) ;
  assign n23106 = ( n11742 & n20483 ) | ( n11742 & n21544 ) | ( n20483 & n21544 ) ;
  assign n23107 = n20014 ^ n4192 ^ n2191 ;
  assign n23108 = ( ~n1781 & n13292 ) | ( ~n1781 & n23107 ) | ( n13292 & n23107 ) ;
  assign n23109 = ( ~n8451 & n20825 ) | ( ~n8451 & n23108 ) | ( n20825 & n23108 ) ;
  assign n23110 = ( ~n9007 & n17174 ) | ( ~n9007 & n21272 ) | ( n17174 & n21272 ) ;
  assign n23111 = ~n8855 & n21723 ;
  assign n23112 = n23111 ^ n13829 ^ 1'b0 ;
  assign n23113 = n17701 | n23031 ;
  assign n23114 = ( n18543 & ~n21932 ) | ( n18543 & n22439 ) | ( ~n21932 & n22439 ) ;
  assign n23115 = n21600 ^ n8722 ^ n2467 ;
  assign n23116 = ( n3247 & ~n3999 ) | ( n3247 & n13251 ) | ( ~n3999 & n13251 ) ;
  assign n23117 = n20518 ^ n12219 ^ n1735 ;
  assign n23120 = ( n1230 & n1508 ) | ( n1230 & n8529 ) | ( n1508 & n8529 ) ;
  assign n23118 = x90 & n8590 ;
  assign n23119 = n23118 ^ n21312 ^ n19964 ;
  assign n23121 = n23120 ^ n23119 ^ 1'b0 ;
  assign n23122 = n16273 & n23121 ;
  assign n23123 = n18784 ^ n1380 ^ 1'b0 ;
  assign n23124 = n10784 | n23123 ;
  assign n23125 = n3838 ^ n1595 ^ n1454 ;
  assign n23126 = n23125 ^ n20807 ^ x50 ;
  assign n23127 = n18019 ^ n2050 ^ x75 ;
  assign n23128 = ( n6531 & ~n20662 ) | ( n6531 & n23127 ) | ( ~n20662 & n23127 ) ;
  assign n23129 = n14603 ^ n10318 ^ n2558 ;
  assign n23130 = n1263 & ~n11563 ;
  assign n23131 = n23130 ^ n18972 ^ 1'b0 ;
  assign n23132 = n23131 ^ n14292 ^ n4746 ;
  assign n23133 = ~n1335 & n11922 ;
  assign n23134 = n23133 ^ n19929 ^ n17059 ;
  assign n23135 = n23134 ^ n9977 ^ 1'b0 ;
  assign n23136 = ( n14386 & n20742 ) | ( n14386 & n23135 ) | ( n20742 & n23135 ) ;
  assign n23137 = n15676 ^ n11433 ^ n4756 ;
  assign n23138 = n13164 ^ n9190 ^ n1470 ;
  assign n23139 = ~n20486 & n23138 ;
  assign n23140 = n23139 ^ n18934 ^ n14886 ;
  assign n23141 = ( n3599 & ~n9597 ) | ( n3599 & n15258 ) | ( ~n9597 & n15258 ) ;
  assign n23142 = n23141 ^ n11024 ^ n5005 ;
  assign n23143 = ( n6662 & n9452 ) | ( n6662 & n23142 ) | ( n9452 & n23142 ) ;
  assign n23144 = n6746 ^ n3572 ^ 1'b0 ;
  assign n23145 = n9511 & n23144 ;
  assign n23146 = n23145 ^ n3681 ^ 1'b0 ;
  assign n23147 = n23143 & ~n23146 ;
  assign n23148 = x60 & ~n12190 ;
  assign n23149 = n7277 & n23148 ;
  assign n23150 = n23149 ^ n1032 ^ 1'b0 ;
  assign n23151 = n15309 | n23150 ;
  assign n23152 = n144 & ~n22518 ;
  assign n23153 = ~n19547 & n23152 ;
  assign n23154 = n23153 ^ n15030 ^ 1'b0 ;
  assign n23155 = n12551 & n23154 ;
  assign n23156 = n17788 ^ n14498 ^ 1'b0 ;
  assign n23157 = ( ~n12219 & n22443 ) | ( ~n12219 & n23156 ) | ( n22443 & n23156 ) ;
  assign n23158 = n18197 ^ n11093 ^ n7739 ;
  assign n23159 = n10411 ^ n6838 ^ n2040 ;
  assign n23160 = n1694 & ~n3887 ;
  assign n23161 = ( n2360 & ~n9517 ) | ( n2360 & n23160 ) | ( ~n9517 & n23160 ) ;
  assign n23162 = n16253 ^ n8032 ^ 1'b0 ;
  assign n23163 = ~n5078 & n5471 ;
  assign n23164 = n13034 & n23163 ;
  assign n23167 = n7819 ^ n2527 ^ 1'b0 ;
  assign n23168 = n12205 | n23167 ;
  assign n23169 = ( n499 & n22160 ) | ( n499 & n23168 ) | ( n22160 & n23168 ) ;
  assign n23165 = n4083 & n19047 ;
  assign n23166 = n23165 ^ x50 ^ 1'b0 ;
  assign n23170 = n23169 ^ n23166 ^ n2897 ;
  assign n23171 = n20185 ^ n7412 ^ n1262 ;
  assign n23172 = n1407 & ~n2928 ;
  assign n23173 = ~x125 & n23172 ;
  assign n23174 = ( n8094 & ~n11285 ) | ( n8094 & n23173 ) | ( ~n11285 & n23173 ) ;
  assign n23175 = ~n3111 & n15735 ;
  assign n23176 = n23175 ^ n10541 ^ 1'b0 ;
  assign n23177 = n14703 | n15406 ;
  assign n23178 = n662 & ~n23177 ;
  assign n23179 = ( n3211 & n8998 ) | ( n3211 & ~n15004 ) | ( n8998 & ~n15004 ) ;
  assign n23180 = ( ~n4656 & n7264 ) | ( ~n4656 & n13524 ) | ( n7264 & n13524 ) ;
  assign n23181 = n9162 ^ n4819 ^ n1925 ;
  assign n23182 = n23181 ^ n19305 ^ n4187 ;
  assign n23183 = ~n4417 & n21114 ;
  assign n23185 = n5979 ^ n1833 ^ 1'b0 ;
  assign n23184 = n10624 ^ n144 ^ 1'b0 ;
  assign n23186 = n23185 ^ n23184 ^ n13674 ;
  assign n23187 = ( n1766 & n16479 ) | ( n1766 & n22638 ) | ( n16479 & n22638 ) ;
  assign n23188 = n20099 ^ n13868 ^ n11742 ;
  assign n23189 = n11823 ^ n7208 ^ n5327 ;
  assign n23190 = n23189 ^ n5717 ^ n4151 ;
  assign n23191 = n7038 ^ n4331 ^ 1'b0 ;
  assign n23192 = ~n23190 & n23191 ;
  assign n23193 = ( n8920 & n13099 ) | ( n8920 & n14689 ) | ( n13099 & n14689 ) ;
  assign n23195 = n22255 ^ n5724 ^ 1'b0 ;
  assign n23196 = ( n4717 & n6772 ) | ( n4717 & ~n23195 ) | ( n6772 & ~n23195 ) ;
  assign n23194 = n3491 & ~n8128 ;
  assign n23197 = n23196 ^ n23194 ^ 1'b0 ;
  assign n23199 = n3464 ^ n812 ^ 1'b0 ;
  assign n23200 = ~n4048 & n23199 ;
  assign n23198 = n2789 ^ n1676 ^ n1222 ;
  assign n23201 = n23200 ^ n23198 ^ n13621 ;
  assign n23202 = ~n5818 & n10867 ;
  assign n23203 = ( n11742 & n22278 ) | ( n11742 & n23202 ) | ( n22278 & n23202 ) ;
  assign n23204 = n23203 ^ n6416 ^ n3992 ;
  assign n23205 = ( n8591 & n23201 ) | ( n8591 & ~n23204 ) | ( n23201 & ~n23204 ) ;
  assign n23206 = ( x66 & n23197 ) | ( x66 & n23205 ) | ( n23197 & n23205 ) ;
  assign n23207 = n11227 ^ n3209 ^ 1'b0 ;
  assign n23208 = ~n6060 & n23207 ;
  assign n23209 = n23208 ^ n16439 ^ 1'b0 ;
  assign n23210 = ( n3148 & ~n3622 ) | ( n3148 & n5443 ) | ( ~n3622 & n5443 ) ;
  assign n23211 = ( n304 & n7318 ) | ( n304 & ~n19834 ) | ( n7318 & ~n19834 ) ;
  assign n23212 = n7962 & ~n11845 ;
  assign n23213 = n23212 ^ x112 ^ 1'b0 ;
  assign n23214 = ( n3034 & n6860 ) | ( n3034 & n18814 ) | ( n6860 & n18814 ) ;
  assign n23215 = n23214 ^ n1887 ^ 1'b0 ;
  assign n23216 = ( ~n11906 & n13112 ) | ( ~n11906 & n23215 ) | ( n13112 & n23215 ) ;
  assign n23217 = ~n23213 & n23216 ;
  assign n23218 = ~n23211 & n23217 ;
  assign n23219 = n23218 ^ n12981 ^ n1042 ;
  assign n23220 = n18514 ^ n15815 ^ n9093 ;
  assign n23221 = n12977 ^ n6257 ^ 1'b0 ;
  assign n23222 = n3146 & ~n23221 ;
  assign n23223 = n19561 ^ n10656 ^ 1'b0 ;
  assign n23224 = n23222 & n23223 ;
  assign n23225 = ~n4141 & n14480 ;
  assign n23226 = n17359 & n23225 ;
  assign n23227 = ( n5176 & ~n11047 ) | ( n5176 & n19971 ) | ( ~n11047 & n19971 ) ;
  assign n23228 = n19740 & n23227 ;
  assign n23229 = n23228 ^ n5001 ^ 1'b0 ;
  assign n23230 = n8627 ^ n2190 ^ 1'b0 ;
  assign n23231 = n1407 & ~n23230 ;
  assign n23232 = n19133 & n23231 ;
  assign n23233 = ( ~n2111 & n3104 ) | ( ~n2111 & n5466 ) | ( n3104 & n5466 ) ;
  assign n23234 = n23233 ^ n20829 ^ n12158 ;
  assign n23235 = ~n2851 & n4029 ;
  assign n23236 = n23235 ^ n20971 ^ 1'b0 ;
  assign n23237 = ( n10767 & ~n12835 ) | ( n10767 & n19492 ) | ( ~n12835 & n19492 ) ;
  assign n23238 = ~n23236 & n23237 ;
  assign n23239 = n10006 ^ n4318 ^ 1'b0 ;
  assign n23240 = ~n6751 & n20051 ;
  assign n23241 = n23240 ^ n20957 ^ 1'b0 ;
  assign n23242 = n23239 | n23241 ;
  assign n23244 = n10475 ^ n6856 ^ n745 ;
  assign n23245 = n23244 ^ n4748 ^ n4207 ;
  assign n23243 = n4511 & n19323 ;
  assign n23246 = n23245 ^ n23243 ^ 1'b0 ;
  assign n23247 = ( ~n10655 & n20021 ) | ( ~n10655 & n21420 ) | ( n20021 & n21420 ) ;
  assign n23248 = n23247 ^ n3322 ^ 1'b0 ;
  assign n23249 = n23246 & n23248 ;
  assign n23251 = n10003 | n14007 ;
  assign n23250 = n22239 ^ n13323 ^ n3453 ;
  assign n23252 = n23251 ^ n23250 ^ 1'b0 ;
  assign n23253 = n15635 & ~n23252 ;
  assign n23254 = ( ~n200 & n7549 ) | ( ~n200 & n8187 ) | ( n7549 & n8187 ) ;
  assign n23255 = ( n13941 & n16808 ) | ( n13941 & n23254 ) | ( n16808 & n23254 ) ;
  assign n23256 = ( ~n1738 & n11128 ) | ( ~n1738 & n12792 ) | ( n11128 & n12792 ) ;
  assign n23257 = ( ~n16979 & n23255 ) | ( ~n16979 & n23256 ) | ( n23255 & n23256 ) ;
  assign n23258 = ( n553 & n1478 ) | ( n553 & ~n8284 ) | ( n1478 & ~n8284 ) ;
  assign n23259 = n1113 & ~n8156 ;
  assign n23260 = ( n10006 & ~n21229 ) | ( n10006 & n23259 ) | ( ~n21229 & n23259 ) ;
  assign n23261 = ( ~n5283 & n9404 ) | ( ~n5283 & n23260 ) | ( n9404 & n23260 ) ;
  assign n23262 = ( n6374 & ~n10880 ) | ( n6374 & n23261 ) | ( ~n10880 & n23261 ) ;
  assign n23263 = n19240 ^ n2645 ^ n435 ;
  assign n23264 = ( n9354 & ~n19502 ) | ( n9354 & n23263 ) | ( ~n19502 & n23263 ) ;
  assign n23265 = n19000 ^ n12023 ^ 1'b0 ;
  assign n23266 = ~n15550 & n23265 ;
  assign n23267 = n10486 ^ n10101 ^ n8574 ;
  assign n23269 = ( n7682 & ~n12311 ) | ( n7682 & n13960 ) | ( ~n12311 & n13960 ) ;
  assign n23270 = ( ~n331 & n17239 ) | ( ~n331 & n23269 ) | ( n17239 & n23269 ) ;
  assign n23268 = n8413 | n21747 ;
  assign n23271 = n23270 ^ n23268 ^ 1'b0 ;
  assign n23272 = ( n2894 & n11605 ) | ( n2894 & n15474 ) | ( n11605 & n15474 ) ;
  assign n23273 = n23272 ^ n10008 ^ n8090 ;
  assign n23276 = ~n1854 & n3334 ;
  assign n23277 = n23276 ^ n9475 ^ 1'b0 ;
  assign n23274 = n3297 ^ n665 ^ x33 ;
  assign n23275 = n23274 ^ n18239 ^ n4617 ;
  assign n23278 = n23277 ^ n23275 ^ n8316 ;
  assign n23279 = n6149 ^ n2163 ^ n1116 ;
  assign n23280 = n23279 ^ n4589 ^ n659 ;
  assign n23281 = n23280 ^ n5537 ^ 1'b0 ;
  assign n23282 = n711 & n7517 ;
  assign n23283 = ~n1545 & n23282 ;
  assign n23284 = n12505 ^ n791 ^ 1'b0 ;
  assign n23285 = ~n23283 & n23284 ;
  assign n23286 = ( n6164 & n9627 ) | ( n6164 & n23285 ) | ( n9627 & n23285 ) ;
  assign n23287 = ~n8088 & n23286 ;
  assign n23288 = n17867 ^ n17605 ^ n11272 ;
  assign n23289 = ( ~n267 & n3052 ) | ( ~n267 & n11051 ) | ( n3052 & n11051 ) ;
  assign n23290 = n14233 ^ n12659 ^ n2830 ;
  assign n23291 = n23290 ^ n3401 ^ n1059 ;
  assign n23292 = n11330 ^ n5234 ^ 1'b0 ;
  assign n23293 = n7929 & ~n23292 ;
  assign n23294 = ~n3966 & n17889 ;
  assign n23295 = n372 & n23294 ;
  assign n23296 = n5980 & ~n16466 ;
  assign n23297 = n23296 ^ n7734 ^ 1'b0 ;
  assign n23298 = ~n11100 & n16566 ;
  assign n23299 = ~n6208 & n23298 ;
  assign n23301 = ( n12583 & n18386 ) | ( n12583 & ~n23141 ) | ( n18386 & ~n23141 ) ;
  assign n23300 = n8142 & ~n13771 ;
  assign n23302 = n23301 ^ n23300 ^ 1'b0 ;
  assign n23303 = ( n6666 & ~n23299 ) | ( n6666 & n23302 ) | ( ~n23299 & n23302 ) ;
  assign n23304 = ( n8599 & n12818 ) | ( n8599 & n18076 ) | ( n12818 & n18076 ) ;
  assign n23305 = ~n1927 & n2312 ;
  assign n23306 = ~n5405 & n23305 ;
  assign n23307 = n15211 & n23306 ;
  assign n23308 = n1494 | n23307 ;
  assign n23309 = ( n2057 & n15772 ) | ( n2057 & n23308 ) | ( n15772 & n23308 ) ;
  assign n23310 = ( n3918 & n11585 ) | ( n3918 & ~n14877 ) | ( n11585 & ~n14877 ) ;
  assign n23311 = ( ~n13804 & n15616 ) | ( ~n13804 & n23310 ) | ( n15616 & n23310 ) ;
  assign n23312 = n7471 ^ n7296 ^ 1'b0 ;
  assign n23313 = n4743 | n23312 ;
  assign n23315 = n6308 ^ n2105 ^ 1'b0 ;
  assign n23316 = n5090 & ~n23315 ;
  assign n23314 = ~n2390 & n3551 ;
  assign n23317 = n23316 ^ n23314 ^ 1'b0 ;
  assign n23318 = n14819 ^ n8351 ^ 1'b0 ;
  assign n23319 = n7466 | n23318 ;
  assign n23320 = n20331 & ~n23319 ;
  assign n23321 = n6737 | n21336 ;
  assign n23322 = ( ~n1260 & n7651 ) | ( ~n1260 & n16953 ) | ( n7651 & n16953 ) ;
  assign n23323 = n23322 ^ n3907 ^ 1'b0 ;
  assign n23324 = n12126 ^ n3401 ^ 1'b0 ;
  assign n23325 = n5687 & n23324 ;
  assign n23326 = n3680 & ~n23325 ;
  assign n23327 = n731 | n5001 ;
  assign n23328 = n3718 & ~n23327 ;
  assign n23329 = n23173 ^ n17800 ^ 1'b0 ;
  assign n23330 = n8356 ^ n6420 ^ 1'b0 ;
  assign n23331 = n9441 | n23330 ;
  assign n23333 = ( n6187 & n11616 ) | ( n6187 & n16225 ) | ( n11616 & n16225 ) ;
  assign n23332 = ( n5557 & ~n9567 ) | ( n5557 & n20669 ) | ( ~n9567 & n20669 ) ;
  assign n23334 = n23333 ^ n23332 ^ n9407 ;
  assign n23335 = n15628 ^ n15572 ^ n5655 ;
  assign n23336 = ( n1404 & ~n3334 ) | ( n1404 & n3892 ) | ( ~n3334 & n3892 ) ;
  assign n23337 = n2183 ^ n355 ^ 1'b0 ;
  assign n23338 = ( n12324 & ~n23336 ) | ( n12324 & n23337 ) | ( ~n23336 & n23337 ) ;
  assign n23339 = ~n2697 & n23338 ;
  assign n23342 = ( n846 & n15749 ) | ( n846 & n20966 ) | ( n15749 & n20966 ) ;
  assign n23340 = n11521 ^ n3787 ^ 1'b0 ;
  assign n23341 = ( x71 & n8216 ) | ( x71 & ~n23340 ) | ( n8216 & ~n23340 ) ;
  assign n23343 = n23342 ^ n23341 ^ n3066 ;
  assign n23344 = n20955 ^ n11631 ^ n8728 ;
  assign n23345 = ( ~n1291 & n5602 ) | ( ~n1291 & n10673 ) | ( n5602 & n10673 ) ;
  assign n23346 = n23345 ^ n4538 ^ 1'b0 ;
  assign n23347 = ( ~n10788 & n13051 ) | ( ~n10788 & n15873 ) | ( n13051 & n15873 ) ;
  assign n23348 = n23346 & n23347 ;
  assign n23349 = n23348 ^ n5594 ^ 1'b0 ;
  assign n23351 = n4859 ^ n3962 ^ n1801 ;
  assign n23350 = n13875 ^ n5533 ^ n827 ;
  assign n23352 = n23351 ^ n23350 ^ n16683 ;
  assign n23353 = n8480 & ~n9223 ;
  assign n23354 = ( n1181 & n11970 ) | ( n1181 & n23353 ) | ( n11970 & n23353 ) ;
  assign n23355 = ( ~n12649 & n13880 ) | ( ~n12649 & n23354 ) | ( n13880 & n23354 ) ;
  assign n23356 = ( n2981 & ~n6576 ) | ( n2981 & n13428 ) | ( ~n6576 & n13428 ) ;
  assign n23359 = ( n7976 & ~n12476 ) | ( n7976 & n19638 ) | ( ~n12476 & n19638 ) ;
  assign n23358 = n13562 | n15964 ;
  assign n23357 = n6919 ^ n5359 ^ n3637 ;
  assign n23360 = n23359 ^ n23358 ^ n23357 ;
  assign n23361 = n13631 ^ n13091 ^ n7243 ;
  assign n23362 = n12996 ^ n10278 ^ n8469 ;
  assign n23363 = ~n5943 & n12304 ;
  assign n23364 = n15646 & n23363 ;
  assign n23365 = n9614 ^ n4025 ^ x8 ;
  assign n23366 = n22784 & n23365 ;
  assign n23367 = ~n19938 & n23366 ;
  assign n23369 = ( ~n325 & n5630 ) | ( ~n325 & n10805 ) | ( n5630 & n10805 ) ;
  assign n23370 = n23369 ^ n10228 ^ n5731 ;
  assign n23368 = ( ~n5153 & n5214 ) | ( ~n5153 & n6964 ) | ( n5214 & n6964 ) ;
  assign n23371 = n23370 ^ n23368 ^ 1'b0 ;
  assign n23372 = n16635 ^ n11749 ^ n2436 ;
  assign n23373 = ( x29 & n684 ) | ( x29 & ~n14165 ) | ( n684 & ~n14165 ) ;
  assign n23374 = n17439 ^ n13624 ^ 1'b0 ;
  assign n23375 = n18283 ^ n11062 ^ n9952 ;
  assign n23376 = n14367 | n16390 ;
  assign n23377 = ( n2482 & n9817 ) | ( n2482 & n15097 ) | ( n9817 & n15097 ) ;
  assign n23378 = n12653 & n23377 ;
  assign n23379 = ( n17166 & n23141 ) | ( n17166 & n23378 ) | ( n23141 & n23378 ) ;
  assign n23380 = n9145 & n17588 ;
  assign n23381 = ( n1576 & ~n1638 ) | ( n1576 & n5612 ) | ( ~n1638 & n5612 ) ;
  assign n23382 = n23381 ^ n18846 ^ n13914 ;
  assign n23383 = n957 | n6098 ;
  assign n23384 = n23383 ^ n4890 ^ 1'b0 ;
  assign n23385 = ( n1896 & ~n1945 ) | ( n1896 & n6507 ) | ( ~n1945 & n6507 ) ;
  assign n23386 = ( n9255 & n13608 ) | ( n9255 & n23385 ) | ( n13608 & n23385 ) ;
  assign n23387 = n10990 ^ n8907 ^ 1'b0 ;
  assign n23388 = ~n23386 & n23387 ;
  assign n23389 = ( n11714 & n23384 ) | ( n11714 & ~n23388 ) | ( n23384 & ~n23388 ) ;
  assign n23390 = n12195 ^ n11322 ^ n2605 ;
  assign n23391 = n6925 & n11882 ;
  assign n23392 = ~n5325 & n23391 ;
  assign n23393 = n9279 ^ n3066 ^ 1'b0 ;
  assign n23394 = n17268 & ~n23393 ;
  assign n23395 = n17630 ^ n6596 ^ n308 ;
  assign n23396 = n23395 ^ n5512 ^ 1'b0 ;
  assign n23397 = ( n11148 & ~n20937 ) | ( n11148 & n21637 ) | ( ~n20937 & n21637 ) ;
  assign n23398 = ~n4051 & n4212 ;
  assign n23399 = ( n12076 & n13923 ) | ( n12076 & n23398 ) | ( n13923 & n23398 ) ;
  assign n23400 = ( n1739 & n4186 ) | ( n1739 & n22547 ) | ( n4186 & n22547 ) ;
  assign n23401 = n2269 & ~n21463 ;
  assign n23402 = n2270 & ~n18756 ;
  assign n23403 = ~n22762 & n23402 ;
  assign n23404 = n5715 | n23403 ;
  assign n23405 = n16629 | n23404 ;
  assign n23406 = n20030 ^ n14006 ^ n2126 ;
  assign n23407 = n23406 ^ n15359 ^ 1'b0 ;
  assign n23408 = n6764 ^ n4666 ^ 1'b0 ;
  assign n23409 = ~n4032 & n23408 ;
  assign n23410 = n17737 ^ n3373 ^ 1'b0 ;
  assign n23411 = n23409 & ~n23410 ;
  assign n23412 = n7141 & n23411 ;
  assign n23413 = ~n23407 & n23412 ;
  assign n23414 = n16816 ^ n7564 ^ 1'b0 ;
  assign n23415 = n1106 | n23414 ;
  assign n23416 = n23415 ^ n13413 ^ n7677 ;
  assign n23420 = ( n1702 & n4459 ) | ( n1702 & n8444 ) | ( n4459 & n8444 ) ;
  assign n23417 = n651 & n19515 ;
  assign n23418 = n19967 & n23417 ;
  assign n23419 = n11047 | n23418 ;
  assign n23421 = n23420 ^ n23419 ^ n14044 ;
  assign n23422 = n5020 ^ n1335 ^ 1'b0 ;
  assign n23423 = ~n8088 & n23422 ;
  assign n23424 = n23423 ^ n16411 ^ n1864 ;
  assign n23425 = ~n11159 & n15766 ;
  assign n23426 = n23425 ^ n13643 ^ n11235 ;
  assign n23427 = n16892 ^ n10535 ^ n8825 ;
  assign n23428 = ~n4429 & n8494 ;
  assign n23429 = ( ~n4587 & n21470 ) | ( ~n4587 & n23428 ) | ( n21470 & n23428 ) ;
  assign n23430 = n6392 ^ n3804 ^ 1'b0 ;
  assign n23431 = n23429 | n23430 ;
  assign n23432 = ~n13818 & n17623 ;
  assign n23433 = n23432 ^ n14789 ^ 1'b0 ;
  assign n23434 = n23433 ^ n6835 ^ 1'b0 ;
  assign n23435 = n7408 | n23434 ;
  assign n23437 = n4349 | n17077 ;
  assign n23438 = n6562 | n23437 ;
  assign n23436 = n3106 & ~n6368 ;
  assign n23439 = n23438 ^ n23436 ^ 1'b0 ;
  assign n23440 = n21885 ^ n12678 ^ n4877 ;
  assign n23441 = ( n11641 & n21926 ) | ( n11641 & n23440 ) | ( n21926 & n23440 ) ;
  assign n23442 = ( ~n7814 & n8825 ) | ( ~n7814 & n12124 ) | ( n8825 & n12124 ) ;
  assign n23443 = n2590 | n15789 ;
  assign n23444 = ( n19549 & n23442 ) | ( n19549 & n23443 ) | ( n23442 & n23443 ) ;
  assign n23445 = ( ~n6396 & n11550 ) | ( ~n6396 & n23444 ) | ( n11550 & n23444 ) ;
  assign n23446 = n16384 ^ n14662 ^ n5371 ;
  assign n23447 = n23446 ^ n21673 ^ n11784 ;
  assign n23448 = ~n1199 & n6201 ;
  assign n23449 = n5586 & n23448 ;
  assign n23450 = n20754 ^ n15328 ^ n3250 ;
  assign n23451 = ( n17145 & ~n18434 ) | ( n17145 & n23450 ) | ( ~n18434 & n23450 ) ;
  assign n23452 = ( n19512 & n23449 ) | ( n19512 & ~n23451 ) | ( n23449 & ~n23451 ) ;
  assign n23453 = n22304 ^ n12759 ^ n5385 ;
  assign n23454 = n23453 ^ n5176 ^ 1'b0 ;
  assign n23455 = ~n12621 & n23454 ;
  assign n23457 = n13805 ^ n13494 ^ n6203 ;
  assign n23458 = ( n8078 & ~n18318 ) | ( n8078 & n23457 ) | ( ~n18318 & n23457 ) ;
  assign n23459 = n23458 ^ n18491 ^ n11540 ;
  assign n23456 = ~n4422 & n10857 ;
  assign n23460 = n23459 ^ n23456 ^ 1'b0 ;
  assign n23461 = ( ~n10835 & n13133 ) | ( ~n10835 & n14402 ) | ( n13133 & n14402 ) ;
  assign n23462 = n3191 | n15228 ;
  assign n23463 = n589 & ~n23462 ;
  assign n23464 = n938 | n7171 ;
  assign n23465 = n23464 ^ n11527 ^ 1'b0 ;
  assign n23466 = ( n6865 & n23463 ) | ( n6865 & ~n23465 ) | ( n23463 & ~n23465 ) ;
  assign n23467 = ~n1987 & n6636 ;
  assign n23468 = ~n9511 & n23467 ;
  assign n23469 = n5784 | n23468 ;
  assign n23470 = n23469 ^ n17884 ^ 1'b0 ;
  assign n23471 = ~n3256 & n8081 ;
  assign n23472 = ~n21233 & n23471 ;
  assign n23473 = n23472 ^ n15049 ^ 1'b0 ;
  assign n23474 = n12717 & n13075 ;
  assign n23475 = ~n11359 & n23474 ;
  assign n23476 = ( n4988 & n22226 ) | ( n4988 & ~n23475 ) | ( n22226 & ~n23475 ) ;
  assign n23477 = ( n1239 & ~n11641 ) | ( n1239 & n15571 ) | ( ~n11641 & n15571 ) ;
  assign n23478 = n23477 ^ n2714 ^ 1'b0 ;
  assign n23479 = ( n19224 & n21983 ) | ( n19224 & ~n23478 ) | ( n21983 & ~n23478 ) ;
  assign n23480 = ( n11515 & n11642 ) | ( n11515 & ~n12702 ) | ( n11642 & ~n12702 ) ;
  assign n23481 = n23480 ^ n18218 ^ n17868 ;
  assign n23482 = ( n5594 & n9630 ) | ( n5594 & ~n14786 ) | ( n9630 & ~n14786 ) ;
  assign n23483 = n23482 ^ n5651 ^ 1'b0 ;
  assign n23484 = n23481 | n23483 ;
  assign n23485 = ~n1421 & n4383 ;
  assign n23486 = n10283 & n23485 ;
  assign n23487 = n2238 & n11735 ;
  assign n23488 = n23487 ^ n9420 ^ 1'b0 ;
  assign n23489 = n16308 | n23488 ;
  assign n23490 = n23486 & ~n23489 ;
  assign n23491 = n20308 ^ n7520 ^ 1'b0 ;
  assign n23492 = n23490 | n23491 ;
  assign n23493 = n19878 ^ n9722 ^ n753 ;
  assign n23494 = n9948 | n10646 ;
  assign n23495 = n23494 ^ n14385 ^ 1'b0 ;
  assign n23496 = x26 & n22161 ;
  assign n23497 = ( n19977 & n23495 ) | ( n19977 & n23496 ) | ( n23495 & n23496 ) ;
  assign n23498 = n23497 ^ n19840 ^ n4252 ;
  assign n23499 = n9314 ^ n7945 ^ 1'b0 ;
  assign n23500 = n3453 & ~n23499 ;
  assign n23501 = ( ~n1404 & n16086 ) | ( ~n1404 & n23500 ) | ( n16086 & n23500 ) ;
  assign n23502 = n23501 ^ n5196 ^ n1020 ;
  assign n23503 = ( ~x63 & n5896 ) | ( ~x63 & n21803 ) | ( n5896 & n21803 ) ;
  assign n23509 = ( n2384 & n8891 ) | ( n2384 & n19482 ) | ( n8891 & n19482 ) ;
  assign n23510 = ( n3742 & n5732 ) | ( n3742 & n23509 ) | ( n5732 & n23509 ) ;
  assign n23504 = ( ~n3068 & n8813 ) | ( ~n3068 & n9355 ) | ( n8813 & n9355 ) ;
  assign n23505 = n1381 & n3118 ;
  assign n23506 = n23505 ^ n4376 ^ 1'b0 ;
  assign n23507 = ( n5784 & n23504 ) | ( n5784 & ~n23506 ) | ( n23504 & ~n23506 ) ;
  assign n23508 = n23507 ^ n21486 ^ n14964 ;
  assign n23511 = n23510 ^ n23508 ^ n2672 ;
  assign n23512 = n23511 ^ n5501 ^ n1883 ;
  assign n23513 = n9386 ^ n2784 ^ n659 ;
  assign n23514 = n7375 ^ n7368 ^ n701 ;
  assign n23515 = n877 & n23514 ;
  assign n23516 = n3281 & n13387 ;
  assign n23517 = n23516 ^ n15604 ^ n12347 ;
  assign n23518 = n10475 ^ n909 ^ 1'b0 ;
  assign n23519 = n23518 ^ n15589 ^ 1'b0 ;
  assign n23520 = ~n23517 & n23519 ;
  assign n23521 = n17518 ^ n16953 ^ 1'b0 ;
  assign n23522 = n16546 | n23521 ;
  assign n23523 = n3835 ^ n2722 ^ n2624 ;
  assign n23524 = ( n11647 & n15885 ) | ( n11647 & n23523 ) | ( n15885 & n23523 ) ;
  assign n23525 = ~n23522 & n23524 ;
  assign n23526 = n12208 & n23525 ;
  assign n23527 = ( ~n3571 & n6234 ) | ( ~n3571 & n18080 ) | ( n6234 & n18080 ) ;
  assign n23528 = n6032 ^ n3185 ^ 1'b0 ;
  assign n23529 = n13393 & ~n23528 ;
  assign n23530 = ( n23310 & n23527 ) | ( n23310 & n23529 ) | ( n23527 & n23529 ) ;
  assign n23531 = n829 & n9539 ;
  assign n23532 = ( n7767 & ~n8961 ) | ( n7767 & n13604 ) | ( ~n8961 & n13604 ) ;
  assign n23533 = ( n312 & n23531 ) | ( n312 & ~n23532 ) | ( n23531 & ~n23532 ) ;
  assign n23534 = n8843 ^ n3219 ^ n195 ;
  assign n23535 = ~n3623 & n14759 ;
  assign n23536 = ( n8785 & n23482 ) | ( n8785 & n23535 ) | ( n23482 & n23535 ) ;
  assign n23537 = n16731 ^ n12409 ^ n8973 ;
  assign n23538 = ~n1545 & n19090 ;
  assign n23539 = n5552 & n9202 ;
  assign n23540 = ( n1483 & ~n6546 ) | ( n1483 & n11157 ) | ( ~n6546 & n11157 ) ;
  assign n23541 = n23540 ^ n8972 ^ n6288 ;
  assign n23542 = n8430 ^ n3938 ^ x55 ;
  assign n23543 = n11000 & n23542 ;
  assign n23544 = ~n23541 & n23543 ;
  assign n23545 = ( n4302 & ~n9966 ) | ( n4302 & n19934 ) | ( ~n9966 & n19934 ) ;
  assign n23546 = n22316 ^ n17019 ^ 1'b0 ;
  assign n23547 = n23546 ^ n12968 ^ 1'b0 ;
  assign n23548 = ~n15759 & n22977 ;
  assign n23549 = ( n5580 & n11738 ) | ( n5580 & n17534 ) | ( n11738 & n17534 ) ;
  assign n23550 = n23549 ^ n21900 ^ n17904 ;
  assign n23551 = ( x44 & n7975 ) | ( x44 & n12867 ) | ( n7975 & n12867 ) ;
  assign n23552 = n17190 & ~n23551 ;
  assign n23553 = ~n9808 & n23552 ;
  assign n23556 = n176 | n2526 ;
  assign n23554 = n1244 & n4629 ;
  assign n23555 = n6427 & n23554 ;
  assign n23557 = n23556 ^ n23555 ^ n862 ;
  assign n23558 = ( n4444 & ~n8443 ) | ( n4444 & n14704 ) | ( ~n8443 & n14704 ) ;
  assign n23559 = ~n858 & n4996 ;
  assign n23560 = n5964 ^ n3057 ^ n201 ;
  assign n23561 = n23560 ^ n19415 ^ n14537 ;
  assign n23570 = n7006 ^ n5147 ^ n4653 ;
  assign n23568 = n9064 ^ n305 ^ 1'b0 ;
  assign n23569 = n23568 ^ n13176 ^ n10974 ;
  assign n23571 = n23570 ^ n23569 ^ n400 ;
  assign n23572 = ~n3272 & n19979 ;
  assign n23573 = ~n23377 & n23572 ;
  assign n23574 = n23571 & ~n23573 ;
  assign n23575 = n23574 ^ n16429 ^ 1'b0 ;
  assign n23562 = ~n484 & n3593 ;
  assign n23563 = n22443 & n23562 ;
  assign n23564 = ( n1259 & n6338 ) | ( n1259 & ~n10950 ) | ( n6338 & ~n10950 ) ;
  assign n23565 = ( n15969 & n23563 ) | ( n15969 & ~n23564 ) | ( n23563 & ~n23564 ) ;
  assign n23566 = n23565 ^ x20 ^ 1'b0 ;
  assign n23567 = ~n16980 & n23566 ;
  assign n23576 = n23575 ^ n23567 ^ 1'b0 ;
  assign n23577 = n8729 & n23576 ;
  assign n23578 = ~n16812 & n23089 ;
  assign n23579 = ( n6118 & n12195 ) | ( n6118 & n19692 ) | ( n12195 & n19692 ) ;
  assign n23580 = n23579 ^ n11745 ^ n6910 ;
  assign n23581 = n10635 | n19144 ;
  assign n23582 = n15397 & ~n23581 ;
  assign n23583 = n23582 ^ n20201 ^ n10041 ;
  assign n23584 = ( n2109 & n2197 ) | ( n2109 & n12925 ) | ( n2197 & n12925 ) ;
  assign n23585 = n9559 ^ n5180 ^ n2044 ;
  assign n23586 = n23585 ^ n7855 ^ n1135 ;
  assign n23588 = ( n1747 & n6277 ) | ( n1747 & ~n19402 ) | ( n6277 & ~n19402 ) ;
  assign n23587 = n1738 & ~n4791 ;
  assign n23589 = n23588 ^ n23587 ^ 1'b0 ;
  assign n23590 = n8133 ^ n1542 ^ 1'b0 ;
  assign n23591 = ( ~n2977 & n23589 ) | ( ~n2977 & n23590 ) | ( n23589 & n23590 ) ;
  assign n23592 = ( n6299 & ~n7448 ) | ( n6299 & n7705 ) | ( ~n7448 & n7705 ) ;
  assign n23593 = n20092 ^ n18387 ^ n7453 ;
  assign n23594 = n19776 & n23593 ;
  assign n23595 = n23592 & n23594 ;
  assign n23596 = ( ~n3671 & n10475 ) | ( ~n3671 & n19316 ) | ( n10475 & n19316 ) ;
  assign n23597 = n6475 ^ n3014 ^ 1'b0 ;
  assign n23598 = n23596 & ~n23597 ;
  assign n23599 = n15749 ^ n6833 ^ 1'b0 ;
  assign n23600 = ~n11303 & n23599 ;
  assign n23601 = ( ~n640 & n3848 ) | ( ~n640 & n23600 ) | ( n3848 & n23600 ) ;
  assign n23602 = n23601 ^ n19142 ^ n10066 ;
  assign n23603 = ( n13210 & n17376 ) | ( n13210 & ~n17681 ) | ( n17376 & ~n17681 ) ;
  assign n23604 = n23603 ^ n12998 ^ n10339 ;
  assign n23605 = n12834 | n19793 ;
  assign n23606 = n11134 | n23605 ;
  assign n23607 = ( n10412 & n10670 ) | ( n10412 & ~n23606 ) | ( n10670 & ~n23606 ) ;
  assign n23608 = ( ~n6208 & n15749 ) | ( ~n6208 & n23607 ) | ( n15749 & n23607 ) ;
  assign n23611 = n15522 ^ n5077 ^ 1'b0 ;
  assign n23609 = n6069 ^ n4077 ^ n3494 ;
  assign n23610 = n14769 | n23609 ;
  assign n23612 = n23611 ^ n23610 ^ n3834 ;
  assign n23613 = n5035 | n17098 ;
  assign n23614 = n23613 ^ n15485 ^ 1'b0 ;
  assign n23615 = n23614 ^ n16857 ^ 1'b0 ;
  assign n23616 = n4762 & ~n17976 ;
  assign n23617 = n23616 ^ n16174 ^ 1'b0 ;
  assign n23618 = ( n3261 & ~n23269 ) | ( n3261 & n23617 ) | ( ~n23269 & n23617 ) ;
  assign n23619 = n2253 & ~n23618 ;
  assign n23620 = n12867 & n23619 ;
  assign n23621 = n22714 ^ n7756 ^ n1082 ;
  assign n23622 = ( n7122 & n10808 ) | ( n7122 & ~n18431 ) | ( n10808 & ~n18431 ) ;
  assign n23623 = ( n11700 & ~n23621 ) | ( n11700 & n23622 ) | ( ~n23621 & n23622 ) ;
  assign n23624 = ( n13872 & n14113 ) | ( n13872 & ~n23623 ) | ( n14113 & ~n23623 ) ;
  assign n23625 = n8074 & n22941 ;
  assign n23626 = n23625 ^ n18452 ^ 1'b0 ;
  assign n23627 = n10111 & n23626 ;
  assign n23629 = ( n10535 & ~n12577 ) | ( n10535 & n21207 ) | ( ~n12577 & n21207 ) ;
  assign n23628 = n16274 ^ n9892 ^ 1'b0 ;
  assign n23630 = n23629 ^ n23628 ^ n6709 ;
  assign n23631 = n15451 ^ n3982 ^ n3033 ;
  assign n23632 = n9792 ^ n4881 ^ 1'b0 ;
  assign n23633 = n17988 ^ n7380 ^ n426 ;
  assign n23634 = n23633 ^ n22291 ^ 1'b0 ;
  assign n23635 = ~n23632 & n23634 ;
  assign n23636 = n23635 ^ n14619 ^ n13391 ;
  assign n23637 = n23636 ^ n1809 ^ 1'b0 ;
  assign n23639 = n6141 ^ n2293 ^ 1'b0 ;
  assign n23638 = n16334 | n21893 ;
  assign n23640 = n23639 ^ n23638 ^ n14710 ;
  assign n23641 = n10670 ^ n9174 ^ 1'b0 ;
  assign n23642 = ~n23640 & n23641 ;
  assign n23643 = n22831 ^ n3001 ^ n1314 ;
  assign n23644 = n18128 ^ n1765 ^ 1'b0 ;
  assign n23645 = n905 & ~n23644 ;
  assign n23646 = n13919 ^ n6903 ^ 1'b0 ;
  assign n23647 = n23645 & ~n23646 ;
  assign n23648 = n23643 & n23647 ;
  assign n23649 = n7605 ^ n5254 ^ 1'b0 ;
  assign n23650 = ( n739 & ~n11568 ) | ( n739 & n23649 ) | ( ~n11568 & n23649 ) ;
  assign n23651 = n5266 ^ n2536 ^ n2029 ;
  assign n23652 = n23651 ^ n3982 ^ 1'b0 ;
  assign n23653 = ~n8529 & n23652 ;
  assign n23654 = n23653 ^ n14745 ^ n365 ;
  assign n23660 = ( x32 & n8946 ) | ( x32 & n13762 ) | ( n8946 & n13762 ) ;
  assign n23655 = n11777 ^ n5252 ^ 1'b0 ;
  assign n23656 = n23655 ^ n4308 ^ n1061 ;
  assign n23657 = n11939 & ~n16807 ;
  assign n23658 = n23656 & n23657 ;
  assign n23659 = n23658 ^ n4192 ^ 1'b0 ;
  assign n23661 = n23660 ^ n23659 ^ n3510 ;
  assign n23662 = n21415 ^ n3285 ^ 1'b0 ;
  assign n23663 = n1757 & ~n2015 ;
  assign n23664 = n23663 ^ n12675 ^ 1'b0 ;
  assign n23665 = n23313 ^ n313 ^ 1'b0 ;
  assign n23666 = ~n15155 & n23665 ;
  assign n23667 = n15811 ^ n13456 ^ n9126 ;
  assign n23668 = n23667 ^ n5307 ^ n3150 ;
  assign n23669 = n7139 ^ n3904 ^ 1'b0 ;
  assign n23670 = ( n3598 & n5949 ) | ( n3598 & n23556 ) | ( n5949 & n23556 ) ;
  assign n23671 = n23670 ^ n10583 ^ n9867 ;
  assign n23672 = ( n16711 & n23669 ) | ( n16711 & n23671 ) | ( n23669 & n23671 ) ;
  assign n23673 = n4318 | n9532 ;
  assign n23674 = n873 & ~n23673 ;
  assign n23675 = n23674 ^ n18293 ^ 1'b0 ;
  assign n23676 = n13335 & ~n23675 ;
  assign n23679 = n7718 ^ n3893 ^ n273 ;
  assign n23677 = n17091 ^ n8808 ^ n4948 ;
  assign n23678 = n23677 ^ n11275 ^ 1'b0 ;
  assign n23680 = n23679 ^ n23678 ^ n4132 ;
  assign n23681 = n1376 | n4181 ;
  assign n23682 = n4922 | n23681 ;
  assign n23683 = n3416 ^ n1277 ^ 1'b0 ;
  assign n23684 = n23682 & n23683 ;
  assign n23685 = ( n19041 & n23680 ) | ( n19041 & n23684 ) | ( n23680 & n23684 ) ;
  assign n23686 = n12453 ^ n7584 ^ n5765 ;
  assign n23687 = n713 & ~n23686 ;
  assign n23688 = n21900 & n23687 ;
  assign n23689 = n3630 | n6134 ;
  assign n23690 = n23689 ^ n20235 ^ 1'b0 ;
  assign n23691 = ( n2275 & ~n18820 ) | ( n2275 & n23690 ) | ( ~n18820 & n23690 ) ;
  assign n23693 = n5294 ^ x126 ^ 1'b0 ;
  assign n23692 = n18062 ^ n6140 ^ n467 ;
  assign n23694 = n23693 ^ n23692 ^ n8328 ;
  assign n23695 = n23694 ^ n4879 ^ 1'b0 ;
  assign n23696 = n6452 ^ n1153 ^ 1'b0 ;
  assign n23697 = n5652 & n23696 ;
  assign n23698 = ( n10130 & n14540 ) | ( n10130 & ~n22862 ) | ( n14540 & ~n22862 ) ;
  assign n23699 = ( n1129 & n18398 ) | ( n1129 & ~n23698 ) | ( n18398 & ~n23698 ) ;
  assign n23700 = ( n1640 & ~n23697 ) | ( n1640 & n23699 ) | ( ~n23697 & n23699 ) ;
  assign n23702 = ( n865 & ~n13168 ) | ( n865 & n17703 ) | ( ~n13168 & n17703 ) ;
  assign n23701 = n17319 ^ n14986 ^ 1'b0 ;
  assign n23703 = n23702 ^ n23701 ^ n13452 ;
  assign n23704 = n11646 ^ n2662 ^ 1'b0 ;
  assign n23705 = n17430 & n23429 ;
  assign n23706 = ( n16495 & n23704 ) | ( n16495 & ~n23705 ) | ( n23704 & ~n23705 ) ;
  assign n23707 = n2901 & ~n11115 ;
  assign n23708 = n23707 ^ n19507 ^ 1'b0 ;
  assign n23709 = n23708 ^ n17819 ^ n1362 ;
  assign n23710 = n20223 & n20930 ;
  assign n23711 = n23710 ^ n15947 ^ 1'b0 ;
  assign n23712 = ~n5167 & n8073 ;
  assign n23713 = n23712 ^ n4664 ^ 1'b0 ;
  assign n23714 = n23713 ^ n348 ^ 1'b0 ;
  assign n23715 = n11468 ^ n7591 ^ n2536 ;
  assign n23716 = ( n7992 & n9528 ) | ( n7992 & ~n18618 ) | ( n9528 & ~n18618 ) ;
  assign n23717 = n23716 ^ n23227 ^ n3317 ;
  assign n23718 = ( ~n1228 & n10124 ) | ( ~n1228 & n17900 ) | ( n10124 & n17900 ) ;
  assign n23719 = n12487 ^ n4377 ^ 1'b0 ;
  assign n23720 = n20084 ^ n9599 ^ 1'b0 ;
  assign n23721 = ~n20946 & n23720 ;
  assign n23722 = n23074 ^ n15037 ^ n14273 ;
  assign n23725 = n1399 & n12697 ;
  assign n23723 = n12807 ^ n10603 ^ n591 ;
  assign n23724 = ( n21393 & n21973 ) | ( n21393 & n23723 ) | ( n21973 & n23723 ) ;
  assign n23726 = n23725 ^ n23724 ^ n16932 ;
  assign n23730 = n7034 ^ n151 ^ 1'b0 ;
  assign n23731 = n480 & ~n23730 ;
  assign n23727 = n3994 ^ n3592 ^ n892 ;
  assign n23728 = n23727 ^ n13538 ^ n8261 ;
  assign n23729 = n23728 ^ n10549 ^ 1'b0 ;
  assign n23732 = n23731 ^ n23729 ^ n6116 ;
  assign n23733 = ( n1668 & ~n10053 ) | ( n1668 & n11303 ) | ( ~n10053 & n11303 ) ;
  assign n23734 = n10579 ^ n6779 ^ n1130 ;
  assign n23735 = ( x15 & ~x94 ) | ( x15 & n9805 ) | ( ~x94 & n9805 ) ;
  assign n23736 = ( n23733 & n23734 ) | ( n23733 & ~n23735 ) | ( n23734 & ~n23735 ) ;
  assign n23737 = n23736 ^ n17616 ^ n16467 ;
  assign n23738 = ( n2292 & n5053 ) | ( n2292 & n8651 ) | ( n5053 & n8651 ) ;
  assign n23739 = ( n5707 & n16439 ) | ( n5707 & ~n23738 ) | ( n16439 & ~n23738 ) ;
  assign n23740 = ~n4447 & n23739 ;
  assign n23741 = n23740 ^ n13040 ^ 1'b0 ;
  assign n23742 = ( n9648 & n17519 ) | ( n9648 & n23741 ) | ( n17519 & n23741 ) ;
  assign n23743 = n8608 ^ n4386 ^ n434 ;
  assign n23744 = n19885 & n23743 ;
  assign n23746 = ( n6114 & n13021 ) | ( n6114 & n19785 ) | ( n13021 & n19785 ) ;
  assign n23745 = n3316 & n17763 ;
  assign n23747 = n23746 ^ n23745 ^ 1'b0 ;
  assign n23748 = ( n9599 & ~n10313 ) | ( n9599 & n20801 ) | ( ~n10313 & n20801 ) ;
  assign n23749 = n7290 | n23748 ;
  assign n23750 = n17665 ^ n14059 ^ n1221 ;
  assign n23751 = n6305 ^ n810 ^ 1'b0 ;
  assign n23752 = n23750 & ~n23751 ;
  assign n23753 = n460 & ~n1587 ;
  assign n23754 = ( ~n3931 & n15387 ) | ( ~n3931 & n15576 ) | ( n15387 & n15576 ) ;
  assign n23755 = n13565 ^ n4202 ^ 1'b0 ;
  assign n23756 = ( ~n4022 & n23754 ) | ( ~n4022 & n23755 ) | ( n23754 & n23755 ) ;
  assign n23757 = n12034 ^ n4269 ^ 1'b0 ;
  assign n23761 = ( ~x32 & n12523 ) | ( ~x32 & n16781 ) | ( n12523 & n16781 ) ;
  assign n23758 = n5716 & ~n16888 ;
  assign n23759 = n23758 ^ n10195 ^ n7029 ;
  assign n23760 = n17172 | n23759 ;
  assign n23762 = n23761 ^ n23760 ^ 1'b0 ;
  assign n23763 = ( n2762 & n3530 ) | ( n2762 & ~n19695 ) | ( n3530 & ~n19695 ) ;
  assign n23764 = ( n1856 & ~n5918 ) | ( n1856 & n23763 ) | ( ~n5918 & n23763 ) ;
  assign n23765 = n23764 ^ n8377 ^ 1'b0 ;
  assign n23766 = n12365 & ~n23765 ;
  assign n23767 = ( n5539 & n6805 ) | ( n5539 & n10701 ) | ( n6805 & n10701 ) ;
  assign n23768 = ( n9126 & n14463 ) | ( n9126 & ~n23767 ) | ( n14463 & ~n23767 ) ;
  assign n23769 = n18938 ^ n8040 ^ n3384 ;
  assign n23770 = n23769 ^ n8278 ^ n931 ;
  assign n23771 = ( n4104 & n23768 ) | ( n4104 & ~n23770 ) | ( n23768 & ~n23770 ) ;
  assign n23772 = n23771 ^ n9831 ^ n3040 ;
  assign n23773 = n10246 | n23772 ;
  assign n23774 = n6181 & ~n23773 ;
  assign n23775 = n7577 ^ n1517 ^ 1'b0 ;
  assign n23776 = n2113 | n23775 ;
  assign n23777 = n4467 & n23776 ;
  assign n23780 = n15631 ^ n2121 ^ n265 ;
  assign n23778 = n18746 ^ n374 ^ 1'b0 ;
  assign n23779 = ~n13673 & n23778 ;
  assign n23781 = n23780 ^ n23779 ^ n13011 ;
  assign n23782 = n7406 ^ n3699 ^ n496 ;
  assign n23783 = n23782 ^ n9746 ^ n4689 ;
  assign n23784 = ( ~n2849 & n11760 ) | ( ~n2849 & n23783 ) | ( n11760 & n23783 ) ;
  assign n23788 = n18592 ^ n6408 ^ 1'b0 ;
  assign n23789 = ~n6427 & n23788 ;
  assign n23785 = n11837 ^ n10568 ^ n4568 ;
  assign n23786 = n5594 & n7768 ;
  assign n23787 = ~n23785 & n23786 ;
  assign n23790 = n23789 ^ n23787 ^ n9672 ;
  assign n23791 = ~n10389 & n23790 ;
  assign n23792 = n9511 ^ n7380 ^ n1261 ;
  assign n23793 = n4862 ^ n4199 ^ 1'b0 ;
  assign n23794 = n23792 & ~n23793 ;
  assign n23795 = n5198 | n12789 ;
  assign n23796 = n23795 ^ n12411 ^ 1'b0 ;
  assign n23797 = n12280 ^ n9200 ^ 1'b0 ;
  assign n23798 = n21103 | n23797 ;
  assign n23799 = n11005 ^ n1195 ^ 1'b0 ;
  assign n23800 = ( ~n9475 & n10919 ) | ( ~n9475 & n18493 ) | ( n10919 & n18493 ) ;
  assign n23801 = n23800 ^ n18823 ^ n10391 ;
  assign n23802 = ( n10486 & n14300 ) | ( n10486 & n17127 ) | ( n14300 & n17127 ) ;
  assign n23803 = n23802 ^ n18623 ^ n15593 ;
  assign n23804 = n6510 ^ n5272 ^ x3 ;
  assign n23805 = n23804 ^ n6574 ^ 1'b0 ;
  assign n23806 = n5284 | n23805 ;
  assign n23807 = n23806 ^ n16683 ^ n3098 ;
  assign n23811 = n4788 | n16938 ;
  assign n23812 = n23811 ^ n4422 ^ 1'b0 ;
  assign n23813 = n23812 ^ n9105 ^ n2738 ;
  assign n23808 = ( ~n6440 & n9536 ) | ( ~n6440 & n9937 ) | ( n9536 & n9937 ) ;
  assign n23809 = n23808 ^ n11684 ^ 1'b0 ;
  assign n23810 = ~n8855 & n23809 ;
  assign n23814 = n23813 ^ n23810 ^ n17618 ;
  assign n23815 = n2588 ^ n2489 ^ 1'b0 ;
  assign n23816 = n17155 & n19948 ;
  assign n23817 = ( n827 & n4095 ) | ( n827 & ~n15017 ) | ( n4095 & ~n15017 ) ;
  assign n23818 = n23817 ^ n8448 ^ n3005 ;
  assign n23819 = n19330 ^ n7202 ^ n1459 ;
  assign n23822 = ( ~n9231 & n15270 ) | ( ~n9231 & n16917 ) | ( n15270 & n16917 ) ;
  assign n23823 = n18044 | n23822 ;
  assign n23824 = n23823 ^ n23245 ^ 1'b0 ;
  assign n23820 = ( n777 & n4353 ) | ( n777 & ~n12565 ) | ( n4353 & ~n12565 ) ;
  assign n23821 = ( n2036 & n11133 ) | ( n2036 & n23820 ) | ( n11133 & n23820 ) ;
  assign n23825 = n23824 ^ n23821 ^ 1'b0 ;
  assign n23826 = n4134 ^ n2846 ^ n562 ;
  assign n23827 = n176 & n23826 ;
  assign n23828 = ( n8315 & n18451 ) | ( n8315 & ~n23827 ) | ( n18451 & ~n23827 ) ;
  assign n23829 = n4719 & n17086 ;
  assign n23830 = n23829 ^ n12612 ^ 1'b0 ;
  assign n23831 = n8823 ^ n8028 ^ n7953 ;
  assign n23832 = n23831 ^ n8516 ^ 1'b0 ;
  assign n23833 = ( n1299 & n1908 ) | ( n1299 & ~n23792 ) | ( n1908 & ~n23792 ) ;
  assign n23834 = n23833 ^ n11915 ^ 1'b0 ;
  assign n23835 = n23834 ^ n15594 ^ 1'b0 ;
  assign n23836 = n6114 & ~n23835 ;
  assign n23837 = n23836 ^ n15498 ^ n11476 ;
  assign n23839 = ( x69 & n9426 ) | ( x69 & ~n13447 ) | ( n9426 & ~n13447 ) ;
  assign n23838 = n23131 ^ n8363 ^ 1'b0 ;
  assign n23840 = n23839 ^ n23838 ^ n17554 ;
  assign n23841 = ( ~n11303 & n11584 ) | ( ~n11303 & n17943 ) | ( n11584 & n17943 ) ;
  assign n23842 = n6130 ^ n1099 ^ x114 ;
  assign n23843 = n13299 ^ n10766 ^ n3376 ;
  assign n23844 = ( n4555 & n8168 ) | ( n4555 & ~n10201 ) | ( n8168 & ~n10201 ) ;
  assign n23845 = n23070 ^ n11063 ^ 1'b0 ;
  assign n23846 = n23844 & n23845 ;
  assign n23847 = ( n1542 & ~n2503 ) | ( n1542 & n7295 ) | ( ~n2503 & n7295 ) ;
  assign n23848 = ~n4720 & n23847 ;
  assign n23849 = ~n8132 & n23848 ;
  assign n23850 = n11237 | n23849 ;
  assign n23851 = n2305 & ~n23850 ;
  assign n23853 = n5962 & n10003 ;
  assign n23854 = ~n12881 & n23853 ;
  assign n23852 = n10559 | n19875 ;
  assign n23855 = n23854 ^ n23852 ^ 1'b0 ;
  assign n23856 = ( n423 & ~n620 ) | ( n423 & n15777 ) | ( ~n620 & n15777 ) ;
  assign n23857 = n21106 & ~n23856 ;
  assign n23864 = ( n1745 & n17224 ) | ( n1745 & ~n18220 ) | ( n17224 & ~n18220 ) ;
  assign n23865 = n23864 ^ n6080 ^ n2973 ;
  assign n23858 = n5549 ^ n5353 ^ 1'b0 ;
  assign n23860 = ~n553 & n16803 ;
  assign n23859 = n15986 ^ n5632 ^ n3130 ;
  assign n23861 = n23860 ^ n23859 ^ 1'b0 ;
  assign n23862 = n23858 & ~n23861 ;
  assign n23863 = ( ~n7459 & n21900 ) | ( ~n7459 & n23862 ) | ( n21900 & n23862 ) ;
  assign n23866 = n23865 ^ n23863 ^ n2546 ;
  assign n23867 = ( ~n265 & n8585 ) | ( ~n265 & n17116 ) | ( n8585 & n17116 ) ;
  assign n23868 = n23867 ^ n2408 ^ 1'b0 ;
  assign n23869 = n20830 ^ n14901 ^ 1'b0 ;
  assign n23870 = n7262 | n23869 ;
  assign n23871 = ( n414 & n7040 ) | ( n414 & ~n12598 ) | ( n7040 & ~n12598 ) ;
  assign n23872 = n17538 ^ n6967 ^ n5520 ;
  assign n23873 = n23872 ^ n21453 ^ n6202 ;
  assign n23874 = ( ~n2449 & n5896 ) | ( ~n2449 & n22693 ) | ( n5896 & n22693 ) ;
  assign n23875 = n23874 ^ n22559 ^ n20844 ;
  assign n23876 = n14269 ^ n6181 ^ n1775 ;
  assign n23879 = n8128 | n17239 ;
  assign n23880 = ( ~n4812 & n8180 ) | ( ~n4812 & n23879 ) | ( n8180 & n23879 ) ;
  assign n23881 = ( n10605 & n18646 ) | ( n10605 & n23880 ) | ( n18646 & n23880 ) ;
  assign n23877 = n15989 ^ n3820 ^ n2658 ;
  assign n23878 = ( n16685 & ~n17273 ) | ( n16685 & n23877 ) | ( ~n17273 & n23877 ) ;
  assign n23882 = n23881 ^ n23878 ^ 1'b0 ;
  assign n23888 = n1476 & n3786 ;
  assign n23883 = n2406 ^ n355 ^ 1'b0 ;
  assign n23884 = n2377 | n23883 ;
  assign n23885 = n14443 ^ n6430 ^ n1148 ;
  assign n23886 = n12030 & n23885 ;
  assign n23887 = n23884 & n23886 ;
  assign n23889 = n23888 ^ n23887 ^ n17778 ;
  assign n23890 = n14467 | n23889 ;
  assign n23891 = n7763 & ~n13011 ;
  assign n23892 = ~n5129 & n23891 ;
  assign n23893 = n23892 ^ n20110 ^ n3354 ;
  assign n23894 = n17000 ^ n15396 ^ n7401 ;
  assign n23895 = n4804 | n23894 ;
  assign n23896 = n5265 & n5843 ;
  assign n23897 = n23896 ^ n2315 ^ 1'b0 ;
  assign n23898 = n16549 ^ n15647 ^ 1'b0 ;
  assign n23899 = ~n23897 & n23898 ;
  assign n23900 = ( n4095 & ~n6428 ) | ( n4095 & n22592 ) | ( ~n6428 & n22592 ) ;
  assign n23901 = ( n6839 & n23899 ) | ( n6839 & ~n23900 ) | ( n23899 & ~n23900 ) ;
  assign n23902 = ( n7370 & n11359 ) | ( n7370 & n23901 ) | ( n11359 & n23901 ) ;
  assign n23903 = n7343 ^ n312 ^ 1'b0 ;
  assign n23904 = ~n13653 & n23903 ;
  assign n23905 = n5979 & n16782 ;
  assign n23906 = n20396 & n23905 ;
  assign n23907 = ( n3617 & n10805 ) | ( n3617 & n21991 ) | ( n10805 & n21991 ) ;
  assign n23908 = n23907 ^ n18335 ^ n9501 ;
  assign n23909 = n10102 ^ n2236 ^ 1'b0 ;
  assign n23910 = ( ~n923 & n5144 ) | ( ~n923 & n12840 ) | ( n5144 & n12840 ) ;
  assign n23911 = n4649 ^ n170 ^ 1'b0 ;
  assign n23912 = n11589 ^ n9717 ^ n1009 ;
  assign n23913 = n23912 ^ n15525 ^ n5253 ;
  assign n23914 = n12270 ^ n9951 ^ 1'b0 ;
  assign n23915 = n13332 ^ n6047 ^ 1'b0 ;
  assign n23916 = ~n19702 & n23915 ;
  assign n23917 = n17943 ^ n4515 ^ 1'b0 ;
  assign n23918 = ( n1478 & ~n6000 ) | ( n1478 & n16310 ) | ( ~n6000 & n16310 ) ;
  assign n23919 = n5272 ^ n4177 ^ n738 ;
  assign n23920 = n23919 ^ n12935 ^ n2054 ;
  assign n23921 = n23920 ^ n12862 ^ n3544 ;
  assign n23922 = n19031 ^ n17530 ^ n2349 ;
  assign n23923 = ( n2348 & n23680 ) | ( n2348 & ~n23922 ) | ( n23680 & ~n23922 ) ;
  assign n23924 = n16654 ^ n6396 ^ n5771 ;
  assign n23925 = n17558 ^ n8726 ^ 1'b0 ;
  assign n23926 = n23924 | n23925 ;
  assign n23927 = n5201 & n12238 ;
  assign n23928 = ~n5243 & n23927 ;
  assign n23929 = ( n18521 & ~n23926 ) | ( n18521 & n23928 ) | ( ~n23926 & n23928 ) ;
  assign n23930 = n19942 ^ n11764 ^ n6324 ;
  assign n23931 = n21879 ^ n3757 ^ 1'b0 ;
  assign n23932 = n7383 | n23931 ;
  assign n23933 = n16274 ^ n10681 ^ n1345 ;
  assign n23934 = n18268 | n23933 ;
  assign n23935 = ~n2271 & n4191 ;
  assign n23936 = n9749 & n23935 ;
  assign n23937 = n1268 & n15877 ;
  assign n23938 = n16111 ^ n13038 ^ 1'b0 ;
  assign n23939 = n19233 ^ n9771 ^ 1'b0 ;
  assign n23943 = n723 & n23120 ;
  assign n23944 = ~n1913 & n23943 ;
  assign n23940 = n3144 & ~n6494 ;
  assign n23941 = ( n13959 & n23120 ) | ( n13959 & n23940 ) | ( n23120 & n23940 ) ;
  assign n23942 = n23941 ^ n2969 ^ 1'b0 ;
  assign n23945 = n23944 ^ n23942 ^ n14196 ;
  assign n23946 = n23033 ^ n9767 ^ n4232 ;
  assign n23947 = n11460 ^ n8350 ^ 1'b0 ;
  assign n23948 = ~n4933 & n23947 ;
  assign n23949 = n5253 & ~n23948 ;
  assign n23950 = ~n3173 & n23949 ;
  assign n23951 = ( n858 & n5507 ) | ( n858 & n8211 ) | ( n5507 & n8211 ) ;
  assign n23952 = n23201 ^ n13321 ^ n12877 ;
  assign n23953 = ( n18019 & ~n23951 ) | ( n18019 & n23952 ) | ( ~n23951 & n23952 ) ;
  assign n23954 = n21635 ^ n20946 ^ n12788 ;
  assign n23955 = n10946 ^ n3881 ^ 1'b0 ;
  assign n23956 = n4417 & ~n23955 ;
  assign n23957 = n23956 ^ n7572 ^ n6413 ;
  assign n23958 = n15248 & n23957 ;
  assign n23959 = n23958 ^ n12588 ^ n1074 ;
  assign n23960 = n7350 & n12548 ;
  assign n23961 = ~n1247 & n23960 ;
  assign n23962 = n3281 | n12643 ;
  assign n23963 = n23962 ^ n11363 ^ 1'b0 ;
  assign n23964 = ~n6215 & n17640 ;
  assign n23965 = n23964 ^ n4857 ^ 1'b0 ;
  assign n23966 = ( ~n23961 & n23963 ) | ( ~n23961 & n23965 ) | ( n23963 & n23965 ) ;
  assign n23967 = n18057 ^ n17835 ^ n16948 ;
  assign n23968 = n23967 ^ n19441 ^ 1'b0 ;
  assign n23973 = n10130 ^ n2780 ^ n1114 ;
  assign n23969 = ~n496 & n11269 ;
  assign n23970 = ( ~n4020 & n15710 ) | ( ~n4020 & n23969 ) | ( n15710 & n23969 ) ;
  assign n23971 = ( n7894 & n8154 ) | ( n7894 & n18905 ) | ( n8154 & n18905 ) ;
  assign n23972 = n23970 | n23971 ;
  assign n23974 = n23973 ^ n23972 ^ 1'b0 ;
  assign n23975 = n1657 & n4265 ;
  assign n23976 = n23975 ^ n10120 ^ 1'b0 ;
  assign n23977 = ( n3173 & n3691 ) | ( n3173 & n7448 ) | ( n3691 & n7448 ) ;
  assign n23978 = ( n581 & ~n3680 ) | ( n581 & n21616 ) | ( ~n3680 & n21616 ) ;
  assign n23979 = n4798 | n11552 ;
  assign n23980 = n23979 ^ n16144 ^ 1'b0 ;
  assign n23981 = ( n6297 & n13479 ) | ( n6297 & n23980 ) | ( n13479 & n23980 ) ;
  assign n23982 = ( n9464 & ~n11488 ) | ( n9464 & n19101 ) | ( ~n11488 & n19101 ) ;
  assign n23983 = n10594 ^ n9346 ^ 1'b0 ;
  assign n23986 = n5313 & n9808 ;
  assign n23987 = n3798 & n23986 ;
  assign n23988 = n20162 & ~n23213 ;
  assign n23989 = n23987 & n23988 ;
  assign n23984 = ~n735 & n14927 ;
  assign n23985 = ~n485 & n23984 ;
  assign n23990 = n23989 ^ n23985 ^ n19112 ;
  assign n23991 = ( n7152 & n11235 ) | ( n7152 & n20862 ) | ( n11235 & n20862 ) ;
  assign n23994 = ( n1454 & n1729 ) | ( n1454 & n6531 ) | ( n1729 & n6531 ) ;
  assign n23992 = x92 & ~n5172 ;
  assign n23993 = ~n23645 & n23992 ;
  assign n23995 = n23994 ^ n23993 ^ 1'b0 ;
  assign n23996 = ( ~n6935 & n8298 ) | ( ~n6935 & n23995 ) | ( n8298 & n23995 ) ;
  assign n23997 = ( n3710 & n23991 ) | ( n3710 & ~n23996 ) | ( n23991 & ~n23996 ) ;
  assign n23998 = n1612 & ~n9558 ;
  assign n23999 = n8966 | n23998 ;
  assign n24000 = n11204 | n23999 ;
  assign n24001 = ( n5359 & ~n14302 ) | ( n5359 & n24000 ) | ( ~n14302 & n24000 ) ;
  assign n24002 = ( ~n3489 & n4101 ) | ( ~n3489 & n24001 ) | ( n4101 & n24001 ) ;
  assign n24003 = ( n3880 & ~n13154 ) | ( n3880 & n24002 ) | ( ~n13154 & n24002 ) ;
  assign n24004 = n5859 & n24003 ;
  assign n24005 = n24004 ^ n14258 ^ 1'b0 ;
  assign n24006 = ( ~n4655 & n8576 ) | ( ~n4655 & n20610 ) | ( n8576 & n20610 ) ;
  assign n24007 = n15783 ^ n2401 ^ n1616 ;
  assign n24008 = ( n6432 & n17542 ) | ( n6432 & n24007 ) | ( n17542 & n24007 ) ;
  assign n24009 = n24008 ^ n19395 ^ n16637 ;
  assign n24010 = n24009 ^ n1258 ^ 1'b0 ;
  assign n24011 = n24006 & n24010 ;
  assign n24012 = n4525 | n10288 ;
  assign n24013 = n24012 ^ n3423 ^ 1'b0 ;
  assign n24014 = n5986 & ~n19861 ;
  assign n24015 = n14753 ^ n7097 ^ n1327 ;
  assign n24016 = n24015 ^ n14627 ^ 1'b0 ;
  assign n24017 = n24014 & ~n24016 ;
  assign n24018 = ( n19842 & ~n24013 ) | ( n19842 & n24017 ) | ( ~n24013 & n24017 ) ;
  assign n24019 = ( n3814 & ~n4000 ) | ( n3814 & n13991 ) | ( ~n4000 & n13991 ) ;
  assign n24020 = n13147 ^ n4957 ^ n2340 ;
  assign n24021 = n24020 ^ n20266 ^ n5438 ;
  assign n24022 = ( n2798 & ~n8469 ) | ( n2798 & n16336 ) | ( ~n8469 & n16336 ) ;
  assign n24023 = n1685 | n18330 ;
  assign n24024 = ( n9672 & n12057 ) | ( n9672 & ~n24023 ) | ( n12057 & ~n24023 ) ;
  assign n24025 = n11460 | n16384 ;
  assign n24026 = n24025 ^ n14762 ^ 1'b0 ;
  assign n24027 = ~n10262 & n10476 ;
  assign n24028 = n322 & ~n3049 ;
  assign n24029 = n24028 ^ n8095 ^ 1'b0 ;
  assign n24030 = n24029 ^ n10954 ^ 1'b0 ;
  assign n24031 = n11656 ^ n6310 ^ 1'b0 ;
  assign n24032 = n24030 | n24031 ;
  assign n24033 = ( ~n4581 & n24027 ) | ( ~n4581 & n24032 ) | ( n24027 & n24032 ) ;
  assign n24034 = n19938 ^ n7922 ^ n7355 ;
  assign n24035 = n1264 ^ n768 ^ 1'b0 ;
  assign n24036 = n9388 | n24035 ;
  assign n24037 = ( n15507 & n19433 ) | ( n15507 & ~n24036 ) | ( n19433 & ~n24036 ) ;
  assign n24038 = ( n21742 & ~n22876 ) | ( n21742 & n24037 ) | ( ~n22876 & n24037 ) ;
  assign n24041 = n13078 ^ n4151 ^ n3269 ;
  assign n24042 = n14059 & n24041 ;
  assign n24043 = ( n3266 & ~n13907 ) | ( n3266 & n24042 ) | ( ~n13907 & n24042 ) ;
  assign n24039 = ( n5233 & ~n8430 ) | ( n5233 & n18049 ) | ( ~n8430 & n18049 ) ;
  assign n24040 = n8284 & ~n24039 ;
  assign n24044 = n24043 ^ n24040 ^ n10449 ;
  assign n24045 = n16716 & n23301 ;
  assign n24046 = n21061 ^ n8681 ^ n7584 ;
  assign n24047 = ( n13463 & ~n24045 ) | ( n13463 & n24046 ) | ( ~n24045 & n24046 ) ;
  assign n24048 = n923 | n21627 ;
  assign n24050 = ( ~n2613 & n6984 ) | ( ~n2613 & n16624 ) | ( n6984 & n16624 ) ;
  assign n24049 = ( ~n11620 & n18503 ) | ( ~n11620 & n21015 ) | ( n18503 & n21015 ) ;
  assign n24051 = n24050 ^ n24049 ^ n15811 ;
  assign n24052 = n2583 & ~n9394 ;
  assign n24053 = n24052 ^ n6530 ^ 1'b0 ;
  assign n24054 = n10229 ^ n9802 ^ n9475 ;
  assign n24055 = n24054 ^ n17097 ^ 1'b0 ;
  assign n24056 = n19199 & n24055 ;
  assign n24057 = ( n4381 & ~n4486 ) | ( n4381 & n11530 ) | ( ~n4486 & n11530 ) ;
  assign n24058 = n13751 ^ n7815 ^ n2759 ;
  assign n24059 = n7351 ^ n4629 ^ 1'b0 ;
  assign n24060 = ( n1748 & n2118 ) | ( n1748 & n24059 ) | ( n2118 & n24059 ) ;
  assign n24061 = n8777 ^ n918 ^ 1'b0 ;
  assign n24062 = ( n24058 & ~n24060 ) | ( n24058 & n24061 ) | ( ~n24060 & n24061 ) ;
  assign n24063 = n23081 ^ n11270 ^ n1476 ;
  assign n24064 = n14323 & n21653 ;
  assign n24065 = ~n24063 & n24064 ;
  assign n24066 = n24065 ^ n14273 ^ n10365 ;
  assign n24067 = ( n10937 & ~n11741 ) | ( n10937 & n14973 ) | ( ~n11741 & n14973 ) ;
  assign n24068 = ( n6413 & ~n12469 ) | ( n6413 & n24067 ) | ( ~n12469 & n24067 ) ;
  assign n24069 = ( ~n3220 & n22426 ) | ( ~n3220 & n24068 ) | ( n22426 & n24068 ) ;
  assign n24070 = n337 & n14046 ;
  assign n24071 = n24070 ^ n19294 ^ n14661 ;
  assign n24072 = n9952 ^ n7275 ^ n5009 ;
  assign n24073 = n9627 & ~n21370 ;
  assign n24074 = n11337 & n24073 ;
  assign n24075 = ( n7412 & ~n8183 ) | ( n7412 & n12770 ) | ( ~n8183 & n12770 ) ;
  assign n24076 = n6247 ^ n143 ^ 1'b0 ;
  assign n24077 = n11159 | n24076 ;
  assign n24078 = n5963 | n24077 ;
  assign n24079 = ~n8653 & n23409 ;
  assign n24080 = n24079 ^ n10282 ^ 1'b0 ;
  assign n24081 = ( n3667 & n12231 ) | ( n3667 & n24080 ) | ( n12231 & n24080 ) ;
  assign n24082 = n12830 | n16905 ;
  assign n24083 = n2900 | n3298 ;
  assign n24084 = ~n14639 & n24083 ;
  assign n24085 = n1287 | n3485 ;
  assign n24086 = n15320 | n24085 ;
  assign n24087 = ( n2605 & n5541 ) | ( n2605 & ~n15697 ) | ( n5541 & ~n15697 ) ;
  assign n24088 = n19434 ^ n4074 ^ 1'b0 ;
  assign n24089 = ( n639 & ~n13480 ) | ( n639 & n24088 ) | ( ~n13480 & n24088 ) ;
  assign n24090 = n12027 & n14973 ;
  assign n24091 = n3443 & n24090 ;
  assign n24092 = n24091 ^ n5509 ^ 1'b0 ;
  assign n24102 = n17452 ^ n13049 ^ n3581 ;
  assign n24101 = n1687 & ~n23247 ;
  assign n24093 = ( x108 & n4405 ) | ( x108 & n8816 ) | ( n4405 & n8816 ) ;
  assign n24094 = n17986 ^ n16216 ^ 1'b0 ;
  assign n24095 = n23153 | n24094 ;
  assign n24096 = n24095 ^ n18691 ^ n13953 ;
  assign n24097 = n8659 ^ n4617 ^ 1'b0 ;
  assign n24098 = ~n1899 & n18025 ;
  assign n24099 = n24097 & n24098 ;
  assign n24100 = ( n24093 & n24096 ) | ( n24093 & n24099 ) | ( n24096 & n24099 ) ;
  assign n24103 = n24102 ^ n24101 ^ n24100 ;
  assign n24104 = n18813 ^ n12173 ^ n2094 ;
  assign n24107 = n23285 ^ n9419 ^ n160 ;
  assign n24105 = n12015 ^ n4437 ^ n703 ;
  assign n24106 = n24105 ^ n9586 ^ n6252 ;
  assign n24108 = n24107 ^ n24106 ^ n6153 ;
  assign n24109 = n13075 & n24003 ;
  assign n24110 = ~n17496 & n24109 ;
  assign n24111 = n12098 ^ n10269 ^ n847 ;
  assign n24112 = ( ~n6324 & n10697 ) | ( ~n6324 & n24111 ) | ( n10697 & n24111 ) ;
  assign n24113 = n24112 ^ n3364 ^ 1'b0 ;
  assign n24114 = n22190 & n24113 ;
  assign n24115 = n16844 ^ n8350 ^ n3652 ;
  assign n24116 = n21854 ^ n18280 ^ n6425 ;
  assign n24117 = ~n18526 & n24116 ;
  assign n24118 = n24115 & n24117 ;
  assign n24120 = n6580 | n17917 ;
  assign n24119 = n15061 ^ n6898 ^ 1'b0 ;
  assign n24121 = n24120 ^ n24119 ^ n6445 ;
  assign n24126 = n12903 ^ n8797 ^ 1'b0 ;
  assign n24127 = n14695 & ~n24126 ;
  assign n24122 = ( n4367 & n10690 ) | ( n4367 & ~n11832 ) | ( n10690 & ~n11832 ) ;
  assign n24123 = n24122 ^ n19380 ^ n8698 ;
  assign n24124 = n15862 | n24123 ;
  assign n24125 = n24124 ^ n15046 ^ 1'b0 ;
  assign n24128 = n24127 ^ n24125 ^ n9296 ;
  assign n24129 = ( ~n6018 & n14148 ) | ( ~n6018 & n16264 ) | ( n14148 & n16264 ) ;
  assign n24130 = n16844 ^ n8170 ^ n4497 ;
  assign n24131 = n5898 & ~n14618 ;
  assign n24132 = ~n24130 & n24131 ;
  assign n24133 = ( n4259 & ~n18451 ) | ( n4259 & n24132 ) | ( ~n18451 & n24132 ) ;
  assign n24134 = ( n5885 & n12697 ) | ( n5885 & ~n24133 ) | ( n12697 & ~n24133 ) ;
  assign n24136 = n13529 ^ n12260 ^ n4914 ;
  assign n24135 = ( n10238 & n13300 ) | ( n10238 & ~n22649 ) | ( n13300 & ~n22649 ) ;
  assign n24137 = n24136 ^ n24135 ^ 1'b0 ;
  assign n24138 = n14560 & ~n16981 ;
  assign n24139 = ~n8385 & n8658 ;
  assign n24140 = n23007 ^ n6498 ^ 1'b0 ;
  assign n24141 = x9 & n243 ;
  assign n24142 = n4037 & n16719 ;
  assign n24143 = n7405 & ~n9395 ;
  assign n24144 = n24142 & n24143 ;
  assign n24145 = ( n2163 & n11508 ) | ( n2163 & ~n24144 ) | ( n11508 & ~n24144 ) ;
  assign n24149 = n5216 | n11494 ;
  assign n24150 = n24149 ^ n18240 ^ 1'b0 ;
  assign n24151 = n4445 & ~n24150 ;
  assign n24146 = n4212 ^ n816 ^ 1'b0 ;
  assign n24147 = n20234 & ~n24146 ;
  assign n24148 = ( ~n4348 & n5877 ) | ( ~n4348 & n24147 ) | ( n5877 & n24147 ) ;
  assign n24152 = n24151 ^ n24148 ^ n16935 ;
  assign n24153 = n19937 ^ n11742 ^ n3276 ;
  assign n24154 = ~n15218 & n24153 ;
  assign n24155 = n20255 ^ n17311 ^ n2878 ;
  assign n24156 = n7246 & ~n22529 ;
  assign n24157 = n24156 ^ n10590 ^ 1'b0 ;
  assign n24158 = ( n12364 & n22372 ) | ( n12364 & n24157 ) | ( n22372 & n24157 ) ;
  assign n24159 = n214 & n3379 ;
  assign n24160 = ( n3765 & ~n17945 ) | ( n3765 & n20201 ) | ( ~n17945 & n20201 ) ;
  assign n24161 = ( n5624 & n24159 ) | ( n5624 & n24160 ) | ( n24159 & n24160 ) ;
  assign n24162 = ( n1910 & ~n8127 ) | ( n1910 & n11789 ) | ( ~n8127 & n11789 ) ;
  assign n24163 = n24162 ^ n995 ^ 1'b0 ;
  assign n24164 = n21036 ^ n1259 ^ 1'b0 ;
  assign n24165 = ~n1067 & n24164 ;
  assign n24166 = n24165 ^ n6125 ^ 1'b0 ;
  assign n24167 = ( n2175 & n4973 ) | ( n2175 & n17340 ) | ( n4973 & n17340 ) ;
  assign n24168 = n5466 & ~n24167 ;
  assign n24169 = n24168 ^ n1573 ^ 1'b0 ;
  assign n24170 = n16351 ^ n3407 ^ 1'b0 ;
  assign n24171 = n13632 & n24170 ;
  assign n24172 = ~n19815 & n24171 ;
  assign n24173 = ~n923 & n17161 ;
  assign n24174 = ~n10267 & n24173 ;
  assign n24175 = ( n7344 & n13248 ) | ( n7344 & n24174 ) | ( n13248 & n24174 ) ;
  assign n24176 = n24175 ^ n10732 ^ n8565 ;
  assign n24177 = ~n4386 & n8985 ;
  assign n24178 = n3073 & n24177 ;
  assign n24179 = n4524 ^ n3761 ^ 1'b0 ;
  assign n24180 = n24178 | n24179 ;
  assign n24181 = n7820 ^ n2745 ^ 1'b0 ;
  assign n24182 = n9689 | n24181 ;
  assign n24183 = ( n723 & n10521 ) | ( n723 & n24182 ) | ( n10521 & n24182 ) ;
  assign n24184 = ( n20329 & ~n24180 ) | ( n20329 & n24183 ) | ( ~n24180 & n24183 ) ;
  assign n24185 = ( n6764 & n8153 ) | ( n6764 & n13983 ) | ( n8153 & n13983 ) ;
  assign n24186 = ( n15439 & ~n15873 ) | ( n15439 & n24185 ) | ( ~n15873 & n24185 ) ;
  assign n24187 = ( n24176 & n24184 ) | ( n24176 & n24186 ) | ( n24184 & n24186 ) ;
  assign n24188 = n21774 ^ n10270 ^ n476 ;
  assign n24189 = ( n7676 & ~n13063 ) | ( n7676 & n24188 ) | ( ~n13063 & n24188 ) ;
  assign n24190 = n9758 & ~n21043 ;
  assign n24191 = n4649 & n24190 ;
  assign n24192 = n24191 ^ n13616 ^ 1'b0 ;
  assign n24193 = n24192 ^ n11700 ^ 1'b0 ;
  assign n24194 = ( x65 & n16724 ) | ( x65 & ~n18239 ) | ( n16724 & ~n18239 ) ;
  assign n24195 = n3553 & n9754 ;
  assign n24196 = ( n1239 & ~n1885 ) | ( n1239 & n4521 ) | ( ~n1885 & n4521 ) ;
  assign n24197 = n24195 | n24196 ;
  assign n24198 = ( n5191 & ~n12650 ) | ( n5191 & n22888 ) | ( ~n12650 & n22888 ) ;
  assign n24199 = ( n19054 & ~n19277 ) | ( n19054 & n24198 ) | ( ~n19277 & n24198 ) ;
  assign n24200 = n14956 ^ n3938 ^ 1'b0 ;
  assign n24201 = n12102 & ~n22894 ;
  assign n24202 = n24201 ^ n13813 ^ 1'b0 ;
  assign n24204 = ( ~n4579 & n6657 ) | ( ~n4579 & n17393 ) | ( n6657 & n17393 ) ;
  assign n24203 = n13212 & ~n13324 ;
  assign n24205 = n24204 ^ n24203 ^ 1'b0 ;
  assign n24206 = n17012 | n21212 ;
  assign n24207 = ( n8011 & n17307 ) | ( n8011 & n24037 ) | ( n17307 & n24037 ) ;
  assign n24208 = n17266 ^ n6525 ^ n3836 ;
  assign n24209 = n24207 | n24208 ;
  assign n24210 = n24209 ^ n20533 ^ n11134 ;
  assign n24211 = n18903 ^ n6268 ^ 1'b0 ;
  assign n24215 = n11304 ^ n5591 ^ n4087 ;
  assign n24216 = ~n5701 & n24215 ;
  assign n24217 = ~n21003 & n24216 ;
  assign n24218 = n24217 ^ n10947 ^ n10100 ;
  assign n24212 = n4531 ^ n455 ^ 1'b0 ;
  assign n24213 = ~n3212 & n24212 ;
  assign n24214 = n1957 & ~n24213 ;
  assign n24219 = n24218 ^ n24214 ^ n18904 ;
  assign n24220 = n16635 ^ n13999 ^ 1'b0 ;
  assign n24221 = n24220 ^ n6756 ^ n801 ;
  assign n24222 = ~n1072 & n7194 ;
  assign n24224 = n6979 | n16357 ;
  assign n24223 = n12860 & n18829 ;
  assign n24225 = n24224 ^ n24223 ^ n14146 ;
  assign n24226 = n24225 ^ n20108 ^ 1'b0 ;
  assign n24227 = n9338 & ~n24226 ;
  assign n24228 = n16157 ^ n4296 ^ 1'b0 ;
  assign n24229 = n1481 & ~n24228 ;
  assign n24230 = n24229 ^ n6072 ^ 1'b0 ;
  assign n24231 = ( x57 & ~n3666 ) | ( x57 & n24230 ) | ( ~n3666 & n24230 ) ;
  assign n24232 = n3647 ^ n620 ^ 1'b0 ;
  assign n24233 = n2954 | n10963 ;
  assign n24234 = n24233 ^ n1972 ^ 1'b0 ;
  assign n24235 = n9343 & n24234 ;
  assign n24236 = ( ~n7385 & n11261 ) | ( ~n7385 & n24235 ) | ( n11261 & n24235 ) ;
  assign n24237 = ~n1322 & n4667 ;
  assign n24238 = ~n20641 & n24237 ;
  assign n24239 = ( ~n8065 & n24236 ) | ( ~n8065 & n24238 ) | ( n24236 & n24238 ) ;
  assign n24240 = ( ~n20233 & n24232 ) | ( ~n20233 & n24239 ) | ( n24232 & n24239 ) ;
  assign n24241 = ( ~n7914 & n9096 ) | ( ~n7914 & n13053 ) | ( n9096 & n13053 ) ;
  assign n24242 = n24241 ^ n19282 ^ n234 ;
  assign n24243 = n1055 & n2457 ;
  assign n24244 = n24243 ^ n7004 ^ 1'b0 ;
  assign n24245 = ~n6645 & n24244 ;
  assign n24246 = n3772 ^ n2440 ^ 1'b0 ;
  assign n24247 = n2085 | n24246 ;
  assign n24248 = n24247 ^ n17761 ^ n9666 ;
  assign n24249 = ~n10455 & n24248 ;
  assign n24250 = n4175 | n14972 ;
  assign n24251 = n21043 ^ n4945 ^ 1'b0 ;
  assign n24252 = n4384 | n24251 ;
  assign n24253 = n24250 & n24252 ;
  assign n24254 = n4845 & ~n5929 ;
  assign n24255 = n24254 ^ n9938 ^ 1'b0 ;
  assign n24256 = n24255 ^ n14718 ^ n2461 ;
  assign n24257 = n13243 ^ n6499 ^ 1'b0 ;
  assign n24258 = ( n1731 & ~n19086 ) | ( n1731 & n19876 ) | ( ~n19086 & n19876 ) ;
  assign n24259 = n15103 ^ n14647 ^ 1'b0 ;
  assign n24260 = n8061 ^ n1331 ^ 1'b0 ;
  assign n24261 = n18065 | n24260 ;
  assign n24262 = ( n148 & n3516 ) | ( n148 & n24261 ) | ( n3516 & n24261 ) ;
  assign n24263 = n12838 & n24262 ;
  assign n24264 = ~n18500 & n24263 ;
  assign n24265 = n10406 & n18293 ;
  assign n24266 = n24265 ^ n13751 ^ 1'b0 ;
  assign n24267 = n8396 & n9723 ;
  assign n24268 = n22424 & n24267 ;
  assign n24269 = n14472 | n24268 ;
  assign n24270 = n4671 | n24269 ;
  assign n24271 = n15816 ^ n8748 ^ 1'b0 ;
  assign n24272 = n9212 & n24271 ;
  assign n24273 = n24272 ^ n23748 ^ n18892 ;
  assign n24274 = n1559 & ~n21692 ;
  assign n24275 = n23207 ^ n8317 ^ n1317 ;
  assign n24276 = n22113 ^ n14729 ^ n8227 ;
  assign n24277 = n5332 & n24276 ;
  assign n24278 = n18003 ^ n4598 ^ n1728 ;
  assign n24279 = n24278 ^ n14102 ^ n13532 ;
  assign n24280 = n4044 & n6418 ;
  assign n24281 = ~n16151 & n24280 ;
  assign n24282 = n705 & ~n8302 ;
  assign n24283 = n24282 ^ n14192 ^ 1'b0 ;
  assign n24284 = n15902 | n24283 ;
  assign n24285 = n24284 ^ n19047 ^ 1'b0 ;
  assign n24289 = n1360 & n9853 ;
  assign n24290 = n24289 ^ n12820 ^ n10350 ;
  assign n24288 = n1380 & n10152 ;
  assign n24286 = n8314 ^ n4190 ^ 1'b0 ;
  assign n24287 = n19575 & ~n24286 ;
  assign n24291 = n24290 ^ n24288 ^ n24287 ;
  assign n24292 = ( ~n17665 & n22644 ) | ( ~n17665 & n23892 ) | ( n22644 & n23892 ) ;
  assign n24293 = n8797 ^ n5876 ^ n797 ;
  assign n24294 = ( n7787 & ~n21593 ) | ( n7787 & n24293 ) | ( ~n21593 & n24293 ) ;
  assign n24295 = ( n2908 & n14620 ) | ( n2908 & ~n24294 ) | ( n14620 & ~n24294 ) ;
  assign n24296 = ( n5695 & n24292 ) | ( n5695 & n24295 ) | ( n24292 & n24295 ) ;
  assign n24297 = ( ~n11541 & n15772 ) | ( ~n11541 & n18067 ) | ( n15772 & n18067 ) ;
  assign n24298 = ( ~n1130 & n2768 ) | ( ~n1130 & n12124 ) | ( n2768 & n12124 ) ;
  assign n24299 = n24298 ^ n6903 ^ 1'b0 ;
  assign n24300 = ( n11504 & n23029 ) | ( n11504 & n24299 ) | ( n23029 & n24299 ) ;
  assign n24301 = ( n2029 & n6451 ) | ( n2029 & n23051 ) | ( n6451 & n23051 ) ;
  assign n24302 = n24301 ^ n9040 ^ n458 ;
  assign n24303 = ( n3747 & n16461 ) | ( n3747 & ~n24302 ) | ( n16461 & ~n24302 ) ;
  assign n24306 = ( n3047 & ~n5618 ) | ( n3047 & n10607 ) | ( ~n5618 & n10607 ) ;
  assign n24304 = n13109 ^ n6539 ^ n4944 ;
  assign n24305 = n24304 ^ n24191 ^ n11963 ;
  assign n24307 = n24306 ^ n24305 ^ n22029 ;
  assign n24308 = ( n2580 & n4008 ) | ( n2580 & n9160 ) | ( n4008 & n9160 ) ;
  assign n24309 = n23785 & n24308 ;
  assign n24310 = n24309 ^ n2070 ^ 1'b0 ;
  assign n24311 = n24310 ^ n13218 ^ n4794 ;
  assign n24312 = n10139 | n21230 ;
  assign n24313 = n22944 ^ n22340 ^ 1'b0 ;
  assign n24314 = ~n24312 & n24313 ;
  assign n24315 = ( n2305 & ~n3390 ) | ( n2305 & n11350 ) | ( ~n3390 & n11350 ) ;
  assign n24316 = ( n2024 & n7036 ) | ( n2024 & ~n24315 ) | ( n7036 & ~n24315 ) ;
  assign n24317 = n17599 ^ n13857 ^ n9244 ;
  assign n24318 = n19971 & ~n22301 ;
  assign n24319 = n24318 ^ n19830 ^ 1'b0 ;
  assign n24320 = n24317 | n24319 ;
  assign n24321 = ( n12499 & n24316 ) | ( n12499 & ~n24320 ) | ( n24316 & ~n24320 ) ;
  assign n24324 = n1110 & n5917 ;
  assign n24325 = n24324 ^ n12649 ^ 1'b0 ;
  assign n24322 = n1665 & ~n8567 ;
  assign n24323 = n24322 ^ n2906 ^ 1'b0 ;
  assign n24326 = n24325 ^ n24323 ^ n19058 ;
  assign n24327 = n9614 ^ n3564 ^ n3428 ;
  assign n24328 = n16865 ^ n1845 ^ 1'b0 ;
  assign n24329 = ( n17195 & n24327 ) | ( n17195 & ~n24328 ) | ( n24327 & ~n24328 ) ;
  assign n24330 = n19039 & n22943 ;
  assign n24331 = n3948 & ~n24330 ;
  assign n24332 = ~n9292 & n24331 ;
  assign n24333 = n880 | n901 ;
  assign n24334 = n24333 ^ n2124 ^ 1'b0 ;
  assign n24335 = n24334 ^ n8888 ^ 1'b0 ;
  assign n24336 = ~n2219 & n24335 ;
  assign n24337 = ( n11177 & n24332 ) | ( n11177 & n24336 ) | ( n24332 & n24336 ) ;
  assign n24338 = n16942 ^ n14379 ^ 1'b0 ;
  assign n24339 = ~n18263 & n19569 ;
  assign n24340 = n24339 ^ n14919 ^ 1'b0 ;
  assign n24341 = ( n10720 & n10909 ) | ( n10720 & n24340 ) | ( n10909 & n24340 ) ;
  assign n24342 = n2260 & n11439 ;
  assign n24343 = ( n486 & ~n8111 ) | ( n486 & n12881 ) | ( ~n8111 & n12881 ) ;
  assign n24344 = ( n1761 & ~n14389 ) | ( n1761 & n24343 ) | ( ~n14389 & n24343 ) ;
  assign n24345 = ( n22738 & n24342 ) | ( n22738 & ~n24344 ) | ( n24342 & ~n24344 ) ;
  assign n24346 = n4729 | n22618 ;
  assign n24347 = n24346 ^ n10138 ^ 1'b0 ;
  assign n24348 = ( ~n1301 & n16193 ) | ( ~n1301 & n16778 ) | ( n16193 & n16778 ) ;
  assign n24349 = n24348 ^ n6675 ^ 1'b0 ;
  assign n24350 = n11871 & ~n24349 ;
  assign n24351 = n18183 ^ n7065 ^ n5222 ;
  assign n24352 = n2714 & ~n24351 ;
  assign n24353 = n3638 | n20854 ;
  assign n24354 = n7200 & ~n24353 ;
  assign n24355 = n15568 & ~n24354 ;
  assign n24356 = n14100 & n24355 ;
  assign n24357 = n24356 ^ n19083 ^ 1'b0 ;
  assign n24358 = n24357 ^ n12312 ^ n8676 ;
  assign n24359 = n24358 ^ n17479 ^ n14627 ;
  assign n24360 = n13475 ^ n11064 ^ n4433 ;
  assign n24361 = n24360 ^ n11861 ^ 1'b0 ;
  assign n24362 = n2582 & n8641 ;
  assign n24363 = n24362 ^ n5890 ^ 1'b0 ;
  assign n24364 = n24363 ^ n11349 ^ n5046 ;
  assign n24365 = n24364 ^ n24165 ^ n23415 ;
  assign n24366 = n18386 ^ n16754 ^ n7847 ;
  assign n24367 = n7225 ^ n867 ^ 1'b0 ;
  assign n24368 = n4222 & n24367 ;
  assign n24369 = ~n6206 & n24368 ;
  assign n24370 = n23804 ^ n9829 ^ n8082 ;
  assign n24371 = ~n2593 & n15612 ;
  assign n24372 = n3188 ^ n3102 ^ n2320 ;
  assign n24373 = n24372 ^ n19767 ^ 1'b0 ;
  assign n24374 = n6951 & ~n24373 ;
  assign n24375 = ( n1805 & n10524 ) | ( n1805 & n24374 ) | ( n10524 & n24374 ) ;
  assign n24376 = ~n3340 & n11963 ;
  assign n24377 = n24376 ^ n14960 ^ 1'b0 ;
  assign n24378 = ( n24371 & ~n24375 ) | ( n24371 & n24377 ) | ( ~n24375 & n24377 ) ;
  assign n24379 = n8356 ^ n6885 ^ 1'b0 ;
  assign n24380 = ( ~n4282 & n8347 ) | ( ~n4282 & n22970 ) | ( n8347 & n22970 ) ;
  assign n24381 = ( n5737 & n24379 ) | ( n5737 & n24380 ) | ( n24379 & n24380 ) ;
  assign n24382 = ( n8981 & n9867 ) | ( n8981 & ~n15301 ) | ( n9867 & ~n15301 ) ;
  assign n24383 = ( ~n3564 & n24122 ) | ( ~n3564 & n24382 ) | ( n24122 & n24382 ) ;
  assign n24384 = ( ~n5416 & n6820 ) | ( ~n5416 & n21528 ) | ( n6820 & n21528 ) ;
  assign n24385 = n11386 & n24384 ;
  assign n24386 = n24385 ^ n23626 ^ 1'b0 ;
  assign n24387 = n18387 ^ n1570 ^ 1'b0 ;
  assign n24388 = n12869 & ~n24387 ;
  assign n24389 = n24388 ^ n10754 ^ n9834 ;
  assign n24390 = n19395 ^ n10415 ^ 1'b0 ;
  assign n24391 = n4184 & ~n24390 ;
  assign n24392 = ~n1659 & n24391 ;
  assign n24393 = n24389 & n24392 ;
  assign n24394 = n16385 ^ n12881 ^ n7937 ;
  assign n24395 = n21377 ^ n6937 ^ 1'b0 ;
  assign n24396 = ~n4606 & n17208 ;
  assign n24397 = ( n2465 & ~n14405 ) | ( n2465 & n14956 ) | ( ~n14405 & n14956 ) ;
  assign n24398 = n24397 ^ n3080 ^ n2370 ;
  assign n24399 = ( n7601 & n7627 ) | ( n7601 & ~n24398 ) | ( n7627 & ~n24398 ) ;
  assign n24402 = n1993 ^ n1483 ^ n186 ;
  assign n24403 = n17851 ^ n6305 ^ 1'b0 ;
  assign n24404 = ~n18095 & n24403 ;
  assign n24405 = ( n8096 & n24402 ) | ( n8096 & ~n24404 ) | ( n24402 & ~n24404 ) ;
  assign n24400 = ( ~n2094 & n4549 ) | ( ~n2094 & n9618 ) | ( n4549 & n9618 ) ;
  assign n24401 = n24400 ^ n17766 ^ n12261 ;
  assign n24406 = n24405 ^ n24401 ^ n18140 ;
  assign n24407 = n2716 & n17540 ;
  assign n24408 = n24407 ^ n14922 ^ 1'b0 ;
  assign n24409 = n24408 ^ n6729 ^ 1'b0 ;
  assign n24410 = ~n7231 & n24409 ;
  assign n24412 = n15320 ^ n14165 ^ n523 ;
  assign n24413 = ~n1569 & n24412 ;
  assign n24411 = n3465 | n12565 ;
  assign n24414 = n24413 ^ n24411 ^ 1'b0 ;
  assign n24417 = n2205 ^ n1967 ^ 1'b0 ;
  assign n24415 = ( n4093 & n6924 ) | ( n4093 & ~n16944 ) | ( n6924 & ~n16944 ) ;
  assign n24416 = ~n18763 & n24415 ;
  assign n24418 = n24417 ^ n24416 ^ 1'b0 ;
  assign n24419 = n3324 & ~n6919 ;
  assign n24420 = n17305 & n24419 ;
  assign n24421 = n24420 ^ n8779 ^ 1'b0 ;
  assign n24426 = n11761 ^ n2621 ^ 1'b0 ;
  assign n24427 = n21728 | n24426 ;
  assign n24428 = n6900 & n24427 ;
  assign n24422 = n5098 & n17041 ;
  assign n24423 = n24422 ^ n3361 ^ 1'b0 ;
  assign n24424 = ( n1639 & ~n2379 ) | ( n1639 & n24423 ) | ( ~n2379 & n24423 ) ;
  assign n24425 = n24424 ^ n12521 ^ 1'b0 ;
  assign n24429 = n24428 ^ n24425 ^ 1'b0 ;
  assign n24431 = ( n4771 & n5786 ) | ( n4771 & n16218 ) | ( n5786 & n16218 ) ;
  assign n24430 = ( n957 & n8954 ) | ( n957 & ~n10559 ) | ( n8954 & ~n10559 ) ;
  assign n24432 = n24431 ^ n24430 ^ 1'b0 ;
  assign n24433 = ( ~n3880 & n11102 ) | ( ~n3880 & n24432 ) | ( n11102 & n24432 ) ;
  assign n24434 = n2044 & ~n7631 ;
  assign n24435 = n3196 ^ n1996 ^ n941 ;
  assign n24436 = ( n8094 & n24434 ) | ( n8094 & n24435 ) | ( n24434 & n24435 ) ;
  assign n24437 = n21667 ^ n13297 ^ n4534 ;
  assign n24438 = ~n18905 & n24437 ;
  assign n24439 = n12335 ^ n6933 ^ x108 ;
  assign n24440 = ( n17241 & n24438 ) | ( n17241 & n24439 ) | ( n24438 & n24439 ) ;
  assign n24441 = n14986 ^ n3543 ^ n1929 ;
  assign n24443 = n12189 ^ n10571 ^ 1'b0 ;
  assign n24442 = n17063 ^ n14016 ^ n13335 ;
  assign n24444 = n24443 ^ n24442 ^ n14083 ;
  assign n24445 = n4437 & ~n5230 ;
  assign n24446 = ~n19835 & n24445 ;
  assign n24447 = n22873 & ~n24446 ;
  assign n24448 = ~n15424 & n15936 ;
  assign n24449 = n24448 ^ n3364 ^ 1'b0 ;
  assign n24450 = n24449 ^ n11618 ^ 1'b0 ;
  assign n24451 = ~n4534 & n24450 ;
  assign n24456 = n6227 & ~n8546 ;
  assign n24457 = n24456 ^ n2165 ^ 1'b0 ;
  assign n24458 = n4831 | n24457 ;
  assign n24459 = n24458 ^ n2031 ^ 1'b0 ;
  assign n24452 = n9817 & ~n14774 ;
  assign n24453 = n8005 & n24452 ;
  assign n24454 = ( ~n4076 & n12256 ) | ( ~n4076 & n24453 ) | ( n12256 & n24453 ) ;
  assign n24455 = ( n22621 & n23333 ) | ( n22621 & ~n24454 ) | ( n23333 & ~n24454 ) ;
  assign n24460 = n24459 ^ n24455 ^ n6167 ;
  assign n24461 = n2977 & n7197 ;
  assign n24462 = n24461 ^ n10598 ^ 1'b0 ;
  assign n24463 = ~n8060 & n24462 ;
  assign n24464 = n24463 ^ n7150 ^ 1'b0 ;
  assign n24465 = n12273 ^ n8557 ^ 1'b0 ;
  assign n24466 = n15949 & n24465 ;
  assign n24467 = ( n24454 & ~n24464 ) | ( n24454 & n24466 ) | ( ~n24464 & n24466 ) ;
  assign n24468 = n14355 ^ n9642 ^ n2688 ;
  assign n24469 = n10048 ^ n1031 ^ 1'b0 ;
  assign n24470 = n7846 ^ n4876 ^ n2805 ;
  assign n24471 = n19768 ^ n10087 ^ 1'b0 ;
  assign n24472 = n24471 ^ n21874 ^ n6123 ;
  assign n24473 = n24472 ^ n18214 ^ 1'b0 ;
  assign n24474 = ( ~n2807 & n8681 ) | ( ~n2807 & n10413 ) | ( n8681 & n10413 ) ;
  assign n24475 = ( ~n202 & n9336 ) | ( ~n202 & n24474 ) | ( n9336 & n24474 ) ;
  assign n24476 = ~n4583 & n10056 ;
  assign n24477 = ~n10329 & n24476 ;
  assign n24478 = n24477 ^ n14080 ^ 1'b0 ;
  assign n24479 = n24475 | n24478 ;
  assign n24480 = ( n7722 & n23433 ) | ( n7722 & n24479 ) | ( n23433 & n24479 ) ;
  assign n24481 = ( ~n4465 & n8346 ) | ( ~n4465 & n18070 ) | ( n8346 & n18070 ) ;
  assign n24482 = n7381 & n24481 ;
  assign n24484 = ( n4330 & ~n5948 ) | ( n4330 & n21867 ) | ( ~n5948 & n21867 ) ;
  assign n24483 = ( n8989 & n11159 ) | ( n8989 & n12257 ) | ( n11159 & n12257 ) ;
  assign n24485 = n24484 ^ n24483 ^ 1'b0 ;
  assign n24486 = n10518 & n24485 ;
  assign n24487 = n24486 ^ n21211 ^ 1'b0 ;
  assign n24488 = n23449 ^ n10545 ^ 1'b0 ;
  assign n24489 = n10203 ^ n2679 ^ 1'b0 ;
  assign n24490 = n14438 & ~n24489 ;
  assign n24491 = n15886 ^ n1538 ^ n974 ;
  assign n24492 = n4973 ^ n1773 ^ n549 ;
  assign n24493 = n24492 ^ n19314 ^ n7182 ;
  assign n24494 = n24493 ^ n21871 ^ n8285 ;
  assign n24495 = n6917 | n23403 ;
  assign n24496 = n20714 & ~n24495 ;
  assign n24497 = x44 & ~n11943 ;
  assign n24498 = ~n2689 & n24497 ;
  assign n24499 = n24496 | n24498 ;
  assign n24500 = ( ~n8458 & n15216 ) | ( ~n8458 & n21984 ) | ( n15216 & n21984 ) ;
  assign n24501 = n1626 & ~n10761 ;
  assign n24502 = n15568 ^ n6952 ^ 1'b0 ;
  assign n24503 = n7807 & ~n24502 ;
  assign n24504 = ( n1334 & n21021 ) | ( n1334 & ~n24503 ) | ( n21021 & ~n24503 ) ;
  assign n24505 = n10327 | n11664 ;
  assign n24506 = n19823 & ~n22084 ;
  assign n24507 = n12894 & n24506 ;
  assign n24508 = n10375 ^ n6988 ^ 1'b0 ;
  assign n24509 = n7449 & n24508 ;
  assign n24515 = ( ~n7127 & n15595 ) | ( ~n7127 & n15811 ) | ( n15595 & n15811 ) ;
  assign n24516 = ( n17304 & n18108 ) | ( n17304 & ~n24515 ) | ( n18108 & ~n24515 ) ;
  assign n24511 = n5180 ^ n3799 ^ n3473 ;
  assign n24510 = ~n10138 & n14085 ;
  assign n24512 = n24511 ^ n24510 ^ 1'b0 ;
  assign n24513 = n15320 & ~n24512 ;
  assign n24514 = ~n13563 & n24513 ;
  assign n24517 = n24516 ^ n24514 ^ 1'b0 ;
  assign n24518 = n15583 ^ n6880 ^ n5488 ;
  assign n24519 = n24518 ^ n3931 ^ 1'b0 ;
  assign n24520 = n22287 ^ n6668 ^ 1'b0 ;
  assign n24521 = n23940 & n24520 ;
  assign n24522 = ( n2886 & n24519 ) | ( n2886 & ~n24521 ) | ( n24519 & ~n24521 ) ;
  assign n24523 = n3197 | n11594 ;
  assign n24524 = n4191 & ~n24523 ;
  assign n24525 = n24524 ^ n22600 ^ 1'b0 ;
  assign n24526 = ( n8816 & ~n9742 ) | ( n8816 & n24525 ) | ( ~n9742 & n24525 ) ;
  assign n24527 = n5725 | n9072 ;
  assign n24528 = x99 & ~n9669 ;
  assign n24529 = n24528 ^ n11840 ^ n6281 ;
  assign n24530 = n2583 & ~n14848 ;
  assign n24531 = n11935 ^ n5681 ^ n5022 ;
  assign n24532 = n13227 ^ n9289 ^ 1'b0 ;
  assign n24533 = ~n24531 & n24532 ;
  assign n24534 = n24533 ^ n524 ^ 1'b0 ;
  assign n24535 = ~n1036 & n1146 ;
  assign n24536 = n11284 ^ n2695 ^ n726 ;
  assign n24537 = ( n6851 & n24535 ) | ( n6851 & ~n24536 ) | ( n24535 & ~n24536 ) ;
  assign n24540 = ( n1947 & n4188 ) | ( n1947 & n10015 ) | ( n4188 & n10015 ) ;
  assign n24538 = ( n2036 & n4778 ) | ( n2036 & n21130 ) | ( n4778 & n21130 ) ;
  assign n24539 = n24538 ^ n8299 ^ 1'b0 ;
  assign n24541 = n24540 ^ n24539 ^ n981 ;
  assign n24542 = n12008 | n17213 ;
  assign n24543 = n13312 & n24542 ;
  assign n24544 = ~n4416 & n24543 ;
  assign n24545 = n24544 ^ n6631 ^ 1'b0 ;
  assign n24546 = ( n3883 & n8029 ) | ( n3883 & ~n13634 ) | ( n8029 & ~n13634 ) ;
  assign n24547 = n24546 ^ n5694 ^ n3778 ;
  assign n24548 = ~n11369 & n17616 ;
  assign n24549 = n24548 ^ n7601 ^ 1'b0 ;
  assign n24550 = n5906 & ~n24549 ;
  assign n24551 = ~n24547 & n24550 ;
  assign n24552 = n1341 | n8746 ;
  assign n24553 = n24552 ^ n6805 ^ 1'b0 ;
  assign n24554 = n24553 ^ n16781 ^ n10549 ;
  assign n24555 = n16604 ^ n9743 ^ 1'b0 ;
  assign n24556 = n24554 & ~n24555 ;
  assign n24560 = ( x25 & n10071 ) | ( x25 & n12429 ) | ( n10071 & n12429 ) ;
  assign n24561 = ( n1919 & n2733 ) | ( n1919 & n4696 ) | ( n2733 & n4696 ) ;
  assign n24562 = ~n13357 & n24561 ;
  assign n24563 = ~n24560 & n24562 ;
  assign n24564 = ( ~n2968 & n11052 ) | ( ~n2968 & n24563 ) | ( n11052 & n24563 ) ;
  assign n24557 = n2306 ^ n1946 ^ 1'b0 ;
  assign n24558 = ( n1048 & n4905 ) | ( n1048 & n24557 ) | ( n4905 & n24557 ) ;
  assign n24559 = n1420 | n24558 ;
  assign n24565 = n24564 ^ n24559 ^ 1'b0 ;
  assign n24566 = n3025 & ~n9670 ;
  assign n24567 = ~n7667 & n14161 ;
  assign n24568 = ~n13665 & n24567 ;
  assign n24569 = n24568 ^ n14073 ^ n8346 ;
  assign n24570 = n24569 ^ n20225 ^ n14230 ;
  assign n24571 = ( ~n4876 & n11318 ) | ( ~n4876 & n14291 ) | ( n11318 & n14291 ) ;
  assign n24572 = n19193 & n24571 ;
  assign n24573 = n24572 ^ n4458 ^ 1'b0 ;
  assign n24574 = n24573 ^ n24112 ^ n6552 ;
  assign n24575 = n1798 | n2068 ;
  assign n24576 = n4079 ^ n3312 ^ n1973 ;
  assign n24577 = n24576 ^ n2308 ^ n2204 ;
  assign n24578 = n24577 ^ n18174 ^ n11529 ;
  assign n24579 = n24578 ^ n20309 ^ 1'b0 ;
  assign n24580 = n16762 & n24579 ;
  assign n24581 = ( ~n8363 & n9694 ) | ( ~n8363 & n24571 ) | ( n9694 & n24571 ) ;
  assign n24582 = ( n5649 & n9662 ) | ( n5649 & n11592 ) | ( n9662 & n11592 ) ;
  assign n24583 = n15194 | n19322 ;
  assign n24584 = n8387 & ~n24583 ;
  assign n24585 = n18216 & n20478 ;
  assign n24586 = n24584 & n24585 ;
  assign n24587 = n24586 ^ n20510 ^ n1189 ;
  assign n24588 = n24582 | n24587 ;
  assign n24589 = n3522 & n3886 ;
  assign n24590 = n24589 ^ n8632 ^ n4491 ;
  assign n24595 = ( n1664 & ~n7610 ) | ( n1664 & n18049 ) | ( ~n7610 & n18049 ) ;
  assign n24596 = n24595 ^ n10566 ^ n6043 ;
  assign n24593 = n18748 ^ n13729 ^ n5212 ;
  assign n24592 = ~n3423 & n16458 ;
  assign n24591 = n20772 ^ n17207 ^ n9551 ;
  assign n24594 = n24593 ^ n24592 ^ n24591 ;
  assign n24597 = n24596 ^ n24594 ^ n3147 ;
  assign n24598 = n23831 ^ n18672 ^ 1'b0 ;
  assign n24599 = n6950 | n7091 ;
  assign n24600 = n24599 ^ n20429 ^ n770 ;
  assign n24601 = n19462 ^ n12978 ^ n5062 ;
  assign n24602 = ( ~n15291 & n16866 ) | ( ~n15291 & n24601 ) | ( n16866 & n24601 ) ;
  assign n24603 = n24298 ^ n18855 ^ n5667 ;
  assign n24604 = n22010 & ~n24603 ;
  assign n24605 = n24604 ^ n24399 ^ 1'b0 ;
  assign n24613 = n18216 ^ n7517 ^ n3580 ;
  assign n24609 = n8679 ^ n342 ^ 1'b0 ;
  assign n24610 = n24609 ^ n9248 ^ n2138 ;
  assign n24608 = ~n3912 & n22272 ;
  assign n24611 = n24610 ^ n24608 ^ 1'b0 ;
  assign n24607 = ( ~n6952 & n11498 ) | ( ~n6952 & n21282 ) | ( n11498 & n21282 ) ;
  assign n24612 = n24611 ^ n24607 ^ n2363 ;
  assign n24614 = n24613 ^ n24612 ^ 1'b0 ;
  assign n24606 = n2454 & n24308 ;
  assign n24615 = n24614 ^ n24606 ^ 1'b0 ;
  assign n24616 = n15300 & n15837 ;
  assign n24617 = n24616 ^ n6548 ^ 1'b0 ;
  assign n24618 = n24617 ^ n7111 ^ n623 ;
  assign n24619 = ( n2775 & n3941 ) | ( n2775 & ~n6639 ) | ( n3941 & ~n6639 ) ;
  assign n24620 = x110 & ~n22238 ;
  assign n24621 = n24619 & n24620 ;
  assign n24622 = x105 & ~n24621 ;
  assign n24623 = ( n3814 & n19424 ) | ( n3814 & ~n21533 ) | ( n19424 & ~n21533 ) ;
  assign n24624 = n24623 ^ n3710 ^ 1'b0 ;
  assign n24625 = ~n784 & n2950 ;
  assign n24626 = n24625 ^ n10664 ^ 1'b0 ;
  assign n24627 = ( n7535 & n11591 ) | ( n7535 & ~n24626 ) | ( n11591 & ~n24626 ) ;
  assign n24628 = n19577 ^ n11814 ^ n10766 ;
  assign n24629 = ~n231 & n13633 ;
  assign n24630 = ( n6685 & n6845 ) | ( n6685 & ~n24629 ) | ( n6845 & ~n24629 ) ;
  assign n24634 = ( ~n189 & n5595 ) | ( ~n189 & n19268 ) | ( n5595 & n19268 ) ;
  assign n24631 = ( n13570 & ~n14272 ) | ( n13570 & n16351 ) | ( ~n14272 & n16351 ) ;
  assign n24632 = ( n8751 & n12840 ) | ( n8751 & n24631 ) | ( n12840 & n24631 ) ;
  assign n24633 = n24632 ^ n23052 ^ n1626 ;
  assign n24635 = n24634 ^ n24633 ^ 1'b0 ;
  assign n24636 = n8080 ^ n6544 ^ n2512 ;
  assign n24637 = ( n6680 & n9101 ) | ( n6680 & ~n24636 ) | ( n9101 & ~n24636 ) ;
  assign n24638 = x73 & n24637 ;
  assign n24639 = n5848 ^ n2635 ^ 1'b0 ;
  assign n24640 = n22950 & ~n24639 ;
  assign n24641 = n10433 & ~n13894 ;
  assign n24642 = n24174 & n24641 ;
  assign n24643 = ( n15164 & n15401 ) | ( n15164 & ~n19767 ) | ( n15401 & ~n19767 ) ;
  assign n24644 = ( ~n2134 & n4743 ) | ( ~n2134 & n21757 ) | ( n4743 & n21757 ) ;
  assign n24645 = n19464 ^ n14562 ^ n4236 ;
  assign n24646 = n14405 ^ n11658 ^ n3220 ;
  assign n24647 = ( n1019 & ~n20893 ) | ( n1019 & n24646 ) | ( ~n20893 & n24646 ) ;
  assign n24648 = n2733 ^ n2535 ^ 1'b0 ;
  assign n24649 = n20889 | n24648 ;
  assign n24650 = ( n3475 & ~n18289 ) | ( n3475 & n18526 ) | ( ~n18289 & n18526 ) ;
  assign n24651 = ( ~n15691 & n16267 ) | ( ~n15691 & n24650 ) | ( n16267 & n24650 ) ;
  assign n24652 = ( n11064 & n11134 ) | ( n11064 & ~n11775 ) | ( n11134 & ~n11775 ) ;
  assign n24653 = ~n18811 & n24652 ;
  assign n24654 = n24653 ^ n1559 ^ 1'b0 ;
  assign n24655 = n20277 & ~n24654 ;
  assign n24657 = n8638 & n9087 ;
  assign n24658 = n24657 ^ n14508 ^ 1'b0 ;
  assign n24656 = n16308 ^ n3996 ^ n1199 ;
  assign n24659 = n24658 ^ n24656 ^ n15576 ;
  assign n24660 = n17411 | n24659 ;
  assign n24661 = ( n1973 & ~n5817 ) | ( n1973 & n12105 ) | ( ~n5817 & n12105 ) ;
  assign n24662 = n24661 ^ n18088 ^ n2430 ;
  assign n24663 = n24023 ^ n5639 ^ 1'b0 ;
  assign n24664 = n24663 ^ n13669 ^ 1'b0 ;
  assign n24665 = n12853 & n14995 ;
  assign n24666 = n24665 ^ n10133 ^ 1'b0 ;
  assign n24667 = n16861 ^ n12316 ^ n6103 ;
  assign n24668 = ~n14230 & n24667 ;
  assign n24669 = n24668 ^ n9075 ^ 1'b0 ;
  assign n24670 = x85 & ~n662 ;
  assign n24671 = n24670 ^ n19386 ^ 1'b0 ;
  assign n24672 = ~n7565 & n9751 ;
  assign n24673 = n24672 ^ n6234 ^ 1'b0 ;
  assign n24677 = n3619 & ~n5485 ;
  assign n24678 = ~n20477 & n24677 ;
  assign n24674 = ( n658 & n5502 ) | ( n658 & ~n18814 ) | ( n5502 & ~n18814 ) ;
  assign n24675 = n24674 ^ n4936 ^ 1'b0 ;
  assign n24676 = n11376 & n24675 ;
  assign n24679 = n24678 ^ n24676 ^ 1'b0 ;
  assign n24680 = n8577 ^ n4710 ^ n2869 ;
  assign n24681 = n24680 ^ n15143 ^ n5201 ;
  assign n24682 = n10688 ^ n2075 ^ 1'b0 ;
  assign n24683 = n9739 | n24682 ;
  assign n24684 = n24683 ^ n11169 ^ n7175 ;
  assign n24685 = n24684 ^ n20691 ^ n7047 ;
  assign n24686 = n9515 ^ n3985 ^ 1'b0 ;
  assign n24687 = n8390 & n24686 ;
  assign n24688 = n24687 ^ n11623 ^ n5942 ;
  assign n24689 = n16811 ^ n10891 ^ n7791 ;
  assign n24690 = n24689 ^ n547 ^ 1'b0 ;
  assign n24691 = n16351 | n24690 ;
  assign n24692 = n9643 ^ n1963 ^ 1'b0 ;
  assign n24693 = n10024 & n24692 ;
  assign n24694 = n9730 ^ n2323 ^ 1'b0 ;
  assign n24695 = ( n3471 & n13573 ) | ( n3471 & n14590 ) | ( n13573 & n14590 ) ;
  assign n24696 = ( n664 & n1605 ) | ( n664 & n15778 ) | ( n1605 & n15778 ) ;
  assign n24697 = ( n10946 & ~n10954 ) | ( n10946 & n24696 ) | ( ~n10954 & n24696 ) ;
  assign n24698 = ( x112 & ~n5238 ) | ( x112 & n24697 ) | ( ~n5238 & n24697 ) ;
  assign n24700 = n13973 ^ n2915 ^ 1'b0 ;
  assign n24699 = ~n8255 & n10869 ;
  assign n24701 = n24700 ^ n24699 ^ 1'b0 ;
  assign n24702 = n20491 ^ n12351 ^ 1'b0 ;
  assign n24703 = n7052 | n24702 ;
  assign n24704 = ~n8743 & n12943 ;
  assign n24705 = n24704 ^ n14613 ^ 1'b0 ;
  assign n24706 = ~n4302 & n4784 ;
  assign n24707 = n17552 ^ n11262 ^ n240 ;
  assign n24708 = n8834 ^ n5775 ^ n1993 ;
  assign n24709 = n9613 | n20801 ;
  assign n24710 = ( n6750 & n17345 ) | ( n6750 & n24709 ) | ( n17345 & n24709 ) ;
  assign n24711 = n24175 ^ n12365 ^ 1'b0 ;
  assign n24712 = n4504 & ~n24711 ;
  assign n24713 = ( n919 & n11574 ) | ( n919 & ~n24712 ) | ( n11574 & ~n24712 ) ;
  assign n24714 = n24713 ^ n20462 ^ n15181 ;
  assign n24715 = ~n10674 & n17711 ;
  assign n24716 = n24715 ^ n9009 ^ n5051 ;
  assign n24717 = n10021 & ~n20160 ;
  assign n24718 = n24717 ^ n11166 ^ n7111 ;
  assign n24719 = n21684 ^ n11842 ^ 1'b0 ;
  assign n24720 = ~n24718 & n24719 ;
  assign n24721 = n13399 ^ n2340 ^ 1'b0 ;
  assign n24722 = n24721 ^ n8792 ^ n6719 ;
  assign n24724 = ( ~n4713 & n10386 ) | ( ~n4713 & n17535 ) | ( n10386 & n17535 ) ;
  assign n24723 = n3500 & ~n23556 ;
  assign n24725 = n24724 ^ n24723 ^ 1'b0 ;
  assign n24726 = n24725 ^ n21798 ^ n7810 ;
  assign n24727 = n17546 ^ n8571 ^ 1'b0 ;
  assign n24728 = n24727 ^ n15016 ^ n7768 ;
  assign n24729 = n24188 & ~n24728 ;
  assign n24730 = n7739 ^ n6088 ^ n4968 ;
  assign n24731 = n23048 ^ n5242 ^ n2319 ;
  assign n24732 = ( n11278 & n24730 ) | ( n11278 & n24731 ) | ( n24730 & n24731 ) ;
  assign n24734 = n6311 ^ n5337 ^ n3848 ;
  assign n24735 = ( n3282 & n4833 ) | ( n3282 & ~n24734 ) | ( n4833 & ~n24734 ) ;
  assign n24733 = ( n1692 & n21635 ) | ( n1692 & ~n23651 ) | ( n21635 & ~n23651 ) ;
  assign n24736 = n24735 ^ n24733 ^ n8479 ;
  assign n24737 = n11293 ^ n10369 ^ 1'b0 ;
  assign n24738 = n23406 | n24737 ;
  assign n24739 = n16191 ^ n9477 ^ 1'b0 ;
  assign n24740 = ~n2105 & n24739 ;
  assign n24741 = ~n24738 & n24740 ;
  assign n24742 = ( n14192 & n24713 ) | ( n14192 & ~n24741 ) | ( n24713 & ~n24741 ) ;
  assign n24743 = n5170 | n13242 ;
  assign n24744 = n5800 & ~n24743 ;
  assign n24745 = n4428 | n17722 ;
  assign n24746 = n24744 & ~n24745 ;
  assign n24747 = ~n13905 & n21178 ;
  assign n24748 = n24747 ^ n1179 ^ 1'b0 ;
  assign n24751 = n14429 ^ n10809 ^ n3434 ;
  assign n24749 = ~n6635 & n15303 ;
  assign n24750 = n24749 ^ n4833 ^ 1'b0 ;
  assign n24752 = n24751 ^ n24750 ^ n6008 ;
  assign n24753 = n17013 ^ n3390 ^ n1496 ;
  assign n24760 = ( ~n3281 & n12735 ) | ( ~n3281 & n21359 ) | ( n12735 & n21359 ) ;
  assign n24758 = n19043 ^ n8623 ^ n1677 ;
  assign n24759 = n9339 | n24758 ;
  assign n24755 = ( n5675 & n9277 ) | ( n5675 & ~n14209 ) | ( n9277 & ~n14209 ) ;
  assign n24756 = n24755 ^ n11579 ^ n5801 ;
  assign n24754 = ~n8548 & n8692 ;
  assign n24757 = n24756 ^ n24754 ^ 1'b0 ;
  assign n24761 = n24760 ^ n24759 ^ n24757 ;
  assign n24762 = n9459 ^ n8918 ^ n916 ;
  assign n24763 = ~n2603 & n24762 ;
  assign n24764 = n3918 & n24763 ;
  assign n24765 = n455 & ~n24764 ;
  assign n24766 = n200 & n649 ;
  assign n24767 = ~n12259 & n24766 ;
  assign n24768 = n24561 ^ n14692 ^ n3698 ;
  assign n24769 = ( n8343 & n24767 ) | ( n8343 & ~n24768 ) | ( n24767 & ~n24768 ) ;
  assign n24770 = n8570 ^ n5981 ^ 1'b0 ;
  assign n24772 = n14264 ^ n9490 ^ 1'b0 ;
  assign n24773 = n19362 | n24772 ;
  assign n24771 = ~n2213 & n12532 ;
  assign n24774 = n24773 ^ n24771 ^ n16550 ;
  assign n24775 = n24774 ^ n11416 ^ 1'b0 ;
  assign n24776 = ~n3825 & n24775 ;
  assign n24778 = ( n2560 & n12520 ) | ( n2560 & ~n12745 ) | ( n12520 & ~n12745 ) ;
  assign n24779 = n24778 ^ n5843 ^ 1'b0 ;
  assign n24777 = ( n11741 & n14802 ) | ( n11741 & ~n18230 ) | ( n14802 & ~n18230 ) ;
  assign n24780 = n24779 ^ n24777 ^ n2118 ;
  assign n24781 = n10210 ^ n8961 ^ n798 ;
  assign n24782 = n4050 ^ n4017 ^ n1820 ;
  assign n24783 = ( ~n13601 & n15772 ) | ( ~n13601 & n24782 ) | ( n15772 & n24782 ) ;
  assign n24784 = ( n2686 & n7949 ) | ( n2686 & ~n11671 ) | ( n7949 & ~n11671 ) ;
  assign n24785 = ( n4384 & n22985 ) | ( n4384 & n24784 ) | ( n22985 & n24784 ) ;
  assign n24786 = n6694 ^ n3268 ^ n1370 ;
  assign n24787 = n8152 & ~n15980 ;
  assign n24788 = n13172 ^ n3779 ^ 1'b0 ;
  assign n24789 = ~n16978 & n24788 ;
  assign n24790 = ~n24787 & n24789 ;
  assign n24791 = n11751 | n24790 ;
  assign n24792 = n24791 ^ n12203 ^ 1'b0 ;
  assign n24793 = n858 & ~n13423 ;
  assign n24797 = ~n2953 & n14521 ;
  assign n24798 = n24797 ^ n1569 ^ 1'b0 ;
  assign n24796 = n1326 | n3581 ;
  assign n24799 = n24798 ^ n24796 ^ n15360 ;
  assign n24794 = ~n3366 & n11063 ;
  assign n24795 = n24794 ^ n22291 ^ 1'b0 ;
  assign n24800 = n24799 ^ n24795 ^ 1'b0 ;
  assign n24801 = x92 & n9977 ;
  assign n24802 = n24800 & n24801 ;
  assign n24803 = n2465 ^ n2305 ^ 1'b0 ;
  assign n24804 = n20702 | n24803 ;
  assign n24805 = ( n7844 & ~n16719 ) | ( n7844 & n24804 ) | ( ~n16719 & n24804 ) ;
  assign n24806 = n9489 ^ n5784 ^ n4687 ;
  assign n24807 = ~n2371 & n14116 ;
  assign n24808 = n1321 | n24807 ;
  assign n24809 = n24808 ^ n6811 ^ 1'b0 ;
  assign n24810 = ~n7262 & n24809 ;
  assign n24811 = ( n14854 & n24806 ) | ( n14854 & ~n24810 ) | ( n24806 & ~n24810 ) ;
  assign n24812 = n3407 & ~n15909 ;
  assign n24813 = n24812 ^ n9220 ^ n2642 ;
  assign n24815 = ( n565 & ~n10311 ) | ( n565 & n15843 ) | ( ~n10311 & n15843 ) ;
  assign n24814 = n2113 & ~n22391 ;
  assign n24816 = n24815 ^ n24814 ^ n5604 ;
  assign n24817 = ( n1832 & ~n6893 ) | ( n1832 & n7906 ) | ( ~n6893 & n7906 ) ;
  assign n24818 = n19983 ^ n4827 ^ 1'b0 ;
  assign n24819 = n7304 & n24818 ;
  assign n24820 = ~n8146 & n24819 ;
  assign n24821 = n11344 & ~n20400 ;
  assign n24822 = ~n11051 & n24821 ;
  assign n24823 = n7426 & ~n16116 ;
  assign n24824 = n24822 & n24823 ;
  assign n24825 = n17676 & ~n24824 ;
  assign n24826 = ~n19165 & n24825 ;
  assign n24827 = n12889 ^ n5658 ^ n1436 ;
  assign n24828 = ( n2409 & n6179 ) | ( n2409 & ~n12710 ) | ( n6179 & ~n12710 ) ;
  assign n24829 = n16229 ^ n14534 ^ n1217 ;
  assign n24830 = ~n3428 & n3937 ;
  assign n24831 = n11785 & n24830 ;
  assign n24832 = ( n3579 & n19457 ) | ( n3579 & n24831 ) | ( n19457 & n24831 ) ;
  assign n24833 = n24832 ^ n12224 ^ 1'b0 ;
  assign n24834 = n13880 & n24833 ;
  assign n24835 = ~n1826 & n24834 ;
  assign n24836 = ~n21879 & n24835 ;
  assign n24837 = n24836 ^ n14481 ^ n8748 ;
  assign n24838 = ( n3199 & n14190 ) | ( n3199 & n23015 ) | ( n14190 & n23015 ) ;
  assign n24839 = n9241 ^ n3503 ^ 1'b0 ;
  assign n24840 = n320 | n24839 ;
  assign n24841 = n725 & ~n24840 ;
  assign n24842 = n24659 ^ n17236 ^ 1'b0 ;
  assign n24843 = n11970 & ~n23118 ;
  assign n24844 = n18184 ^ n14598 ^ n1826 ;
  assign n24845 = n24844 ^ n19933 ^ n330 ;
  assign n24846 = n22309 ^ n7038 ^ 1'b0 ;
  assign n24847 = n1554 | n6427 ;
  assign n24848 = n24847 ^ n21894 ^ n17284 ;
  assign n24849 = n14480 & n20474 ;
  assign n24850 = n8072 ^ n6524 ^ n934 ;
  assign n24851 = ( n6955 & n10304 ) | ( n6955 & n24850 ) | ( n10304 & n24850 ) ;
  assign n24852 = ~n759 & n24851 ;
  assign n24853 = n24852 ^ n12740 ^ 1'b0 ;
  assign n24854 = n24853 ^ n16656 ^ 1'b0 ;
  assign n24855 = n24854 ^ n8540 ^ n3816 ;
  assign n24856 = n7518 ^ n5225 ^ n5135 ;
  assign n24857 = n15890 | n24856 ;
  assign n24858 = n8666 | n24857 ;
  assign n24859 = n24858 ^ n18962 ^ 1'b0 ;
  assign n24860 = n7617 & ~n17253 ;
  assign n24861 = n24859 & n24860 ;
  assign n24862 = n19357 ^ n6441 ^ 1'b0 ;
  assign n24863 = ~n17671 & n24862 ;
  assign n24864 = ( ~n3181 & n8205 ) | ( ~n3181 & n15631 ) | ( n8205 & n15631 ) ;
  assign n24865 = n15770 | n16229 ;
  assign n24866 = ~n24864 & n24865 ;
  assign n24867 = ~n12796 & n13609 ;
  assign n24868 = ( ~n1443 & n5269 ) | ( ~n1443 & n13659 ) | ( n5269 & n13659 ) ;
  assign n24869 = n2264 ^ n1351 ^ 1'b0 ;
  assign n24870 = ( n6617 & n14010 ) | ( n6617 & n24869 ) | ( n14010 & n24869 ) ;
  assign n24871 = ( n18842 & ~n24868 ) | ( n18842 & n24870 ) | ( ~n24868 & n24870 ) ;
  assign n24872 = n2729 ^ n1130 ^ n328 ;
  assign n24876 = n5448 ^ n4592 ^ n2707 ;
  assign n24874 = n4401 ^ x16 ^ 1'b0 ;
  assign n24873 = ~n1013 & n7814 ;
  assign n24875 = n24874 ^ n24873 ^ 1'b0 ;
  assign n24877 = n24876 ^ n24875 ^ n13539 ;
  assign n24878 = ( n4056 & n9955 ) | ( n4056 & n18534 ) | ( n9955 & n18534 ) ;
  assign n24879 = n24878 ^ n15719 ^ n12884 ;
  assign n24880 = ( n7351 & ~n24877 ) | ( n7351 & n24879 ) | ( ~n24877 & n24879 ) ;
  assign n24881 = ( n2796 & n12877 ) | ( n2796 & n14135 ) | ( n12877 & n14135 ) ;
  assign n24882 = n7262 ^ n6123 ^ 1'b0 ;
  assign n24883 = n24882 ^ n11134 ^ n1172 ;
  assign n24884 = n8478 & ~n13352 ;
  assign n24885 = n11564 & n24884 ;
  assign n24886 = n21855 ^ n1120 ^ 1'b0 ;
  assign n24887 = ~n13948 & n24886 ;
  assign n24890 = ( n6343 & n6675 ) | ( n6343 & ~n7678 ) | ( n6675 & ~n7678 ) ;
  assign n24888 = ( n4314 & n5103 ) | ( n4314 & n21425 ) | ( n5103 & n21425 ) ;
  assign n24889 = n24888 ^ n11480 ^ n6189 ;
  assign n24891 = n24890 ^ n24889 ^ n6418 ;
  assign n24892 = n13284 & n24891 ;
  assign n24893 = n24892 ^ n9316 ^ 1'b0 ;
  assign n24894 = n1180 & n9126 ;
  assign n24895 = ( n4074 & ~n10955 ) | ( n4074 & n24894 ) | ( ~n10955 & n24894 ) ;
  assign n24896 = ( n329 & n2109 ) | ( n329 & n4841 ) | ( n2109 & n4841 ) ;
  assign n24897 = ( n15121 & n21767 ) | ( n15121 & n24896 ) | ( n21767 & n24896 ) ;
  assign n24898 = n17406 ^ n12923 ^ n6087 ;
  assign n24899 = ( n5241 & n9674 ) | ( n5241 & n12566 ) | ( n9674 & n12566 ) ;
  assign n24900 = ( n17906 & n24898 ) | ( n17906 & ~n24899 ) | ( n24898 & ~n24899 ) ;
  assign n24901 = ( ~n24895 & n24897 ) | ( ~n24895 & n24900 ) | ( n24897 & n24900 ) ;
  assign n24902 = n4615 | n19241 ;
  assign n24903 = n7929 & ~n24902 ;
  assign n24904 = n7493 ^ n2585 ^ n572 ;
  assign n24905 = ( ~n9173 & n17206 ) | ( ~n9173 & n18561 ) | ( n17206 & n18561 ) ;
  assign n24906 = n17781 ^ n4037 ^ n1480 ;
  assign n24907 = n24034 ^ n7810 ^ 1'b0 ;
  assign n24908 = n14015 & n24907 ;
  assign n24909 = n5136 & n16159 ;
  assign n24910 = n14196 & n24909 ;
  assign n24913 = n9001 & ~n12894 ;
  assign n24914 = n24913 ^ n15408 ^ 1'b0 ;
  assign n24911 = n11250 & ~n17870 ;
  assign n24912 = ~n5593 & n24911 ;
  assign n24915 = n24914 ^ n24912 ^ 1'b0 ;
  assign n24916 = ( n1215 & ~n9034 ) | ( n1215 & n19924 ) | ( ~n9034 & n19924 ) ;
  assign n24917 = n9921 & ~n22029 ;
  assign n24918 = n1906 & n24917 ;
  assign n24919 = ( n974 & n2142 ) | ( n974 & n24918 ) | ( n2142 & n24918 ) ;
  assign n24920 = n20251 ^ n2963 ^ n2676 ;
  assign n24921 = n24920 ^ n19926 ^ n3495 ;
  assign n24922 = n19906 ^ n10996 ^ n8923 ;
  assign n24923 = ( n2210 & n14123 ) | ( n2210 & ~n24922 ) | ( n14123 & ~n24922 ) ;
  assign n24924 = ~n5389 & n7718 ;
  assign n24925 = n24924 ^ n17295 ^ 1'b0 ;
  assign n24926 = n964 | n24578 ;
  assign n24927 = n2049 | n4470 ;
  assign n24928 = n21203 ^ n4072 ^ n2184 ;
  assign n24929 = n1783 ^ x88 ^ 1'b0 ;
  assign n24930 = n6382 ^ n6267 ^ n2625 ;
  assign n24931 = n7058 ^ n5774 ^ 1'b0 ;
  assign n24932 = n13019 ^ n3965 ^ n1517 ;
  assign n24933 = ( n17012 & n24931 ) | ( n17012 & n24932 ) | ( n24931 & n24932 ) ;
  assign n24934 = n2580 ^ n2294 ^ x123 ;
  assign n24935 = n24934 ^ n17843 ^ n8853 ;
  assign n24936 = n21562 ^ n981 ^ 1'b0 ;
  assign n24937 = n16984 ^ n2586 ^ 1'b0 ;
  assign n24938 = ~n2537 & n24937 ;
  assign n24939 = n6576 & n24938 ;
  assign n24940 = n7944 & n24939 ;
  assign n24941 = n18840 ^ n4190 ^ 1'b0 ;
  assign n24942 = n18075 ^ n7174 ^ 1'b0 ;
  assign n24943 = ~n24941 & n24942 ;
  assign n24944 = n6363 ^ n6044 ^ n1603 ;
  assign n24945 = ~n6167 & n24944 ;
  assign n24946 = n11651 ^ n3070 ^ 1'b0 ;
  assign n24947 = n15995 ^ n4438 ^ n2145 ;
  assign n24948 = n3878 | n20765 ;
  assign n24949 = n18306 | n24948 ;
  assign n24950 = n21152 ^ n12612 ^ 1'b0 ;
  assign n24951 = n24949 & ~n24950 ;
  assign n24952 = n7722 ^ n4948 ^ 1'b0 ;
  assign n24953 = ( ~n8146 & n24951 ) | ( ~n8146 & n24952 ) | ( n24951 & n24952 ) ;
  assign n24954 = n22165 ^ n6893 ^ 1'b0 ;
  assign n24955 = ( n549 & n9728 ) | ( n549 & ~n11337 ) | ( n9728 & ~n11337 ) ;
  assign n24956 = n24955 ^ n12526 ^ 1'b0 ;
  assign n24957 = ~n1331 & n24956 ;
  assign n24958 = n24957 ^ n4095 ^ n663 ;
  assign n24960 = n3404 ^ n417 ^ 1'b0 ;
  assign n24959 = n7061 & n11834 ;
  assign n24961 = n24960 ^ n24959 ^ n14254 ;
  assign n24962 = n5021 ^ n1895 ^ 1'b0 ;
  assign n24963 = n4902 & ~n24962 ;
  assign n24964 = n24963 ^ n21153 ^ n15151 ;
  assign n24965 = n19243 ^ n15541 ^ n14540 ;
  assign n24966 = n7489 ^ n3838 ^ 1'b0 ;
  assign n24967 = n12050 & ~n24966 ;
  assign n24968 = n15200 ^ n2852 ^ n1569 ;
  assign n24969 = n24968 ^ n3207 ^ n477 ;
  assign n24970 = n15622 ^ n2733 ^ 1'b0 ;
  assign n24971 = n18440 | n24970 ;
  assign n24972 = n24971 ^ n12182 ^ 1'b0 ;
  assign n24973 = n21871 ^ n12380 ^ n2280 ;
  assign n24974 = n14373 ^ n12616 ^ n10190 ;
  assign n24975 = n11807 ^ n7223 ^ 1'b0 ;
  assign n24976 = n1421 | n24975 ;
  assign n24979 = n14070 ^ n6043 ^ n837 ;
  assign n24980 = ( ~n5698 & n8255 ) | ( ~n5698 & n24979 ) | ( n8255 & n24979 ) ;
  assign n24977 = ~n1207 & n12722 ;
  assign n24978 = n24977 ^ n2893 ^ 1'b0 ;
  assign n24981 = n24980 ^ n24978 ^ 1'b0 ;
  assign n24982 = ( n4115 & ~n12129 ) | ( n4115 & n12935 ) | ( ~n12129 & n12935 ) ;
  assign n24983 = ( ~n5629 & n9493 ) | ( ~n5629 & n9749 ) | ( n9493 & n9749 ) ;
  assign n24984 = n16148 ^ n322 ^ 1'b0 ;
  assign n24985 = ( n12504 & n16577 ) | ( n12504 & ~n24984 ) | ( n16577 & ~n24984 ) ;
  assign n24986 = n6657 ^ n2362 ^ n755 ;
  assign n24987 = ( ~n4429 & n10317 ) | ( ~n4429 & n24986 ) | ( n10317 & n24986 ) ;
  assign n24988 = ( n15804 & n24105 ) | ( n15804 & n24987 ) | ( n24105 & n24987 ) ;
  assign n24989 = n24988 ^ n22295 ^ n14533 ;
  assign n24990 = n24989 ^ n11095 ^ 1'b0 ;
  assign n24992 = ( n7823 & n9062 ) | ( n7823 & ~n23792 ) | ( n9062 & ~n23792 ) ;
  assign n24991 = n7380 & n10048 ;
  assign n24993 = n24992 ^ n24991 ^ 1'b0 ;
  assign n24994 = n24993 ^ n13278 ^ n3221 ;
  assign n24995 = n365 & ~n13730 ;
  assign n24996 = n4053 & n24995 ;
  assign n24997 = n22136 ^ n10831 ^ n5862 ;
  assign n24998 = ( n1134 & ~n24996 ) | ( n1134 & n24997 ) | ( ~n24996 & n24997 ) ;
  assign n24999 = n8718 ^ n5150 ^ n2317 ;
  assign n25000 = n12754 ^ n3712 ^ 1'b0 ;
  assign n25001 = ( n3552 & ~n13827 ) | ( n3552 & n25000 ) | ( ~n13827 & n25000 ) ;
  assign n25002 = n9761 | n25001 ;
  assign n25003 = n24999 & ~n25002 ;
  assign n25004 = n1867 & ~n4438 ;
  assign n25005 = n25004 ^ n8402 ^ 1'b0 ;
  assign n25006 = n1145 & ~n17089 ;
  assign n25007 = n25005 & n25006 ;
  assign n25008 = ( n6461 & n8233 ) | ( n6461 & ~n8305 ) | ( n8233 & ~n8305 ) ;
  assign n25009 = n10616 ^ n2733 ^ 1'b0 ;
  assign n25010 = ( ~n6676 & n13241 ) | ( ~n6676 & n25009 ) | ( n13241 & n25009 ) ;
  assign n25011 = ( ~n7368 & n25008 ) | ( ~n7368 & n25010 ) | ( n25008 & n25010 ) ;
  assign n25012 = ( ~n5347 & n18386 ) | ( ~n5347 & n20964 ) | ( n18386 & n20964 ) ;
  assign n25013 = n21690 ^ n7421 ^ n5464 ;
  assign n25014 = ( ~n23510 & n25012 ) | ( ~n23510 & n25013 ) | ( n25012 & n25013 ) ;
  assign n25015 = n18535 ^ n14820 ^ 1'b0 ;
  assign n25016 = n25015 ^ n3580 ^ n2912 ;
  assign n25017 = n17715 ^ n6287 ^ n392 ;
  assign n25018 = n1052 & ~n15282 ;
  assign n25019 = n628 & ~n5272 ;
  assign n25020 = n25019 ^ n12380 ^ 1'b0 ;
  assign n25021 = ( n4124 & n20252 ) | ( n4124 & ~n25020 ) | ( n20252 & ~n25020 ) ;
  assign n25022 = n25021 ^ n6377 ^ 1'b0 ;
  assign n25024 = n4422 | n6623 ;
  assign n25025 = n14523 | n25024 ;
  assign n25023 = n22163 ^ n16227 ^ n16140 ;
  assign n25026 = n25025 ^ n25023 ^ n10551 ;
  assign n25027 = ( n3188 & ~n5202 ) | ( n3188 & n11878 ) | ( ~n5202 & n11878 ) ;
  assign n25028 = n25027 ^ n2893 ^ 1'b0 ;
  assign n25032 = ( n3474 & n5655 ) | ( n3474 & ~n12089 ) | ( n5655 & ~n12089 ) ;
  assign n25030 = ( n782 & n16086 ) | ( n782 & n16194 ) | ( n16086 & n16194 ) ;
  assign n25031 = n25030 ^ n19966 ^ n6667 ;
  assign n25029 = n12316 ^ n2441 ^ 1'b0 ;
  assign n25033 = n25032 ^ n25031 ^ n25029 ;
  assign n25034 = n25033 ^ n19549 ^ n2653 ;
  assign n25035 = ( n2072 & n9163 ) | ( n2072 & ~n14214 ) | ( n9163 & ~n14214 ) ;
  assign n25036 = n24330 ^ n16458 ^ n681 ;
  assign n25037 = n13413 ^ n6376 ^ 1'b0 ;
  assign n25038 = n15322 ^ n9670 ^ 1'b0 ;
  assign n25039 = n8309 | n25038 ;
  assign n25040 = n3984 ^ n2822 ^ 1'b0 ;
  assign n25041 = n25039 | n25040 ;
  assign n25042 = n21307 & ~n25041 ;
  assign n25043 = n20221 ^ n5369 ^ 1'b0 ;
  assign n25044 = n2454 & ~n25043 ;
  assign n25045 = ( n754 & ~n1013 ) | ( n754 & n9951 ) | ( ~n1013 & n9951 ) ;
  assign n25046 = n25045 ^ n9446 ^ n5822 ;
  assign n25047 = n23095 & n25046 ;
  assign n25048 = ( n1031 & n14859 ) | ( n1031 & n25047 ) | ( n14859 & n25047 ) ;
  assign n25049 = n25048 ^ n14673 ^ n1958 ;
  assign n25050 = n25044 & ~n25049 ;
  assign n25052 = n1945 | n4972 ;
  assign n25051 = n12635 & n18553 ;
  assign n25053 = n25052 ^ n25051 ^ 1'b0 ;
  assign n25054 = n25050 | n25053 ;
  assign n25055 = ( n10962 & n15010 ) | ( n10962 & ~n20634 ) | ( n15010 & ~n20634 ) ;
  assign n25056 = ( ~n620 & n18890 ) | ( ~n620 & n25055 ) | ( n18890 & n25055 ) ;
  assign n25057 = ( n2798 & n17589 ) | ( n2798 & ~n24247 ) | ( n17589 & ~n24247 ) ;
  assign n25058 = n25057 ^ n19293 ^ n728 ;
  assign n25059 = n25058 ^ n1228 ^ 1'b0 ;
  assign n25060 = ( n4285 & ~n17856 ) | ( n4285 & n20579 ) | ( ~n17856 & n20579 ) ;
  assign n25061 = n5545 ^ n3524 ^ n1744 ;
  assign n25062 = n827 & ~n2965 ;
  assign n25065 = ( n3952 & n4879 ) | ( n3952 & n14740 ) | ( n4879 & n14740 ) ;
  assign n25063 = n11698 ^ n11241 ^ n535 ;
  assign n25064 = n5930 & ~n25063 ;
  assign n25066 = n25065 ^ n25064 ^ 1'b0 ;
  assign n25067 = n25066 ^ n5996 ^ n5359 ;
  assign n25068 = ~n5009 & n25067 ;
  assign n25069 = ~n25062 & n25068 ;
  assign n25070 = ( n14134 & ~n17262 ) | ( n14134 & n19294 ) | ( ~n17262 & n19294 ) ;
  assign n25071 = n6111 ^ n1975 ^ n1273 ;
  assign n25072 = n25071 ^ n16943 ^ n11939 ;
  assign n25073 = ( ~n7836 & n24122 ) | ( ~n7836 & n25072 ) | ( n24122 & n25072 ) ;
  assign n25074 = n3452 ^ n3237 ^ 1'b0 ;
  assign n25075 = n25074 ^ n15501 ^ n2827 ;
  assign n25076 = n25075 ^ n16595 ^ n6527 ;
  assign n25077 = n16413 ^ n424 ^ 1'b0 ;
  assign n25078 = n25076 & ~n25077 ;
  assign n25079 = n8884 & n25078 ;
  assign n25080 = ( n19760 & ~n24356 ) | ( n19760 & n25079 ) | ( ~n24356 & n25079 ) ;
  assign n25081 = n16911 ^ n7120 ^ n4903 ;
  assign n25082 = ( ~n15472 & n16488 ) | ( ~n15472 & n24192 ) | ( n16488 & n24192 ) ;
  assign n25083 = n13991 ^ n5742 ^ 1'b0 ;
  assign n25084 = n23160 & n25083 ;
  assign n25085 = ( n16552 & n25082 ) | ( n16552 & ~n25084 ) | ( n25082 & ~n25084 ) ;
  assign n25086 = ~n485 & n18392 ;
  assign n25087 = ~n3882 & n7061 ;
  assign n25088 = n17384 & n25087 ;
  assign n25089 = n11923 & ~n12923 ;
  assign n25090 = n25089 ^ n17711 ^ 1'b0 ;
  assign n25091 = n25090 ^ n12366 ^ 1'b0 ;
  assign n25092 = ~n25088 & n25091 ;
  assign n25093 = ( ~n2994 & n3097 ) | ( ~n2994 & n21243 ) | ( n3097 & n21243 ) ;
  assign n25094 = ~n303 & n11832 ;
  assign n25095 = n25093 & n25094 ;
  assign n25096 = ( n6107 & ~n9972 ) | ( n6107 & n16255 ) | ( ~n9972 & n16255 ) ;
  assign n25097 = n22573 ^ n3427 ^ n2889 ;
  assign n25098 = n15775 & n25097 ;
  assign n25099 = n25096 & n25098 ;
  assign n25100 = n23971 ^ n17688 ^ n3851 ;
  assign n25101 = n25100 ^ n14338 ^ 1'b0 ;
  assign n25102 = ~n1999 & n25101 ;
  assign n25103 = n24408 ^ n8535 ^ n6337 ;
  assign n25104 = n20811 ^ n176 ^ 1'b0 ;
  assign n25105 = ( n3861 & ~n4240 ) | ( n3861 & n16050 ) | ( ~n4240 & n16050 ) ;
  assign n25106 = n25105 ^ n11306 ^ n1034 ;
  assign n25107 = ( ~n9928 & n13490 ) | ( ~n9928 & n14277 ) | ( n13490 & n14277 ) ;
  assign n25108 = n3309 & n5912 ;
  assign n25109 = x32 & n12161 ;
  assign n25110 = ( n394 & ~n7630 ) | ( n394 & n25109 ) | ( ~n7630 & n25109 ) ;
  assign n25111 = ( n2016 & ~n2800 ) | ( n2016 & n7740 ) | ( ~n2800 & n7740 ) ;
  assign n25112 = ( n4303 & ~n4926 ) | ( n4303 & n25111 ) | ( ~n4926 & n25111 ) ;
  assign n25113 = n15813 | n25112 ;
  assign n25114 = n14967 ^ n12288 ^ 1'b0 ;
  assign n25115 = n19314 & n25114 ;
  assign n25116 = n6787 | n13392 ;
  assign n25117 = n13610 & ~n25116 ;
  assign n25118 = n7344 & n13634 ;
  assign n25119 = n25118 ^ n9279 ^ 1'b0 ;
  assign n25120 = n25119 ^ n4050 ^ 1'b0 ;
  assign n25121 = n13893 ^ n1039 ^ 1'b0 ;
  assign n25122 = n16295 | n25121 ;
  assign n25123 = n19475 ^ n3576 ^ 1'b0 ;
  assign n25124 = n11252 & ~n25123 ;
  assign n25125 = n22200 & n24553 ;
  assign n25126 = n25125 ^ n9481 ^ 1'b0 ;
  assign n25127 = ( n13554 & ~n25124 ) | ( n13554 & n25126 ) | ( ~n25124 & n25126 ) ;
  assign n25128 = ( n21048 & n25122 ) | ( n21048 & ~n25127 ) | ( n25122 & ~n25127 ) ;
  assign n25129 = ( ~n384 & n4815 ) | ( ~n384 & n15515 ) | ( n4815 & n15515 ) ;
  assign n25130 = ( n3617 & ~n8491 ) | ( n3617 & n25129 ) | ( ~n8491 & n25129 ) ;
  assign n25131 = n4971 | n11540 ;
  assign n25132 = n25131 ^ n23265 ^ 1'b0 ;
  assign n25133 = n25132 ^ n21811 ^ n20187 ;
  assign n25134 = n17478 ^ n13313 ^ 1'b0 ;
  assign n25135 = n6525 | n25134 ;
  assign n25136 = n11792 | n14061 ;
  assign n25137 = n25136 ^ n20498 ^ n1635 ;
  assign n25138 = n7860 & ~n25137 ;
  assign n25139 = ( n3315 & n15555 ) | ( n3315 & n24364 ) | ( n15555 & n24364 ) ;
  assign n25140 = n5232 ^ n2376 ^ n1621 ;
  assign n25141 = n15766 ^ n12753 ^ n3946 ;
  assign n25142 = ( n2215 & n25140 ) | ( n2215 & ~n25141 ) | ( n25140 & ~n25141 ) ;
  assign n25143 = n25142 ^ n23057 ^ n7088 ;
  assign n25146 = n2973 ^ n2222 ^ n1952 ;
  assign n25145 = n19008 ^ n4674 ^ 1'b0 ;
  assign n25144 = n22395 ^ n417 ^ 1'b0 ;
  assign n25147 = n25146 ^ n25145 ^ n25144 ;
  assign n25148 = ( ~n371 & n5228 ) | ( ~n371 & n13157 ) | ( n5228 & n13157 ) ;
  assign n25149 = n20622 & ~n25148 ;
  assign n25150 = ( n2392 & n15613 ) | ( n2392 & ~n21191 ) | ( n15613 & ~n21191 ) ;
  assign n25151 = ( ~n2671 & n21268 ) | ( ~n2671 & n25150 ) | ( n21268 & n25150 ) ;
  assign n25152 = n1880 & ~n10636 ;
  assign n25153 = ~n14862 & n25152 ;
  assign n25154 = n11871 ^ n9567 ^ n509 ;
  assign n25155 = ( n496 & ~n18761 ) | ( n496 & n25154 ) | ( ~n18761 & n25154 ) ;
  assign n25157 = n13967 ^ n1562 ^ n201 ;
  assign n25156 = n16245 ^ n13969 ^ n2102 ;
  assign n25158 = n25157 ^ n25156 ^ 1'b0 ;
  assign n25159 = ( n25153 & n25155 ) | ( n25153 & n25158 ) | ( n25155 & n25158 ) ;
  assign n25160 = n13924 ^ n8547 ^ n7551 ;
  assign n25161 = n1183 | n25160 ;
  assign n25162 = n9028 | n25161 ;
  assign n25163 = n25162 ^ n20481 ^ 1'b0 ;
  assign n25164 = ~n25159 & n25163 ;
  assign n25165 = ( n2901 & ~n4015 ) | ( n2901 & n4120 ) | ( ~n4015 & n4120 ) ;
  assign n25166 = n25165 ^ n11975 ^ 1'b0 ;
  assign n25167 = n15978 ^ n8702 ^ 1'b0 ;
  assign n25168 = n1911 & ~n25167 ;
  assign n25169 = n25168 ^ n15907 ^ 1'b0 ;
  assign n25170 = n238 & n10358 ;
  assign n25171 = ~n14220 & n25170 ;
  assign n25172 = n7592 & n25171 ;
  assign n25173 = n11837 ^ n10092 ^ n994 ;
  assign n25174 = n25173 ^ n16436 ^ n5851 ;
  assign n25175 = n4968 ^ n3748 ^ n3642 ;
  assign n25176 = n22151 ^ n5024 ^ 1'b0 ;
  assign n25177 = ( n898 & n5148 ) | ( n898 & ~n5753 ) | ( n5148 & ~n5753 ) ;
  assign n25178 = ( n6150 & n20484 ) | ( n6150 & ~n25177 ) | ( n20484 & ~n25177 ) ;
  assign n25179 = ( n6931 & n22131 ) | ( n6931 & n25178 ) | ( n22131 & n25178 ) ;
  assign n25180 = ( n7220 & ~n12913 ) | ( n7220 & n25179 ) | ( ~n12913 & n25179 ) ;
  assign n25181 = ( ~n9317 & n14378 ) | ( ~n9317 & n18366 ) | ( n14378 & n18366 ) ;
  assign n25182 = n4666 & ~n17019 ;
  assign n25183 = ~n25181 & n25182 ;
  assign n25184 = n6859 & ~n23755 ;
  assign n25185 = n25184 ^ n21747 ^ 1'b0 ;
  assign n25186 = n13914 ^ n13415 ^ n245 ;
  assign n25187 = n3917 | n21973 ;
  assign n25188 = n19942 ^ n7357 ^ 1'b0 ;
  assign n25189 = n2713 | n25188 ;
  assign n25190 = n25189 ^ n13956 ^ 1'b0 ;
  assign n25191 = n24938 ^ n23704 ^ n18950 ;
  assign n25192 = n11258 ^ n6434 ^ 1'b0 ;
  assign n25193 = n24384 & ~n25192 ;
  assign n25194 = n2868 | n9942 ;
  assign n25195 = n25194 ^ n9287 ^ 1'b0 ;
  assign n25196 = n21204 ^ n6823 ^ x63 ;
  assign n25197 = n3117 | n5692 ;
  assign n25198 = n25197 ^ n15905 ^ 1'b0 ;
  assign n25199 = ( n209 & n12278 ) | ( n209 & ~n25198 ) | ( n12278 & ~n25198 ) ;
  assign n25200 = n19142 ^ n18846 ^ n7961 ;
  assign n25201 = n4448 ^ n613 ^ 1'b0 ;
  assign n25202 = n5080 & ~n10340 ;
  assign n25203 = n25202 ^ n4752 ^ 1'b0 ;
  assign n25204 = ( n10916 & n13608 ) | ( n10916 & ~n16136 ) | ( n13608 & ~n16136 ) ;
  assign n25205 = n25204 ^ n5997 ^ 1'b0 ;
  assign n25206 = n25205 ^ n23679 ^ n10340 ;
  assign n25207 = ~n6697 & n11749 ;
  assign n25208 = n25207 ^ n9821 ^ 1'b0 ;
  assign n25209 = n11624 & n13104 ;
  assign n25210 = n25209 ^ n16138 ^ 1'b0 ;
  assign n25211 = ( ~n22370 & n25208 ) | ( ~n22370 & n25210 ) | ( n25208 & n25210 ) ;
  assign n25212 = n4712 & n4738 ;
  assign n25213 = n25212 ^ n12943 ^ n4263 ;
  assign n25214 = x111 & n25213 ;
  assign n25215 = n1648 | n6547 ;
  assign n25216 = n10176 & ~n25215 ;
  assign n25217 = n23803 ^ n453 ^ 1'b0 ;
  assign n25218 = n18032 & ~n25217 ;
  assign n25219 = n23731 ^ n2971 ^ 1'b0 ;
  assign n25220 = n9434 & ~n25219 ;
  assign n25221 = ( n11536 & n13830 ) | ( n11536 & n25220 ) | ( n13830 & n25220 ) ;
  assign n25222 = n3705 & n25221 ;
  assign n25223 = n25222 ^ n17946 ^ 1'b0 ;
  assign n25224 = n8339 & n13643 ;
  assign n25225 = n18185 ^ n16220 ^ n9942 ;
  assign n25228 = n24725 ^ n1531 ^ 1'b0 ;
  assign n25226 = n22409 ^ n14840 ^ n3525 ;
  assign n25227 = ~n4790 & n25226 ;
  assign n25229 = n25228 ^ n25227 ^ 1'b0 ;
  assign n25230 = ( n15550 & n24328 ) | ( n15550 & n25229 ) | ( n24328 & n25229 ) ;
  assign n25231 = ( ~x62 & n7059 ) | ( ~x62 & n19207 ) | ( n7059 & n19207 ) ;
  assign n25232 = ( ~n2889 & n7914 ) | ( ~n2889 & n14067 ) | ( n7914 & n14067 ) ;
  assign n25233 = ( n8958 & n25231 ) | ( n8958 & n25232 ) | ( n25231 & n25232 ) ;
  assign n25234 = n23195 ^ n9658 ^ n8144 ;
  assign n25235 = n13998 | n25234 ;
  assign n25236 = n25235 ^ n14059 ^ 1'b0 ;
  assign n25237 = n25236 ^ n13437 ^ n9261 ;
  assign n25239 = ( ~n902 & n4031 ) | ( ~n902 & n22031 ) | ( n4031 & n22031 ) ;
  assign n25240 = n25239 ^ n5087 ^ 1'b0 ;
  assign n25238 = n2147 | n21133 ;
  assign n25241 = n25240 ^ n25238 ^ 1'b0 ;
  assign n25242 = n9934 ^ x41 ^ 1'b0 ;
  assign n25243 = ~n25241 & n25242 ;
  assign n25244 = n4948 ^ n4784 ^ 1'b0 ;
  assign n25245 = ( n2504 & n6538 ) | ( n2504 & n25244 ) | ( n6538 & n25244 ) ;
  assign n25246 = n24586 ^ n17450 ^ n4217 ;
  assign n25247 = n9412 ^ n7702 ^ n6333 ;
  assign n25248 = n19101 & ~n22289 ;
  assign n25249 = n25247 & n25248 ;
  assign n25250 = ( ~n2454 & n25246 ) | ( ~n2454 & n25249 ) | ( n25246 & n25249 ) ;
  assign n25251 = n13743 ^ n2931 ^ 1'b0 ;
  assign n25252 = n14664 ^ n8878 ^ n667 ;
  assign n25253 = n5909 ^ n1899 ^ 1'b0 ;
  assign n25254 = n14088 & n25253 ;
  assign n25255 = n2842 & ~n4814 ;
  assign n25256 = ~n5090 & n25255 ;
  assign n25257 = n24955 ^ n21767 ^ n15352 ;
  assign n25258 = n21692 ^ n7564 ^ 1'b0 ;
  assign n25259 = n7996 & ~n25258 ;
  assign n25260 = n25259 ^ n21608 ^ n1685 ;
  assign n25261 = n18813 ^ n8809 ^ n5731 ;
  assign n25262 = n21267 ^ n18891 ^ 1'b0 ;
  assign n25263 = ( ~n19758 & n25261 ) | ( ~n19758 & n25262 ) | ( n25261 & n25262 ) ;
  assign n25264 = n14115 ^ n14113 ^ 1'b0 ;
  assign n25265 = ( n10900 & n12340 ) | ( n10900 & n13147 ) | ( n12340 & n13147 ) ;
  assign n25266 = n394 & ~n3460 ;
  assign n25267 = n24095 | n25266 ;
  assign n25268 = ( ~n2514 & n3247 ) | ( ~n2514 & n13122 ) | ( n3247 & n13122 ) ;
  assign n25269 = ( n3537 & ~n3991 ) | ( n3537 & n25268 ) | ( ~n3991 & n25268 ) ;
  assign n25270 = n2047 | n3629 ;
  assign n25271 = n25269 & ~n25270 ;
  assign n25272 = ( n8742 & n9696 ) | ( n8742 & n23621 ) | ( n9696 & n23621 ) ;
  assign n25273 = n8981 & n25272 ;
  assign n25274 = ( ~n8307 & n13815 ) | ( ~n8307 & n14006 ) | ( n13815 & n14006 ) ;
  assign n25275 = ( n19683 & n20530 ) | ( n19683 & n25274 ) | ( n20530 & n25274 ) ;
  assign n25276 = n25275 ^ n14148 ^ n9758 ;
  assign n25277 = ~n4109 & n25276 ;
  assign n25278 = n25277 ^ n10693 ^ 1'b0 ;
  assign n25279 = n7834 | n12094 ;
  assign n25280 = n11448 & ~n25279 ;
  assign n25281 = n25280 ^ n16184 ^ n2541 ;
  assign n25282 = n25281 ^ n7404 ^ n870 ;
  assign n25283 = n22637 ^ n3674 ^ 1'b0 ;
  assign n25284 = ~n25282 & n25283 ;
  assign n25285 = n21402 ^ n13331 ^ 1'b0 ;
  assign n25286 = n1174 | n25285 ;
  assign n25287 = n21371 ^ n19264 ^ n1543 ;
  assign n25288 = n25287 ^ n12208 ^ n2942 ;
  assign n25289 = ( n5897 & ~n25286 ) | ( n5897 & n25288 ) | ( ~n25286 & n25288 ) ;
  assign n25290 = n20545 ^ n19668 ^ n4805 ;
  assign n25291 = n15993 ^ n3309 ^ 1'b0 ;
  assign n25292 = n23564 & n25291 ;
  assign n25293 = n5243 & ~n14946 ;
  assign n25294 = ~n8944 & n25293 ;
  assign n25295 = ( n269 & ~n6302 ) | ( n269 & n25294 ) | ( ~n6302 & n25294 ) ;
  assign n25298 = n9897 | n12449 ;
  assign n25299 = n11448 & ~n25298 ;
  assign n25296 = n9202 | n14425 ;
  assign n25297 = n25296 ^ n22211 ^ n15864 ;
  assign n25300 = n25299 ^ n25297 ^ n1264 ;
  assign n25301 = n9334 ^ n715 ^ 1'b0 ;
  assign n25302 = ~n14598 & n25301 ;
  assign n25303 = ( n2780 & n10469 ) | ( n2780 & ~n24045 ) | ( n10469 & ~n24045 ) ;
  assign n25304 = n7378 | n25303 ;
  assign n25305 = n5311 | n25304 ;
  assign n25306 = n5878 & n23416 ;
  assign n25307 = n20390 ^ n8082 ^ n5757 ;
  assign n25308 = ( n3041 & ~n4567 ) | ( n3041 & n5310 ) | ( ~n4567 & n5310 ) ;
  assign n25309 = n25308 ^ n14130 ^ 1'b0 ;
  assign n25310 = n11304 ^ n3470 ^ n1335 ;
  assign n25311 = n25310 ^ n9919 ^ n9167 ;
  assign n25312 = n2645 & ~n7087 ;
  assign n25313 = ~n25239 & n25312 ;
  assign n25314 = n25313 ^ n14820 ^ n4801 ;
  assign n25317 = n1626 & ~n3285 ;
  assign n25318 = n25317 ^ n2243 ^ 1'b0 ;
  assign n25315 = n3310 ^ n1861 ^ 1'b0 ;
  assign n25316 = n4967 | n25315 ;
  assign n25319 = n25318 ^ n25316 ^ n5358 ;
  assign n25320 = ( ~n2169 & n16550 ) | ( ~n2169 & n25319 ) | ( n16550 & n25319 ) ;
  assign n25321 = n25320 ^ n18138 ^ 1'b0 ;
  assign n25322 = n25321 ^ n24787 ^ n18739 ;
  assign n25324 = n3212 | n8342 ;
  assign n25323 = ( ~n17737 & n17860 ) | ( ~n17737 & n21738 ) | ( n17860 & n21738 ) ;
  assign n25325 = n25324 ^ n25323 ^ n2214 ;
  assign n25326 = n25325 ^ n25088 ^ 1'b0 ;
  assign n25327 = n2242 & n19221 ;
  assign n25328 = ~n10418 & n25327 ;
  assign n25329 = n23699 ^ n2536 ^ 1'b0 ;
  assign n25330 = n15110 ^ n2875 ^ n767 ;
  assign n25331 = n25330 ^ n3340 ^ 1'b0 ;
  assign n25332 = ~n5793 & n15411 ;
  assign n25333 = ~n25331 & n25332 ;
  assign n25334 = ( n2353 & ~n4873 ) | ( n2353 & n11512 ) | ( ~n4873 & n11512 ) ;
  assign n25335 = n25334 ^ n13357 ^ n7479 ;
  assign n25336 = ( n5859 & n6098 ) | ( n5859 & ~n17169 ) | ( n6098 & ~n17169 ) ;
  assign n25337 = n850 & n7359 ;
  assign n25338 = ~n5918 & n12296 ;
  assign n25339 = ~n4992 & n10132 ;
  assign n25340 = n25339 ^ n6939 ^ 1'b0 ;
  assign n25341 = n25340 ^ n5722 ^ 1'b0 ;
  assign n25342 = n25338 & n25341 ;
  assign n25343 = n25337 | n25342 ;
  assign n25344 = n25336 & n25343 ;
  assign n25345 = n6645 | n24453 ;
  assign n25346 = ( ~n1484 & n21147 ) | ( ~n1484 & n21658 ) | ( n21147 & n21658 ) ;
  assign n25347 = ( n5800 & ~n15324 ) | ( n5800 & n25346 ) | ( ~n15324 & n25346 ) ;
  assign n25348 = n23592 ^ n10311 ^ n640 ;
  assign n25349 = n25348 ^ n10739 ^ n820 ;
  assign n25350 = ( ~n1967 & n12011 ) | ( ~n1967 & n25349 ) | ( n12011 & n25349 ) ;
  assign n25351 = n8133 & ~n13239 ;
  assign n25352 = n2800 & n25351 ;
  assign n25353 = n24405 ^ x38 ^ 1'b0 ;
  assign n25354 = ~n25352 & n25353 ;
  assign n25355 = n25354 ^ n5390 ^ 1'b0 ;
  assign n25356 = n22251 & n25355 ;
  assign n25357 = n8646 & n25023 ;
  assign n25358 = ~n24959 & n25357 ;
  assign n25359 = n23169 ^ n12354 ^ n11627 ;
  assign n25360 = n25359 ^ n8090 ^ 1'b0 ;
  assign n25361 = ~n18462 & n25360 ;
  assign n25362 = ~n13941 & n25361 ;
  assign n25363 = n3768 | n4948 ;
  assign n25364 = n1414 & ~n25363 ;
  assign n25365 = ( n14299 & n17350 ) | ( n14299 & ~n25364 ) | ( n17350 & ~n25364 ) ;
  assign n25366 = n25365 ^ n16969 ^ 1'b0 ;
  assign n25367 = ~n6082 & n19815 ;
  assign n25368 = n25367 ^ n14646 ^ n8234 ;
  assign n25369 = ( n3536 & ~n10968 ) | ( n3536 & n25368 ) | ( ~n10968 & n25368 ) ;
  assign n25376 = n3939 | n4634 ;
  assign n25377 = n9860 | n25376 ;
  assign n25378 = n25377 ^ n3100 ^ 1'b0 ;
  assign n25371 = n1735 | n10202 ;
  assign n25372 = n6826 & ~n25371 ;
  assign n25373 = ( n509 & n12980 ) | ( n509 & n25372 ) | ( n12980 & n25372 ) ;
  assign n25374 = n25373 ^ n6864 ^ 1'b0 ;
  assign n25370 = ( n7159 & ~n13439 ) | ( n7159 & n19862 ) | ( ~n13439 & n19862 ) ;
  assign n25375 = n25374 ^ n25370 ^ 1'b0 ;
  assign n25379 = n25378 ^ n25375 ^ n8056 ;
  assign n25380 = ( n18709 & n25369 ) | ( n18709 & ~n25379 ) | ( n25369 & ~n25379 ) ;
  assign n25381 = ( x1 & n8890 ) | ( x1 & ~n15963 ) | ( n8890 & ~n15963 ) ;
  assign n25382 = n19159 ^ n10557 ^ n1703 ;
  assign n25383 = n7091 & ~n10276 ;
  assign n25384 = ~n11150 & n14323 ;
  assign n25385 = n25384 ^ n17725 ^ 1'b0 ;
  assign n25386 = n5801 & ~n23116 ;
  assign n25387 = n25386 ^ n7384 ^ 1'b0 ;
  assign n25388 = ( n870 & n3384 ) | ( n870 & ~n3973 ) | ( n3384 & ~n3973 ) ;
  assign n25389 = n1064 & ~n25388 ;
  assign n25390 = ~n13051 & n25389 ;
  assign n25391 = ( n2842 & ~n3300 ) | ( n2842 & n7343 ) | ( ~n3300 & n7343 ) ;
  assign n25392 = n8946 & n25391 ;
  assign n25393 = n25390 & n25392 ;
  assign n25394 = n9871 & n25393 ;
  assign n25395 = n25394 ^ n10784 ^ n1563 ;
  assign n25396 = n25395 ^ n16267 ^ n9497 ;
  assign n25397 = n10801 ^ n5604 ^ 1'b0 ;
  assign n25398 = n4199 ^ n275 ^ 1'b0 ;
  assign n25399 = n20792 & n23639 ;
  assign n25400 = n25399 ^ n9037 ^ 1'b0 ;
  assign n25401 = ( n5662 & n25398 ) | ( n5662 & ~n25400 ) | ( n25398 & ~n25400 ) ;
  assign n25402 = ( n5243 & n5740 ) | ( n5243 & n9220 ) | ( n5740 & n9220 ) ;
  assign n25403 = ( ~n4154 & n4872 ) | ( ~n4154 & n7388 ) | ( n4872 & n7388 ) ;
  assign n25404 = n25403 ^ n19427 ^ 1'b0 ;
  assign n25405 = n13122 ^ n8393 ^ n2733 ;
  assign n25406 = n10643 ^ n1048 ^ 1'b0 ;
  assign n25407 = n25405 & ~n25406 ;
  assign n25408 = n24363 ^ n22115 ^ 1'b0 ;
  assign n25409 = ( n2957 & n15703 ) | ( n2957 & n16120 ) | ( n15703 & n16120 ) ;
  assign n25410 = n7454 ^ n4742 ^ n141 ;
  assign n25411 = ( n6887 & n10416 ) | ( n6887 & ~n25410 ) | ( n10416 & ~n25410 ) ;
  assign n25412 = ~n8214 & n11819 ;
  assign n25413 = ~n11743 & n18739 ;
  assign n25414 = ( n6507 & n20499 ) | ( n6507 & ~n25413 ) | ( n20499 & ~n25413 ) ;
  assign n25415 = n24367 ^ n16338 ^ n7176 ;
  assign n25416 = ( ~n1288 & n15644 ) | ( ~n1288 & n25415 ) | ( n15644 & n25415 ) ;
  assign n25417 = ( x8 & n6215 ) | ( x8 & ~n25416 ) | ( n6215 & ~n25416 ) ;
  assign n25418 = n4458 & n9052 ;
  assign n25419 = ( ~n1120 & n7569 ) | ( ~n1120 & n15173 ) | ( n7569 & n15173 ) ;
  assign n25420 = n15110 & n16566 ;
  assign n25421 = ( n25418 & n25419 ) | ( n25418 & n25420 ) | ( n25419 & n25420 ) ;
  assign n25422 = n12960 ^ n1956 ^ 1'b0 ;
  assign n25423 = n23299 ^ n5491 ^ 1'b0 ;
  assign n25424 = n9599 & n25423 ;
  assign n25425 = ( ~n13865 & n25422 ) | ( ~n13865 & n25424 ) | ( n25422 & n25424 ) ;
  assign n25426 = n21334 ^ n16693 ^ n15218 ;
  assign n25427 = n25426 ^ n20248 ^ n12206 ;
  assign n25428 = n25427 ^ n9297 ^ 1'b0 ;
  assign n25429 = n9247 & ~n25428 ;
  assign n25433 = ( n10307 & n14266 ) | ( n10307 & ~n15686 ) | ( n14266 & ~n15686 ) ;
  assign n25430 = n953 | n7313 ;
  assign n25431 = n7412 | n25430 ;
  assign n25432 = n10272 & n25431 ;
  assign n25434 = n25433 ^ n25432 ^ 1'b0 ;
  assign n25435 = n7185 & n7874 ;
  assign n25436 = ~n16379 & n25435 ;
  assign n25437 = ( n14998 & ~n16155 ) | ( n14998 & n25436 ) | ( ~n16155 & n25436 ) ;
  assign n25438 = ~n20855 & n25437 ;
  assign n25439 = n25438 ^ n16993 ^ 1'b0 ;
  assign n25440 = n2372 | n25439 ;
  assign n25441 = n11458 ^ n6844 ^ n5381 ;
  assign n25442 = n25441 ^ n16275 ^ n12174 ;
  assign n25443 = ( n4810 & n12132 ) | ( n4810 & n24093 ) | ( n12132 & n24093 ) ;
  assign n25444 = n25443 ^ n12560 ^ n2080 ;
  assign n25445 = ( n2844 & n9549 ) | ( n2844 & n19370 ) | ( n9549 & n19370 ) ;
  assign n25446 = n25445 ^ n13236 ^ n10979 ;
  assign n25447 = n23725 ^ n23078 ^ n7957 ;
  assign n25448 = ~n1082 & n3998 ;
  assign n25449 = n25334 ^ n9630 ^ n744 ;
  assign n25450 = n15487 | n25449 ;
  assign n25451 = ( ~n3354 & n25448 ) | ( ~n3354 & n25450 ) | ( n25448 & n25450 ) ;
  assign n25452 = n15103 ^ n413 ^ 1'b0 ;
  assign n25453 = n13421 | n25452 ;
  assign n25454 = n15823 ^ n3999 ^ 1'b0 ;
  assign n25455 = ~n10181 & n25454 ;
  assign n25456 = n19990 ^ n19142 ^ n11015 ;
  assign n25457 = ( n1501 & n14336 ) | ( n1501 & ~n24278 ) | ( n14336 & ~n24278 ) ;
  assign n25459 = ( ~n755 & n2811 ) | ( ~n755 & n18814 ) | ( n2811 & n18814 ) ;
  assign n25460 = ~n17014 & n25459 ;
  assign n25461 = ~n20464 & n25460 ;
  assign n25462 = ( n5344 & n7785 ) | ( n5344 & ~n25461 ) | ( n7785 & ~n25461 ) ;
  assign n25463 = n25462 ^ n25025 ^ n13483 ;
  assign n25458 = ( ~n1395 & n8292 ) | ( ~n1395 & n15314 ) | ( n8292 & n15314 ) ;
  assign n25464 = n25463 ^ n25458 ^ n12263 ;
  assign n25465 = n4932 ^ x81 ^ 1'b0 ;
  assign n25466 = ( n5062 & ~n13218 ) | ( n5062 & n25340 ) | ( ~n13218 & n25340 ) ;
  assign n25467 = n25466 ^ n4730 ^ 1'b0 ;
  assign n25468 = n17886 ^ n13314 ^ n5746 ;
  assign n25469 = ( ~n1422 & n12055 ) | ( ~n1422 & n25468 ) | ( n12055 & n25468 ) ;
  assign n25470 = n6832 ^ n5621 ^ 1'b0 ;
  assign n25474 = n3347 ^ n3321 ^ 1'b0 ;
  assign n25475 = n7906 | n25474 ;
  assign n25471 = ( ~n5313 & n8432 ) | ( ~n5313 & n21973 ) | ( n8432 & n21973 ) ;
  assign n25472 = n25471 ^ n24070 ^ 1'b0 ;
  assign n25473 = n14200 | n25472 ;
  assign n25476 = n25475 ^ n25473 ^ n17949 ;
  assign n25477 = n5689 ^ n5591 ^ n4014 ;
  assign n25478 = ( n8038 & ~n23250 ) | ( n8038 & n25477 ) | ( ~n23250 & n25477 ) ;
  assign n25479 = n21500 ^ n16155 ^ n13578 ;
  assign n25480 = n15320 ^ n1907 ^ 1'b0 ;
  assign n25481 = n25480 ^ n10383 ^ 1'b0 ;
  assign n25482 = n25481 ^ n19441 ^ n7859 ;
  assign n25483 = n19830 | n25482 ;
  assign n25484 = n12009 ^ n8082 ^ 1'b0 ;
  assign n25485 = n232 & ~n25484 ;
  assign n25486 = ( n1676 & n3050 ) | ( n1676 & ~n3399 ) | ( n3050 & ~n3399 ) ;
  assign n25487 = n220 | n25486 ;
  assign n25488 = n25485 | n25487 ;
  assign n25489 = n4346 ^ n3503 ^ n1819 ;
  assign n25490 = n9402 ^ n2779 ^ 1'b0 ;
  assign n25491 = n25489 | n25490 ;
  assign n25492 = n17276 ^ n7759 ^ n3815 ;
  assign n25493 = ( n21984 & n25491 ) | ( n21984 & n25492 ) | ( n25491 & n25492 ) ;
  assign n25494 = n14784 ^ n3935 ^ 1'b0 ;
  assign n25495 = n4784 & ~n25494 ;
  assign n25496 = n15953 ^ n14819 ^ n10023 ;
  assign n25497 = n25495 | n25496 ;
  assign n25498 = n12816 ^ n10767 ^ n8730 ;
  assign n25499 = ( n21879 & n25051 ) | ( n21879 & n25498 ) | ( n25051 & n25498 ) ;
  assign n25500 = n14937 ^ n3516 ^ n176 ;
  assign n25501 = n21924 ^ n18398 ^ 1'b0 ;
  assign n25502 = ~n7118 & n25501 ;
  assign n25503 = ~n13916 & n25502 ;
  assign n25504 = n10140 | n14117 ;
  assign n25505 = n5117 & ~n18728 ;
  assign n25506 = n25504 & n25505 ;
  assign n25507 = ~n3511 & n24938 ;
  assign n25508 = n782 | n14378 ;
  assign n25509 = n6120 & ~n25508 ;
  assign n25510 = n12011 ^ n5346 ^ 1'b0 ;
  assign n25511 = n25510 ^ n20074 ^ n11478 ;
  assign n25512 = n7202 & ~n10955 ;
  assign n25513 = n25512 ^ n8555 ^ 1'b0 ;
  assign n25514 = ( ~n2639 & n3935 ) | ( ~n2639 & n25513 ) | ( n3935 & n25513 ) ;
  assign n25515 = n17500 ^ n3651 ^ 1'b0 ;
  assign n25516 = ( ~n5658 & n8760 ) | ( ~n5658 & n13319 ) | ( n8760 & n13319 ) ;
  assign n25517 = n2276 & n16076 ;
  assign n25518 = n25517 ^ n11937 ^ 1'b0 ;
  assign n25519 = ~n1912 & n13260 ;
  assign n25520 = n25519 ^ n20596 ^ 1'b0 ;
  assign n25521 = ( ~n5209 & n6434 ) | ( ~n5209 & n9200 ) | ( n6434 & n9200 ) ;
  assign n25522 = n22413 ^ n16062 ^ n4015 ;
  assign n25523 = ( n8126 & ~n25521 ) | ( n8126 & n25522 ) | ( ~n25521 & n25522 ) ;
  assign n25524 = n13144 ^ n406 ^ 1'b0 ;
  assign n25525 = n25523 | n25524 ;
  assign n25526 = n25525 ^ n4568 ^ n2097 ;
  assign n25528 = n7920 ^ n3766 ^ 1'b0 ;
  assign n25529 = ~n22779 & n25528 ;
  assign n25527 = ( n667 & n5539 ) | ( n667 & ~n7806 ) | ( n5539 & ~n7806 ) ;
  assign n25530 = n25529 ^ n25527 ^ n6960 ;
  assign n25531 = n14880 ^ n4844 ^ 1'b0 ;
  assign n25532 = n20729 ^ n15900 ^ n3478 ;
  assign n25533 = n8863 | n10484 ;
  assign n25534 = n25532 | n25533 ;
  assign n25535 = ( n21326 & n25531 ) | ( n21326 & n25534 ) | ( n25531 & n25534 ) ;
  assign n25536 = ~n5499 & n6430 ;
  assign n25537 = n17458 ^ n15979 ^ n6057 ;
  assign n25538 = ( ~n2057 & n25536 ) | ( ~n2057 & n25537 ) | ( n25536 & n25537 ) ;
  assign n25539 = ( n885 & n1619 ) | ( n885 & n5287 ) | ( n1619 & n5287 ) ;
  assign n25540 = ( ~n545 & n6052 ) | ( ~n545 & n25539 ) | ( n6052 & n25539 ) ;
  assign n25541 = n11988 | n25540 ;
  assign n25542 = n10498 ^ n8559 ^ n5969 ;
  assign n25543 = n6139 | n6179 ;
  assign n25544 = n24175 & ~n25543 ;
  assign n25545 = n25104 ^ n11568 ^ 1'b0 ;
  assign n25546 = n21079 & ~n25545 ;
  assign n25547 = n1788 ^ n1378 ^ 1'b0 ;
  assign n25548 = ~n15259 & n25547 ;
  assign n25549 = ~n900 & n20061 ;
  assign n25550 = n3357 & n25549 ;
  assign n25551 = ( n18331 & ~n24595 ) | ( n18331 & n25550 ) | ( ~n24595 & n25550 ) ;
  assign n25555 = n14943 ^ n13417 ^ n8433 ;
  assign n25553 = n9389 & ~n12983 ;
  assign n25554 = n10962 & n25553 ;
  assign n25552 = ( ~n9659 & n12613 ) | ( ~n9659 & n24767 ) | ( n12613 & n24767 ) ;
  assign n25556 = n25555 ^ n25554 ^ n25552 ;
  assign n25557 = n20985 ^ n2315 ^ 1'b0 ;
  assign n25560 = ( n3641 & n7994 ) | ( n3641 & ~n9863 ) | ( n7994 & ~n9863 ) ;
  assign n25558 = ( n2534 & ~n3295 ) | ( n2534 & n12176 ) | ( ~n3295 & n12176 ) ;
  assign n25559 = n25558 ^ n19642 ^ n1538 ;
  assign n25561 = n25560 ^ n25559 ^ n728 ;
  assign n25562 = n25561 ^ n15211 ^ n5615 ;
  assign n25563 = n5125 ^ n1314 ^ 1'b0 ;
  assign n25564 = ( n8409 & ~n18019 ) | ( n8409 & n25563 ) | ( ~n18019 & n25563 ) ;
  assign n25565 = n12004 ^ n6368 ^ 1'b0 ;
  assign n25566 = ( n6537 & ~n18330 ) | ( n6537 & n22687 ) | ( ~n18330 & n22687 ) ;
  assign n25567 = n5368 | n8869 ;
  assign n25568 = n25566 | n25567 ;
  assign n25569 = n21067 ^ n16965 ^ n226 ;
  assign n25570 = n1399 & ~n9906 ;
  assign n25571 = ~n25569 & n25570 ;
  assign n25572 = n2429 & ~n13811 ;
  assign n25573 = n20499 & n25572 ;
  assign n25574 = n25573 ^ n14148 ^ n12717 ;
  assign n25575 = n16548 ^ n12781 ^ n9480 ;
  assign n25576 = ( n3661 & ~n11503 ) | ( n3661 & n18108 ) | ( ~n11503 & n18108 ) ;
  assign n25577 = ( n7059 & n9555 ) | ( n7059 & n15587 ) | ( n9555 & n15587 ) ;
  assign n25578 = ( ~n241 & n1267 ) | ( ~n241 & n8374 ) | ( n1267 & n8374 ) ;
  assign n25579 = n5421 ^ n3352 ^ n967 ;
  assign n25580 = n20283 ^ n7938 ^ 1'b0 ;
  assign n25581 = ~n25579 & n25580 ;
  assign n25582 = n25581 ^ n13845 ^ 1'b0 ;
  assign n25583 = n15231 ^ n4731 ^ n729 ;
  assign n25584 = ( n17843 & ~n25582 ) | ( n17843 & n25583 ) | ( ~n25582 & n25583 ) ;
  assign n25585 = ( ~n3066 & n6033 ) | ( ~n3066 & n25584 ) | ( n6033 & n25584 ) ;
  assign n25586 = n6058 & n20059 ;
  assign n25587 = ( n1695 & n6631 ) | ( n1695 & n9291 ) | ( n6631 & n9291 ) ;
  assign n25588 = ( n3535 & n4600 ) | ( n3535 & ~n12565 ) | ( n4600 & ~n12565 ) ;
  assign n25589 = n25588 ^ n2331 ^ n912 ;
  assign n25590 = ( ~n2372 & n9326 ) | ( ~n2372 & n25589 ) | ( n9326 & n25589 ) ;
  assign n25591 = n25590 ^ n16155 ^ 1'b0 ;
  assign n25592 = n25587 & n25591 ;
  assign n25593 = n2705 & n25287 ;
  assign n25594 = n25593 ^ n12764 ^ n6742 ;
  assign n25595 = n25594 ^ n9410 ^ 1'b0 ;
  assign n25596 = n12569 ^ n8257 ^ n3192 ;
  assign n25597 = n25596 ^ n11505 ^ n10383 ;
  assign n25598 = n25597 ^ n24357 ^ 1'b0 ;
  assign n25599 = ( ~n6158 & n25595 ) | ( ~n6158 & n25598 ) | ( n25595 & n25598 ) ;
  assign n25600 = n25599 ^ n13365 ^ 1'b0 ;
  assign n25601 = n15773 | n25600 ;
  assign n25602 = n14647 ^ n4746 ^ n3146 ;
  assign n25604 = n18398 ^ n12973 ^ n9079 ;
  assign n25603 = ( x108 & ~n11776 ) | ( x108 & n20170 ) | ( ~n11776 & n20170 ) ;
  assign n25605 = n25604 ^ n25603 ^ n4014 ;
  assign n25606 = n19069 ^ n3328 ^ 1'b0 ;
  assign n25607 = n14232 & ~n25606 ;
  assign n25608 = n342 & n25607 ;
  assign n25609 = n22515 ^ n3270 ^ 1'b0 ;
  assign n25610 = ~n8810 & n25609 ;
  assign n25611 = ( n679 & n17518 ) | ( n679 & n25610 ) | ( n17518 & n25610 ) ;
  assign n25612 = n23255 ^ n19541 ^ n16861 ;
  assign n25613 = n8896 ^ n6228 ^ n1736 ;
  assign n25614 = ( n3853 & ~n14860 ) | ( n3853 & n25613 ) | ( ~n14860 & n25613 ) ;
  assign n25615 = ~n1045 & n4044 ;
  assign n25616 = n21015 & n25615 ;
  assign n25617 = n13450 ^ n11225 ^ n3197 ;
  assign n25618 = n25617 ^ n20263 ^ 1'b0 ;
  assign n25619 = n1793 | n7868 ;
  assign n25620 = n25618 & ~n25619 ;
  assign n25621 = ( n2500 & ~n16790 ) | ( n2500 & n17055 ) | ( ~n16790 & n17055 ) ;
  assign n25622 = n12934 | n25621 ;
  assign n25623 = ( n3738 & n8352 ) | ( n3738 & ~n22370 ) | ( n8352 & ~n22370 ) ;
  assign n25624 = n17207 ^ n8672 ^ 1'b0 ;
  assign n25625 = n17739 ^ n13981 ^ n9998 ;
  assign n25626 = n12845 | n25625 ;
  assign n25627 = n3546 & ~n9919 ;
  assign n25628 = n8152 ^ n5562 ^ n1079 ;
  assign n25629 = n10050 & n17351 ;
  assign n25630 = n25629 ^ n15769 ^ n2863 ;
  assign n25631 = n25628 | n25630 ;
  assign n25632 = ~n6573 & n13729 ;
  assign n25633 = n25632 ^ n6639 ^ 1'b0 ;
  assign n25634 = ( n7445 & ~n7703 ) | ( n7445 & n15474 ) | ( ~n7703 & n15474 ) ;
  assign n25635 = n25634 ^ n22176 ^ 1'b0 ;
  assign n25636 = n4435 & n11516 ;
  assign n25637 = n25636 ^ n24049 ^ 1'b0 ;
  assign n25638 = ( n11121 & n11211 ) | ( n11121 & ~n13664 ) | ( n11211 & ~n13664 ) ;
  assign n25639 = n9355 & ~n14819 ;
  assign n25640 = n25639 ^ n1587 ^ 1'b0 ;
  assign n25641 = ( n17484 & ~n25638 ) | ( n17484 & n25640 ) | ( ~n25638 & n25640 ) ;
  assign n25642 = ( n1470 & ~n19081 ) | ( n1470 & n19673 ) | ( ~n19081 & n19673 ) ;
  assign n25643 = n20261 ^ n17280 ^ n6325 ;
  assign n25644 = n15808 ^ n11886 ^ n8133 ;
  assign n25645 = ~n8787 & n9046 ;
  assign n25646 = n25645 ^ n19849 ^ 1'b0 ;
  assign n25647 = n1009 & n4987 ;
  assign n25648 = ( n9153 & n18779 ) | ( n9153 & n19209 ) | ( n18779 & n19209 ) ;
  assign n25649 = n12522 ^ n11383 ^ n4214 ;
  assign n25650 = n24464 ^ n19262 ^ 1'b0 ;
  assign n25651 = n17872 | n21219 ;
  assign n25652 = n25651 ^ n18149 ^ 1'b0 ;
  assign n25653 = n25652 ^ n13109 ^ 1'b0 ;
  assign n25654 = n3887 & n6018 ;
  assign n25655 = n25364 ^ n8413 ^ 1'b0 ;
  assign n25656 = n2762 & n25655 ;
  assign n25657 = ( n6838 & ~n25654 ) | ( n6838 & n25656 ) | ( ~n25654 & n25656 ) ;
  assign n25658 = n25653 & ~n25657 ;
  assign n25659 = n11613 ^ n8210 ^ 1'b0 ;
  assign n25660 = ~n9986 & n21521 ;
  assign n25661 = ~n5020 & n25660 ;
  assign n25662 = ( n3975 & ~n20616 ) | ( n3975 & n25661 ) | ( ~n20616 & n25661 ) ;
  assign n25663 = n14233 | n18153 ;
  assign n25664 = ( n5477 & n7041 ) | ( n5477 & n25663 ) | ( n7041 & n25663 ) ;
  assign n25665 = n25664 ^ n22236 ^ 1'b0 ;
  assign n25666 = n744 & n25665 ;
  assign n25667 = n16862 & n25666 ;
  assign n25669 = n6721 & ~n19585 ;
  assign n25670 = n25669 ^ n15917 ^ 1'b0 ;
  assign n25668 = ~n8055 & n11137 ;
  assign n25671 = n25670 ^ n25668 ^ 1'b0 ;
  assign n25672 = ( n9344 & ~n15260 ) | ( n9344 & n21005 ) | ( ~n15260 & n21005 ) ;
  assign n25673 = n25672 ^ n9544 ^ n6057 ;
  assign n25674 = n8104 ^ n3090 ^ 1'b0 ;
  assign n25675 = n25674 ^ n13550 ^ n1610 ;
  assign n25677 = n3007 | n4438 ;
  assign n25676 = n20664 ^ n15051 ^ n12903 ;
  assign n25678 = n25677 ^ n25676 ^ n592 ;
  assign n25679 = n16643 ^ n15525 ^ n6182 ;
  assign n25680 = n25679 ^ n639 ^ 1'b0 ;
  assign n25681 = ~n3021 & n23510 ;
  assign n25682 = n25681 ^ n7371 ^ 1'b0 ;
  assign n25683 = n4187 | n23216 ;
  assign n25684 = n9057 ^ n3798 ^ 1'b0 ;
  assign n25685 = ( ~n4919 & n9007 ) | ( ~n4919 & n16127 ) | ( n9007 & n16127 ) ;
  assign n25686 = n25685 ^ n7598 ^ n4220 ;
  assign n25687 = n25686 ^ n22135 ^ n20971 ;
  assign n25688 = n2621 | n23488 ;
  assign n25689 = ~n1773 & n21855 ;
  assign n25690 = n12895 & n25689 ;
  assign n25691 = n14716 ^ n7575 ^ 1'b0 ;
  assign n25692 = ~n14472 & n14792 ;
  assign n25693 = n25691 & n25692 ;
  assign n25694 = ( ~n8067 & n8440 ) | ( ~n8067 & n19196 ) | ( n8440 & n19196 ) ;
  assign n25695 = ( n4860 & ~n11577 ) | ( n4860 & n25694 ) | ( ~n11577 & n25694 ) ;
  assign n25696 = ( ~n1573 & n11756 ) | ( ~n1573 & n25695 ) | ( n11756 & n25695 ) ;
  assign n25697 = ( n6649 & n7975 ) | ( n6649 & n15798 ) | ( n7975 & n15798 ) ;
  assign n25698 = n24344 ^ n8690 ^ n4035 ;
  assign n25699 = n20888 ^ n18569 ^ 1'b0 ;
  assign n25700 = n16297 ^ n16236 ^ n3014 ;
  assign n25701 = n7860 ^ n6411 ^ n1570 ;
  assign n25702 = n25701 ^ n16741 ^ 1'b0 ;
  assign n25703 = n13815 ^ n12134 ^ n6337 ;
  assign n25704 = n23817 ^ n4650 ^ 1'b0 ;
  assign n25705 = n7912 ^ n6311 ^ n1838 ;
  assign n25706 = n25705 ^ n17599 ^ n17354 ;
  assign n25707 = n25706 ^ n8854 ^ n5993 ;
  assign n25708 = n7100 ^ n5494 ^ n2884 ;
  assign n25709 = ( ~n4230 & n25226 ) | ( ~n4230 & n25708 ) | ( n25226 & n25708 ) ;
  assign n25710 = n13594 & n22465 ;
  assign n25711 = n1517 | n12928 ;
  assign n25712 = n25711 ^ n5402 ^ 1'b0 ;
  assign n25713 = ( ~n1743 & n4342 ) | ( ~n1743 & n9249 ) | ( n4342 & n9249 ) ;
  assign n25714 = n23087 | n25713 ;
  assign n25715 = n25712 & ~n25714 ;
  assign n25716 = n10271 & ~n25159 ;
  assign n25717 = n16500 & ~n23419 ;
  assign n25718 = ( n1390 & n1624 ) | ( n1390 & n14429 ) | ( n1624 & n14429 ) ;
  assign n25719 = n25718 ^ n21116 ^ 1'b0 ;
  assign n25721 = n8853 ^ n7076 ^ n3805 ;
  assign n25720 = n2099 | n2167 ;
  assign n25722 = n25721 ^ n25720 ^ n2907 ;
  assign n25723 = n11500 ^ n10670 ^ 1'b0 ;
  assign n25737 = n10561 ^ n7680 ^ n7427 ;
  assign n25731 = ( ~n2488 & n3486 ) | ( ~n2488 & n15593 ) | ( n3486 & n15593 ) ;
  assign n25729 = n6535 & n6656 ;
  assign n25730 = ~n1592 & n25729 ;
  assign n25732 = n25731 ^ n25730 ^ n22040 ;
  assign n25733 = n10280 | n12616 ;
  assign n25734 = n25733 ^ n7869 ^ 1'b0 ;
  assign n25735 = n1544 | n25734 ;
  assign n25736 = n25732 | n25735 ;
  assign n25727 = ( n1617 & n7854 ) | ( n1617 & n23346 ) | ( n7854 & n23346 ) ;
  assign n25725 = n7098 & ~n21657 ;
  assign n25726 = n25725 ^ n13144 ^ n7685 ;
  assign n25724 = n3178 ^ n225 ^ 1'b0 ;
  assign n25728 = n25727 ^ n25726 ^ n25724 ;
  assign n25738 = n25737 ^ n25736 ^ n25728 ;
  assign n25739 = n15960 ^ n8143 ^ 1'b0 ;
  assign n25740 = ~n3090 & n15898 ;
  assign n25741 = n9977 ^ n8488 ^ n2328 ;
  assign n25742 = ~n24815 & n25741 ;
  assign n25743 = ~n16576 & n25742 ;
  assign n25744 = n8046 ^ n5079 ^ 1'b0 ;
  assign n25745 = n25743 | n25744 ;
  assign n25746 = n22505 ^ n17473 ^ n8182 ;
  assign n25747 = x77 & n5409 ;
  assign n25748 = n25747 ^ n12734 ^ n173 ;
  assign n25749 = n24040 ^ n21704 ^ n6261 ;
  assign n25750 = n8531 ^ n2717 ^ 1'b0 ;
  assign n25751 = ( n2948 & n13814 ) | ( n2948 & ~n25750 ) | ( n13814 & ~n25750 ) ;
  assign n25752 = n22733 ^ n15034 ^ n7555 ;
  assign n25753 = ( n2779 & n4234 ) | ( n2779 & n9124 ) | ( n4234 & n9124 ) ;
  assign n25754 = ~n928 & n25753 ;
  assign n25755 = n25754 ^ n7576 ^ 1'b0 ;
  assign n25756 = ( n4886 & ~n5416 ) | ( n4886 & n12904 ) | ( ~n5416 & n12904 ) ;
  assign n25757 = n25756 ^ n13233 ^ 1'b0 ;
  assign n25758 = n13290 ^ n179 ^ 1'b0 ;
  assign n25759 = n12335 & n25758 ;
  assign n25760 = n9262 | n17397 ;
  assign n25761 = n7515 | n25760 ;
  assign n25762 = n25761 ^ n21545 ^ 1'b0 ;
  assign n25763 = n25759 & n25762 ;
  assign n25764 = n14923 ^ n14757 ^ n3040 ;
  assign n25765 = ( n7537 & n12737 ) | ( n7537 & n15171 ) | ( n12737 & n15171 ) ;
  assign n25766 = ( n418 & ~n1883 ) | ( n418 & n11824 ) | ( ~n1883 & n11824 ) ;
  assign n25767 = ( n14278 & n15033 ) | ( n14278 & n25766 ) | ( n15033 & n25766 ) ;
  assign n25768 = n25767 ^ n12325 ^ 1'b0 ;
  assign n25769 = n25765 & ~n25768 ;
  assign n25770 = ( ~n10554 & n12656 ) | ( ~n10554 & n25769 ) | ( n12656 & n25769 ) ;
  assign n25771 = n2970 | n5553 ;
  assign n25772 = n25771 ^ n19150 ^ n14437 ;
  assign n25773 = ( n4934 & ~n8888 ) | ( n4934 & n16230 ) | ( ~n8888 & n16230 ) ;
  assign n25774 = n24875 ^ n9297 ^ 1'b0 ;
  assign n25775 = ~n7108 & n25774 ;
  assign n25776 = n25775 ^ n10406 ^ n10123 ;
  assign n25777 = n22840 ^ n22295 ^ n4264 ;
  assign n25778 = n7296 | n19612 ;
  assign n25779 = ~n12050 & n25778 ;
  assign n25780 = ~n931 & n15976 ;
  assign n25781 = n25780 ^ n18151 ^ 1'b0 ;
  assign n25782 = ~n14351 & n21778 ;
  assign n25783 = n25782 ^ n25603 ^ 1'b0 ;
  assign n25784 = n12622 ^ n934 ^ 1'b0 ;
  assign n25785 = ( n12768 & n17670 ) | ( n12768 & ~n24564 ) | ( n17670 & ~n24564 ) ;
  assign n25786 = n17875 ^ n11568 ^ n275 ;
  assign n25787 = n25786 ^ n6684 ^ n4873 ;
  assign n25788 = ( ~n5068 & n9588 ) | ( ~n5068 & n13762 ) | ( n9588 & n13762 ) ;
  assign n25789 = ( n4585 & n5283 ) | ( n4585 & n5421 ) | ( n5283 & n5421 ) ;
  assign n25790 = n25789 ^ n13767 ^ 1'b0 ;
  assign n25791 = n1466 & ~n18171 ;
  assign n25792 = ~n18005 & n25791 ;
  assign n25797 = ( ~n2125 & n7607 ) | ( ~n2125 & n8443 ) | ( n7607 & n8443 ) ;
  assign n25794 = n3151 | n5442 ;
  assign n25795 = n15570 | n25794 ;
  assign n25793 = ( n4356 & n4556 ) | ( n4356 & n24119 ) | ( n4556 & n24119 ) ;
  assign n25796 = n25795 ^ n25793 ^ n9327 ;
  assign n25798 = n25797 ^ n25796 ^ n11260 ;
  assign n25799 = ~n8748 & n25798 ;
  assign n25800 = n25799 ^ n15894 ^ 1'b0 ;
  assign n25802 = ( n1965 & n14444 ) | ( n1965 & n19365 ) | ( n14444 & n19365 ) ;
  assign n25801 = n3458 & ~n6935 ;
  assign n25803 = n25802 ^ n25801 ^ 1'b0 ;
  assign n25804 = n4858 & n10384 ;
  assign n25805 = ( n16042 & ~n23888 ) | ( n16042 & n25804 ) | ( ~n23888 & n25804 ) ;
  assign n25806 = n12288 ^ n3996 ^ 1'b0 ;
  assign n25807 = n2747 | n6038 ;
  assign n25808 = n25807 ^ n15140 ^ 1'b0 ;
  assign n25809 = n25808 ^ n6334 ^ n3035 ;
  assign n25810 = n4774 & n25809 ;
  assign n25811 = n25810 ^ n21054 ^ n18433 ;
  assign n25812 = n10551 ^ n3864 ^ n3309 ;
  assign n25813 = ( n14184 & n15063 ) | ( n14184 & n25812 ) | ( n15063 & n25812 ) ;
  assign n25814 = ( x22 & n459 ) | ( x22 & ~n20908 ) | ( n459 & ~n20908 ) ;
  assign n25817 = n1112 & ~n16510 ;
  assign n25815 = n16298 ^ n3060 ^ 1'b0 ;
  assign n25816 = n3005 & ~n25815 ;
  assign n25818 = n25817 ^ n25816 ^ 1'b0 ;
  assign n25819 = ( n1095 & ~n2458 ) | ( n1095 & n5377 ) | ( ~n2458 & n5377 ) ;
  assign n25820 = n13241 ^ n5199 ^ 1'b0 ;
  assign n25821 = n25819 & ~n25820 ;
  assign n25822 = ( n3401 & ~n5263 ) | ( n3401 & n10441 ) | ( ~n5263 & n10441 ) ;
  assign n25823 = n25822 ^ n19686 ^ n15824 ;
  assign n25824 = n21179 ^ n11313 ^ n4456 ;
  assign n25825 = n25587 ^ n17291 ^ 1'b0 ;
  assign n25826 = ( n1739 & ~n8876 ) | ( n1739 & n18213 ) | ( ~n8876 & n18213 ) ;
  assign n25827 = ( n14445 & ~n17284 ) | ( n14445 & n25826 ) | ( ~n17284 & n25826 ) ;
  assign n25828 = n3387 & ~n12469 ;
  assign n25829 = n25828 ^ n3520 ^ 1'b0 ;
  assign n25830 = n9802 & n20681 ;
  assign n25831 = n24940 ^ n23570 ^ 1'b0 ;
  assign n25832 = n17695 | n25831 ;
  assign n25833 = ( ~n2780 & n5142 ) | ( ~n2780 & n20941 ) | ( n5142 & n20941 ) ;
  assign n25834 = ~n3063 & n8625 ;
  assign n25835 = n25833 & n25834 ;
  assign n25836 = n7962 & ~n10959 ;
  assign n25837 = n1176 & n25836 ;
  assign n25838 = n23793 ^ n14634 ^ 1'b0 ;
  assign n25839 = n186 | n25838 ;
  assign n25840 = n25839 ^ n20008 ^ 1'b0 ;
  assign n25841 = ~n25837 & n25840 ;
  assign n25842 = ( n5689 & ~n5774 ) | ( n5689 & n11270 ) | ( ~n5774 & n11270 ) ;
  assign n25843 = n7501 ^ n7396 ^ n5644 ;
  assign n25844 = ( n5827 & ~n7721 ) | ( n5827 & n25843 ) | ( ~n7721 & n25843 ) ;
  assign n25845 = ~n602 & n9766 ;
  assign n25846 = n25845 ^ n18958 ^ n17429 ;
  assign n25847 = n25846 ^ n5887 ^ 1'b0 ;
  assign n25848 = n25593 ^ n22809 ^ n18406 ;
  assign n25852 = ~n1625 & n6448 ;
  assign n25849 = n6281 ^ n1152 ^ 1'b0 ;
  assign n25850 = n17704 & n25849 ;
  assign n25851 = n25850 ^ n22414 ^ n19751 ;
  assign n25853 = n25852 ^ n25851 ^ n1525 ;
  assign n25854 = n25021 ^ n13649 ^ 1'b0 ;
  assign n25855 = n17945 ^ n13134 ^ n3568 ;
  assign n25856 = n2384 | n14854 ;
  assign n25857 = n14748 ^ n6771 ^ n1084 ;
  assign n25858 = n25857 ^ n24918 ^ x14 ;
  assign n25859 = ~n447 & n25858 ;
  assign n25860 = n25859 ^ n6077 ^ 1'b0 ;
  assign n25861 = ( n10878 & n25856 ) | ( n10878 & ~n25860 ) | ( n25856 & ~n25860 ) ;
  assign n25862 = n11580 ^ n3304 ^ n1508 ;
  assign n25863 = n21627 ^ n17897 ^ 1'b0 ;
  assign n25864 = ( n23425 & ~n24619 ) | ( n23425 & n25863 ) | ( ~n24619 & n25863 ) ;
  assign n25865 = n3665 & ~n12030 ;
  assign n25866 = n25865 ^ n14254 ^ n5166 ;
  assign n25867 = n15606 ^ n12768 ^ n1031 ;
  assign n25868 = ( n10627 & n10684 ) | ( n10627 & n25867 ) | ( n10684 & n25867 ) ;
  assign n25869 = n1735 | n25868 ;
  assign n25870 = n10459 & ~n25869 ;
  assign n25871 = n843 & n17028 ;
  assign n25872 = ~n13833 & n25871 ;
  assign n25873 = n25872 ^ n10699 ^ n9835 ;
  assign n25874 = ( n8962 & ~n19908 ) | ( n8962 & n23443 ) | ( ~n19908 & n23443 ) ;
  assign n25875 = n25874 ^ n18185 ^ n1813 ;
  assign n25876 = n13256 ^ n8317 ^ 1'b0 ;
  assign n25877 = n12027 ^ n5827 ^ n3988 ;
  assign n25878 = n22574 ^ n15496 ^ n12613 ;
  assign n25879 = n6910 ^ n3816 ^ 1'b0 ;
  assign n25880 = n25879 ^ n3461 ^ 1'b0 ;
  assign n25881 = n1295 & n20028 ;
  assign n25882 = n4358 & n25881 ;
  assign n25883 = n19834 ^ n16568 ^ n4302 ;
  assign n25884 = n17575 ^ n17288 ^ 1'b0 ;
  assign n25885 = n19078 ^ n405 ^ 1'b0 ;
  assign n25886 = n25884 & n25885 ;
  assign n25887 = ( ~n7427 & n25883 ) | ( ~n7427 & n25886 ) | ( n25883 & n25886 ) ;
  assign n25888 = n15349 ^ n9900 ^ n8077 ;
  assign n25889 = ( n2202 & n14278 ) | ( n2202 & ~n18763 ) | ( n14278 & ~n18763 ) ;
  assign n25890 = n25889 ^ n6267 ^ n1612 ;
  assign n25891 = n25890 ^ n3040 ^ n2283 ;
  assign n25892 = ( n2792 & ~n5535 ) | ( n2792 & n25891 ) | ( ~n5535 & n25891 ) ;
  assign n25893 = ~n1959 & n10767 ;
  assign n25894 = ( n10058 & n12392 ) | ( n10058 & ~n25664 ) | ( n12392 & ~n25664 ) ;
  assign n25895 = n1278 & n21012 ;
  assign n25896 = n14402 & n25895 ;
  assign n25902 = n21465 & n22518 ;
  assign n25897 = ~n6020 & n22128 ;
  assign n25898 = ( n4833 & n6000 ) | ( n4833 & n25897 ) | ( n6000 & n25897 ) ;
  assign n25899 = ~n6307 & n25898 ;
  assign n25900 = n25899 ^ n4109 ^ 1'b0 ;
  assign n25901 = n5222 & n25900 ;
  assign n25903 = n25902 ^ n25901 ^ 1'b0 ;
  assign n25904 = n3907 ^ n2804 ^ 1'b0 ;
  assign n25905 = ~n5556 & n25904 ;
  assign n25906 = n1568 & ~n1862 ;
  assign n25907 = n21243 ^ n19310 ^ n12354 ;
  assign n25908 = ( n8670 & n16440 ) | ( n8670 & n25907 ) | ( n16440 & n25907 ) ;
  assign n25909 = n8164 ^ n4298 ^ n1646 ;
  assign n25910 = ( n8234 & n22061 ) | ( n8234 & n25909 ) | ( n22061 & n25909 ) ;
  assign n25911 = n25910 ^ n6874 ^ n1563 ;
  assign n25912 = n23831 ^ n7045 ^ n5089 ;
  assign n25913 = n25912 ^ n4647 ^ 1'b0 ;
  assign n25914 = n5927 | n25913 ;
  assign n25915 = ( n10212 & ~n25911 ) | ( n10212 & n25914 ) | ( ~n25911 & n25914 ) ;
  assign n25916 = n12385 ^ n526 ^ 1'b0 ;
  assign n25917 = ( ~n16715 & n18291 ) | ( ~n16715 & n25916 ) | ( n18291 & n25916 ) ;
  assign n25918 = n3790 ^ n851 ^ 1'b0 ;
  assign n25919 = n7236 & ~n25918 ;
  assign n25922 = n20871 ^ n13063 ^ n1981 ;
  assign n25920 = n24116 ^ n15993 ^ 1'b0 ;
  assign n25921 = n16716 & ~n25920 ;
  assign n25923 = n25922 ^ n25921 ^ 1'b0 ;
  assign n25925 = ( n1363 & n8892 ) | ( n1363 & n24731 ) | ( n8892 & n24731 ) ;
  assign n25924 = n11438 ^ n6541 ^ 1'b0 ;
  assign n25926 = n25925 ^ n25924 ^ n11818 ;
  assign n25927 = n498 & ~n7047 ;
  assign n25928 = ( n6525 & n12755 ) | ( n6525 & ~n25927 ) | ( n12755 & ~n25927 ) ;
  assign n25929 = n25928 ^ n24294 ^ n5071 ;
  assign n25930 = n25929 ^ n3045 ^ n2707 ;
  assign n25933 = n19797 ^ n6381 ^ n535 ;
  assign n25934 = n16038 | n25933 ;
  assign n25931 = ( n1453 & n2054 ) | ( n1453 & ~n11769 ) | ( n2054 & ~n11769 ) ;
  assign n25932 = ( n3864 & ~n24367 ) | ( n3864 & n25931 ) | ( ~n24367 & n25931 ) ;
  assign n25935 = n25934 ^ n25932 ^ n10719 ;
  assign n25936 = n25427 ^ n25000 ^ n17557 ;
  assign n25938 = ( n3770 & n11948 ) | ( n3770 & n16580 ) | ( n11948 & n16580 ) ;
  assign n25937 = n862 | n4461 ;
  assign n25939 = n25938 ^ n25937 ^ 1'b0 ;
  assign n25941 = n18314 ^ n14649 ^ n9925 ;
  assign n25940 = ~n426 & n6118 ;
  assign n25942 = n25941 ^ n25940 ^ 1'b0 ;
  assign n25943 = n11370 | n12351 ;
  assign n25944 = n9780 ^ n705 ^ 1'b0 ;
  assign n25945 = ~n12805 & n25944 ;
  assign n25946 = n9258 | n25945 ;
  assign n25947 = n10298 ^ n789 ^ 1'b0 ;
  assign n25948 = n4517 & ~n4862 ;
  assign n25949 = ~n11161 & n25948 ;
  assign n25950 = n14144 ^ n1254 ^ 1'b0 ;
  assign n25951 = ( ~n2593 & n19910 ) | ( ~n2593 & n25950 ) | ( n19910 & n25950 ) ;
  assign n25952 = ( x3 & ~n695 ) | ( x3 & n3611 ) | ( ~n695 & n3611 ) ;
  assign n25953 = n18065 ^ n1569 ^ 1'b0 ;
  assign n25954 = n5906 & n25953 ;
  assign n25955 = ~n4877 & n25954 ;
  assign n25956 = ( n18005 & n25952 ) | ( n18005 & ~n25955 ) | ( n25952 & ~n25955 ) ;
  assign n25957 = n20371 & n25956 ;
  assign n25958 = n8056 & n25957 ;
  assign n25959 = n25958 ^ n3747 ^ 1'b0 ;
  assign n25960 = ( n16502 & n21539 ) | ( n16502 & ~n25959 ) | ( n21539 & ~n25959 ) ;
  assign n25961 = ( n4607 & n7915 ) | ( n4607 & ~n20003 ) | ( n7915 & ~n20003 ) ;
  assign n25962 = ( n5226 & ~n16055 ) | ( n5226 & n25961 ) | ( ~n16055 & n25961 ) ;
  assign n25963 = n25962 ^ n18075 ^ n9262 ;
  assign n25973 = ( n773 & n11258 ) | ( n773 & ~n20327 ) | ( n11258 & ~n20327 ) ;
  assign n25971 = ~n1302 & n14584 ;
  assign n25972 = ~n17534 & n25971 ;
  assign n25974 = n25973 ^ n25972 ^ n3043 ;
  assign n25964 = n4021 & n8978 ;
  assign n25965 = n5877 ^ n4761 ^ n2515 ;
  assign n25966 = n4357 & n25965 ;
  assign n25967 = n15879 & n25966 ;
  assign n25968 = n25967 ^ n4191 ^ n217 ;
  assign n25969 = n25968 ^ n25573 ^ n8019 ;
  assign n25970 = ( n16041 & n25964 ) | ( n16041 & n25969 ) | ( n25964 & n25969 ) ;
  assign n25975 = n25974 ^ n25970 ^ n19202 ;
  assign n25976 = n12520 ^ n6187 ^ 1'b0 ;
  assign n25977 = n25976 ^ n8930 ^ n4710 ;
  assign n25978 = n22180 ^ n17720 ^ n8207 ;
  assign n25979 = ( n15993 & n25977 ) | ( n15993 & n25978 ) | ( n25977 & n25978 ) ;
  assign n25980 = n16784 ^ n14862 ^ n4798 ;
  assign n25981 = ( n8698 & n22131 ) | ( n8698 & ~n25980 ) | ( n22131 & ~n25980 ) ;
  assign n25982 = n3437 ^ n1883 ^ n1747 ;
  assign n25983 = n25982 ^ n1332 ^ 1'b0 ;
  assign n25984 = n6406 ^ n5419 ^ 1'b0 ;
  assign n25985 = n25984 ^ n2716 ^ 1'b0 ;
  assign n25986 = n25983 | n25985 ;
  assign n25987 = n8263 ^ n5915 ^ 1'b0 ;
  assign n25988 = n2970 | n24767 ;
  assign n25989 = n5155 | n25988 ;
  assign n25990 = n10078 ^ n7675 ^ n1359 ;
  assign n25991 = n25990 ^ n16485 ^ n11920 ;
  assign n25992 = ~n20820 & n25991 ;
  assign n25993 = n13264 & n16232 ;
  assign n25994 = n3825 | n10986 ;
  assign n25995 = ( ~n22715 & n25993 ) | ( ~n22715 & n25994 ) | ( n25993 & n25994 ) ;
  assign n25997 = n11199 ^ n8715 ^ n7547 ;
  assign n25996 = n2236 & n4035 ;
  assign n25998 = n25997 ^ n25996 ^ n23532 ;
  assign n25999 = ( n738 & n3657 ) | ( n738 & n8147 ) | ( n3657 & n8147 ) ;
  assign n26000 = n25999 ^ n14111 ^ 1'b0 ;
  assign n26001 = n19066 ^ n2592 ^ 1'b0 ;
  assign n26002 = n26000 | n26001 ;
  assign n26003 = n13338 ^ n1519 ^ n553 ;
  assign n26004 = n26003 ^ n7695 ^ 1'b0 ;
  assign n26005 = n22357 | n26004 ;
  assign n26006 = ~n1403 & n20578 ;
  assign n26007 = ( n19595 & ~n26005 ) | ( n19595 & n26006 ) | ( ~n26005 & n26006 ) ;
  assign n26008 = ( n1028 & n2090 ) | ( n1028 & n4880 ) | ( n2090 & n4880 ) ;
  assign n26009 = n10238 ^ n6198 ^ 1'b0 ;
  assign n26010 = n16732 & n26009 ;
  assign n26011 = ~n26008 & n26010 ;
  assign n26012 = ( x104 & n17327 ) | ( x104 & ~n26011 ) | ( n17327 & ~n26011 ) ;
  assign n26013 = n5108 ^ n3622 ^ 1'b0 ;
  assign n26014 = ( ~n3242 & n12618 ) | ( ~n3242 & n19647 ) | ( n12618 & n19647 ) ;
  assign n26015 = ( x9 & ~n14272 ) | ( x9 & n25701 ) | ( ~n14272 & n25701 ) ;
  assign n26016 = ~n3156 & n3986 ;
  assign n26017 = ( ~n10549 & n14869 ) | ( ~n10549 & n24576 ) | ( n14869 & n24576 ) ;
  assign n26018 = ( n6656 & n9895 ) | ( n6656 & ~n12768 ) | ( n9895 & ~n12768 ) ;
  assign n26019 = n26018 ^ n8463 ^ 1'b0 ;
  assign n26020 = ( ~n7015 & n18859 ) | ( ~n7015 & n20824 ) | ( n18859 & n20824 ) ;
  assign n26021 = ( n1462 & n11748 ) | ( n1462 & ~n12786 ) | ( n11748 & ~n12786 ) ;
  assign n26022 = n18581 ^ n12325 ^ n475 ;
  assign n26023 = ( n3784 & n4305 ) | ( n3784 & n26022 ) | ( n4305 & n26022 ) ;
  assign n26024 = n18516 ^ n6966 ^ n2978 ;
  assign n26025 = n26024 ^ n17727 ^ 1'b0 ;
  assign n26026 = n23649 ^ n7144 ^ 1'b0 ;
  assign n26031 = ( n1254 & n5439 ) | ( n1254 & ~n25652 ) | ( n5439 & ~n25652 ) ;
  assign n26028 = ( n9538 & n11351 ) | ( n9538 & ~n18591 ) | ( n11351 & ~n18591 ) ;
  assign n26029 = n2145 & n26028 ;
  assign n26030 = ~n25529 & n26029 ;
  assign n26032 = n26031 ^ n26030 ^ n4396 ;
  assign n26033 = n26032 ^ n16246 ^ 1'b0 ;
  assign n26027 = n4197 | n15557 ;
  assign n26034 = n26033 ^ n26027 ^ 1'b0 ;
  assign n26035 = x62 | n5177 ;
  assign n26036 = n13532 & ~n26035 ;
  assign n26037 = ( n7268 & ~n13061 ) | ( n7268 & n13355 ) | ( ~n13061 & n13355 ) ;
  assign n26038 = n9261 | n12682 ;
  assign n26039 = n26038 ^ n11657 ^ n1118 ;
  assign n26041 = ( n1559 & n8486 ) | ( n1559 & n8672 ) | ( n8486 & n8672 ) ;
  assign n26040 = ( ~n4495 & n9542 ) | ( ~n4495 & n15589 ) | ( n9542 & n15589 ) ;
  assign n26042 = n26041 ^ n26040 ^ n19818 ;
  assign n26043 = ~n4988 & n9917 ;
  assign n26044 = n18154 & ~n26043 ;
  assign n26048 = n14753 ^ n6494 ^ n3569 ;
  assign n26045 = ( n4872 & n6888 ) | ( n4872 & n13088 ) | ( n6888 & n13088 ) ;
  assign n26046 = ( n5470 & n15255 ) | ( n5470 & n26045 ) | ( n15255 & n26045 ) ;
  assign n26047 = n16476 & n26046 ;
  assign n26049 = n26048 ^ n26047 ^ 1'b0 ;
  assign n26050 = ( n1188 & ~n12476 ) | ( n1188 & n26049 ) | ( ~n12476 & n26049 ) ;
  assign n26051 = n14759 ^ n10111 ^ n8617 ;
  assign n26052 = n26051 ^ n5101 ^ n2294 ;
  assign n26053 = ( n26044 & ~n26050 ) | ( n26044 & n26052 ) | ( ~n26050 & n26052 ) ;
  assign n26054 = n13371 ^ n11392 ^ n7060 ;
  assign n26055 = n26054 ^ n18720 ^ n2852 ;
  assign n26056 = n11894 ^ n1973 ^ 1'b0 ;
  assign n26057 = n26056 ^ n15776 ^ n3079 ;
  assign n26058 = n15595 ^ n3188 ^ n947 ;
  assign n26059 = n26058 ^ n18457 ^ 1'b0 ;
  assign n26060 = n14360 & ~n16804 ;
  assign n26061 = n26060 ^ n24715 ^ 1'b0 ;
  assign n26062 = n3141 & ~n11996 ;
  assign n26063 = n24029 ^ n9409 ^ n6744 ;
  assign n26064 = n26063 ^ n2816 ^ 1'b0 ;
  assign n26065 = n14902 ^ n13404 ^ 1'b0 ;
  assign n26066 = n14555 & ~n18686 ;
  assign n26067 = n19990 ^ n12874 ^ n609 ;
  assign n26068 = n26067 ^ n24133 ^ n11568 ;
  assign n26069 = n19447 ^ n13002 ^ n10929 ;
  assign n26070 = n14077 ^ n13940 ^ 1'b0 ;
  assign n26071 = n26069 & ~n26070 ;
  assign n26072 = n9481 ^ n3619 ^ n331 ;
  assign n26073 = n4189 & ~n25419 ;
  assign n26074 = ~n4278 & n26073 ;
  assign n26075 = ( n10512 & n11079 ) | ( n10512 & ~n26074 ) | ( n11079 & ~n26074 ) ;
  assign n26076 = n26072 & ~n26075 ;
  assign n26077 = ~n17842 & n26076 ;
  assign n26078 = ( n3516 & n5822 ) | ( n3516 & ~n11160 ) | ( n5822 & ~n11160 ) ;
  assign n26079 = n20533 ^ n5870 ^ 1'b0 ;
  assign n26080 = n26078 & n26079 ;
  assign n26081 = n14307 ^ n6645 ^ 1'b0 ;
  assign n26082 = n3541 & n26081 ;
  assign n26083 = n14287 | n14402 ;
  assign n26084 = n14486 | n26083 ;
  assign n26085 = n2688 ^ n524 ^ 1'b0 ;
  assign n26086 = n26084 & n26085 ;
  assign n26087 = n26086 ^ n830 ^ 1'b0 ;
  assign n26088 = ( ~n17249 & n18536 ) | ( ~n17249 & n26087 ) | ( n18536 & n26087 ) ;
  assign n26089 = n22344 ^ n17135 ^ n15220 ;
  assign n26090 = n26089 ^ n23885 ^ n1932 ;
  assign n26091 = n23200 ^ n9744 ^ 1'b0 ;
  assign n26092 = n25226 ^ n15350 ^ n13773 ;
  assign n26093 = n26092 ^ n23638 ^ n13964 ;
  assign n26094 = n724 ^ n183 ^ 1'b0 ;
  assign n26095 = n13822 & n26094 ;
  assign n26096 = n26095 ^ n1925 ^ 1'b0 ;
  assign n26097 = n26096 ^ n7404 ^ n6087 ;
  assign n26098 = n10413 ^ n4441 ^ 1'b0 ;
  assign n26099 = n26098 ^ n21232 ^ 1'b0 ;
  assign n26100 = ~n12985 & n26099 ;
  assign n26101 = n25694 ^ n4788 ^ n1967 ;
  assign n26102 = n21688 & n22926 ;
  assign n26103 = n26101 & n26102 ;
  assign n26105 = n5197 ^ n3006 ^ 1'b0 ;
  assign n26106 = n1011 & ~n26105 ;
  assign n26104 = n8655 | n18771 ;
  assign n26107 = n26106 ^ n26104 ^ 1'b0 ;
  assign n26109 = ~n9405 & n10573 ;
  assign n26110 = ( ~n6697 & n17036 ) | ( ~n6697 & n26109 ) | ( n17036 & n26109 ) ;
  assign n26111 = n26110 ^ n11538 ^ n9819 ;
  assign n26108 = n18944 ^ n15028 ^ n12101 ;
  assign n26112 = n26111 ^ n26108 ^ n5232 ;
  assign n26113 = n17443 ^ n12753 ^ n5361 ;
  assign n26114 = n9208 & ~n9983 ;
  assign n26115 = n26114 ^ n8984 ^ 1'b0 ;
  assign n26116 = n13773 ^ n7157 ^ n6229 ;
  assign n26117 = n26116 ^ n13381 ^ n9779 ;
  assign n26118 = n26117 ^ n1461 ^ 1'b0 ;
  assign n26119 = n19340 ^ n18127 ^ n12792 ;
  assign n26120 = n21156 ^ n9521 ^ 1'b0 ;
  assign n26121 = n26120 ^ n16274 ^ n16166 ;
  assign n26122 = n15455 ^ n1829 ^ 1'b0 ;
  assign n26123 = n11775 & ~n26122 ;
  assign n26124 = ~n15934 & n20012 ;
  assign n26125 = n6181 & n26124 ;
  assign n26126 = ( n6654 & ~n8535 ) | ( n6654 & n10920 ) | ( ~n8535 & n10920 ) ;
  assign n26127 = ~n5987 & n14190 ;
  assign n26128 = n26127 ^ n14562 ^ 1'b0 ;
  assign n26129 = n8426 & ~n15387 ;
  assign n26130 = n26129 ^ n9821 ^ 1'b0 ;
  assign n26131 = ( n7299 & n16520 ) | ( n7299 & ~n26130 ) | ( n16520 & ~n26130 ) ;
  assign n26132 = n26131 ^ n19977 ^ n1294 ;
  assign n26133 = ( ~n12273 & n26128 ) | ( ~n12273 & n26132 ) | ( n26128 & n26132 ) ;
  assign n26134 = n14438 ^ n13172 ^ n10127 ;
  assign n26135 = n26134 ^ n8268 ^ 1'b0 ;
  assign n26138 = ( n4153 & ~n6202 ) | ( n4153 & n7359 ) | ( ~n6202 & n7359 ) ;
  assign n26136 = n22267 ^ n15423 ^ n488 ;
  assign n26137 = ( n7512 & ~n12802 ) | ( n7512 & n26136 ) | ( ~n12802 & n26136 ) ;
  assign n26139 = n26138 ^ n26137 ^ n12438 ;
  assign n26140 = n333 & n7316 ;
  assign n26141 = n3915 & n26140 ;
  assign n26142 = n26141 ^ n10904 ^ n10022 ;
  assign n26143 = ( n3716 & n25051 ) | ( n3716 & ~n26142 ) | ( n25051 & ~n26142 ) ;
  assign n26144 = n23670 ^ n9658 ^ n1428 ;
  assign n26149 = n12200 ^ n8263 ^ 1'b0 ;
  assign n26150 = n26149 ^ n20324 ^ n15948 ;
  assign n26148 = n19034 ^ n14448 ^ n11348 ;
  assign n26145 = n563 | n5547 ;
  assign n26146 = n26145 ^ n3385 ^ 1'b0 ;
  assign n26147 = ( n4174 & n18372 ) | ( n4174 & ~n26146 ) | ( n18372 & ~n26146 ) ;
  assign n26151 = n26150 ^ n26148 ^ n26147 ;
  assign n26152 = n8855 | n13606 ;
  assign n26153 = n5616 | n26152 ;
  assign n26154 = n10449 | n20865 ;
  assign n26155 = n26154 ^ n8903 ^ 1'b0 ;
  assign n26156 = n18345 | n20982 ;
  assign n26157 = n10903 & ~n26156 ;
  assign n26158 = n2433 | n17090 ;
  assign n26159 = n5086 | n26158 ;
  assign n26160 = n17542 ^ n5106 ^ n2087 ;
  assign n26161 = n8871 & ~n26160 ;
  assign n26162 = n2448 & n26161 ;
  assign n26163 = ( n7016 & n7056 ) | ( n7016 & n26162 ) | ( n7056 & n26162 ) ;
  assign n26164 = n18603 & ~n26163 ;
  assign n26165 = n26164 ^ n1300 ^ 1'b0 ;
  assign n26166 = n26165 ^ n17316 ^ n1078 ;
  assign n26167 = ( n5131 & n26159 ) | ( n5131 & ~n26166 ) | ( n26159 & ~n26166 ) ;
  assign n26168 = n20584 ^ n11966 ^ n716 ;
  assign n26169 = n26168 ^ n22802 ^ n14380 ;
  assign n26170 = n9167 ^ n3301 ^ 1'b0 ;
  assign n26171 = n10843 | n26170 ;
  assign n26172 = ( ~n6984 & n20112 ) | ( ~n6984 & n26171 ) | ( n20112 & n26171 ) ;
  assign n26173 = n14389 ^ n6978 ^ 1'b0 ;
  assign n26174 = n25924 & n26173 ;
  assign n26176 = ~n9323 & n12050 ;
  assign n26175 = n9292 & ~n16995 ;
  assign n26177 = n26176 ^ n26175 ^ 1'b0 ;
  assign n26178 = n5113 | n7582 ;
  assign n26179 = ( n1911 & ~n3078 ) | ( n1911 & n13889 ) | ( ~n3078 & n13889 ) ;
  assign n26180 = ( n5578 & ~n12319 ) | ( n5578 & n18755 ) | ( ~n12319 & n18755 ) ;
  assign n26181 = ( n12290 & ~n26179 ) | ( n12290 & n26180 ) | ( ~n26179 & n26180 ) ;
  assign n26182 = ( n10828 & ~n26178 ) | ( n10828 & n26181 ) | ( ~n26178 & n26181 ) ;
  assign n26183 = n11177 ^ n7304 ^ n7014 ;
  assign n26184 = ~n5876 & n24986 ;
  assign n26185 = ( n857 & n26183 ) | ( n857 & n26184 ) | ( n26183 & n26184 ) ;
  assign n26191 = n18713 ^ n1719 ^ 1'b0 ;
  assign n26192 = n2819 | n26191 ;
  assign n26193 = n3039 | n26192 ;
  assign n26189 = n1989 & n19424 ;
  assign n26190 = n10152 & n26189 ;
  assign n26186 = ~n3689 & n11026 ;
  assign n26187 = n26186 ^ n8923 ^ 1'b0 ;
  assign n26188 = ~n8682 & n26187 ;
  assign n26194 = n26193 ^ n26190 ^ n26188 ;
  assign n26195 = ( ~n6135 & n18881 ) | ( ~n6135 & n25236 ) | ( n18881 & n25236 ) ;
  assign n26196 = n9813 ^ n4771 ^ n1151 ;
  assign n26197 = n12544 & n26196 ;
  assign n26203 = ( ~n4989 & n6492 ) | ( ~n4989 & n15449 ) | ( n6492 & n15449 ) ;
  assign n26198 = ( n340 & ~n1543 ) | ( n340 & n22541 ) | ( ~n1543 & n22541 ) ;
  assign n26199 = n10311 & ~n26198 ;
  assign n26200 = n26199 ^ n1027 ^ 1'b0 ;
  assign n26201 = n26200 ^ n5108 ^ n573 ;
  assign n26202 = n9358 & n26201 ;
  assign n26204 = n26203 ^ n26202 ^ 1'b0 ;
  assign n26205 = n24849 ^ n4202 ^ 1'b0 ;
  assign n26206 = n2094 | n26205 ;
  assign n26207 = ( ~n1921 & n19156 ) | ( ~n1921 & n19501 ) | ( n19156 & n19501 ) ;
  assign n26208 = n26207 ^ n20322 ^ n15183 ;
  assign n26209 = n19109 & ~n26208 ;
  assign n26210 = n7591 & n26209 ;
  assign n26211 = n5095 ^ n2156 ^ 1'b0 ;
  assign n26212 = ( n14580 & ~n21427 ) | ( n14580 & n26211 ) | ( ~n21427 & n26211 ) ;
  assign n26213 = n26212 ^ n8072 ^ n4627 ;
  assign n26214 = ( n11433 & n20786 ) | ( n11433 & ~n21106 ) | ( n20786 & ~n21106 ) ;
  assign n26217 = n6535 ^ n3393 ^ 1'b0 ;
  assign n26218 = n25521 | n26217 ;
  assign n26215 = n1339 | n11184 ;
  assign n26216 = n26215 ^ n14571 ^ 1'b0 ;
  assign n26219 = n26218 ^ n26216 ^ n3603 ;
  assign n26220 = n20821 ^ n20305 ^ n18390 ;
  assign n26221 = ( n18735 & n26188 ) | ( n18735 & n26220 ) | ( n26188 & n26220 ) ;
  assign n26222 = n6118 ^ n3270 ^ n1207 ;
  assign n26223 = n1951 | n6662 ;
  assign n26224 = ( n1518 & n3582 ) | ( n1518 & ~n12159 ) | ( n3582 & ~n12159 ) ;
  assign n26225 = n26224 ^ n7892 ^ 1'b0 ;
  assign n26226 = ~n17354 & n26225 ;
  assign n26227 = ( n224 & n20867 ) | ( n224 & ~n26226 ) | ( n20867 & ~n26226 ) ;
  assign n26228 = n13414 ^ n11837 ^ n10294 ;
  assign n26229 = n26228 ^ n5774 ^ 1'b0 ;
  assign n26230 = n925 | n26229 ;
  assign n26231 = n9178 ^ n870 ^ 1'b0 ;
  assign n26232 = n8351 & ~n26231 ;
  assign n26233 = n18855 & n26232 ;
  assign n26234 = n10254 & n26233 ;
  assign n26235 = ( n1360 & ~n3194 ) | ( n1360 & n3977 ) | ( ~n3194 & n3977 ) ;
  assign n26236 = n9797 & n18744 ;
  assign n26237 = n26236 ^ n2286 ^ n1808 ;
  assign n26238 = ( n7580 & ~n9856 ) | ( n7580 & n18995 ) | ( ~n9856 & n18995 ) ;
  assign n26239 = ( n12615 & n16776 ) | ( n12615 & n26238 ) | ( n16776 & n26238 ) ;
  assign n26240 = n16099 ^ n15210 ^ n13825 ;
  assign n26241 = n26240 ^ n6268 ^ 1'b0 ;
  assign n26242 = n11722 ^ n9338 ^ n8806 ;
  assign n26243 = ( n3382 & n24328 ) | ( n3382 & ~n26242 ) | ( n24328 & ~n26242 ) ;
  assign n26244 = n11243 & n21766 ;
  assign n26245 = ( n12544 & n20843 ) | ( n12544 & ~n26244 ) | ( n20843 & ~n26244 ) ;
  assign n26246 = n2882 & n21118 ;
  assign n26247 = n17188 & n26246 ;
  assign n26248 = n16370 & ~n26247 ;
  assign n26249 = n409 | n26248 ;
  assign n26250 = n17895 ^ n16729 ^ n4103 ;
  assign n26251 = n26250 ^ n20650 ^ 1'b0 ;
  assign n26252 = n8442 & n26251 ;
  assign n26253 = n21712 & n26252 ;
  assign n26254 = n2846 ^ n1277 ^ 1'b0 ;
  assign n26255 = ~n201 & n23244 ;
  assign n26256 = n26255 ^ n5855 ^ 1'b0 ;
  assign n26257 = n9680 & ~n26256 ;
  assign n26258 = ( ~n20766 & n26254 ) | ( ~n20766 & n26257 ) | ( n26254 & n26257 ) ;
  assign n26259 = n23211 ^ n3353 ^ 1'b0 ;
  assign n26260 = ( n14405 & n14453 ) | ( n14405 & n14720 ) | ( n14453 & n14720 ) ;
  assign n26261 = ( ~n8065 & n16031 ) | ( ~n8065 & n26260 ) | ( n16031 & n26260 ) ;
  assign n26262 = n26261 ^ n10010 ^ n8982 ;
  assign n26263 = n16637 ^ n6086 ^ n4240 ;
  assign n26264 = n648 & ~n10383 ;
  assign n26265 = ~n13756 & n26264 ;
  assign n26266 = ( n1007 & n13894 ) | ( n1007 & n24204 ) | ( n13894 & n24204 ) ;
  assign n26267 = ( n6403 & n26265 ) | ( n6403 & ~n26266 ) | ( n26265 & ~n26266 ) ;
  assign n26268 = n14030 ^ n9776 ^ n3598 ;
  assign n26269 = n5116 ^ n4394 ^ 1'b0 ;
  assign n26270 = ~n6580 & n26269 ;
  assign n26274 = ( n5442 & n11555 ) | ( n5442 & ~n12353 ) | ( n11555 & ~n12353 ) ;
  assign n26271 = n16495 ^ n8827 ^ n6153 ;
  assign n26272 = n3928 & ~n26271 ;
  assign n26273 = n26272 ^ n7948 ^ 1'b0 ;
  assign n26275 = n26274 ^ n26273 ^ n22084 ;
  assign n26276 = n11907 ^ n3788 ^ 1'b0 ;
  assign n26277 = n26276 ^ n6957 ^ n681 ;
  assign n26278 = ~n3156 & n11505 ;
  assign n26279 = n2396 | n8223 ;
  assign n26280 = n4926 & ~n26279 ;
  assign n26281 = ( ~n21015 & n26278 ) | ( ~n21015 & n26280 ) | ( n26278 & n26280 ) ;
  assign n26282 = n3055 | n7909 ;
  assign n26283 = n26282 ^ n25039 ^ 1'b0 ;
  assign n26284 = n26283 ^ n17826 ^ n2724 ;
  assign n26285 = n5975 & n26284 ;
  assign n26286 = n24578 ^ n9895 ^ n8388 ;
  assign n26287 = n3912 | n16429 ;
  assign n26289 = n6358 & n10925 ;
  assign n26290 = n26289 ^ n5748 ^ n4058 ;
  assign n26288 = ~n2789 & n23810 ;
  assign n26291 = n26290 ^ n26288 ^ 1'b0 ;
  assign n26292 = n16744 ^ n10697 ^ n2999 ;
  assign n26293 = ~n12765 & n16867 ;
  assign n26294 = ~n26292 & n26293 ;
  assign n26295 = n941 | n5522 ;
  assign n26296 = n26295 ^ n8543 ^ 1'b0 ;
  assign n26297 = ( n880 & n2260 ) | ( n880 & ~n26296 ) | ( n2260 & ~n26296 ) ;
  assign n26298 = n26297 ^ n2023 ^ 1'b0 ;
  assign n26299 = n26298 ^ n19222 ^ n8827 ;
  assign n26300 = ( n6084 & n26294 ) | ( n6084 & ~n26299 ) | ( n26294 & ~n26299 ) ;
  assign n26301 = n17017 ^ n12795 ^ n4291 ;
  assign n26302 = n26301 ^ n19346 ^ 1'b0 ;
  assign n26305 = n10357 ^ n2176 ^ 1'b0 ;
  assign n26306 = ~n375 & n26305 ;
  assign n26307 = n26306 ^ n2507 ^ n1343 ;
  assign n26308 = n26307 ^ n25220 ^ 1'b0 ;
  assign n26303 = n9015 ^ n6956 ^ n345 ;
  assign n26304 = n26303 ^ n5112 ^ 1'b0 ;
  assign n26309 = n26308 ^ n26304 ^ n2733 ;
  assign n26310 = ( n4376 & ~n8060 ) | ( n4376 & n16726 ) | ( ~n8060 & n16726 ) ;
  assign n26312 = ~n624 & n7821 ;
  assign n26313 = n26312 ^ n7375 ^ n2169 ;
  assign n26311 = n16328 | n20468 ;
  assign n26314 = n26313 ^ n26311 ^ 1'b0 ;
  assign n26315 = n3746 ^ n3456 ^ 1'b0 ;
  assign n26316 = n921 & n26315 ;
  assign n26317 = n26316 ^ n312 ^ 1'b0 ;
  assign n26318 = n23171 ^ n14129 ^ 1'b0 ;
  assign n26319 = n4879 & ~n6215 ;
  assign n26320 = n22538 & n26319 ;
  assign n26323 = ~n8235 & n15421 ;
  assign n26321 = n18511 ^ n3848 ^ 1'b0 ;
  assign n26322 = n13297 & ~n26321 ;
  assign n26324 = n26323 ^ n26322 ^ n12575 ;
  assign n26325 = ( n8923 & n18362 ) | ( n8923 & n24796 ) | ( n18362 & n24796 ) ;
  assign n26328 = n22562 ^ n6525 ^ 1'b0 ;
  assign n26326 = ~n668 & n19983 ;
  assign n26327 = n25232 & n26326 ;
  assign n26329 = n26328 ^ n26327 ^ n26184 ;
  assign n26330 = n23161 ^ n13919 ^ n9128 ;
  assign n26331 = n12246 ^ n2107 ^ 1'b0 ;
  assign n26332 = n12781 | n26331 ;
  assign n26333 = ~n9352 & n25961 ;
  assign n26334 = n6779 ^ n5955 ^ 1'b0 ;
  assign n26335 = n8257 & n26334 ;
  assign n26336 = n2954 ^ n998 ^ 1'b0 ;
  assign n26337 = ~n13249 & n26336 ;
  assign n26338 = ~n26335 & n26337 ;
  assign n26339 = ( n4588 & ~n20328 ) | ( n4588 & n23912 ) | ( ~n20328 & n23912 ) ;
  assign n26340 = n10257 & ~n11915 ;
  assign n26341 = n26339 & n26340 ;
  assign n26342 = n10875 | n26341 ;
  assign n26343 = n14882 ^ n4374 ^ 1'b0 ;
  assign n26344 = ~n703 & n26343 ;
  assign n26345 = ~n16209 & n26344 ;
  assign n26346 = n26345 ^ n3427 ^ 1'b0 ;
  assign n26347 = n24525 ^ n22132 ^ 1'b0 ;
  assign n26348 = n5416 ^ n3096 ^ 1'b0 ;
  assign n26349 = n26348 ^ n20918 ^ n5504 ;
  assign n26350 = n26349 ^ n2733 ^ x100 ;
  assign n26351 = n13097 ^ n11965 ^ n8067 ;
  assign n26352 = ( n12447 & n15686 ) | ( n12447 & n26351 ) | ( n15686 & n26351 ) ;
  assign n26353 = n1755 | n12402 ;
  assign n26354 = n6161 | n26353 ;
  assign n26355 = n24070 ^ n8166 ^ 1'b0 ;
  assign n26356 = n11978 ^ n8868 ^ 1'b0 ;
  assign n26357 = n4073 & n10001 ;
  assign n26358 = n8953 ^ n6955 ^ n2625 ;
  assign n26359 = ~n1557 & n26358 ;
  assign n26360 = n26359 ^ n6145 ^ 1'b0 ;
  assign n26361 = n6014 & ~n6284 ;
  assign n26362 = ~n7367 & n26361 ;
  assign n26363 = n13545 ^ n2605 ^ 1'b0 ;
  assign n26364 = ~n11028 & n26363 ;
  assign n26369 = n10857 ^ n5329 ^ 1'b0 ;
  assign n26370 = ~n18080 & n26369 ;
  assign n26371 = n6548 | n26370 ;
  assign n26365 = ( n1517 & n9856 ) | ( n1517 & ~n16426 ) | ( n9856 & ~n16426 ) ;
  assign n26366 = n2660 | n12911 ;
  assign n26367 = n26365 | n26366 ;
  assign n26368 = n10491 & n26367 ;
  assign n26372 = n26371 ^ n26368 ^ 1'b0 ;
  assign n26373 = ( n26362 & n26364 ) | ( n26362 & ~n26372 ) | ( n26364 & ~n26372 ) ;
  assign n26374 = n26373 ^ n21854 ^ n12926 ;
  assign n26375 = ( n738 & ~n11646 ) | ( n738 & n18203 ) | ( ~n11646 & n18203 ) ;
  assign n26376 = n4092 & ~n10212 ;
  assign n26377 = n26376 ^ n13286 ^ 1'b0 ;
  assign n26378 = n26377 ^ n24609 ^ n15187 ;
  assign n26379 = n26378 ^ n8856 ^ n7700 ;
  assign n26383 = n457 & n8651 ;
  assign n26384 = ~n1867 & n26383 ;
  assign n26382 = ( n2860 & ~n9658 ) | ( n2860 & n18797 ) | ( ~n9658 & n18797 ) ;
  assign n26380 = ( n5817 & n12552 ) | ( n5817 & ~n23149 ) | ( n12552 & ~n23149 ) ;
  assign n26381 = n26380 ^ n763 ^ 1'b0 ;
  assign n26385 = n26384 ^ n26382 ^ n26381 ;
  assign n26386 = ( n11482 & n13104 ) | ( n11482 & ~n17535 ) | ( n13104 & ~n17535 ) ;
  assign n26387 = ~n16100 & n17319 ;
  assign n26388 = n26386 & n26387 ;
  assign n26389 = n2992 & ~n18301 ;
  assign n26390 = n3714 & n26389 ;
  assign n26391 = ( ~n1210 & n2495 ) | ( ~n1210 & n17770 ) | ( n2495 & n17770 ) ;
  assign n26392 = n2733 ^ n1931 ^ 1'b0 ;
  assign n26393 = n26392 ^ n22902 ^ n4259 ;
  assign n26394 = n10148 ^ n3037 ^ 1'b0 ;
  assign n26395 = ~n18711 & n26394 ;
  assign n26396 = n26395 ^ n10162 ^ 1'b0 ;
  assign n26397 = n2667 & ~n7689 ;
  assign n26398 = n26397 ^ n3056 ^ 1'b0 ;
  assign n26399 = n26398 ^ n2805 ^ n1515 ;
  assign n26400 = ( n9902 & n15278 ) | ( n9902 & ~n23769 ) | ( n15278 & ~n23769 ) ;
  assign n26401 = ( n20571 & n23440 ) | ( n20571 & ~n23660 ) | ( n23440 & ~n23660 ) ;
  assign n26402 = n22052 ^ n7783 ^ 1'b0 ;
  assign n26403 = n16270 & n26402 ;
  assign n26404 = n26403 ^ n15772 ^ n2429 ;
  assign n26405 = n26404 ^ n16560 ^ n1566 ;
  assign n26406 = n2053 & n8989 ;
  assign n26407 = ~n4502 & n26406 ;
  assign n26408 = x41 & ~n7400 ;
  assign n26409 = n6740 | n26408 ;
  assign n26410 = n4610 ^ n3897 ^ n3073 ;
  assign n26412 = n11763 ^ n6572 ^ 1'b0 ;
  assign n26411 = ( n8343 & ~n19342 ) | ( n8343 & n22295 ) | ( ~n19342 & n22295 ) ;
  assign n26413 = n26412 ^ n26411 ^ n19704 ;
  assign n26414 = ( n21276 & ~n26410 ) | ( n21276 & n26413 ) | ( ~n26410 & n26413 ) ;
  assign n26415 = ( n2366 & n5987 ) | ( n2366 & n17934 ) | ( n5987 & n17934 ) ;
  assign n26416 = n18597 ^ n17526 ^ 1'b0 ;
  assign n26417 = ~n5178 & n7089 ;
  assign n26418 = n3805 & n26417 ;
  assign n26419 = ( x29 & ~n1987 ) | ( x29 & n26418 ) | ( ~n1987 & n26418 ) ;
  assign n26420 = n15843 & n26419 ;
  assign n26421 = n4994 ^ n4280 ^ 1'b0 ;
  assign n26422 = n9886 & ~n26421 ;
  assign n26423 = ~n22859 & n26422 ;
  assign n26424 = n17086 & ~n26423 ;
  assign n26425 = ~n25857 & n26424 ;
  assign n26426 = n8340 ^ n8277 ^ n4396 ;
  assign n26427 = ~n12427 & n23365 ;
  assign n26428 = ~n3159 & n26427 ;
  assign n26429 = ~n26426 & n26428 ;
  assign n26430 = n8897 & n11142 ;
  assign n26431 = n26430 ^ n23006 ^ 1'b0 ;
  assign n26432 = ( n3659 & ~n10581 ) | ( n3659 & n16600 ) | ( ~n10581 & n16600 ) ;
  assign n26433 = n6187 ^ n602 ^ 1'b0 ;
  assign n26434 = n8548 ^ n3729 ^ 1'b0 ;
  assign n26435 = ( ~n2547 & n26433 ) | ( ~n2547 & n26434 ) | ( n26433 & n26434 ) ;
  assign n26436 = ( n838 & n6130 ) | ( n838 & n10639 ) | ( n6130 & n10639 ) ;
  assign n26437 = n26436 ^ n1868 ^ n1714 ;
  assign n26438 = ~n1750 & n18802 ;
  assign n26439 = n26438 ^ n25607 ^ 1'b0 ;
  assign n26440 = ~n13494 & n25084 ;
  assign n26441 = n5327 & n10164 ;
  assign n26442 = n26441 ^ n524 ^ 1'b0 ;
  assign n26444 = n6014 & ~n22632 ;
  assign n26445 = n5656 & n26444 ;
  assign n26446 = ( ~n7154 & n9803 ) | ( ~n7154 & n26445 ) | ( n9803 & n26445 ) ;
  assign n26443 = n17185 ^ n8950 ^ n5421 ;
  assign n26447 = n26446 ^ n26443 ^ n2336 ;
  assign n26448 = n26447 ^ n17267 ^ 1'b0 ;
  assign n26449 = ( n12755 & n13119 ) | ( n12755 & ~n20578 ) | ( n13119 & ~n20578 ) ;
  assign n26450 = n19875 ^ n3428 ^ n3193 ;
  assign n26451 = n26450 ^ n2760 ^ n1565 ;
  assign n26452 = n17511 & ~n22760 ;
  assign n26453 = n26452 ^ n1251 ^ 1'b0 ;
  assign n26454 = ( n1397 & n9943 ) | ( n1397 & ~n26453 ) | ( n9943 & ~n26453 ) ;
  assign n26455 = ( n22695 & n23294 ) | ( n22695 & ~n26454 ) | ( n23294 & ~n26454 ) ;
  assign n26456 = n16801 ^ n13327 ^ n12320 ;
  assign n26457 = n26456 ^ n12467 ^ 1'b0 ;
  assign n26458 = n10465 ^ n5202 ^ n1336 ;
  assign n26459 = ( n8927 & n11089 ) | ( n8927 & n26458 ) | ( n11089 & n26458 ) ;
  assign n26460 = ( ~n3885 & n18256 ) | ( ~n3885 & n20501 ) | ( n18256 & n20501 ) ;
  assign n26461 = n26460 ^ n22596 ^ n5639 ;
  assign n26462 = n23203 ^ n7582 ^ n3941 ;
  assign n26463 = n19316 ^ n13147 ^ n6058 ;
  assign n26464 = n26463 ^ n4360 ^ 1'b0 ;
  assign n26465 = ~n26462 & n26464 ;
  assign n26466 = n4041 ^ n2112 ^ 1'b0 ;
  assign n26467 = n3563 & ~n26466 ;
  assign n26468 = n26467 ^ n13337 ^ 1'b0 ;
  assign n26471 = n1040 | n1722 ;
  assign n26472 = n11760 & ~n26471 ;
  assign n26469 = ( n4255 & n14237 ) | ( n4255 & ~n19375 ) | ( n14237 & ~n19375 ) ;
  assign n26470 = ( n4490 & ~n22937 ) | ( n4490 & n26469 ) | ( ~n22937 & n26469 ) ;
  assign n26473 = n26472 ^ n26470 ^ n1721 ;
  assign n26474 = n26473 ^ n16881 ^ n2296 ;
  assign n26475 = n12387 ^ n2047 ^ 1'b0 ;
  assign n26476 = n9833 | n26475 ;
  assign n26477 = n3769 & ~n26476 ;
  assign n26478 = n26474 & n26477 ;
  assign n26479 = ( n2136 & n18516 ) | ( n2136 & n20361 ) | ( n18516 & n20361 ) ;
  assign n26480 = ( n3238 & n12756 ) | ( n3238 & n19459 ) | ( n12756 & n19459 ) ;
  assign n26481 = n12163 ^ n5808 ^ 1'b0 ;
  assign n26484 = ( n4278 & ~n12895 ) | ( n4278 & n14232 ) | ( ~n12895 & n14232 ) ;
  assign n26482 = n8315 ^ n4101 ^ n403 ;
  assign n26483 = ( n10557 & ~n16062 ) | ( n10557 & n26482 ) | ( ~n16062 & n26482 ) ;
  assign n26485 = n26484 ^ n26483 ^ n15110 ;
  assign n26486 = n2884 & n20545 ;
  assign n26487 = n21302 ^ n12626 ^ n2392 ;
  assign n26488 = n8208 ^ n962 ^ 1'b0 ;
  assign n26489 = n26488 ^ n22768 ^ 1'b0 ;
  assign n26490 = ~n405 & n6664 ;
  assign n26491 = n25872 & n26490 ;
  assign n26492 = n22894 ^ n8082 ^ 1'b0 ;
  assign n26493 = ~n26491 & n26492 ;
  assign n26494 = ( n3286 & n5808 ) | ( n3286 & ~n10594 ) | ( n5808 & ~n10594 ) ;
  assign n26495 = n12159 & ~n26494 ;
  assign n26496 = n9588 ^ n2128 ^ n846 ;
  assign n26497 = n3205 | n6231 ;
  assign n26498 = n12429 & ~n26497 ;
  assign n26499 = n16253 ^ n1031 ^ 1'b0 ;
  assign n26500 = ( n6386 & n26498 ) | ( n6386 & n26499 ) | ( n26498 & n26499 ) ;
  assign n26501 = ( n11837 & n22135 ) | ( n11837 & ~n24223 ) | ( n22135 & ~n24223 ) ;
  assign n26502 = n19036 ^ n16676 ^ n4738 ;
  assign n26503 = ( n3055 & n20509 ) | ( n3055 & n26502 ) | ( n20509 & n26502 ) ;
  assign n26504 = ( n3919 & n5843 ) | ( n3919 & n7384 ) | ( n5843 & n7384 ) ;
  assign n26505 = n26504 ^ n20821 ^ 1'b0 ;
  assign n26506 = n4205 | n12164 ;
  assign n26507 = n16277 & ~n26506 ;
  assign n26508 = n26507 ^ n11586 ^ n1465 ;
  assign n26509 = n14156 ^ n3160 ^ 1'b0 ;
  assign n26510 = n10892 ^ n6781 ^ n2523 ;
  assign n26511 = ~n3063 & n26510 ;
  assign n26512 = n26509 & n26511 ;
  assign n26513 = n7424 | n13473 ;
  assign n26514 = n26513 ^ n5784 ^ 1'b0 ;
  assign n26515 = ( n3415 & n6511 ) | ( n3415 & ~n21299 ) | ( n6511 & ~n21299 ) ;
  assign n26516 = ( n13954 & n25349 ) | ( n13954 & n26515 ) | ( n25349 & n26515 ) ;
  assign n26517 = ( ~n365 & n12961 ) | ( ~n365 & n26516 ) | ( n12961 & n26516 ) ;
  assign n26518 = ( ~n5689 & n8425 ) | ( ~n5689 & n8853 ) | ( n8425 & n8853 ) ;
  assign n26519 = n18581 & n26518 ;
  assign n26520 = ( ~n1114 & n4954 ) | ( ~n1114 & n10595 ) | ( n4954 & n10595 ) ;
  assign n26521 = n22926 & ~n26520 ;
  assign n26522 = n9065 ^ n670 ^ 1'b0 ;
  assign n26523 = n10058 | n26522 ;
  assign n26524 = n2029 | n16022 ;
  assign n26525 = n26524 ^ n13736 ^ 1'b0 ;
  assign n26526 = n6785 | n25401 ;
  assign n26527 = n26526 ^ n10664 ^ 1'b0 ;
  assign n26528 = n1189 & ~n5065 ;
  assign n26529 = ( n3871 & n7175 ) | ( n3871 & ~n11736 ) | ( n7175 & ~n11736 ) ;
  assign n26530 = n26529 ^ n10640 ^ n5801 ;
  assign n26531 = n26530 ^ n19414 ^ n13337 ;
  assign n26532 = n6369 & n12869 ;
  assign n26533 = ~n9506 & n26532 ;
  assign n26534 = n26533 ^ n17725 ^ n2680 ;
  assign n26535 = ( ~n5155 & n8652 ) | ( ~n5155 & n26534 ) | ( n8652 & n26534 ) ;
  assign n26536 = ( n17249 & ~n20664 ) | ( n17249 & n21620 ) | ( ~n20664 & n21620 ) ;
  assign n26537 = ( n1241 & n3065 ) | ( n1241 & n22312 ) | ( n3065 & n22312 ) ;
  assign n26538 = n26537 ^ n10261 ^ 1'b0 ;
  assign n26539 = n20162 ^ n8146 ^ n926 ;
  assign n26540 = n25877 ^ n11780 ^ 1'b0 ;
  assign n26541 = n13623 & ~n26540 ;
  assign n26542 = n17727 & ~n24298 ;
  assign n26543 = n3825 & n26542 ;
  assign n26544 = n13444 | n26543 ;
  assign n26545 = n26544 ^ n1363 ^ 1'b0 ;
  assign n26546 = n25954 ^ n905 ^ 1'b0 ;
  assign n26549 = n1927 | n15701 ;
  assign n26550 = n14605 & ~n26549 ;
  assign n26547 = n11942 | n15162 ;
  assign n26548 = n9032 & ~n26547 ;
  assign n26551 = n26550 ^ n26548 ^ n4236 ;
  assign n26552 = n22474 ^ n12646 ^ n4867 ;
  assign n26553 = ( n1645 & ~n1696 ) | ( n1645 & n4148 ) | ( ~n1696 & n4148 ) ;
  assign n26554 = ~n24751 & n26553 ;
  assign n26555 = ~n25244 & n26554 ;
  assign n26556 = ( n2665 & ~n22082 ) | ( n2665 & n26555 ) | ( ~n22082 & n26555 ) ;
  assign n26557 = n6653 ^ n5308 ^ n4156 ;
  assign n26558 = n2946 | n26557 ;
  assign n26559 = n275 | n8058 ;
  assign n26560 = n26559 ^ n15633 ^ n12560 ;
  assign n26561 = ( ~n3392 & n4314 ) | ( ~n3392 & n14128 ) | ( n4314 & n14128 ) ;
  assign n26562 = ( n7272 & n26560 ) | ( n7272 & n26561 ) | ( n26560 & n26561 ) ;
  assign n26563 = n26562 ^ n4660 ^ 1'b0 ;
  assign n26564 = n3322 | n26563 ;
  assign n26565 = n3022 & ~n23360 ;
  assign n26566 = ~n6602 & n9687 ;
  assign n26567 = n26566 ^ x35 ^ 1'b0 ;
  assign n26568 = n7144 | n26567 ;
  assign n26569 = n26568 ^ n261 ^ 1'b0 ;
  assign n26570 = ( ~n6975 & n12983 ) | ( ~n6975 & n18618 ) | ( n12983 & n18618 ) ;
  assign n26571 = x121 | n12570 ;
  assign n26572 = n19881 ^ n17946 ^ n277 ;
  assign n26573 = ( n3939 & n13452 ) | ( n3939 & ~n16918 ) | ( n13452 & ~n16918 ) ;
  assign n26577 = ( ~n3680 & n7511 ) | ( ~n3680 & n20104 ) | ( n7511 & n20104 ) ;
  assign n26574 = n24334 ^ n6382 ^ n5899 ;
  assign n26575 = n26574 ^ n23007 ^ 1'b0 ;
  assign n26576 = n23205 & ~n26575 ;
  assign n26578 = n26577 ^ n26576 ^ n584 ;
  assign n26579 = ~n8630 & n25473 ;
  assign n26580 = n22634 ^ n9682 ^ 1'b0 ;
  assign n26581 = n4699 | n26580 ;
  assign n26582 = n26581 ^ n18664 ^ n8739 ;
  assign n26583 = ( ~n1594 & n13660 ) | ( ~n1594 & n20430 ) | ( n13660 & n20430 ) ;
  assign n26584 = n26583 ^ n4349 ^ 1'b0 ;
  assign n26585 = n26584 ^ n26315 ^ n25459 ;
  assign n26586 = ( n12354 & n18785 ) | ( n12354 & ~n25815 ) | ( n18785 & ~n25815 ) ;
  assign n26587 = ( n7161 & ~n7220 ) | ( n7161 & n9532 ) | ( ~n7220 & n9532 ) ;
  assign n26588 = n26587 ^ n19720 ^ n8235 ;
  assign n26589 = ( ~x78 & n2851 ) | ( ~x78 & n9547 ) | ( n2851 & n9547 ) ;
  assign n26590 = n26589 ^ n4352 ^ 1'b0 ;
  assign n26591 = n26590 ^ n20383 ^ 1'b0 ;
  assign n26592 = n894 & ~n2345 ;
  assign n26593 = n26592 ^ n6346 ^ 1'b0 ;
  assign n26594 = n26593 ^ n17509 ^ n7923 ;
  assign n26597 = ~n4750 & n5797 ;
  assign n26598 = n26597 ^ n12643 ^ 1'b0 ;
  assign n26595 = ~n4721 & n10886 ;
  assign n26596 = n26595 ^ n18065 ^ 1'b0 ;
  assign n26599 = n26598 ^ n26596 ^ n14734 ;
  assign n26600 = n26599 ^ n22861 ^ n15877 ;
  assign n26601 = ( n5081 & n6734 ) | ( n5081 & n8583 ) | ( n6734 & n8583 ) ;
  assign n26602 = n11058 ^ n7239 ^ n4598 ;
  assign n26603 = ( ~n7945 & n26601 ) | ( ~n7945 & n26602 ) | ( n26601 & n26602 ) ;
  assign n26604 = n26603 ^ n18956 ^ 1'b0 ;
  assign n26605 = n15583 ^ n4664 ^ 1'b0 ;
  assign n26606 = n10244 & n26605 ;
  assign n26607 = n26606 ^ n4306 ^ n1309 ;
  assign n26608 = ( n21881 & n22491 ) | ( n21881 & n26607 ) | ( n22491 & n26607 ) ;
  assign n26609 = n26608 ^ n12096 ^ 1'b0 ;
  assign n26610 = n22623 ^ n16650 ^ 1'b0 ;
  assign n26611 = n13782 ^ n10403 ^ 1'b0 ;
  assign n26612 = n26610 & ~n26611 ;
  assign n26613 = n12985 | n25418 ;
  assign n26614 = n26613 ^ n3390 ^ 1'b0 ;
  assign n26615 = n13693 ^ n905 ^ 1'b0 ;
  assign n26616 = n17565 & ~n26615 ;
  assign n26617 = n5406 & n6056 ;
  assign n26618 = n26617 ^ n861 ^ 1'b0 ;
  assign n26619 = ( n440 & n11889 ) | ( n440 & ~n26618 ) | ( n11889 & ~n26618 ) ;
  assign n26620 = n18204 | n24980 ;
  assign n26621 = ~n1474 & n4268 ;
  assign n26622 = n26620 & n26621 ;
  assign n26623 = ( n11894 & ~n22919 ) | ( n11894 & n26622 ) | ( ~n22919 & n26622 ) ;
  assign n26624 = ( ~n6731 & n7758 ) | ( ~n6731 & n12457 ) | ( n7758 & n12457 ) ;
  assign n26626 = ( ~n3364 & n5373 ) | ( ~n3364 & n15133 ) | ( n5373 & n15133 ) ;
  assign n26625 = n1480 & n21312 ;
  assign n26627 = n26626 ^ n26625 ^ 1'b0 ;
  assign n26628 = ( n240 & n6649 ) | ( n240 & ~n10242 ) | ( n6649 & ~n10242 ) ;
  assign n26629 = ( n7626 & n26627 ) | ( n7626 & ~n26628 ) | ( n26627 & ~n26628 ) ;
  assign n26630 = n10339 ^ n5054 ^ n4380 ;
  assign n26631 = ( ~n22132 & n22467 ) | ( ~n22132 & n26630 ) | ( n22467 & n26630 ) ;
  assign n26632 = n6543 ^ n733 ^ 1'b0 ;
  assign n26633 = n545 & ~n26632 ;
  assign n26634 = n20878 ^ n9246 ^ n6465 ;
  assign n26635 = n26634 ^ n16627 ^ 1'b0 ;
  assign n26636 = n16874 | n26635 ;
  assign n26637 = n25471 ^ n22640 ^ n5527 ;
  assign n26638 = n26242 ^ n16635 ^ n8276 ;
  assign n26639 = n13335 ^ n4815 ^ n1861 ;
  assign n26640 = n26639 ^ n9424 ^ 1'b0 ;
  assign n26641 = n6549 & ~n26640 ;
  assign n26642 = ( n17526 & n26638 ) | ( n17526 & n26641 ) | ( n26638 & n26641 ) ;
  assign n26643 = n25922 ^ n17245 ^ 1'b0 ;
  assign n26644 = n18273 ^ n12068 ^ n6685 ;
  assign n26645 = n25944 ^ n14485 ^ 1'b0 ;
  assign n26649 = n2528 ^ x50 ^ 1'b0 ;
  assign n26650 = n1703 | n26649 ;
  assign n26651 = n26650 ^ n19072 ^ n4675 ;
  assign n26646 = n11666 & ~n12544 ;
  assign n26647 = n26646 ^ n4792 ^ 1'b0 ;
  assign n26648 = ~n8548 & n26647 ;
  assign n26652 = n26651 ^ n26648 ^ 1'b0 ;
  assign n26653 = n1055 ^ n372 ^ 1'b0 ;
  assign n26654 = n5077 | n26653 ;
  assign n26655 = ( n12802 & ~n23839 ) | ( n12802 & n26654 ) | ( ~n23839 & n26654 ) ;
  assign n26656 = n24634 ^ n22626 ^ 1'b0 ;
  assign n26657 = ~n371 & n23222 ;
  assign n26659 = ( ~n1523 & n8152 ) | ( ~n1523 & n11862 ) | ( n8152 & n11862 ) ;
  assign n26658 = n13462 ^ n5537 ^ n3619 ;
  assign n26660 = n26659 ^ n26658 ^ n11742 ;
  assign n26661 = n14424 ^ n2801 ^ n236 ;
  assign n26662 = ~n15937 & n26661 ;
  assign n26663 = n26662 ^ n10665 ^ 1'b0 ;
  assign n26664 = n26663 ^ n5365 ^ 1'b0 ;
  assign n26665 = n21669 & ~n26664 ;
  assign n26666 = n24540 ^ n15484 ^ n12400 ;
  assign n26667 = n11885 ^ n908 ^ 1'b0 ;
  assign n26668 = n26666 & n26667 ;
  assign n26669 = ~n11470 & n26668 ;
  assign n26670 = n26669 ^ n9010 ^ 1'b0 ;
  assign n26671 = ( n13705 & n21918 ) | ( n13705 & ~n22040 ) | ( n21918 & ~n22040 ) ;
  assign n26673 = n17904 ^ n15963 ^ n2077 ;
  assign n26672 = ( ~n15721 & n18144 ) | ( ~n15721 & n21147 ) | ( n18144 & n21147 ) ;
  assign n26674 = n26673 ^ n26672 ^ n22190 ;
  assign n26675 = n12392 ^ n8221 ^ n6548 ;
  assign n26676 = n11578 ^ n7243 ^ n3880 ;
  assign n26677 = ( n23357 & n26675 ) | ( n23357 & ~n26676 ) | ( n26675 & ~n26676 ) ;
  assign n26678 = ( ~n8277 & n10611 ) | ( ~n8277 & n18892 ) | ( n10611 & n18892 ) ;
  assign n26679 = n20811 ^ n3381 ^ n1480 ;
  assign n26680 = n3853 ^ n2459 ^ 1'b0 ;
  assign n26681 = n26680 ^ n20209 ^ 1'b0 ;
  assign n26682 = ~n26679 & n26681 ;
  assign n26683 = n2705 & n26682 ;
  assign n26684 = ( n3718 & ~n26678 ) | ( n3718 & n26683 ) | ( ~n26678 & n26683 ) ;
  assign n26685 = n22635 ^ n16205 ^ n11699 ;
  assign n26686 = ( ~n19897 & n21935 ) | ( ~n19897 & n22230 ) | ( n21935 & n22230 ) ;
  assign n26687 = ~n2070 & n25761 ;
  assign n26688 = n26687 ^ n1019 ^ 1'b0 ;
  assign n26689 = ~n16817 & n26688 ;
  assign n26690 = n4421 ^ n3935 ^ 1'b0 ;
  assign n26691 = ( n3192 & ~n21567 ) | ( n3192 & n26690 ) | ( ~n21567 & n26690 ) ;
  assign n26692 = n15924 | n26691 ;
  assign n26693 = n26692 ^ n13770 ^ 1'b0 ;
  assign n26694 = n17213 ^ n4581 ^ 1'b0 ;
  assign n26695 = n7115 | n26694 ;
  assign n26696 = n14220 & ~n26695 ;
  assign n26697 = n6452 & n26696 ;
  assign n26698 = ( n5670 & ~n8704 ) | ( n5670 & n26697 ) | ( ~n8704 & n26697 ) ;
  assign n26700 = n11091 ^ n10518 ^ n4421 ;
  assign n26699 = n24795 ^ n5317 ^ n4520 ;
  assign n26701 = n26700 ^ n26699 ^ n10639 ;
  assign n26702 = ~n2928 & n4398 ;
  assign n26703 = n26702 ^ n23336 ^ 1'b0 ;
  assign n26704 = n26703 ^ n12529 ^ 1'b0 ;
  assign n26705 = n26704 ^ x61 ^ 1'b0 ;
  assign n26706 = ( n8309 & n9542 ) | ( n8309 & n11341 ) | ( n9542 & n11341 ) ;
  assign n26707 = ( ~n7780 & n9148 ) | ( ~n7780 & n13843 ) | ( n9148 & n13843 ) ;
  assign n26712 = n16389 ^ n861 ^ 1'b0 ;
  assign n26711 = n23088 ^ n16127 ^ n3211 ;
  assign n26708 = ~n8565 & n9121 ;
  assign n26709 = n20172 & n26708 ;
  assign n26710 = n26709 ^ n24540 ^ n20493 ;
  assign n26713 = n26712 ^ n26711 ^ n26710 ;
  assign n26714 = n3898 | n5714 ;
  assign n26715 = n3190 & ~n26714 ;
  assign n26716 = n26715 ^ n24560 ^ n7545 ;
  assign n26717 = n26716 ^ n8121 ^ n3641 ;
  assign n26718 = ~n1334 & n12762 ;
  assign n26719 = ~n7202 & n26718 ;
  assign n26720 = ~n1871 & n16332 ;
  assign n26721 = n23555 & n26720 ;
  assign n26722 = n11376 ^ n5372 ^ 1'b0 ;
  assign n26723 = n4179 & ~n4997 ;
  assign n26724 = n26723 ^ n3478 ^ 1'b0 ;
  assign n26725 = n10581 ^ n3425 ^ n2884 ;
  assign n26726 = n6073 | n26725 ;
  assign n26727 = n26726 ^ n1573 ^ 1'b0 ;
  assign n26728 = ( n15288 & n24633 ) | ( n15288 & n26727 ) | ( n24633 & n26727 ) ;
  assign n26731 = n20730 ^ n12143 ^ n1490 ;
  assign n26729 = n6605 ^ n883 ^ 1'b0 ;
  assign n26730 = n20484 & ~n26729 ;
  assign n26732 = n26731 ^ n26730 ^ n194 ;
  assign n26733 = ( ~n5778 & n24247 ) | ( ~n5778 & n24302 ) | ( n24247 & n24302 ) ;
  assign n26734 = n26733 ^ n8765 ^ 1'b0 ;
  assign n26735 = n22896 ^ n22812 ^ n20381 ;
  assign n26736 = n26734 | n26735 ;
  assign n26737 = ( n818 & n4412 ) | ( n818 & n14720 ) | ( n4412 & n14720 ) ;
  assign n26738 = n9671 ^ n4001 ^ n1399 ;
  assign n26739 = ( n6034 & n17208 ) | ( n6034 & ~n26738 ) | ( n17208 & ~n26738 ) ;
  assign n26740 = n26739 ^ n25679 ^ n2801 ;
  assign n26741 = n23878 ^ n16573 ^ n13589 ;
  assign n26742 = n6252 | n26741 ;
  assign n26743 = n26740 | n26742 ;
  assign n26745 = n14225 ^ n9628 ^ n1810 ;
  assign n26744 = n6221 & ~n9347 ;
  assign n26746 = n26745 ^ n26744 ^ 1'b0 ;
  assign n26747 = n24663 ^ n19576 ^ n12024 ;
  assign n26748 = n16293 & n20613 ;
  assign n26749 = n4744 & n8429 ;
  assign n26750 = n15376 & n26749 ;
  assign n26751 = ( n15300 & n19793 ) | ( n15300 & ~n26750 ) | ( n19793 & ~n26750 ) ;
  assign n26752 = ( ~n8830 & n15159 ) | ( ~n8830 & n23570 ) | ( n15159 & n23570 ) ;
  assign n26753 = n23653 ^ n5405 ^ 1'b0 ;
  assign n26754 = n6631 ^ n829 ^ 1'b0 ;
  assign n26755 = n26754 ^ n15974 ^ n9177 ;
  assign n26756 = ~n542 & n4483 ;
  assign n26757 = n14120 ^ n13415 ^ 1'b0 ;
  assign n26758 = n26756 & ~n26757 ;
  assign n26759 = n17686 ^ n8136 ^ 1'b0 ;
  assign n26762 = ( n1758 & ~n6899 ) | ( n1758 & n20361 ) | ( ~n6899 & n20361 ) ;
  assign n26760 = n767 & n5180 ;
  assign n26761 = ~n23443 & n26760 ;
  assign n26763 = n26762 ^ n26761 ^ n12539 ;
  assign n26764 = n21267 ^ n10861 ^ 1'b0 ;
  assign n26765 = n23555 | n26764 ;
  assign n26766 = ( n5497 & n19139 ) | ( n5497 & n19896 ) | ( n19139 & n19896 ) ;
  assign n26767 = ( n14368 & n25303 ) | ( n14368 & ~n25378 ) | ( n25303 & ~n25378 ) ;
  assign n26768 = n22720 ^ n8015 ^ n1361 ;
  assign n26769 = ~n22380 & n26768 ;
  assign n26770 = n15248 & n26769 ;
  assign n26771 = n14376 ^ n7298 ^ 1'b0 ;
  assign n26772 = n12323 & n26771 ;
  assign n26773 = ( n4228 & n10069 ) | ( n4228 & ~n23767 ) | ( n10069 & ~n23767 ) ;
  assign n26774 = n13766 ^ n11086 ^ 1'b0 ;
  assign n26775 = ~n4647 & n26774 ;
  assign n26776 = n15623 | n26775 ;
  assign n26777 = n6083 & ~n6874 ;
  assign n26778 = n26777 ^ n5367 ^ 1'b0 ;
  assign n26779 = ~n4750 & n26778 ;
  assign n26780 = ~n13456 & n26779 ;
  assign n26781 = ( n1617 & n26553 ) | ( n1617 & ~n26780 ) | ( n26553 & ~n26780 ) ;
  assign n26782 = n19179 ^ n4079 ^ 1'b0 ;
  assign n26783 = n20293 & ~n26782 ;
  assign n26784 = ( ~n13741 & n13744 ) | ( ~n13741 & n26783 ) | ( n13744 & n26783 ) ;
  assign n26785 = ( ~n13639 & n14582 ) | ( ~n13639 & n19391 ) | ( n14582 & n19391 ) ;
  assign n26786 = n2491 | n26785 ;
  assign n26787 = n10909 | n26786 ;
  assign n26788 = ( n141 & n4095 ) | ( n141 & n26787 ) | ( n4095 & n26787 ) ;
  assign n26789 = n17579 ^ n2306 ^ 1'b0 ;
  assign n26790 = n26788 | n26789 ;
  assign n26791 = n19385 ^ n17475 ^ n6183 ;
  assign n26792 = n22190 ^ n7110 ^ n6865 ;
  assign n26794 = n22398 ^ n12000 ^ n10845 ;
  assign n26793 = n16908 ^ n8450 ^ n216 ;
  assign n26795 = n26794 ^ n26793 ^ n2777 ;
  assign n26796 = ( n11087 & ~n22867 ) | ( n11087 & n23501 ) | ( ~n22867 & n23501 ) ;
  assign n26797 = ( n12553 & n15101 ) | ( n12553 & ~n20108 ) | ( n15101 & ~n20108 ) ;
  assign n26798 = n26797 ^ n20352 ^ n15877 ;
  assign n26799 = ( n14486 & n17788 ) | ( n14486 & ~n24751 ) | ( n17788 & ~n24751 ) ;
  assign n26800 = n13134 ^ n11640 ^ 1'b0 ;
  assign n26801 = n13589 & n26800 ;
  assign n26802 = ~n9935 & n14897 ;
  assign n26803 = n8561 ^ n3916 ^ n2160 ;
  assign n26804 = n7976 & ~n24790 ;
  assign n26805 = ~n26803 & n26804 ;
  assign n26806 = n24247 ^ n10676 ^ n4927 ;
  assign n26807 = ( n8547 & n18073 ) | ( n8547 & ~n24665 ) | ( n18073 & ~n24665 ) ;
  assign n26811 = n8651 ^ n3131 ^ x124 ;
  assign n26808 = n19522 ^ n15893 ^ n15379 ;
  assign n26809 = n26808 ^ n17822 ^ n2308 ;
  assign n26810 = n26809 ^ n11172 ^ n2108 ;
  assign n26812 = n26811 ^ n26810 ^ n12386 ;
  assign n26813 = n15593 ^ n13695 ^ 1'b0 ;
  assign n26814 = n4081 & n26813 ;
  assign n26815 = ( ~n3437 & n23215 ) | ( ~n3437 & n26814 ) | ( n23215 & n26814 ) ;
  assign n26816 = ( n11985 & n24268 ) | ( n11985 & n26815 ) | ( n24268 & n26815 ) ;
  assign n26817 = n6236 | n11899 ;
  assign n26818 = n2752 & ~n12735 ;
  assign n26819 = n15464 & n26147 ;
  assign n26820 = n2166 | n6191 ;
  assign n26821 = x102 & ~n26820 ;
  assign n26822 = ( ~n7068 & n10343 ) | ( ~n7068 & n18569 ) | ( n10343 & n18569 ) ;
  assign n26823 = n7511 ^ n5589 ^ 1'b0 ;
  assign n26824 = n11193 ^ n5657 ^ n1560 ;
  assign n26825 = n4770 ^ n2132 ^ n1667 ;
  assign n26826 = n3096 & ~n26825 ;
  assign n26827 = ~n2887 & n26826 ;
  assign n26828 = n26827 ^ n9477 ^ n206 ;
  assign n26829 = ( ~n20635 & n26824 ) | ( ~n20635 & n26828 ) | ( n26824 & n26828 ) ;
  assign n26830 = n21942 ^ n10191 ^ n3735 ;
  assign n26831 = n26830 ^ n22562 ^ 1'b0 ;
  assign n26832 = ( n20462 & n21653 ) | ( n20462 & n26831 ) | ( n21653 & n26831 ) ;
  assign n26833 = n26832 ^ n23702 ^ x92 ;
  assign n26834 = n11613 ^ n3078 ^ 1'b0 ;
  assign n26835 = ( ~n8931 & n21821 ) | ( ~n8931 & n26834 ) | ( n21821 & n26834 ) ;
  assign n26836 = n2555 & ~n13171 ;
  assign n26837 = n26836 ^ n13753 ^ 1'b0 ;
  assign n26838 = n12585 ^ n187 ^ 1'b0 ;
  assign n26839 = n12602 & n26838 ;
  assign n26840 = ~n11943 & n26839 ;
  assign n26841 = n14246 & n26840 ;
  assign n26842 = n18804 ^ n5866 ^ 1'b0 ;
  assign n26843 = ( n19747 & ~n23971 ) | ( n19747 & n26842 ) | ( ~n23971 & n26842 ) ;
  assign n26844 = n11348 ^ n3587 ^ 1'b0 ;
  assign n26845 = ( n7641 & ~n19189 ) | ( n7641 & n26844 ) | ( ~n19189 & n26844 ) ;
  assign n26846 = n22009 ^ n3554 ^ 1'b0 ;
  assign n26847 = n9989 ^ n1553 ^ 1'b0 ;
  assign n26848 = ( n21133 & n21202 ) | ( n21133 & ~n26847 ) | ( n21202 & ~n26847 ) ;
  assign n26849 = n21993 ^ n20544 ^ n4882 ;
  assign n26850 = n23319 ^ n12418 ^ n3184 ;
  assign n26851 = ( n967 & n10526 ) | ( n967 & ~n12950 ) | ( n10526 & ~n12950 ) ;
  assign n26852 = ( n26849 & ~n26850 ) | ( n26849 & n26851 ) | ( ~n26850 & n26851 ) ;
  assign n26853 = ( ~n1755 & n10149 ) | ( ~n1755 & n10959 ) | ( n10149 & n10959 ) ;
  assign n26854 = n26853 ^ n11033 ^ n7625 ;
  assign n26855 = n26854 ^ n13479 ^ 1'b0 ;
  assign n26856 = ~n15040 & n26855 ;
  assign n26857 = ~n15306 & n22845 ;
  assign n26858 = n26857 ^ n17817 ^ 1'b0 ;
  assign n26859 = n22789 ^ n20381 ^ 1'b0 ;
  assign n26860 = n26858 & ~n26859 ;
  assign n26861 = n3666 & ~n17560 ;
  assign n26862 = n26861 ^ n6974 ^ 1'b0 ;
  assign n26863 = n15586 | n26862 ;
  assign n26864 = n5910 & ~n26863 ;
  assign n26865 = n16630 & n16714 ;
  assign n26866 = n26865 ^ n9628 ^ n6237 ;
  assign n26867 = ~n4357 & n26866 ;
  assign n26868 = ( n17311 & ~n23133 ) | ( n17311 & n24869 ) | ( ~n23133 & n24869 ) ;
  assign n26869 = n1048 | n18703 ;
  assign n26870 = ( n3002 & ~n3421 ) | ( n3002 & n17448 ) | ( ~n3421 & n17448 ) ;
  assign n26871 = ( n7185 & n26038 ) | ( n7185 & n26870 ) | ( n26038 & n26870 ) ;
  assign n26872 = ( n22368 & n23356 ) | ( n22368 & n26871 ) | ( n23356 & n26871 ) ;
  assign n26873 = n13134 ^ n11651 ^ n192 ;
  assign n26874 = n26873 ^ n16374 ^ n3217 ;
  assign n26875 = n26874 ^ n21051 ^ n11126 ;
  assign n26876 = n26875 ^ n18347 ^ 1'b0 ;
  assign n26877 = n16867 & ~n23470 ;
  assign n26878 = n26877 ^ n26476 ^ 1'b0 ;
  assign n26879 = n17120 | n23500 ;
  assign n26882 = n22052 ^ n18484 ^ n6411 ;
  assign n26880 = n21481 ^ n9375 ^ 1'b0 ;
  assign n26881 = n3267 & ~n26880 ;
  assign n26883 = n26882 ^ n26881 ^ n9180 ;
  assign n26884 = n26879 & n26883 ;
  assign n26885 = ~n1422 & n26884 ;
  assign n26886 = n17043 & ~n25378 ;
  assign n26887 = n26886 ^ n2606 ^ 1'b0 ;
  assign n26888 = n16530 ^ n6621 ^ 1'b0 ;
  assign n26889 = n26888 ^ n16782 ^ 1'b0 ;
  assign n26890 = n24054 ^ n1479 ^ n1152 ;
  assign n26891 = ~n1687 & n12328 ;
  assign n26892 = n26891 ^ n18566 ^ 1'b0 ;
  assign n26893 = ( ~n3874 & n5419 ) | ( ~n3874 & n26892 ) | ( n5419 & n26892 ) ;
  assign n26894 = ( n2943 & n13923 ) | ( n2943 & ~n19950 ) | ( n13923 & ~n19950 ) ;
  assign n26897 = n14450 ^ n6923 ^ n6721 ;
  assign n26895 = n20202 ^ n19942 ^ n10901 ;
  assign n26896 = n26895 ^ n11764 ^ n4855 ;
  assign n26898 = n26897 ^ n26896 ^ n26251 ;
  assign n26899 = ( ~n12433 & n23754 ) | ( ~n12433 & n25815 ) | ( n23754 & n25815 ) ;
  assign n26900 = ( n2219 & ~n2305 ) | ( n2219 & n15325 ) | ( ~n2305 & n15325 ) ;
  assign n26902 = n26534 ^ n15901 ^ n10754 ;
  assign n26901 = n11686 & n26668 ;
  assign n26903 = n26902 ^ n26901 ^ 1'b0 ;
  assign n26905 = n21118 ^ n16283 ^ 1'b0 ;
  assign n26904 = n13433 | n19079 ;
  assign n26906 = n26905 ^ n26904 ^ 1'b0 ;
  assign n26907 = ~n14414 & n20419 ;
  assign n26908 = n26907 ^ n26627 ^ 1'b0 ;
  assign n26913 = n15390 ^ n11169 ^ n4951 ;
  assign n26909 = ( n3391 & n3486 ) | ( n3391 & ~n9296 ) | ( n3486 & ~n9296 ) ;
  assign n26910 = ( n5769 & ~n15345 ) | ( n5769 & n26909 ) | ( ~n15345 & n26909 ) ;
  assign n26911 = ~n977 & n2832 ;
  assign n26912 = ~n26910 & n26911 ;
  assign n26914 = n26913 ^ n26912 ^ n3881 ;
  assign n26915 = n5932 & n15238 ;
  assign n26916 = n26915 ^ n14556 ^ 1'b0 ;
  assign n26917 = n26916 ^ n7211 ^ n3055 ;
  assign n26918 = n16457 ^ n13450 ^ n4214 ;
  assign n26919 = n25588 ^ n8203 ^ 1'b0 ;
  assign n26920 = n10792 & n26919 ;
  assign n26921 = n10206 & ~n10564 ;
  assign n26922 = ~n4511 & n26921 ;
  assign n26923 = n8663 & ~n9532 ;
  assign n26924 = n1038 & n26923 ;
  assign n26925 = n2463 & n10898 ;
  assign n26926 = n26924 & n26925 ;
  assign n26927 = ( n9860 & n20117 ) | ( n9860 & n21306 ) | ( n20117 & n21306 ) ;
  assign n26928 = ( n6114 & ~n22303 ) | ( n6114 & n26927 ) | ( ~n22303 & n26927 ) ;
  assign n26929 = n18699 ^ n5241 ^ n624 ;
  assign n26930 = n26583 ^ n20319 ^ n1895 ;
  assign n26931 = n8534 ^ n4340 ^ n3778 ;
  assign n26932 = ~n15924 & n26931 ;
  assign n26933 = n10738 & n26932 ;
  assign n26934 = n26933 ^ n22201 ^ n4164 ;
  assign n26935 = n19403 ^ n4350 ^ 1'b0 ;
  assign n26936 = n3390 | n26935 ;
  assign n26937 = ~n11243 & n21540 ;
  assign n26938 = n26937 ^ n9210 ^ 1'b0 ;
  assign n26939 = n21511 & ~n26938 ;
  assign n26940 = n20676 ^ n12085 ^ 1'b0 ;
  assign n26941 = n18065 | n26940 ;
  assign n26942 = ( n11695 & n15766 ) | ( n11695 & ~n17866 ) | ( n15766 & ~n17866 ) ;
  assign n26943 = n26942 ^ n13982 ^ n11225 ;
  assign n26944 = n1584 & n26454 ;
  assign n26945 = ( n10560 & ~n23919 ) | ( n10560 & n26488 ) | ( ~n23919 & n26488 ) ;
  assign n26946 = ~n2157 & n21765 ;
  assign n26947 = ( n6812 & ~n22564 ) | ( n6812 & n26946 ) | ( ~n22564 & n26946 ) ;
  assign n26948 = n15940 & ~n17526 ;
  assign n26949 = n17911 ^ n10313 ^ 1'b0 ;
  assign n26950 = n20551 ^ n6503 ^ n4910 ;
  assign n26951 = n711 & n4139 ;
  assign n26952 = n26951 ^ n4294 ^ 1'b0 ;
  assign n26953 = n9511 & n26952 ;
  assign n26954 = n26953 ^ n1839 ^ 1'b0 ;
  assign n26955 = ( n14791 & ~n21356 ) | ( n14791 & n26954 ) | ( ~n21356 & n26954 ) ;
  assign n26956 = n23575 ^ n6087 ^ n2844 ;
  assign n26957 = n2011 ^ n774 ^ 1'b0 ;
  assign n26958 = ( ~n3122 & n14517 ) | ( ~n3122 & n26957 ) | ( n14517 & n26957 ) ;
  assign n26959 = n21680 & n26739 ;
  assign n26960 = ( n13790 & n26958 ) | ( n13790 & n26959 ) | ( n26958 & n26959 ) ;
  assign n26961 = ( n721 & n10640 ) | ( n721 & ~n14212 ) | ( n10640 & ~n14212 ) ;
  assign n26962 = n19928 ^ n15020 ^ n1079 ;
  assign n26963 = n26962 ^ n17947 ^ 1'b0 ;
  assign n26964 = ( n2602 & ~n3850 ) | ( n2602 & n9458 ) | ( ~n3850 & n9458 ) ;
  assign n26965 = ( n12053 & ~n13727 ) | ( n12053 & n26964 ) | ( ~n13727 & n26964 ) ;
  assign n26966 = n4839 & n8669 ;
  assign n26967 = n26966 ^ n11690 ^ n2360 ;
  assign n26968 = ~n22615 & n26967 ;
  assign n26969 = n19223 ^ n8002 ^ 1'b0 ;
  assign n26970 = n24484 ^ n4765 ^ 1'b0 ;
  assign n26971 = n26969 & ~n26970 ;
  assign n26972 = n16527 ^ n12778 ^ 1'b0 ;
  assign n26973 = n17332 ^ n11574 ^ n5737 ;
  assign n26974 = n13325 ^ n6645 ^ n1515 ;
  assign n26975 = n20276 & n26974 ;
  assign n26976 = n8446 & n26975 ;
  assign n26977 = ( n13324 & n16462 ) | ( n13324 & ~n26976 ) | ( n16462 & ~n26976 ) ;
  assign n26978 = n24807 ^ n14963 ^ n1971 ;
  assign n26979 = n25369 ^ n9937 ^ n8752 ;
  assign n26980 = ~n517 & n26820 ;
  assign n26981 = ( n3254 & ~n3453 ) | ( n3254 & n25316 ) | ( ~n3453 & n25316 ) ;
  assign n26982 = n5583 & ~n11283 ;
  assign n26983 = n6736 ^ n6709 ^ 1'b0 ;
  assign n26984 = n8261 & n26983 ;
  assign n26985 = n1663 | n23369 ;
  assign n26986 = n26985 ^ n8632 ^ 1'b0 ;
  assign n26987 = n7361 & ~n20407 ;
  assign n26988 = n26987 ^ n5048 ^ 1'b0 ;
  assign n26989 = n19943 & ~n26479 ;
  assign n26990 = n26989 ^ n15728 ^ 1'b0 ;
  assign n26991 = n26988 & ~n26990 ;
  assign n26992 = n18401 ^ n14173 ^ n7262 ;
  assign n26993 = n13312 ^ n10513 ^ 1'b0 ;
  assign n26994 = n14923 & ~n17953 ;
  assign n26995 = n3404 & n26994 ;
  assign n26996 = n26995 ^ n25359 ^ n21063 ;
  assign n26997 = n26996 ^ n7766 ^ 1'b0 ;
  assign n26998 = ( n23443 & n26993 ) | ( n23443 & n26997 ) | ( n26993 & n26997 ) ;
  assign n26999 = ( n3432 & n7465 ) | ( n3432 & n15697 ) | ( n7465 & n15697 ) ;
  assign n27000 = n7171 ^ n1948 ^ x127 ;
  assign n27001 = n27000 ^ n2488 ^ 1'b0 ;
  assign n27002 = n27001 ^ n18767 ^ n3146 ;
  assign n27003 = n17737 ^ n5389 ^ 1'b0 ;
  assign n27004 = n5332 | n27003 ;
  assign n27005 = n27004 ^ n17158 ^ n3679 ;
  assign n27006 = n27005 ^ n10440 ^ n3197 ;
  assign n27007 = n13875 ^ n9732 ^ n2640 ;
  assign n27008 = n18698 ^ n4061 ^ 1'b0 ;
  assign n27009 = n14791 | n21815 ;
  assign n27010 = ~n5048 & n8335 ;
  assign n27011 = n2372 & n27010 ;
  assign n27012 = n22678 ^ n848 ^ n603 ;
  assign n27013 = ( n6258 & ~n27011 ) | ( n6258 & n27012 ) | ( ~n27011 & n27012 ) ;
  assign n27014 = n8992 & n16248 ;
  assign n27015 = n27014 ^ n3080 ^ 1'b0 ;
  assign n27016 = ( ~n7429 & n18619 ) | ( ~n7429 & n22663 ) | ( n18619 & n22663 ) ;
  assign n27017 = n3054 & n27016 ;
  assign n27018 = ~n10587 & n27017 ;
  assign n27019 = ( n12457 & ~n20993 ) | ( n12457 & n23201 ) | ( ~n20993 & n23201 ) ;
  assign n27020 = ( n3823 & ~n4943 ) | ( n3823 & n12278 ) | ( ~n4943 & n12278 ) ;
  assign n27021 = ( n25109 & n25424 ) | ( n25109 & ~n27020 ) | ( n25424 & ~n27020 ) ;
  assign n27022 = ~n6272 & n11111 ;
  assign n27023 = ~n2509 & n27022 ;
  assign n27024 = n8728 ^ n3816 ^ n664 ;
  assign n27025 = ( n11806 & n27023 ) | ( n11806 & ~n27024 ) | ( n27023 & ~n27024 ) ;
  assign n27026 = n15940 ^ n9427 ^ n1637 ;
  assign n27027 = n10855 ^ n8116 ^ n7724 ;
  assign n27028 = n20289 ^ n2280 ^ 1'b0 ;
  assign n27029 = n2585 & ~n27028 ;
  assign n27030 = ( n3785 & n4560 ) | ( n3785 & ~n20516 ) | ( n4560 & ~n20516 ) ;
  assign n27031 = n2733 & ~n19114 ;
  assign n27032 = ~n27030 & n27031 ;
  assign n27033 = ( n11742 & n13896 ) | ( n11742 & n14001 ) | ( n13896 & n14001 ) ;
  assign n27034 = n27033 ^ n11482 ^ 1'b0 ;
  assign n27035 = n2408 & n27034 ;
  assign n27036 = ( n8344 & n9095 ) | ( n8344 & n24634 ) | ( n9095 & n24634 ) ;
  assign n27037 = ( ~n1498 & n11065 ) | ( ~n1498 & n23509 ) | ( n11065 & n23509 ) ;
  assign n27038 = n19026 ^ n12653 ^ n8633 ;
  assign n27039 = ( n967 & n21715 ) | ( n967 & n27038 ) | ( n21715 & n27038 ) ;
  assign n27040 = n21733 ^ n15256 ^ 1'b0 ;
  assign n27042 = ( n2324 & n3725 ) | ( n2324 & n3786 ) | ( n3725 & n3786 ) ;
  assign n27041 = n13482 | n19585 ;
  assign n27043 = n27042 ^ n27041 ^ n19764 ;
  assign n27044 = ( ~n5719 & n9933 ) | ( ~n5719 & n13920 ) | ( n9933 & n13920 ) ;
  assign n27045 = n1647 | n27044 ;
  assign n27046 = n7823 | n10253 ;
  assign n27047 = n12615 ^ n2311 ^ 1'b0 ;
  assign n27048 = ( n15412 & ~n25075 ) | ( n15412 & n27047 ) | ( ~n25075 & n27047 ) ;
  assign n27051 = n12681 | n23944 ;
  assign n27052 = n27051 ^ n20086 ^ 1'b0 ;
  assign n27049 = n21867 ^ n4680 ^ 1'b0 ;
  assign n27050 = n14092 | n27049 ;
  assign n27053 = n27052 ^ n27050 ^ n4396 ;
  assign n27054 = n15676 ^ n11204 ^ 1'b0 ;
  assign n27055 = n8469 ^ n6864 ^ n5787 ;
  assign n27056 = n11222 ^ n9919 ^ n698 ;
  assign n27057 = n9738 & ~n19816 ;
  assign n27058 = n27057 ^ n16157 ^ 1'b0 ;
  assign n27059 = ( n25436 & n27056 ) | ( n25436 & ~n27058 ) | ( n27056 & ~n27058 ) ;
  assign n27060 = n27059 ^ n16345 ^ n13915 ;
  assign n27061 = ~n11170 & n27060 ;
  assign n27062 = ( n22056 & n27055 ) | ( n22056 & ~n27061 ) | ( n27055 & ~n27061 ) ;
  assign n27063 = ( ~n5586 & n7059 ) | ( ~n5586 & n13021 ) | ( n7059 & n13021 ) ;
  assign n27064 = ~n12057 & n22155 ;
  assign n27065 = n24656 ^ n9645 ^ n4545 ;
  assign n27066 = n10973 | n27065 ;
  assign n27067 = n12824 | n23849 ;
  assign n27068 = n24149 & ~n27067 ;
  assign n27069 = n13480 & n18820 ;
  assign n27070 = ~n8695 & n27069 ;
  assign n27071 = n15135 ^ n7524 ^ 1'b0 ;
  assign n27072 = ~n27070 & n27071 ;
  assign n27073 = n22025 ^ n12945 ^ 1'b0 ;
  assign n27074 = n27061 ^ n24122 ^ n8992 ;
  assign n27075 = ( n6772 & ~n11139 ) | ( n6772 & n12030 ) | ( ~n11139 & n12030 ) ;
  assign n27076 = n12489 ^ n2345 ^ n469 ;
  assign n27077 = n27076 ^ n23769 ^ n11448 ;
  assign n27078 = ~n1865 & n19123 ;
  assign n27079 = n2070 & n27078 ;
  assign n27080 = ~n13295 & n27079 ;
  assign n27081 = n6946 | n9637 ;
  assign n27082 = n19878 | n27081 ;
  assign n27083 = n22937 & ~n25282 ;
  assign n27084 = n27083 ^ n20632 ^ 1'b0 ;
  assign n27085 = n6942 ^ n3456 ^ 1'b0 ;
  assign n27086 = n7479 ^ n1482 ^ n979 ;
  assign n27087 = n9354 ^ n197 ^ 1'b0 ;
  assign n27088 = n16131 & n18532 ;
  assign n27089 = n27088 ^ n16281 ^ 1'b0 ;
  assign n27090 = n27089 ^ n2007 ^ 1'b0 ;
  assign n27091 = ~n2005 & n27090 ;
  assign n27092 = n8864 ^ n5882 ^ 1'b0 ;
  assign n27093 = n21402 ^ n1013 ^ 1'b0 ;
  assign n27094 = n27092 & ~n27093 ;
  assign n27095 = n20481 ^ n7249 ^ n1781 ;
  assign n27096 = n27095 ^ n12509 ^ n6633 ;
  assign n27097 = n23759 ^ n11460 ^ n5694 ;
  assign n27098 = ( ~n3220 & n19810 ) | ( ~n3220 & n27097 ) | ( n19810 & n27097 ) ;
  assign n27099 = n11189 ^ n3778 ^ n3301 ;
  assign n27100 = n27099 ^ n18034 ^ n14233 ;
  assign n27101 = n7738 ^ n2098 ^ 1'b0 ;
  assign n27102 = n23860 ^ n7445 ^ 1'b0 ;
  assign n27103 = ( n5318 & ~n17002 ) | ( n5318 & n21642 ) | ( ~n17002 & n21642 ) ;
  assign n27104 = n3364 & n27103 ;
  assign n27107 = n19648 ^ n4279 ^ n1966 ;
  assign n27108 = n19495 & ~n27107 ;
  assign n27105 = n18511 ^ n339 ^ n187 ;
  assign n27106 = ~n23536 & n27105 ;
  assign n27109 = n27108 ^ n27106 ^ 1'b0 ;
  assign n27110 = n12196 ^ n5496 ^ n576 ;
  assign n27111 = n22635 & ~n27110 ;
  assign n27112 = n13054 ^ n9081 ^ n5100 ;
  assign n27113 = n6355 ^ n1808 ^ 1'b0 ;
  assign n27114 = n4971 | n27113 ;
  assign n27115 = n22163 ^ n4758 ^ 1'b0 ;
  assign n27116 = n14067 | n27115 ;
  assign n27117 = n27114 | n27116 ;
  assign n27118 = n13893 ^ n7176 ^ n2516 ;
  assign n27119 = ( n2630 & n12248 ) | ( n2630 & n27118 ) | ( n12248 & n27118 ) ;
  assign n27120 = ( x121 & ~n7943 ) | ( x121 & n22395 ) | ( ~n7943 & n22395 ) ;
  assign n27121 = n27120 ^ n24294 ^ n10194 ;
  assign n27123 = n5595 & ~n12139 ;
  assign n27124 = n27123 ^ n131 ^ 1'b0 ;
  assign n27122 = n10684 ^ n10355 ^ 1'b0 ;
  assign n27125 = n27124 ^ n27122 ^ x102 ;
  assign n27126 = ( ~n2716 & n14078 ) | ( ~n2716 & n19040 ) | ( n14078 & n19040 ) ;
  assign n27127 = ( ~n4820 & n27125 ) | ( ~n4820 & n27126 ) | ( n27125 & n27126 ) ;
  assign n27128 = ( ~n226 & n1989 ) | ( ~n226 & n13895 ) | ( n1989 & n13895 ) ;
  assign n27129 = ~n8708 & n14139 ;
  assign n27130 = n27129 ^ n12489 ^ 1'b0 ;
  assign n27131 = ( ~n4222 & n5021 ) | ( ~n4222 & n18185 ) | ( n5021 & n18185 ) ;
  assign n27132 = ( n2639 & n4349 ) | ( n2639 & ~n27131 ) | ( n4349 & ~n27131 ) ;
  assign n27133 = n27132 ^ n15838 ^ 1'b0 ;
  assign n27134 = n10290 ^ n429 ^ 1'b0 ;
  assign n27138 = ( ~x62 & n7260 ) | ( ~x62 & n12546 ) | ( n7260 & n12546 ) ;
  assign n27136 = n9867 | n18645 ;
  assign n27137 = n27136 ^ n12525 ^ 1'b0 ;
  assign n27135 = n25360 ^ n15405 ^ n14658 ;
  assign n27139 = n27138 ^ n27137 ^ n27135 ;
  assign n27140 = n5971 | n7915 ;
  assign n27141 = n16491 & ~n27140 ;
  assign n27142 = n27141 ^ n19091 ^ 1'b0 ;
  assign n27143 = n22316 ^ n10901 ^ 1'b0 ;
  assign n27146 = n6238 & n16966 ;
  assign n27145 = ( n12150 & ~n25313 ) | ( n12150 & n26335 ) | ( ~n25313 & n26335 ) ;
  assign n27144 = n5526 & ~n15824 ;
  assign n27147 = n27146 ^ n27145 ^ n27144 ;
  assign n27148 = ( n3343 & ~n15311 ) | ( n3343 & n21442 ) | ( ~n15311 & n21442 ) ;
  assign n27149 = n27148 ^ n26330 ^ n16816 ;
  assign n27150 = n1931 | n13996 ;
  assign n27151 = n27150 ^ n2279 ^ 1'b0 ;
  assign n27152 = n2909 | n27151 ;
  assign n27153 = n796 & ~n7766 ;
  assign n27154 = ~n3146 & n27153 ;
  assign n27155 = ( n2515 & ~n7576 ) | ( n2515 & n18992 ) | ( ~n7576 & n18992 ) ;
  assign n27156 = n27155 ^ n13702 ^ 1'b0 ;
  assign n27157 = n9416 | n27156 ;
  assign n27158 = n16623 ^ n9293 ^ 1'b0 ;
  assign n27159 = ~n27157 & n27158 ;
  assign n27160 = ( n6130 & n7200 ) | ( n6130 & ~n8260 ) | ( n7200 & ~n8260 ) ;
  assign n27161 = ~n9819 & n27160 ;
  assign n27162 = ( ~n17463 & n21470 ) | ( ~n17463 & n22434 ) | ( n21470 & n22434 ) ;
  assign n27163 = ( ~n15306 & n22559 ) | ( ~n15306 & n26543 ) | ( n22559 & n26543 ) ;
  assign n27164 = ( ~n933 & n12993 ) | ( ~n933 & n16339 ) | ( n12993 & n16339 ) ;
  assign n27165 = n27164 ^ n10223 ^ 1'b0 ;
  assign n27166 = n12969 | n13829 ;
  assign n27167 = ( n2792 & ~n4053 ) | ( n2792 & n14862 ) | ( ~n4053 & n14862 ) ;
  assign n27168 = n23378 ^ n21135 ^ n10460 ;
  assign n27169 = n27168 ^ n4392 ^ 1'b0 ;
  assign n27170 = n19282 ^ n4880 ^ 1'b0 ;
  assign n27171 = n27169 & n27170 ;
  assign n27172 = n14935 | n18412 ;
  assign n27173 = n27172 ^ n780 ^ 1'b0 ;
  assign n27174 = ( n4810 & n9261 ) | ( n4810 & n21232 ) | ( n9261 & n21232 ) ;
  assign n27175 = n27174 ^ n3586 ^ 1'b0 ;
  assign n27176 = n6083 ^ x118 ^ 1'b0 ;
  assign n27177 = ( n11693 & n16096 ) | ( n11693 & ~n27176 ) | ( n16096 & ~n27176 ) ;
  assign n27178 = ( n15454 & ~n18319 ) | ( n15454 & n23596 ) | ( ~n18319 & n23596 ) ;
  assign n27181 = ( n6386 & n15139 ) | ( n6386 & ~n17800 ) | ( n15139 & ~n17800 ) ;
  assign n27182 = n11140 & ~n27181 ;
  assign n27179 = n20015 ^ n14885 ^ n7469 ;
  assign n27180 = n11888 | n27179 ;
  assign n27183 = n27182 ^ n27180 ^ n16494 ;
  assign n27186 = n23743 ^ n13390 ^ n6912 ;
  assign n27184 = n7474 ^ n812 ^ 1'b0 ;
  assign n27185 = n27184 ^ n13773 ^ n3389 ;
  assign n27187 = n27186 ^ n27185 ^ n13297 ;
  assign n27190 = n1418 & n6018 ;
  assign n27191 = n6828 & n27190 ;
  assign n27189 = n16673 ^ n4915 ^ n1267 ;
  assign n27192 = n27191 ^ n27189 ^ n15406 ;
  assign n27188 = ( ~n13381 & n13547 ) | ( ~n13381 & n19478 ) | ( n13547 & n19478 ) ;
  assign n27193 = n27192 ^ n27188 ^ n26854 ;
  assign n27194 = n27193 ^ n11234 ^ n9988 ;
  assign n27195 = n20729 ^ n2501 ^ 1'b0 ;
  assign n27196 = n6586 | n27195 ;
  assign n27198 = n22125 ^ n5780 ^ n4474 ;
  assign n27197 = ~n20711 & n25965 ;
  assign n27199 = n27198 ^ n27197 ^ 1'b0 ;
  assign n27200 = n26862 ^ n12490 ^ n2617 ;
  assign n27201 = n390 & n21461 ;
  assign n27202 = ( n7844 & ~n14394 ) | ( n7844 & n27201 ) | ( ~n14394 & n27201 ) ;
  assign n27203 = ( n6872 & n12522 ) | ( n6872 & n19411 ) | ( n12522 & n19411 ) ;
  assign n27204 = ( n16152 & n27148 ) | ( n16152 & ~n27203 ) | ( n27148 & ~n27203 ) ;
  assign n27205 = n27204 ^ n18990 ^ n12118 ;
  assign n27206 = n7779 & ~n12380 ;
  assign n27207 = ( n319 & ~n11687 ) | ( n319 & n17307 ) | ( ~n11687 & n17307 ) ;
  assign n27213 = n6914 ^ n425 ^ 1'b0 ;
  assign n27208 = n11511 & ~n15451 ;
  assign n27209 = n8771 | n18251 ;
  assign n27210 = n27209 ^ n17218 ^ 1'b0 ;
  assign n27211 = ~n27208 & n27210 ;
  assign n27212 = n27211 ^ n1496 ^ 1'b0 ;
  assign n27214 = n27213 ^ n27212 ^ n7377 ;
  assign n27215 = n8279 & ~n9966 ;
  assign n27216 = ~n14815 & n27215 ;
  assign n27217 = n1600 | n17077 ;
  assign n27218 = n27217 ^ n11772 ^ 1'b0 ;
  assign n27219 = ( n2930 & n6251 ) | ( n2930 & ~n18181 ) | ( n6251 & ~n18181 ) ;
  assign n27220 = ~n1643 & n27219 ;
  assign n27221 = n6305 ^ n5097 ^ n629 ;
  assign n27225 = n860 | n7622 ;
  assign n27224 = ( ~n2380 & n2620 ) | ( ~n2380 & n4921 ) | ( n2620 & n4921 ) ;
  assign n27222 = n11849 ^ n5264 ^ n1969 ;
  assign n27223 = ~n15012 & n27222 ;
  assign n27226 = n27225 ^ n27224 ^ n27223 ;
  assign n27227 = ( n1040 & n27221 ) | ( n1040 & n27226 ) | ( n27221 & n27226 ) ;
  assign n27228 = ( n6610 & ~n15014 ) | ( n6610 & n16939 ) | ( ~n15014 & n16939 ) ;
  assign n27229 = n2250 | n7418 ;
  assign n27230 = n27229 ^ n23626 ^ 1'b0 ;
  assign n27231 = n16282 ^ n2470 ^ n1097 ;
  assign n27232 = ( ~n4344 & n13646 ) | ( ~n4344 & n27231 ) | ( n13646 & n27231 ) ;
  assign n27233 = n27232 ^ n22761 ^ n20022 ;
  assign n27234 = n27230 & n27233 ;
  assign n27235 = n27234 ^ n14303 ^ n7311 ;
  assign n27236 = n5466 ^ x112 ^ 1'b0 ;
  assign n27237 = ~n4748 & n27236 ;
  assign n27238 = ~n3858 & n6546 ;
  assign n27239 = ~n10641 & n27238 ;
  assign n27240 = n5419 & n7651 ;
  assign n27241 = n27239 & n27240 ;
  assign n27242 = ( ~n10223 & n23998 ) | ( ~n10223 & n27241 ) | ( n23998 & n27241 ) ;
  assign n27243 = n27237 & n27242 ;
  assign n27244 = ~n9760 & n9766 ;
  assign n27245 = ( n8154 & n21597 ) | ( n8154 & ~n27244 ) | ( n21597 & ~n27244 ) ;
  assign n27246 = n4585 ^ n4354 ^ 1'b0 ;
  assign n27247 = ~n3950 & n27246 ;
  assign n27248 = n27247 ^ n24721 ^ 1'b0 ;
  assign n27250 = n3891 & n12077 ;
  assign n27251 = n27250 ^ n4797 ^ 1'b0 ;
  assign n27249 = n2232 & ~n19465 ;
  assign n27252 = n27251 ^ n27249 ^ 1'b0 ;
  assign n27253 = n15983 ^ n7139 ^ n3671 ;
  assign n27254 = ( ~n8834 & n11509 ) | ( ~n8834 & n14209 ) | ( n11509 & n14209 ) ;
  assign n27255 = n11851 ^ n7230 ^ 1'b0 ;
  assign n27256 = ~n7605 & n27255 ;
  assign n27257 = ( n7323 & n11939 ) | ( n7323 & ~n27256 ) | ( n11939 & ~n27256 ) ;
  assign n27258 = n20821 | n24067 ;
  assign n27259 = ( n1167 & n7152 ) | ( n1167 & ~n16098 ) | ( n7152 & ~n16098 ) ;
  assign n27260 = n2518 & n22501 ;
  assign n27261 = ~n27259 & n27260 ;
  assign n27262 = n22691 & ~n26959 ;
  assign n27263 = n21827 | n27262 ;
  assign n27264 = n27263 ^ n1486 ^ 1'b0 ;
  assign n27265 = ~n7909 & n18456 ;
  assign n27266 = n3834 & n23368 ;
  assign n27267 = ( n3916 & n7277 ) | ( n3916 & n10087 ) | ( n7277 & n10087 ) ;
  assign n27268 = n17332 | n23083 ;
  assign n27269 = n11355 | n27268 ;
  assign n27270 = n27269 ^ n12471 ^ n6602 ;
  assign n27271 = n25480 ^ n4040 ^ n3516 ;
  assign n27272 = ( n5882 & n5963 ) | ( n5882 & ~n10152 ) | ( n5963 & ~n10152 ) ;
  assign n27273 = n27272 ^ n23143 ^ 1'b0 ;
  assign n27274 = ( n3102 & ~n3934 ) | ( n3102 & n27273 ) | ( ~n3934 & n27273 ) ;
  assign n27275 = n5790 & ~n11333 ;
  assign n27276 = n27275 ^ n13953 ^ 1'b0 ;
  assign n27277 = n10450 ^ n1163 ^ n928 ;
  assign n27278 = n27277 ^ n7707 ^ 1'b0 ;
  assign n27279 = n1081 | n9148 ;
  assign n27280 = n20061 | n27279 ;
  assign n27281 = n10583 ^ n9156 ^ n2851 ;
  assign n27282 = ( n4623 & n10096 ) | ( n4623 & n22802 ) | ( n10096 & n22802 ) ;
  assign n27283 = n27282 ^ n21035 ^ x50 ;
  assign n27284 = ( n3427 & n20974 ) | ( n3427 & ~n24344 ) | ( n20974 & ~n24344 ) ;
  assign n27285 = n20439 ^ n5886 ^ 1'b0 ;
  assign n27286 = n22546 & ~n27285 ;
  assign n27287 = ( ~n24725 & n27284 ) | ( ~n24725 & n27286 ) | ( n27284 & n27286 ) ;
  assign n27288 = ( n224 & n2198 ) | ( n224 & n26111 ) | ( n2198 & n26111 ) ;
  assign n27289 = n10142 & ~n19129 ;
  assign n27290 = n27289 ^ n12340 ^ 1'b0 ;
  assign n27291 = n5509 | n27290 ;
  assign n27292 = n27291 ^ n24070 ^ 1'b0 ;
  assign n27293 = n14533 & ~n16213 ;
  assign n27294 = n27293 ^ n8748 ^ 1'b0 ;
  assign n27295 = ( n11079 & n12030 ) | ( n11079 & n12042 ) | ( n12030 & n12042 ) ;
  assign n27296 = n27295 ^ n9281 ^ 1'b0 ;
  assign n27297 = n13736 & n27296 ;
  assign n27298 = ( n1280 & n5932 ) | ( n1280 & ~n8590 ) | ( n5932 & ~n8590 ) ;
  assign n27299 = ~n25117 & n27298 ;
  assign n27300 = n27299 ^ x112 ^ 1'b0 ;
  assign n27301 = n16213 ^ n2693 ^ n1651 ;
  assign n27302 = n27301 ^ n17542 ^ n7900 ;
  assign n27303 = n3556 | n4015 ;
  assign n27304 = n8028 | n11169 ;
  assign n27305 = n27304 ^ n17450 ^ n13999 ;
  assign n27306 = n6365 & ~n25461 ;
  assign n27307 = n8123 & n27306 ;
  assign n27308 = ~n11501 & n14025 ;
  assign n27309 = n11543 & n27308 ;
  assign n27310 = n1377 & n12553 ;
  assign n27311 = n2749 & n5726 ;
  assign n27312 = n4459 ^ n2497 ^ 1'b0 ;
  assign n27313 = n27311 | n27312 ;
  assign n27314 = n8561 ^ n6208 ^ 1'b0 ;
  assign n27315 = ~n27313 & n27314 ;
  assign n27317 = n6092 & n24041 ;
  assign n27318 = n27317 ^ n19275 ^ 1'b0 ;
  assign n27316 = n6765 | n21837 ;
  assign n27319 = n27318 ^ n27316 ^ 1'b0 ;
  assign n27320 = n23763 ^ n2697 ^ 1'b0 ;
  assign n27321 = ( ~n24759 & n27319 ) | ( ~n24759 & n27320 ) | ( n27319 & n27320 ) ;
  assign n27323 = n2800 ^ n1462 ^ 1'b0 ;
  assign n27324 = n12545 ^ n4877 ^ n3983 ;
  assign n27325 = ( n12659 & n27323 ) | ( n12659 & n27324 ) | ( n27323 & n27324 ) ;
  assign n27322 = n5435 & n12027 ;
  assign n27326 = n27325 ^ n27322 ^ n13656 ;
  assign n27327 = n4900 & n14001 ;
  assign n27328 = ( n2762 & n3894 ) | ( n2762 & n5233 ) | ( n3894 & n5233 ) ;
  assign n27329 = n24832 ^ n21593 ^ n1404 ;
  assign n27330 = x6 & ~n24845 ;
  assign n27331 = ~n27329 & n27330 ;
  assign n27332 = n19148 ^ n2113 ^ 1'b0 ;
  assign n27333 = n23611 & n27332 ;
  assign n27334 = ~n159 & n24968 ;
  assign n27335 = n11731 & n27334 ;
  assign n27336 = n3198 & ~n13617 ;
  assign n27337 = n27336 ^ n23899 ^ 1'b0 ;
  assign n27338 = n18437 ^ n11602 ^ n1050 ;
  assign n27339 = n26046 ^ n15079 ^ n2356 ;
  assign n27340 = n27339 ^ n16627 ^ n4098 ;
  assign n27341 = ( n2740 & n8530 ) | ( n2740 & n21338 ) | ( n8530 & n21338 ) ;
  assign n27342 = n7443 & ~n12071 ;
  assign n27343 = ~n163 & n8429 ;
  assign n27344 = n25828 & n27343 ;
  assign n27345 = n12394 ^ n8642 ^ 1'b0 ;
  assign n27346 = n1993 & n27345 ;
  assign n27347 = n7722 | n26101 ;
  assign n27348 = n27347 ^ n1199 ^ 1'b0 ;
  assign n27353 = n20810 ^ n8758 ^ n6666 ;
  assign n27354 = n27353 ^ n7543 ^ 1'b0 ;
  assign n27355 = n27354 ^ n25510 ^ n7053 ;
  assign n27350 = n10796 ^ n9309 ^ n5560 ;
  assign n27349 = n21051 ^ n578 ^ 1'b0 ;
  assign n27351 = n27350 ^ n27349 ^ n6859 ;
  assign n27352 = ~n9556 & n27351 ;
  assign n27356 = n27355 ^ n27352 ^ 1'b0 ;
  assign n27357 = ( n10761 & n14150 ) | ( n10761 & n24043 ) | ( n14150 & n24043 ) ;
  assign n27358 = ( n18410 & ~n19232 ) | ( n18410 & n22683 ) | ( ~n19232 & n22683 ) ;
  assign n27359 = n27358 ^ n22319 ^ n11757 ;
  assign n27360 = ( n2370 & n3658 ) | ( n2370 & ~n11291 ) | ( n3658 & ~n11291 ) ;
  assign n27361 = n27360 ^ n9132 ^ n1947 ;
  assign n27362 = ( ~n158 & n10328 ) | ( ~n158 & n27361 ) | ( n10328 & n27361 ) ;
  assign n27363 = ( n5078 & ~n6102 ) | ( n5078 & n7461 ) | ( ~n6102 & n7461 ) ;
  assign n27364 = ( n6395 & n19233 ) | ( n6395 & ~n27363 ) | ( n19233 & ~n27363 ) ;
  assign n27365 = n27364 ^ n24342 ^ n2758 ;
  assign n27366 = n17455 ^ n14183 ^ 1'b0 ;
  assign n27367 = n27366 ^ n7634 ^ n6509 ;
  assign n27368 = ~n6192 & n12024 ;
  assign n27369 = n20739 & n27368 ;
  assign n27370 = ( n2761 & ~n17643 ) | ( n2761 & n23081 ) | ( ~n17643 & n23081 ) ;
  assign n27371 = n27370 ^ n4710 ^ 1'b0 ;
  assign n27372 = ~n1479 & n27371 ;
  assign n27373 = ( n6314 & ~n9933 ) | ( n6314 & n27372 ) | ( ~n9933 & n27372 ) ;
  assign n27374 = ( n293 & ~n7160 ) | ( n293 & n15532 ) | ( ~n7160 & n15532 ) ;
  assign n27375 = n14020 ^ n6681 ^ n4229 ;
  assign n27376 = n17207 & n17922 ;
  assign n27377 = n27376 ^ n22627 ^ n20258 ;
  assign n27378 = n27377 ^ n11505 ^ 1'b0 ;
  assign n27385 = ( n12818 & n13738 ) | ( n12818 & n17317 ) | ( n13738 & n17317 ) ;
  assign n27386 = n27385 ^ n26924 ^ n2856 ;
  assign n27383 = n3862 & ~n17429 ;
  assign n27384 = ~n13051 & n27383 ;
  assign n27379 = n19441 | n22455 ;
  assign n27380 = n2392 & ~n27379 ;
  assign n27381 = n27380 ^ n5415 ^ n2069 ;
  assign n27382 = ( n6341 & n9177 ) | ( n6341 & ~n27381 ) | ( n9177 & ~n27381 ) ;
  assign n27387 = n27386 ^ n27384 ^ n27382 ;
  assign n27388 = n13410 ^ n2077 ^ 1'b0 ;
  assign n27389 = n18983 ^ n13600 ^ 1'b0 ;
  assign n27390 = ~n6698 & n27389 ;
  assign n27391 = n16440 ^ n16106 ^ n13603 ;
  assign n27392 = ( n27388 & n27390 ) | ( n27388 & n27391 ) | ( n27390 & n27391 ) ;
  assign n27394 = n6476 ^ n4679 ^ n869 ;
  assign n27393 = n10225 ^ n9087 ^ 1'b0 ;
  assign n27395 = n27394 ^ n27393 ^ n1295 ;
  assign n27398 = n20321 ^ n7224 ^ x97 ;
  assign n27396 = n17372 ^ n4821 ^ n1424 ;
  assign n27397 = n6067 | n27396 ;
  assign n27399 = n27398 ^ n27397 ^ 1'b0 ;
  assign n27400 = ~n18512 & n26673 ;
  assign n27401 = n27400 ^ n19515 ^ 1'b0 ;
  assign n27402 = n15552 ^ n865 ^ 1'b0 ;
  assign n27403 = n13095 | n27402 ;
  assign n27404 = ( n3443 & ~n23998 ) | ( n3443 & n27403 ) | ( ~n23998 & n27403 ) ;
  assign n27405 = n27404 ^ n26756 ^ 1'b0 ;
  assign n27406 = n8398 | n27405 ;
  assign n27407 = n4495 & ~n15016 ;
  assign n27408 = n27407 ^ n10483 ^ 1'b0 ;
  assign n27409 = n27408 ^ n1348 ^ n913 ;
  assign n27410 = n3905 | n23952 ;
  assign n27411 = n27409 | n27410 ;
  assign n27412 = ( ~n15194 & n16778 ) | ( ~n15194 & n20601 ) | ( n16778 & n20601 ) ;
  assign n27413 = n4890 & ~n8198 ;
  assign n27414 = ( ~n3948 & n4069 ) | ( ~n3948 & n27413 ) | ( n4069 & n27413 ) ;
  assign n27415 = n26280 ^ n8260 ^ 1'b0 ;
  assign n27416 = ( n13762 & n27414 ) | ( n13762 & n27415 ) | ( n27414 & n27415 ) ;
  assign n27417 = n801 ^ n753 ^ 1'b0 ;
  assign n27418 = ( n14151 & ~n17768 ) | ( n14151 & n20426 ) | ( ~n17768 & n20426 ) ;
  assign n27419 = n7537 & ~n25394 ;
  assign n27420 = n20609 & n27419 ;
  assign n27421 = n20641 ^ n16136 ^ n6573 ;
  assign n27422 = n27421 ^ n11625 ^ 1'b0 ;
  assign n27423 = n6672 & n18885 ;
  assign n27424 = n2569 & ~n18813 ;
  assign n27425 = n27424 ^ n15378 ^ n1591 ;
  assign n27426 = ( n2400 & ~n6474 ) | ( n2400 & n9841 ) | ( ~n6474 & n9841 ) ;
  assign n27427 = ( n11140 & n17192 ) | ( n11140 & n23009 ) | ( n17192 & n23009 ) ;
  assign n27428 = ( n1583 & ~n3094 ) | ( n1583 & n5444 ) | ( ~n3094 & n5444 ) ;
  assign n27429 = n27428 ^ n16020 ^ 1'b0 ;
  assign n27430 = ~n7198 & n27429 ;
  assign n27431 = n7884 & ~n8973 ;
  assign n27432 = ~n5707 & n27431 ;
  assign n27433 = n4914 & ~n20686 ;
  assign n27434 = n24185 & n27433 ;
  assign n27435 = n22024 & n27434 ;
  assign n27436 = n12343 ^ n11199 ^ n7493 ;
  assign n27437 = n25364 & ~n27436 ;
  assign n27438 = n488 & n18881 ;
  assign n27439 = ( ~n23555 & n24790 ) | ( ~n23555 & n27438 ) | ( n24790 & n27438 ) ;
  assign n27440 = n18612 ^ n8214 ^ n6104 ;
  assign n27441 = n15282 ^ n7913 ^ 1'b0 ;
  assign n27442 = n9490 | n27441 ;
  assign n27443 = n27442 ^ n12612 ^ n10190 ;
  assign n27444 = n4156 ^ n3053 ^ n3036 ;
  assign n27445 = n27444 ^ n8571 ^ n3820 ;
  assign n27446 = n27445 ^ n14446 ^ n4742 ;
  assign n27447 = n27446 ^ n23459 ^ n6018 ;
  assign n27448 = ~n18373 & n19447 ;
  assign n27449 = ~n798 & n27448 ;
  assign n27450 = n4830 | n17906 ;
  assign n27451 = n4832 & ~n27450 ;
  assign n27452 = n9544 ^ n8972 ^ 1'b0 ;
  assign n27453 = ( n18393 & n18957 ) | ( n18393 & ~n27452 ) | ( n18957 & ~n27452 ) ;
  assign n27454 = n27453 ^ n2008 ^ 1'b0 ;
  assign n27455 = n1955 & n27454 ;
  assign n27456 = n15726 ^ n4888 ^ 1'b0 ;
  assign n27457 = x117 & ~n27456 ;
  assign n27458 = ( n1487 & n24001 ) | ( n1487 & ~n27457 ) | ( n24001 & ~n27457 ) ;
  assign n27459 = n10824 ^ n10720 ^ n10466 ;
  assign n27460 = n27459 ^ n22667 ^ n4078 ;
  assign n27461 = n3489 ^ n2936 ^ n2825 ;
  assign n27462 = n27461 ^ n8756 ^ n2823 ;
  assign n27463 = n27462 ^ n23614 ^ n9826 ;
  assign n27464 = n23545 ^ n20089 ^ 1'b0 ;
  assign n27465 = n6073 | n27464 ;
  assign n27466 = ( n3746 & ~n15777 ) | ( n3746 & n19402 ) | ( ~n15777 & n19402 ) ;
  assign n27467 = n22685 ^ n8588 ^ n4348 ;
  assign n27468 = n13296 ^ n11637 ^ 1'b0 ;
  assign n27469 = ( n3376 & n27467 ) | ( n3376 & ~n27468 ) | ( n27467 & ~n27468 ) ;
  assign n27471 = ~n4246 & n7112 ;
  assign n27472 = ~n3029 & n27471 ;
  assign n27473 = n27472 ^ n14501 ^ n13624 ;
  assign n27470 = ( n4007 & n8479 ) | ( n4007 & n21902 ) | ( n8479 & n21902 ) ;
  assign n27474 = n27473 ^ n27470 ^ n22475 ;
  assign n27475 = ~n14120 & n15836 ;
  assign n27476 = n6271 & n27475 ;
  assign n27477 = n6246 & ~n27476 ;
  assign n27478 = n3327 | n13522 ;
  assign n27479 = n3957 & ~n27478 ;
  assign n27480 = n27479 ^ n8292 ^ n7338 ;
  assign n27481 = ( n1568 & n9497 ) | ( n1568 & n19698 ) | ( n9497 & n19698 ) ;
  assign n27482 = n27481 ^ n23216 ^ n12615 ;
  assign n27484 = n1295 & ~n1444 ;
  assign n27485 = n27484 ^ n5022 ^ 1'b0 ;
  assign n27483 = n13398 | n26654 ;
  assign n27486 = n27485 ^ n27483 ^ 1'b0 ;
  assign n27487 = n13038 ^ n7290 ^ n1342 ;
  assign n27488 = n27487 ^ n6676 ^ 1'b0 ;
  assign n27492 = ( n371 & n4294 ) | ( n371 & ~n6446 ) | ( n4294 & ~n6446 ) ;
  assign n27489 = n12172 & ~n12699 ;
  assign n27490 = n27489 ^ n22936 ^ n1913 ;
  assign n27491 = n27183 & ~n27490 ;
  assign n27493 = n27492 ^ n27491 ^ 1'b0 ;
  assign n27494 = ( n11213 & n15237 ) | ( n11213 & ~n15885 ) | ( n15237 & ~n15885 ) ;
  assign n27495 = n25046 ^ n14290 ^ n883 ;
  assign n27496 = n4797 & ~n13473 ;
  assign n27497 = n7205 ^ n2851 ^ n2706 ;
  assign n27498 = n20237 ^ n17327 ^ 1'b0 ;
  assign n27499 = n11895 & ~n24633 ;
  assign n27500 = n18502 & n27499 ;
  assign n27501 = ( ~n27497 & n27498 ) | ( ~n27497 & n27500 ) | ( n27498 & n27500 ) ;
  assign n27502 = n2090 | n2514 ;
  assign n27503 = n12831 & ~n27502 ;
  assign n27504 = n16195 & ~n27503 ;
  assign n27505 = n1048 & ~n14983 ;
  assign n27506 = ( ~n5857 & n13143 ) | ( ~n5857 & n26050 ) | ( n13143 & n26050 ) ;
  assign n27507 = ( n11553 & n22768 ) | ( n11553 & n27506 ) | ( n22768 & n27506 ) ;
  assign n27508 = ( n3998 & ~n15823 ) | ( n3998 & n27507 ) | ( ~n15823 & n27507 ) ;
  assign n27509 = ( n1268 & ~n10858 ) | ( n1268 & n11718 ) | ( ~n10858 & n11718 ) ;
  assign n27510 = ~n8020 & n20230 ;
  assign n27511 = n27509 & ~n27510 ;
  assign n27512 = n3535 | n27511 ;
  assign n27513 = n195 | n27512 ;
  assign n27514 = n27513 ^ n26299 ^ n12760 ;
  assign n27515 = n12771 ^ n3573 ^ n293 ;
  assign n27516 = n15565 ^ n10713 ^ 1'b0 ;
  assign n27517 = n27515 & n27516 ;
  assign n27518 = n20462 ^ n2899 ^ 1'b0 ;
  assign n27519 = n27518 ^ n16495 ^ n7811 ;
  assign n27520 = n27517 & ~n27519 ;
  assign n27522 = n1532 & ~n17527 ;
  assign n27523 = n27522 ^ n3263 ^ 1'b0 ;
  assign n27524 = ~n26727 & n27523 ;
  assign n27525 = n27524 ^ n7610 ^ 1'b0 ;
  assign n27521 = ( n2530 & n21801 ) | ( n2530 & n22287 ) | ( n21801 & n22287 ) ;
  assign n27526 = n27525 ^ n27521 ^ 1'b0 ;
  assign n27527 = n24496 ^ x26 ^ 1'b0 ;
  assign n27528 = n4389 | n27527 ;
  assign n27529 = ~n2923 & n19036 ;
  assign n27530 = n21420 & n27529 ;
  assign n27531 = n17307 ^ n9708 ^ n4723 ;
  assign n27532 = n27531 ^ n11880 ^ n1032 ;
  assign n27533 = n27532 ^ n24496 ^ n2955 ;
  assign n27534 = n21750 ^ n5695 ^ n3673 ;
  assign n27535 = n21226 & n27534 ;
  assign n27536 = n140 & n10888 ;
  assign n27537 = n1399 & n20355 ;
  assign n27538 = n27537 ^ n4917 ^ 1'b0 ;
  assign n27539 = ~n17054 & n27538 ;
  assign n27540 = n27539 ^ n25727 ^ 1'b0 ;
  assign n27541 = ( n5539 & n20941 ) | ( n5539 & n27540 ) | ( n20941 & n27540 ) ;
  assign n27542 = ( n10413 & ~n16419 ) | ( n10413 & n20319 ) | ( ~n16419 & n20319 ) ;
  assign n27543 = n27542 ^ n26261 ^ n15845 ;
  assign n27544 = n21539 ^ n3368 ^ n2328 ;
  assign n27545 = n4879 ^ n218 ^ 1'b0 ;
  assign n27546 = n9306 & n27545 ;
  assign n27547 = n5563 | n12545 ;
  assign n27548 = n27547 ^ n11925 ^ 1'b0 ;
  assign n27549 = n27548 ^ n10139 ^ 1'b0 ;
  assign n27550 = n23985 | n27549 ;
  assign n27551 = n26138 ^ n23012 ^ 1'b0 ;
  assign n27552 = n20863 & ~n23338 ;
  assign n27553 = n27552 ^ n18866 ^ n16436 ;
  assign n27554 = n27553 ^ n14090 ^ 1'b0 ;
  assign n27555 = n7343 | n24587 ;
  assign n27556 = n16555 ^ n9760 ^ n7582 ;
  assign n27557 = n2774 & ~n15664 ;
  assign n27558 = n13981 & n27557 ;
  assign n27559 = n9941 | n27558 ;
  assign n27560 = n27556 & ~n27559 ;
  assign n27561 = n27560 ^ n7490 ^ 1'b0 ;
  assign n27562 = n26507 ^ n19028 ^ n9506 ;
  assign n27563 = n20982 ^ n19357 ^ n14695 ;
  assign n27566 = ~n13800 & n17169 ;
  assign n27564 = ( n5937 & ~n17479 ) | ( n5937 & n20412 ) | ( ~n17479 & n20412 ) ;
  assign n27565 = n19817 & ~n27564 ;
  assign n27567 = n27566 ^ n27565 ^ 1'b0 ;
  assign n27569 = ~n5058 & n15318 ;
  assign n27570 = n27569 ^ n8728 ^ 1'b0 ;
  assign n27568 = n2196 | n23446 ;
  assign n27571 = n27570 ^ n27568 ^ 1'b0 ;
  assign n27572 = ( n2963 & n11654 ) | ( n2963 & n12250 ) | ( n11654 & n12250 ) ;
  assign n27573 = n16244 ^ n3730 ^ 1'b0 ;
  assign n27574 = n4344 & ~n27573 ;
  assign n27575 = n27574 ^ n20512 ^ n14472 ;
  assign n27576 = n27575 ^ n22223 ^ n2852 ;
  assign n27577 = n17661 ^ n12730 ^ n10422 ;
  assign n27578 = n11756 ^ n9149 ^ n170 ;
  assign n27579 = n27578 ^ n10233 ^ 1'b0 ;
  assign n27580 = ~n3357 & n27579 ;
  assign n27581 = ~n6208 & n27580 ;
  assign n27582 = ( n1709 & ~n4976 ) | ( n1709 & n12546 ) | ( ~n4976 & n12546 ) ;
  assign n27583 = n6575 & n27582 ;
  assign n27584 = n15187 ^ n3677 ^ n1268 ;
  assign n27585 = n10424 ^ n6222 ^ n5623 ;
  assign n27586 = ( n15435 & n18049 ) | ( n15435 & ~n27585 ) | ( n18049 & ~n27585 ) ;
  assign n27587 = n19276 ^ n10280 ^ 1'b0 ;
  assign n27588 = ~n12903 & n27587 ;
  assign n27589 = n4267 & ~n14625 ;
  assign n27590 = n860 & ~n27589 ;
  assign n27591 = n6083 & ~n14656 ;
  assign n27592 = ~n6182 & n27591 ;
  assign n27593 = ( ~n6868 & n7746 ) | ( ~n6868 & n19263 ) | ( n7746 & n19263 ) ;
  assign n27594 = n27593 ^ n6162 ^ n4725 ;
  assign n27595 = n27592 | n27594 ;
  assign n27596 = n2695 & ~n4269 ;
  assign n27597 = ( n6071 & ~n18892 ) | ( n6071 & n27596 ) | ( ~n18892 & n27596 ) ;
  assign n27598 = ( n5734 & n7854 ) | ( n5734 & n27597 ) | ( n7854 & n27597 ) ;
  assign n27599 = n26289 ^ n1610 ^ 1'b0 ;
  assign n27600 = n15405 ^ n1339 ^ n959 ;
  assign n27601 = ( n11884 & n27599 ) | ( n11884 & ~n27600 ) | ( n27599 & ~n27600 ) ;
  assign n27602 = n8435 & n15730 ;
  assign n27603 = n27602 ^ n20412 ^ 1'b0 ;
  assign n27604 = n27603 ^ n6396 ^ n2892 ;
  assign n27605 = ( ~n1044 & n1291 ) | ( ~n1044 & n1738 ) | ( n1291 & n1738 ) ;
  assign n27606 = n23388 ^ n14874 ^ n6664 ;
  assign n27607 = ( n9559 & ~n27605 ) | ( n9559 & n27606 ) | ( ~n27605 & n27606 ) ;
  assign n27608 = n10381 ^ n5421 ^ 1'b0 ;
  assign n27609 = n6271 | n27608 ;
  assign n27610 = n16252 ^ n12730 ^ n10484 ;
  assign n27611 = ( n16911 & n27609 ) | ( n16911 & n27610 ) | ( n27609 & n27610 ) ;
  assign n27612 = n27611 ^ n16515 ^ n8082 ;
  assign n27613 = n27612 ^ n10261 ^ n3283 ;
  assign n27614 = n10432 ^ n5390 ^ n3843 ;
  assign n27615 = n14198 & ~n27614 ;
  assign n27616 = n25374 & n27615 ;
  assign n27617 = n18522 ^ n15873 ^ 1'b0 ;
  assign n27618 = ~n27616 & n27617 ;
  assign n27619 = n19318 ^ n13924 ^ 1'b0 ;
  assign n27620 = n5180 & n27619 ;
  assign n27621 = ~n5160 & n27620 ;
  assign n27622 = n27621 ^ n8566 ^ 1'b0 ;
  assign n27623 = n4732 & n9641 ;
  assign n27624 = n1009 | n21654 ;
  assign n27625 = n27624 ^ n10104 ^ 1'b0 ;
  assign n27626 = n11247 ^ n6669 ^ 1'b0 ;
  assign n27627 = n16502 ^ n15775 ^ n4775 ;
  assign n27628 = n24574 ^ n17872 ^ n6407 ;
  assign n27629 = ( n5945 & n10959 ) | ( n5945 & ~n12901 ) | ( n10959 & ~n12901 ) ;
  assign n27630 = n27629 ^ n13996 ^ 1'b0 ;
  assign n27631 = ( n5385 & n18387 ) | ( n5385 & n27630 ) | ( n18387 & n27630 ) ;
  assign n27632 = n4622 & ~n13139 ;
  assign n27633 = n27632 ^ n17834 ^ 1'b0 ;
  assign n27634 = n27633 ^ n18763 ^ n5750 ;
  assign n27635 = n27634 ^ n18612 ^ n18266 ;
  assign n27637 = n11243 & n12583 ;
  assign n27638 = n2050 & n27637 ;
  assign n27636 = n14237 ^ n5289 ^ n3169 ;
  assign n27639 = n27638 ^ n27636 ^ n12980 ;
  assign n27640 = n27639 ^ n23279 ^ n646 ;
  assign n27641 = ( n12540 & n19293 ) | ( n12540 & ~n23728 ) | ( n19293 & ~n23728 ) ;
  assign n27642 = n27641 ^ n21454 ^ n1917 ;
  assign n27643 = n1468 & ~n16685 ;
  assign n27644 = ~n22383 & n27643 ;
  assign n27646 = ~n7487 & n11413 ;
  assign n27647 = n6179 & n27646 ;
  assign n27645 = n11624 & ~n11708 ;
  assign n27648 = n27647 ^ n27645 ^ 1'b0 ;
  assign n27649 = n25328 ^ n16214 ^ n16124 ;
  assign n27650 = ( n3902 & n20494 ) | ( n3902 & ~n23254 ) | ( n20494 & ~n23254 ) ;
  assign n27651 = n27650 ^ n24223 ^ n12384 ;
  assign n27652 = n24637 ^ n20865 ^ n7082 ;
  assign n27653 = ( n1101 & ~n12674 ) | ( n1101 & n16291 ) | ( ~n12674 & n16291 ) ;
  assign n27654 = n27472 ^ n14819 ^ 1'b0 ;
  assign n27655 = n4624 ^ n859 ^ 1'b0 ;
  assign n27659 = n3934 & n5981 ;
  assign n27660 = n12944 & n27659 ;
  assign n27656 = n6187 ^ n190 ^ 1'b0 ;
  assign n27657 = ( n5664 & ~n6466 ) | ( n5664 & n22907 ) | ( ~n6466 & n22907 ) ;
  assign n27658 = ( n5100 & ~n27656 ) | ( n5100 & n27657 ) | ( ~n27656 & n27657 ) ;
  assign n27661 = n27660 ^ n27658 ^ n26178 ;
  assign n27662 = ~n12914 & n22529 ;
  assign n27663 = n3014 ^ n1977 ^ 1'b0 ;
  assign n27665 = ( n3572 & n7813 ) | ( n3572 & ~n13908 ) | ( n7813 & ~n13908 ) ;
  assign n27664 = n17915 ^ n6773 ^ n5062 ;
  assign n27666 = n27665 ^ n27664 ^ n12762 ;
  assign n27667 = n27666 ^ n4789 ^ n3093 ;
  assign n27668 = n12118 ^ n10350 ^ n3779 ;
  assign n27669 = ( ~n14479 & n18443 ) | ( ~n14479 & n27668 ) | ( n18443 & n27668 ) ;
  assign n27670 = n27428 ^ n13942 ^ n7845 ;
  assign n27671 = n7678 ^ n5367 ^ n5315 ;
  assign n27672 = ( n2707 & n2733 ) | ( n2707 & ~n4175 ) | ( n2733 & ~n4175 ) ;
  assign n27673 = n27672 ^ n13956 ^ n13457 ;
  assign n27674 = ( n15336 & ~n18386 ) | ( n15336 & n22259 ) | ( ~n18386 & n22259 ) ;
  assign n27675 = n11970 ^ n7493 ^ n4264 ;
  assign n27676 = n27675 ^ n3494 ^ n2902 ;
  assign n27677 = ~n18905 & n27676 ;
  assign n27679 = n9701 ^ n9430 ^ n1501 ;
  assign n27680 = n27679 ^ n10903 ^ n7498 ;
  assign n27678 = n1301 | n1876 ;
  assign n27681 = n27680 ^ n27678 ^ 1'b0 ;
  assign n27682 = n27681 ^ n16634 ^ 1'b0 ;
  assign n27683 = n3730 | n27682 ;
  assign n27684 = n5740 ^ n1210 ^ 1'b0 ;
  assign n27685 = n27684 ^ n15791 ^ n5485 ;
  assign n27686 = n27685 ^ n11126 ^ 1'b0 ;
  assign n27687 = n23746 ^ n9389 ^ 1'b0 ;
  assign n27688 = n27687 ^ n14551 ^ x59 ;
  assign n27689 = n10575 ^ n10251 ^ n4422 ;
  assign n27690 = n27689 ^ n25513 ^ n21900 ;
  assign n27691 = ~n5462 & n7888 ;
  assign n27692 = n27691 ^ n7916 ^ 1'b0 ;
  assign n27693 = n11662 & ~n27692 ;
  assign n27694 = ( n4056 & n16861 ) | ( n4056 & n27693 ) | ( n16861 & n27693 ) ;
  assign n27695 = ~n1948 & n27694 ;
  assign n27696 = x74 & n4476 ;
  assign n27697 = n14373 & n27696 ;
  assign n27698 = n27697 ^ n9767 ^ n5569 ;
  assign n27699 = ~n4827 & n11586 ;
  assign n27700 = ( n8943 & n21130 ) | ( n8943 & n27699 ) | ( n21130 & n27699 ) ;
  assign n27701 = n5180 ^ n1971 ^ n1869 ;
  assign n27702 = n27701 ^ n10504 ^ n8030 ;
  assign n27703 = n1645 | n11629 ;
  assign n27704 = n12142 | n27703 ;
  assign n27705 = n4164 ^ n1706 ^ n525 ;
  assign n27706 = n27705 ^ n11486 ^ n1982 ;
  assign n27707 = n27706 ^ n10708 ^ n8539 ;
  assign n27708 = n26892 ^ n25129 ^ n9173 ;
  assign n27713 = n23844 ^ n21943 ^ 1'b0 ;
  assign n27711 = ( ~n4300 & n9863 ) | ( ~n4300 & n10566 ) | ( n9863 & n10566 ) ;
  assign n27712 = n27711 ^ n16538 ^ n7135 ;
  assign n27709 = n5922 ^ n840 ^ 1'b0 ;
  assign n27710 = n17755 | n27709 ;
  assign n27714 = n27713 ^ n27712 ^ n27710 ;
  assign n27715 = n26510 ^ n10397 ^ n538 ;
  assign n27716 = ( n7457 & n11112 ) | ( n7457 & n23265 ) | ( n11112 & n23265 ) ;
  assign n27717 = ( n3935 & n9084 ) | ( n3935 & ~n27716 ) | ( n9084 & ~n27716 ) ;
  assign n27718 = n2213 | n22184 ;
  assign n27719 = ( n10545 & n27717 ) | ( n10545 & n27718 ) | ( n27717 & n27718 ) ;
  assign n27720 = n22626 ^ n21711 ^ n15363 ;
  assign n27721 = n19116 ^ n16612 ^ n15610 ;
  assign n27722 = n27721 ^ n6832 ^ n4415 ;
  assign n27723 = n6208 & n27722 ;
  assign n27724 = ~n5444 & n27723 ;
  assign n27725 = n11781 & ~n14278 ;
  assign n27726 = n27725 ^ n21747 ^ 1'b0 ;
  assign n27727 = n13908 & ~n27726 ;
  assign n27729 = ( n300 & ~n2526 ) | ( n300 & n4354 ) | ( ~n2526 & n4354 ) ;
  assign n27730 = n27729 ^ n21654 ^ n12150 ;
  assign n27728 = ~n9411 & n13284 ;
  assign n27731 = n27730 ^ n27728 ^ 1'b0 ;
  assign n27732 = n22163 ^ n20513 ^ n4736 ;
  assign n27733 = n21701 ^ n19434 ^ n9600 ;
  assign n27734 = n26218 ^ n2216 ^ 1'b0 ;
  assign n27735 = ( n8223 & n27733 ) | ( n8223 & n27734 ) | ( n27733 & n27734 ) ;
  assign n27736 = ( ~n475 & n567 ) | ( ~n475 & n19126 ) | ( n567 & n19126 ) ;
  assign n27737 = n19799 ^ n3528 ^ n3428 ;
  assign n27741 = ( n342 & ~n3333 ) | ( n342 & n10436 ) | ( ~n3333 & n10436 ) ;
  assign n27738 = n17915 ^ n15847 ^ n10847 ;
  assign n27739 = n27738 ^ n17232 ^ 1'b0 ;
  assign n27740 = n18303 & ~n27739 ;
  assign n27742 = n27741 ^ n27740 ^ n9565 ;
  assign n27743 = n5906 | n27742 ;
  assign n27745 = ( n9678 & n15276 ) | ( n9678 & n20909 ) | ( n15276 & n20909 ) ;
  assign n27744 = n11044 | n18878 ;
  assign n27746 = n27745 ^ n27744 ^ 1'b0 ;
  assign n27747 = n1335 & n24798 ;
  assign n27748 = n27747 ^ n18739 ^ 1'b0 ;
  assign n27749 = n24233 ^ n9965 ^ n9942 ;
  assign n27750 = n27749 ^ n12545 ^ n10884 ;
  assign n27751 = ( n9167 & n11922 ) | ( n9167 & ~n12337 ) | ( n11922 & ~n12337 ) ;
  assign n27752 = n25884 ^ n18500 ^ n1925 ;
  assign n27753 = ( n6476 & n27751 ) | ( n6476 & ~n27752 ) | ( n27751 & ~n27752 ) ;
  assign n27754 = ( n3511 & ~n4850 ) | ( n3511 & n11163 ) | ( ~n4850 & n11163 ) ;
  assign n27755 = n25789 ^ n11051 ^ n6592 ;
  assign n27756 = n26306 ^ n25839 ^ n6103 ;
  assign n27757 = n21341 ^ n19117 ^ n12315 ;
  assign n27758 = n27757 ^ n22029 ^ n17917 ;
  assign n27764 = ( n2058 & ~n18068 ) | ( n2058 & n24822 ) | ( ~n18068 & n24822 ) ;
  assign n27760 = ( ~n811 & n4570 ) | ( ~n811 & n21590 ) | ( n4570 & n21590 ) ;
  assign n27761 = ( n2151 & ~n16166 ) | ( n2151 & n27760 ) | ( ~n16166 & n27760 ) ;
  assign n27759 = n8117 | n15439 ;
  assign n27762 = n27761 ^ n27759 ^ 1'b0 ;
  assign n27763 = n3615 & ~n27762 ;
  assign n27765 = n27764 ^ n27763 ^ 1'b0 ;
  assign n27766 = n15919 ^ n5647 ^ 1'b0 ;
  assign n27767 = ( n11859 & ~n12227 ) | ( n11859 & n16012 ) | ( ~n12227 & n16012 ) ;
  assign n27768 = ~n23326 & n27767 ;
  assign n27769 = n27768 ^ n5758 ^ 1'b0 ;
  assign n27770 = ~n2957 & n11365 ;
  assign n27771 = n27770 ^ n7741 ^ 1'b0 ;
  assign n27772 = n14077 ^ n3022 ^ 1'b0 ;
  assign n27773 = n21407 ^ n18691 ^ n18425 ;
  assign n27774 = n24889 ^ n17958 ^ n5215 ;
  assign n27775 = n27774 ^ n20967 ^ 1'b0 ;
  assign n27776 = ( n18797 & n27773 ) | ( n18797 & ~n27775 ) | ( n27773 & ~n27775 ) ;
  assign n27777 = n25941 ^ n4972 ^ 1'b0 ;
  assign n27778 = ( n7747 & n16936 ) | ( n7747 & ~n27777 ) | ( n16936 & ~n27777 ) ;
  assign n27779 = n3126 | n3796 ;
  assign n27780 = ( n8482 & n13886 ) | ( n8482 & n27779 ) | ( n13886 & n27779 ) ;
  assign n27781 = ( ~n19013 & n24680 ) | ( ~n19013 & n27780 ) | ( n24680 & n27780 ) ;
  assign n27782 = ~n13395 & n21244 ;
  assign n27783 = n9379 & n20340 ;
  assign n27784 = n27782 & n27783 ;
  assign n27785 = ( n12465 & ~n19277 ) | ( n12465 & n27784 ) | ( ~n19277 & n27784 ) ;
  assign n27788 = ~n199 & n14414 ;
  assign n27789 = ~n12755 & n27788 ;
  assign n27786 = n8667 | n17535 ;
  assign n27787 = n27786 ^ n545 ^ 1'b0 ;
  assign n27790 = n27789 ^ n27787 ^ 1'b0 ;
  assign n27791 = ~n6510 & n7100 ;
  assign n27792 = ~n15003 & n27791 ;
  assign n27793 = n14703 ^ n7182 ^ 1'b0 ;
  assign n27794 = n6218 & ~n27793 ;
  assign n27795 = n13557 ^ n11055 ^ 1'b0 ;
  assign n27796 = n12323 & ~n27795 ;
  assign n27798 = n6537 ^ n3681 ^ n1953 ;
  assign n27797 = ~n14177 & n17371 ;
  assign n27799 = n27798 ^ n27797 ^ 1'b0 ;
  assign n27800 = n14841 ^ n9021 ^ n6406 ;
  assign n27801 = n27800 ^ n15759 ^ n6128 ;
  assign n27802 = n21802 ^ n14423 ^ n3427 ;
  assign n27803 = ( ~x27 & n27801 ) | ( ~x27 & n27802 ) | ( n27801 & n27802 ) ;
  assign n27804 = ( n2832 & n4973 ) | ( n2832 & ~n21022 ) | ( n4973 & ~n21022 ) ;
  assign n27805 = ~n4342 & n20926 ;
  assign n27806 = ( ~n5928 & n9907 ) | ( ~n5928 & n14226 ) | ( n9907 & n14226 ) ;
  assign n27807 = n27806 ^ n24354 ^ n15184 ;
  assign n27808 = n27807 ^ n24208 ^ n3278 ;
  assign n27809 = ~n3184 & n4441 ;
  assign n27810 = ( n8931 & ~n21144 ) | ( n8931 & n27809 ) | ( ~n21144 & n27809 ) ;
  assign n27811 = ~n13038 & n27810 ;
  assign n27812 = ( n9323 & ~n25761 ) | ( n9323 & n27811 ) | ( ~n25761 & n27811 ) ;
  assign n27813 = n10439 ^ n4806 ^ 1'b0 ;
  assign n27814 = n20626 ^ n7358 ^ 1'b0 ;
  assign n27815 = n27814 ^ n22505 ^ 1'b0 ;
  assign n27816 = n4602 | n27815 ;
  assign n27817 = n16945 ^ n5731 ^ n2862 ;
  assign n27818 = n25599 ^ n8289 ^ n7953 ;
  assign n27819 = n3528 | n10176 ;
  assign n27820 = n27819 ^ n4229 ^ 1'b0 ;
  assign n27821 = n27820 ^ n20992 ^ n2301 ;
  assign n27822 = n4155 & ~n9261 ;
  assign n27823 = ( n6159 & n12594 ) | ( n6159 & n27822 ) | ( n12594 & n27822 ) ;
  assign n27824 = ~n23678 & n27823 ;
  assign n27825 = ( ~n459 & n9885 ) | ( ~n459 & n10305 ) | ( n9885 & n10305 ) ;
  assign n27826 = ( n11255 & ~n20240 ) | ( n11255 & n27825 ) | ( ~n20240 & n27825 ) ;
  assign n27827 = n23686 ^ n11443 ^ n8764 ;
  assign n27828 = n27827 ^ n22654 ^ n15479 ;
  assign n27829 = n3499 & n4046 ;
  assign n27830 = n27829 ^ n13031 ^ 1'b0 ;
  assign n27831 = n27830 ^ n12110 ^ n7651 ;
  assign n27832 = n21871 | n27831 ;
  assign n27833 = n4755 | n27832 ;
  assign n27834 = n10514 | n15824 ;
  assign n27835 = n15729 & ~n27834 ;
  assign n27836 = n27835 ^ n1562 ^ n812 ;
  assign n27837 = n18953 ^ n9812 ^ 1'b0 ;
  assign n27838 = ~n1967 & n27837 ;
  assign n27839 = n27838 ^ n15162 ^ n4067 ;
  assign n27840 = n21017 ^ n17943 ^ n9119 ;
  assign n27841 = n4209 & ~n15691 ;
  assign n27842 = ( n6963 & n10838 ) | ( n6963 & ~n27841 ) | ( n10838 & ~n27841 ) ;
  assign n27843 = n17020 & n27842 ;
  assign n27844 = n27843 ^ n26966 ^ n7169 ;
  assign n27845 = n12215 ^ n8833 ^ n1910 ;
  assign n27846 = n26924 ^ n11764 ^ 1'b0 ;
  assign n27847 = n18389 & n27846 ;
  assign n27848 = n18885 & n27847 ;
  assign n27849 = ( n11339 & n11355 ) | ( n11339 & n22742 ) | ( n11355 & n22742 ) ;
  assign n27850 = n12594 ^ n8676 ^ 1'b0 ;
  assign n27851 = ( ~n16171 & n17179 ) | ( ~n16171 & n25653 ) | ( n17179 & n25653 ) ;
  assign n27852 = ( n27388 & ~n27850 ) | ( n27388 & n27851 ) | ( ~n27850 & n27851 ) ;
  assign n27853 = n2504 & n3324 ;
  assign n27854 = ~n1857 & n27853 ;
  assign n27855 = n27854 ^ x123 ^ 1'b0 ;
  assign n27856 = n22395 ^ n15387 ^ n12149 ;
  assign n27857 = n11121 ^ n7780 ^ n5718 ;
  assign n27858 = ~n1467 & n2393 ;
  assign n27859 = n27858 ^ n21701 ^ 1'b0 ;
  assign n27860 = ( ~n1181 & n5800 ) | ( ~n1181 & n27859 ) | ( n5800 & n27859 ) ;
  assign n27861 = ( n9282 & n26180 ) | ( n9282 & ~n27213 ) | ( n26180 & ~n27213 ) ;
  assign n27862 = n23785 ^ n6216 ^ n2516 ;
  assign n27863 = n27861 & n27862 ;
  assign n27864 = n6399 | n23828 ;
  assign n27865 = n19259 ^ n6946 ^ 1'b0 ;
  assign n27866 = ~n5194 & n27865 ;
  assign n27867 = n27866 ^ n16451 ^ 1'b0 ;
  assign n27868 = n3898 & ~n15995 ;
  assign n27869 = n27868 ^ n18255 ^ 1'b0 ;
  assign n27870 = n20203 & ~n25587 ;
  assign n27871 = n27870 ^ n17651 ^ 1'b0 ;
  assign n27872 = ( n15508 & n25529 ) | ( n15508 & ~n27871 ) | ( n25529 & ~n27871 ) ;
  assign n27873 = ( ~n7157 & n10328 ) | ( ~n7157 & n26814 ) | ( n10328 & n26814 ) ;
  assign n27874 = n15016 ^ n4491 ^ 1'b0 ;
  assign n27875 = ( ~n745 & n12892 ) | ( ~n745 & n20380 ) | ( n12892 & n20380 ) ;
  assign n27876 = n27875 ^ n23639 ^ n745 ;
  assign n27877 = ( ~n857 & n23527 ) | ( ~n857 & n27876 ) | ( n23527 & n27876 ) ;
  assign n27878 = n6024 & ~n22708 ;
  assign n27879 = ~n27838 & n27878 ;
  assign n27880 = n27879 ^ n25552 ^ n9850 ;
  assign n27881 = ( n5978 & ~n8485 ) | ( n5978 & n25720 ) | ( ~n8485 & n25720 ) ;
  assign n27882 = n3364 ^ n1610 ^ 1'b0 ;
  assign n27883 = n27881 | n27882 ;
  assign n27884 = n1929 ^ n1454 ^ 1'b0 ;
  assign n27885 = ~n11794 & n27884 ;
  assign n27886 = n1888 & n21021 ;
  assign n27887 = n27886 ^ n10280 ^ 1'b0 ;
  assign n27888 = ( ~n2321 & n5765 ) | ( ~n2321 & n7792 ) | ( n5765 & n7792 ) ;
  assign n27889 = n9934 ^ n8503 ^ n551 ;
  assign n27890 = n901 | n3990 ;
  assign n27891 = n8531 & ~n27890 ;
  assign n27892 = n27891 ^ n669 ^ 1'b0 ;
  assign n27893 = ( n15216 & n25437 ) | ( n15216 & ~n27892 ) | ( n25437 & ~n27892 ) ;
  assign n27894 = n8756 | n14515 ;
  assign n27895 = ( n20351 & ~n27689 ) | ( n20351 & n27894 ) | ( ~n27689 & n27894 ) ;
  assign n27896 = ( ~n2823 & n7857 ) | ( ~n2823 & n9070 ) | ( n7857 & n9070 ) ;
  assign n27897 = n6558 & ~n27896 ;
  assign n27898 = ~n4642 & n10758 ;
  assign n27899 = ~n17108 & n17225 ;
  assign n27900 = n27898 & n27899 ;
  assign n27901 = n27900 ^ n21330 ^ n19293 ;
  assign n27902 = n21249 ^ n3835 ^ 1'b0 ;
  assign n27903 = n6295 & ~n27741 ;
  assign n27904 = ~n7994 & n27903 ;
  assign n27905 = ( n616 & n8076 ) | ( n616 & ~n11867 ) | ( n8076 & ~n11867 ) ;
  assign n27906 = n4361 & ~n4923 ;
  assign n27907 = ( n7103 & n8032 ) | ( n7103 & ~n27906 ) | ( n8032 & ~n27906 ) ;
  assign n27908 = n4622 & ~n4723 ;
  assign n27909 = n27908 ^ n27155 ^ 1'b0 ;
  assign n27910 = ( n6750 & n10651 ) | ( n6750 & ~n27909 ) | ( n10651 & ~n27909 ) ;
  assign n27911 = ( ~n8355 & n25154 ) | ( ~n8355 & n26581 ) | ( n25154 & n26581 ) ;
  assign n27912 = n10867 ^ n5086 ^ n1455 ;
  assign n27913 = n27912 ^ n13011 ^ n1425 ;
  assign n27914 = ( n5943 & n6859 ) | ( n5943 & ~n8967 ) | ( n6859 & ~n8967 ) ;
  assign n27915 = n7726 & n17566 ;
  assign n27916 = n7783 ^ n2271 ^ 1'b0 ;
  assign n27917 = n9641 | n27916 ;
  assign n27918 = ~n2005 & n22193 ;
  assign n27919 = n17807 & n27918 ;
  assign n27920 = n8425 ^ n7429 ^ 1'b0 ;
  assign n27921 = n5681 | n14921 ;
  assign n27922 = n27921 ^ n2140 ^ 1'b0 ;
  assign n27923 = ( n19561 & n23260 ) | ( n19561 & ~n25496 ) | ( n23260 & ~n25496 ) ;
  assign n27924 = n22586 ^ n15847 ^ n670 ;
  assign n27925 = n5415 ^ n4531 ^ n4529 ;
  assign n27926 = n27925 ^ n22693 ^ n12500 ;
  assign n27927 = n27926 ^ n12726 ^ 1'b0 ;
  assign n27928 = n3817 & ~n16385 ;
  assign n27929 = n27928 ^ n8450 ^ 1'b0 ;
  assign n27930 = n10565 & n27929 ;
  assign n27931 = n11819 & n27930 ;
  assign n27932 = n1635 & n23545 ;
  assign n27933 = n27932 ^ n13362 ^ 1'b0 ;
  assign n27934 = n9352 | n25804 ;
  assign n27935 = n27934 ^ n3712 ^ 1'b0 ;
  assign n27936 = ( n6464 & ~n13466 ) | ( n6464 & n27935 ) | ( ~n13466 & n27935 ) ;
  assign n27937 = n10391 ^ n4067 ^ n256 ;
  assign n27938 = ( n7280 & n27810 ) | ( n7280 & n27937 ) | ( n27810 & n27937 ) ;
  assign n27939 = ( ~n3069 & n9411 ) | ( ~n3069 & n9904 ) | ( n9411 & n9904 ) ;
  assign n27940 = n2404 | n3057 ;
  assign n27941 = ( n11419 & n27939 ) | ( n11419 & ~n27940 ) | ( n27939 & ~n27940 ) ;
  assign n27942 = n27941 ^ n21101 ^ n3559 ;
  assign n27943 = n26712 & n27814 ;
  assign n27944 = ( ~n4790 & n5501 ) | ( ~n4790 & n11232 ) | ( n5501 & n11232 ) ;
  assign n27947 = n23693 ^ n3399 ^ 1'b0 ;
  assign n27945 = n25721 ^ n19767 ^ n1535 ;
  assign n27946 = n27945 ^ n12678 ^ n3259 ;
  assign n27948 = n27947 ^ n27946 ^ n8153 ;
  assign n27949 = n5813 ^ n2457 ^ n1967 ;
  assign n27950 = n27949 ^ n19365 ^ 1'b0 ;
  assign n27953 = ( n407 & n1702 ) | ( n407 & ~n5462 ) | ( n1702 & ~n5462 ) ;
  assign n27951 = n3551 & n10161 ;
  assign n27952 = n27951 ^ n4866 ^ 1'b0 ;
  assign n27954 = n27953 ^ n27952 ^ n25957 ;
  assign n27958 = n27438 ^ n12366 ^ n1575 ;
  assign n27955 = n7647 ^ n2256 ^ 1'b0 ;
  assign n27956 = n5706 & n27955 ;
  assign n27957 = ( n7458 & ~n20331 ) | ( n7458 & n27956 ) | ( ~n20331 & n27956 ) ;
  assign n27959 = n27958 ^ n27957 ^ n26785 ;
  assign n27961 = n1550 & ~n8567 ;
  assign n27962 = ( n2935 & n3982 ) | ( n2935 & ~n27961 ) | ( n3982 & ~n27961 ) ;
  assign n27960 = ~n9999 & n23570 ;
  assign n27963 = n27962 ^ n27960 ^ 1'b0 ;
  assign n27964 = ( n17224 & n27146 ) | ( n17224 & n27963 ) | ( n27146 & n27963 ) ;
  assign n27965 = n5394 & n27808 ;
  assign n27966 = ~n6658 & n27965 ;
  assign n27968 = ( n9567 & n16595 ) | ( n9567 & n19433 ) | ( n16595 & n19433 ) ;
  assign n27969 = ~n7932 & n27968 ;
  assign n27967 = ~n426 & n8263 ;
  assign n27970 = n27969 ^ n27967 ^ 1'b0 ;
  assign n27972 = n2050 | n4544 ;
  assign n27973 = n27972 ^ n1261 ^ 1'b0 ;
  assign n27974 = n27973 ^ n24674 ^ n17558 ;
  assign n27971 = n8961 & n19747 ;
  assign n27975 = n27974 ^ n27971 ^ 1'b0 ;
  assign n27976 = ( n258 & ~n14679 ) | ( n258 & n17548 ) | ( ~n14679 & n17548 ) ;
  assign n27977 = n15928 ^ n4412 ^ 1'b0 ;
  assign n27978 = ( n894 & n6967 ) | ( n894 & ~n27977 ) | ( n6967 & ~n27977 ) ;
  assign n27979 = ( n11285 & n26831 ) | ( n11285 & n27978 ) | ( n26831 & n27978 ) ;
  assign n27980 = n2017 | n27979 ;
  assign n27981 = n27976 & ~n27980 ;
  assign n27982 = n4513 | n27981 ;
  assign n27983 = n27982 ^ n20723 ^ 1'b0 ;
  assign n27984 = ( ~n293 & n5947 ) | ( ~n293 & n9222 ) | ( n5947 & n9222 ) ;
  assign n27985 = ( n12612 & n25287 ) | ( n12612 & ~n27984 ) | ( n25287 & ~n27984 ) ;
  assign n27986 = ( x125 & n16441 ) | ( x125 & ~n27985 ) | ( n16441 & ~n27985 ) ;
  assign n27987 = ( n343 & n4670 ) | ( n343 & ~n27986 ) | ( n4670 & ~n27986 ) ;
  assign n27988 = n10405 ^ n7199 ^ 1'b0 ;
  assign n27989 = n12555 & n27988 ;
  assign n27990 = ( ~n411 & n25461 ) | ( ~n411 & n27989 ) | ( n25461 & n27989 ) ;
  assign n27991 = n7848 ^ n5943 ^ 1'b0 ;
  assign n27992 = ( ~n7152 & n15246 ) | ( ~n7152 & n27991 ) | ( n15246 & n27991 ) ;
  assign n27993 = ( n464 & ~n12583 ) | ( n464 & n27992 ) | ( ~n12583 & n27992 ) ;
  assign n27994 = ( n14260 & n20204 ) | ( n14260 & ~n22911 ) | ( n20204 & ~n22911 ) ;
  assign n27995 = n17618 ^ n4632 ^ 1'b0 ;
  assign n27996 = ( n7935 & n21016 ) | ( n7935 & ~n27995 ) | ( n21016 & ~n27995 ) ;
  assign n27997 = ~n7250 & n19681 ;
  assign n27998 = n6113 & n27997 ;
  assign n27999 = ( n3239 & n11605 ) | ( n3239 & n27998 ) | ( n11605 & n27998 ) ;
  assign n28000 = n27095 | n27999 ;
  assign n28001 = n668 & n2412 ;
  assign n28002 = ( ~n15727 & n15754 ) | ( ~n15727 & n21984 ) | ( n15754 & n21984 ) ;
  assign n28003 = n6760 & n28002 ;
  assign n28004 = ~n28001 & n28003 ;
  assign n28005 = n4996 & n6759 ;
  assign n28006 = n28005 ^ n5116 ^ 1'b0 ;
  assign n28007 = n12143 & ~n28006 ;
  assign n28008 = n14678 & n28007 ;
  assign n28009 = n7133 ^ n1266 ^ 1'b0 ;
  assign n28010 = ~n28008 & n28009 ;
  assign n28011 = n19671 ^ n12686 ^ 1'b0 ;
  assign n28012 = n2653 ^ n1349 ^ 1'b0 ;
  assign n28013 = n3382 & n28012 ;
  assign n28014 = ( n25561 & ~n26910 ) | ( n25561 & n28013 ) | ( ~n26910 & n28013 ) ;
  assign n28015 = ( n1626 & n11635 ) | ( n1626 & ~n21211 ) | ( n11635 & ~n21211 ) ;
  assign n28016 = n15361 ^ n5220 ^ 1'b0 ;
  assign n28017 = ( ~n10609 & n18703 ) | ( ~n10609 & n19798 ) | ( n18703 & n19798 ) ;
  assign n28018 = n20226 ^ n4145 ^ n517 ;
  assign n28019 = n12027 ^ n4894 ^ n3337 ;
  assign n28020 = n14160 ^ n9117 ^ 1'b0 ;
  assign n28021 = n13439 & ~n28020 ;
  assign n28022 = ( n15148 & n20426 ) | ( n15148 & ~n28021 ) | ( n20426 & ~n28021 ) ;
  assign n28023 = n13765 | n28022 ;
  assign n28024 = n7746 | n28023 ;
  assign n28025 = ~n8136 & n17426 ;
  assign n28026 = ~n11261 & n20870 ;
  assign n28030 = ( n3307 & ~n5477 ) | ( n3307 & n19196 ) | ( ~n5477 & n19196 ) ;
  assign n28031 = n28030 ^ n19439 ^ n13052 ;
  assign n28032 = x101 & ~n28031 ;
  assign n28027 = n638 | n14501 ;
  assign n28028 = n28027 ^ n12634 ^ 1'b0 ;
  assign n28029 = n17593 & ~n28028 ;
  assign n28033 = n28032 ^ n28029 ^ 1'b0 ;
  assign n28034 = n22700 ^ n16762 ^ 1'b0 ;
  assign n28035 = ( ~n4614 & n4926 ) | ( ~n4614 & n4980 ) | ( n4926 & n4980 ) ;
  assign n28036 = ( n7084 & ~n9911 ) | ( n7084 & n28035 ) | ( ~n9911 & n28035 ) ;
  assign n28037 = n28036 ^ n4197 ^ 1'b0 ;
  assign n28038 = ( n21391 & ~n27211 ) | ( n21391 & n28037 ) | ( ~n27211 & n28037 ) ;
  assign n28041 = n9508 ^ n9354 ^ n8469 ;
  assign n28039 = n7955 & ~n11807 ;
  assign n28040 = n28039 ^ n4931 ^ 1'b0 ;
  assign n28042 = n28041 ^ n28040 ^ n24740 ;
  assign n28043 = n22789 ^ n13641 ^ 1'b0 ;
  assign n28044 = n11528 ^ n11447 ^ n8057 ;
  assign n28045 = n3104 & n8939 ;
  assign n28046 = n28045 ^ n16650 ^ 1'b0 ;
  assign n28047 = ( n4019 & ~n8846 ) | ( n4019 & n28046 ) | ( ~n8846 & n28046 ) ;
  assign n28048 = n28047 ^ n10681 ^ n9593 ;
  assign n28049 = ( n261 & ~n6661 ) | ( n261 & n15206 ) | ( ~n6661 & n15206 ) ;
  assign n28050 = n8546 ^ n1644 ^ n591 ;
  assign n28051 = n28050 ^ n21453 ^ n6645 ;
  assign n28052 = ( n5699 & n22863 ) | ( n5699 & n24315 ) | ( n22863 & n24315 ) ;
  assign n28053 = ( n4209 & ~n19136 ) | ( n4209 & n28052 ) | ( ~n19136 & n28052 ) ;
  assign n28054 = ( n2412 & ~n28051 ) | ( n2412 & n28053 ) | ( ~n28051 & n28053 ) ;
  assign n28055 = n9405 | n19669 ;
  assign n28056 = n17718 & ~n28055 ;
  assign n28057 = n28056 ^ n11961 ^ n4202 ;
  assign n28058 = ( n28049 & n28054 ) | ( n28049 & ~n28057 ) | ( n28054 & ~n28057 ) ;
  assign n28059 = n21035 ^ n18964 ^ n9178 ;
  assign n28060 = ( ~n1441 & n23518 ) | ( ~n1441 & n28059 ) | ( n23518 & n28059 ) ;
  assign n28061 = n28060 ^ n15914 ^ 1'b0 ;
  assign n28062 = n20910 & ~n28061 ;
  assign n28065 = n25874 ^ n11260 ^ n490 ;
  assign n28063 = ( n3291 & n6868 ) | ( n3291 & n21558 ) | ( n6868 & n21558 ) ;
  assign n28064 = n2232 & ~n28063 ;
  assign n28066 = n28065 ^ n28064 ^ 1'b0 ;
  assign n28067 = n12369 ^ n5573 ^ 1'b0 ;
  assign n28068 = ~n25268 & n28067 ;
  assign n28069 = n2343 & ~n9546 ;
  assign n28070 = n28069 ^ n16867 ^ 1'b0 ;
  assign n28071 = n10010 | n28070 ;
  assign n28072 = ( x121 & n5259 ) | ( x121 & ~n17479 ) | ( n5259 & ~n17479 ) ;
  assign n28073 = ( ~n1460 & n18721 ) | ( ~n1460 & n21821 ) | ( n18721 & n21821 ) ;
  assign n28074 = ( ~n15749 & n15962 ) | ( ~n15749 & n19332 ) | ( n15962 & n19332 ) ;
  assign n28075 = n14566 ^ n13490 ^ 1'b0 ;
  assign n28076 = n19327 & ~n23169 ;
  assign n28077 = ~n28075 & n28076 ;
  assign n28078 = n24955 ^ n3286 ^ 1'b0 ;
  assign n28079 = n7193 & ~n28078 ;
  assign n28084 = n19597 ^ n7858 ^ 1'b0 ;
  assign n28082 = ( ~n2474 & n5236 ) | ( ~n2474 & n16253 ) | ( n5236 & n16253 ) ;
  assign n28083 = ( x52 & n1638 ) | ( x52 & n28082 ) | ( n1638 & n28082 ) ;
  assign n28080 = n8970 ^ n6158 ^ n1173 ;
  assign n28081 = n28080 ^ n10132 ^ n2031 ;
  assign n28085 = n28084 ^ n28083 ^ n28081 ;
  assign n28086 = n11512 ^ n11270 ^ n603 ;
  assign n28087 = n28086 ^ n16531 ^ n2847 ;
  assign n28088 = n973 & n1090 ;
  assign n28089 = n28088 ^ n3193 ^ 1'b0 ;
  assign n28094 = n8981 ^ n6239 ^ n6031 ;
  assign n28090 = n11090 ^ n10133 ^ 1'b0 ;
  assign n28091 = ~n3714 & n28090 ;
  assign n28092 = ( ~n10142 & n13391 ) | ( ~n10142 & n28091 ) | ( n13391 & n28091 ) ;
  assign n28093 = n28092 ^ n7923 ^ 1'b0 ;
  assign n28095 = n28094 ^ n28093 ^ n2930 ;
  assign n28096 = ( n12909 & n28089 ) | ( n12909 & ~n28095 ) | ( n28089 & ~n28095 ) ;
  assign n28097 = n17949 | n18880 ;
  assign n28098 = ~n8205 & n16838 ;
  assign n28099 = ( ~n11883 & n21571 ) | ( ~n11883 & n28098 ) | ( n21571 & n28098 ) ;
  assign n28100 = ( n5910 & n6531 ) | ( n5910 & n7104 ) | ( n6531 & n7104 ) ;
  assign n28101 = n18805 ^ n15726 ^ n6118 ;
  assign n28103 = n2907 | n19832 ;
  assign n28104 = n28103 ^ n26598 ^ 1'b0 ;
  assign n28102 = n16652 & ~n18321 ;
  assign n28105 = n28104 ^ n28102 ^ 1'b0 ;
  assign n28106 = n2412 & n20076 ;
  assign n28107 = n1884 & n28106 ;
  assign n28108 = n25237 & ~n28107 ;
  assign n28109 = n28105 & n28108 ;
  assign n28110 = n15046 & ~n18660 ;
  assign n28111 = n28110 ^ n4907 ^ 1'b0 ;
  assign n28112 = ~n24044 & n28111 ;
  assign n28113 = ~n5769 & n28112 ;
  assign n28114 = ( n4623 & n8730 ) | ( n4623 & ~n9550 ) | ( n8730 & ~n9550 ) ;
  assign n28115 = n11243 ^ n7690 ^ n320 ;
  assign n28116 = ( n4934 & n6599 ) | ( n4934 & ~n10364 ) | ( n6599 & ~n10364 ) ;
  assign n28117 = n12537 ^ n12385 ^ 1'b0 ;
  assign n28118 = n24293 | n28117 ;
  assign n28119 = ( ~n2891 & n28116 ) | ( ~n2891 & n28118 ) | ( n28116 & n28118 ) ;
  assign n28120 = ( n6537 & n13811 ) | ( n6537 & n22815 ) | ( n13811 & n22815 ) ;
  assign n28121 = n28120 ^ n22871 ^ n5046 ;
  assign n28122 = ~n4617 & n9309 ;
  assign n28126 = n2535 | n6598 ;
  assign n28127 = n7688 | n28126 ;
  assign n28123 = n5039 ^ n529 ^ 1'b0 ;
  assign n28124 = n8654 | n28123 ;
  assign n28125 = n28124 ^ n22285 ^ n5527 ;
  assign n28128 = n28127 ^ n28125 ^ 1'b0 ;
  assign n28129 = n7414 & ~n24563 ;
  assign n28130 = n28129 ^ n21467 ^ 1'b0 ;
  assign n28131 = n19746 ^ n4834 ^ 1'b0 ;
  assign n28132 = ~n27585 & n28131 ;
  assign n28133 = n9179 ^ n6054 ^ n1370 ;
  assign n28134 = n24283 | n26476 ;
  assign n28135 = n28134 ^ n21037 ^ 1'b0 ;
  assign n28136 = n20476 & ~n28135 ;
  assign n28137 = ~n28133 & n28136 ;
  assign n28138 = ~n280 & n18660 ;
  assign n28139 = n17272 ^ n13123 ^ n6657 ;
  assign n28140 = n28139 ^ n20252 ^ n18187 ;
  assign n28142 = ( n2653 & n3297 ) | ( n2653 & ~n7420 ) | ( n3297 & ~n7420 ) ;
  assign n28141 = n16210 ^ n13352 ^ n9776 ;
  assign n28143 = n28142 ^ n28141 ^ n9432 ;
  assign n28144 = ~n3229 & n13134 ;
  assign n28145 = ~n15873 & n28144 ;
  assign n28146 = n10462 ^ n6080 ^ 1'b0 ;
  assign n28147 = n25933 | n28146 ;
  assign n28148 = ( n24432 & ~n28145 ) | ( n24432 & n28147 ) | ( ~n28145 & n28147 ) ;
  assign n28149 = n28148 ^ n24515 ^ n2443 ;
  assign n28150 = n13786 ^ n9482 ^ 1'b0 ;
  assign n28151 = n18724 ^ n9682 ^ n2393 ;
  assign n28152 = ( ~n14078 & n22929 ) | ( ~n14078 & n28151 ) | ( n22929 & n28151 ) ;
  assign n28153 = n7178 & n21318 ;
  assign n28154 = n5987 | n13095 ;
  assign n28155 = n26603 & ~n28154 ;
  assign n28156 = ( n1703 & n8615 ) | ( n1703 & ~n11698 ) | ( n8615 & ~n11698 ) ;
  assign n28157 = n25943 ^ n13780 ^ 1'b0 ;
  assign n28158 = n28156 | n28157 ;
  assign n28159 = n12524 ^ n8210 ^ n3592 ;
  assign n28160 = n10612 ^ n3914 ^ n1421 ;
  assign n28161 = n271 & n28160 ;
  assign n28162 = ~n9896 & n28161 ;
  assign n28163 = n25369 & ~n28162 ;
  assign n28164 = ( n1157 & n5108 ) | ( n1157 & n26499 ) | ( n5108 & n26499 ) ;
  assign n28165 = n28164 ^ n18933 ^ n10627 ;
  assign n28166 = n25737 ^ n13506 ^ n5932 ;
  assign n28167 = ( n11597 & n12023 ) | ( n11597 & ~n24631 ) | ( n12023 & ~n24631 ) ;
  assign n28168 = n16402 & n28167 ;
  assign n28169 = n28168 ^ n3852 ^ 1'b0 ;
  assign n28170 = n28169 ^ n10966 ^ n7749 ;
  assign n28171 = n20436 ^ n6591 ^ n1421 ;
  assign n28172 = n13205 | n16171 ;
  assign n28173 = n28172 ^ n24824 ^ 1'b0 ;
  assign n28174 = n1913 & n6024 ;
  assign n28175 = n28174 ^ n12478 ^ 1'b0 ;
  assign n28176 = ( n10798 & n13429 ) | ( n10798 & n15276 ) | ( n13429 & n15276 ) ;
  assign n28177 = n28176 ^ n10822 ^ 1'b0 ;
  assign n28178 = n28175 & ~n28177 ;
  assign n28179 = n8220 & n15655 ;
  assign n28181 = ( ~n4797 & n5090 ) | ( ~n4797 & n23353 ) | ( n5090 & n23353 ) ;
  assign n28180 = n1787 & n8053 ;
  assign n28182 = n28181 ^ n28180 ^ 1'b0 ;
  assign n28183 = ( n7922 & ~n12498 ) | ( n7922 & n28182 ) | ( ~n12498 & n28182 ) ;
  assign n28184 = n28183 ^ n16470 ^ 1'b0 ;
  assign n28185 = n24457 | n28184 ;
  assign n28186 = n28185 ^ n27056 ^ n6215 ;
  assign n28187 = ( ~n1601 & n4110 ) | ( ~n1601 & n11258 ) | ( n4110 & n11258 ) ;
  assign n28188 = ( ~n9101 & n11062 ) | ( ~n9101 & n28187 ) | ( n11062 & n28187 ) ;
  assign n28189 = n10422 ^ n2323 ^ n583 ;
  assign n28190 = n8400 ^ n2370 ^ 1'b0 ;
  assign n28191 = ~n16494 & n28190 ;
  assign n28192 = ( n1759 & n2775 ) | ( n1759 & n28191 ) | ( n2775 & n28191 ) ;
  assign n28193 = n17917 ^ n9936 ^ n6293 ;
  assign n28194 = ( n4406 & ~n28192 ) | ( n4406 & n28193 ) | ( ~n28192 & n28193 ) ;
  assign n28195 = ( n8297 & n13554 ) | ( n8297 & ~n22672 ) | ( n13554 & ~n22672 ) ;
  assign n28196 = n10403 | n12218 ;
  assign n28197 = n12464 | n28196 ;
  assign n28198 = ( ~n4307 & n14812 ) | ( ~n4307 & n28197 ) | ( n14812 & n28197 ) ;
  assign n28199 = n18921 ^ n17251 ^ n14020 ;
  assign n28200 = ( n567 & ~n607 ) | ( n567 & n20061 ) | ( ~n607 & n20061 ) ;
  assign n28201 = n17610 & ~n28200 ;
  assign n28202 = n10652 ^ n2099 ^ 1'b0 ;
  assign n28203 = n28202 ^ n10460 ^ n6401 ;
  assign n28204 = ( n6330 & n8096 ) | ( n6330 & n11325 ) | ( n8096 & n11325 ) ;
  assign n28205 = n10545 ^ n6911 ^ n4652 ;
  assign n28206 = n3302 ^ n2280 ^ n387 ;
  assign n28207 = n3272 | n16849 ;
  assign n28208 = n28207 ^ n10619 ^ 1'b0 ;
  assign n28209 = n23827 ^ n15176 ^ n1109 ;
  assign n28210 = n9895 | n28209 ;
  assign n28211 = n9393 | n28210 ;
  assign n28212 = n5316 ^ n3089 ^ 1'b0 ;
  assign n28213 = n5986 & n28212 ;
  assign n28214 = ( n7091 & n15451 ) | ( n7091 & n20169 ) | ( n15451 & n20169 ) ;
  assign n28215 = ( ~n13485 & n14108 ) | ( ~n13485 & n14196 ) | ( n14108 & n14196 ) ;
  assign n28219 = n2630 & n3108 ;
  assign n28216 = n3065 & ~n5424 ;
  assign n28217 = n28216 ^ n6566 ^ 1'b0 ;
  assign n28218 = n13667 & n28217 ;
  assign n28220 = n28219 ^ n28218 ^ n22491 ;
  assign n28221 = n17278 ^ n13996 ^ n6529 ;
  assign n28222 = n13824 ^ n5249 ^ n2665 ;
  assign n28223 = n24697 ^ n10634 ^ n9019 ;
  assign n28224 = n14135 ^ n9107 ^ n3055 ;
  assign n28225 = n28224 ^ n21392 ^ 1'b0 ;
  assign n28226 = n13192 | n28225 ;
  assign n28227 = n28226 ^ n22439 ^ 1'b0 ;
  assign n28228 = n293 & n28227 ;
  assign n28229 = ~n896 & n12676 ;
  assign n28230 = n28229 ^ n8604 ^ 1'b0 ;
  assign n28240 = n20361 & ~n26700 ;
  assign n28231 = n8929 & n23919 ;
  assign n28232 = n28231 ^ n8393 ^ 1'b0 ;
  assign n28233 = n28232 ^ n13643 ^ 1'b0 ;
  assign n28234 = n555 | n954 ;
  assign n28235 = ( n10008 & n16887 ) | ( n10008 & n28234 ) | ( n16887 & n28234 ) ;
  assign n28236 = n17433 ^ n5049 ^ 1'b0 ;
  assign n28237 = ( n20076 & n28235 ) | ( n20076 & n28236 ) | ( n28235 & n28236 ) ;
  assign n28238 = ( ~n19310 & n28233 ) | ( ~n19310 & n28237 ) | ( n28233 & n28237 ) ;
  assign n28239 = ~n20294 & n28238 ;
  assign n28241 = n28240 ^ n28239 ^ 1'b0 ;
  assign n28242 = n21009 ^ n9344 ^ 1'b0 ;
  assign n28243 = n6402 ^ n4697 ^ n1692 ;
  assign n28244 = ( n7413 & ~n28063 ) | ( n7413 & n28243 ) | ( ~n28063 & n28243 ) ;
  assign n28245 = ( ~n10618 & n14203 ) | ( ~n10618 & n23181 ) | ( n14203 & n23181 ) ;
  assign n28246 = n867 | n20926 ;
  assign n28247 = n28246 ^ n19597 ^ n12595 ;
  assign n28248 = n28247 ^ n11537 ^ n7546 ;
  assign n28249 = n15164 ^ n2398 ^ n469 ;
  assign n28250 = ( n234 & ~n22644 ) | ( n234 & n28249 ) | ( ~n22644 & n28249 ) ;
  assign n28251 = n28250 ^ n2732 ^ 1'b0 ;
  assign n28252 = ~n19945 & n28251 ;
  assign n28253 = n8069 ^ n7173 ^ n870 ;
  assign n28254 = n12648 & n20535 ;
  assign n28255 = n28254 ^ n5000 ^ 1'b0 ;
  assign n28256 = ( n2077 & n12593 ) | ( n2077 & n28255 ) | ( n12593 & n28255 ) ;
  assign n28257 = ( n5124 & n12938 ) | ( n5124 & n22917 ) | ( n12938 & n22917 ) ;
  assign n28258 = n28257 ^ n6927 ^ n6905 ;
  assign n28259 = n1640 & n7937 ;
  assign n28260 = ~n541 & n28259 ;
  assign n28261 = n11886 | n21047 ;
  assign n28262 = n847 & ~n28261 ;
  assign n28263 = n28260 | n28262 ;
  assign n28264 = n11713 ^ n7748 ^ 1'b0 ;
  assign n28265 = ( ~n3515 & n7296 ) | ( ~n3515 & n16602 ) | ( n7296 & n16602 ) ;
  assign n28266 = ( n3569 & n12752 ) | ( n3569 & ~n22160 ) | ( n12752 & ~n22160 ) ;
  assign n28267 = ( n7317 & n28265 ) | ( n7317 & n28266 ) | ( n28265 & n28266 ) ;
  assign n28268 = n17795 ^ n2014 ^ 1'b0 ;
  assign n28269 = ( n661 & n14869 ) | ( n661 & ~n27182 ) | ( n14869 & ~n27182 ) ;
  assign n28270 = n10409 & ~n28269 ;
  assign n28271 = ~n6951 & n28270 ;
  assign n28272 = ~n729 & n3910 ;
  assign n28273 = n28272 ^ n1289 ^ 1'b0 ;
  assign n28274 = ( n3070 & ~n3697 ) | ( n3070 & n11789 ) | ( ~n3697 & n11789 ) ;
  assign n28275 = n28274 ^ n20452 ^ n18434 ;
  assign n28276 = ( n16063 & n28273 ) | ( n16063 & ~n28275 ) | ( n28273 & ~n28275 ) ;
  assign n28282 = n20811 ^ n9518 ^ 1'b0 ;
  assign n28283 = n158 | n28282 ;
  assign n28277 = ~n11853 & n16030 ;
  assign n28278 = n3747 & n12599 ;
  assign n28279 = n28278 ^ n7959 ^ 1'b0 ;
  assign n28280 = ( ~n4066 & n28277 ) | ( ~n4066 & n28279 ) | ( n28277 & n28279 ) ;
  assign n28281 = ( ~n4967 & n22513 ) | ( ~n4967 & n28280 ) | ( n22513 & n28280 ) ;
  assign n28284 = n28283 ^ n28281 ^ n1133 ;
  assign n28285 = n8780 ^ n3220 ^ 1'b0 ;
  assign n28286 = n19841 & n28285 ;
  assign n28287 = ( ~n3752 & n3794 ) | ( ~n3752 & n18686 ) | ( n3794 & n18686 ) ;
  assign n28288 = ( n18823 & ~n24932 ) | ( n18823 & n27697 ) | ( ~n24932 & n27697 ) ;
  assign n28289 = ( n23486 & n23739 ) | ( n23486 & n25534 ) | ( n23739 & n25534 ) ;
  assign n28290 = ( ~n6167 & n6458 ) | ( ~n6167 & n8342 ) | ( n6458 & n8342 ) ;
  assign n28291 = ( n5108 & n11686 ) | ( n5108 & n15677 ) | ( n11686 & n15677 ) ;
  assign n28292 = n28291 ^ n28083 ^ 1'b0 ;
  assign n28293 = n21046 & ~n28292 ;
  assign n28294 = n28293 ^ n6181 ^ n5999 ;
  assign n28295 = n28294 ^ n17259 ^ 1'b0 ;
  assign n28296 = ~n28290 & n28295 ;
  assign n28297 = n15981 & ~n23161 ;
  assign n28298 = ~n6120 & n14685 ;
  assign n28299 = n15507 & n28298 ;
  assign n28300 = ( n6737 & n8404 ) | ( n6737 & n28299 ) | ( n8404 & n28299 ) ;
  assign n28301 = n6277 & ~n28300 ;
  assign n28302 = n28301 ^ n7297 ^ 1'b0 ;
  assign n28303 = ( n9133 & ~n9612 ) | ( n9133 & n13309 ) | ( ~n9612 & n13309 ) ;
  assign n28304 = n24513 ^ n17002 ^ n9466 ;
  assign n28305 = n18107 & ~n20249 ;
  assign n28306 = ~n9998 & n28305 ;
  assign n28307 = ( ~n4389 & n5910 ) | ( ~n4389 & n28306 ) | ( n5910 & n28306 ) ;
  assign n28308 = n25008 ^ n6525 ^ n1720 ;
  assign n28309 = n15008 ^ n7986 ^ n1912 ;
  assign n28310 = n11797 & ~n22536 ;
  assign n28311 = n9832 & n28310 ;
  assign n28312 = ( n28308 & ~n28309 ) | ( n28308 & n28311 ) | ( ~n28309 & n28311 ) ;
  assign n28313 = n16544 ^ n9581 ^ 1'b0 ;
  assign n28314 = ~n16819 & n28313 ;
  assign n28315 = n12841 ^ n8253 ^ n5846 ;
  assign n28316 = ( ~n8050 & n28314 ) | ( ~n8050 & n28315 ) | ( n28314 & n28315 ) ;
  assign n28317 = n19686 ^ n9951 ^ 1'b0 ;
  assign n28318 = n1963 & n14762 ;
  assign n28319 = ~n28317 & n28318 ;
  assign n28320 = n28319 ^ n10057 ^ n671 ;
  assign n28321 = n8984 ^ n2209 ^ 1'b0 ;
  assign n28322 = ~n10270 & n28321 ;
  assign n28323 = n22876 ^ n9090 ^ 1'b0 ;
  assign n28324 = n28322 & ~n28323 ;
  assign n28325 = n8227 & ~n14785 ;
  assign n28326 = n28325 ^ n4954 ^ 1'b0 ;
  assign n28327 = n26496 ^ n23629 ^ 1'b0 ;
  assign n28328 = ~n28326 & n28327 ;
  assign n28329 = ~n5015 & n8486 ;
  assign n28330 = ~n9013 & n28329 ;
  assign n28331 = ( n2578 & ~n3133 ) | ( n2578 & n6416 ) | ( ~n3133 & n6416 ) ;
  assign n28332 = ~n28330 & n28331 ;
  assign n28333 = n4230 & n11734 ;
  assign n28334 = n28333 ^ n3983 ^ 1'b0 ;
  assign n28335 = n6749 | n28334 ;
  assign n28336 = n26208 & ~n28335 ;
  assign n28337 = n28336 ^ n12699 ^ n3946 ;
  assign n28338 = n25910 ^ n5604 ^ x18 ;
  assign n28339 = n12300 & ~n28338 ;
  assign n28340 = n508 | n15949 ;
  assign n28341 = n5559 | n7161 ;
  assign n28342 = n2636 ^ n2483 ^ n2249 ;
  assign n28343 = n28342 ^ n5391 ^ x35 ;
  assign n28344 = n28343 ^ n26606 ^ n6714 ;
  assign n28345 = ( n12010 & n24338 ) | ( n12010 & ~n28344 ) | ( n24338 & ~n28344 ) ;
  assign n28346 = n28341 & n28345 ;
  assign n28347 = ~n1755 & n2278 ;
  assign n28348 = n15741 & n28347 ;
  assign n28349 = n28348 ^ n19944 ^ n15040 ;
  assign n28350 = n6946 ^ n1893 ^ n342 ;
  assign n28351 = n14481 | n22881 ;
  assign n28352 = n16209 | n28351 ;
  assign n28353 = n1061 & n17178 ;
  assign n28354 = ( n3196 & n5778 ) | ( n3196 & ~n8243 ) | ( n5778 & ~n8243 ) ;
  assign n28355 = n28354 ^ n9460 ^ n8594 ;
  assign n28356 = n28355 ^ n8073 ^ n3279 ;
  assign n28357 = ( n8780 & n14839 ) | ( n8780 & n19275 ) | ( n14839 & n19275 ) ;
  assign n28359 = n597 & n12648 ;
  assign n28360 = n28359 ^ n6797 ^ 1'b0 ;
  assign n28358 = n14377 ^ n7279 ^ 1'b0 ;
  assign n28361 = n28360 ^ n28358 ^ n24320 ;
  assign n28362 = ( n3104 & n5865 ) | ( n3104 & ~n19853 ) | ( n5865 & ~n19853 ) ;
  assign n28363 = ( ~n1069 & n3074 ) | ( ~n1069 & n20221 ) | ( n3074 & n20221 ) ;
  assign n28364 = ( n1109 & ~n17332 ) | ( n1109 & n28363 ) | ( ~n17332 & n28363 ) ;
  assign n28365 = ( ~n2221 & n7301 ) | ( ~n2221 & n28083 ) | ( n7301 & n28083 ) ;
  assign n28370 = n2882 ^ n1738 ^ 1'b0 ;
  assign n28366 = n6661 ^ n3820 ^ 1'b0 ;
  assign n28367 = n6125 | n28366 ;
  assign n28368 = n28367 ^ n12697 ^ n12366 ;
  assign n28369 = ~n5937 & n28368 ;
  assign n28371 = n28370 ^ n28369 ^ 1'b0 ;
  assign n28372 = n2740 ^ n2176 ^ x102 ;
  assign n28373 = n28372 ^ n8139 ^ n4475 ;
  assign n28374 = ~n17243 & n28373 ;
  assign n28375 = n28374 ^ n26092 ^ 1'b0 ;
  assign n28376 = n16775 ^ n11878 ^ n2581 ;
  assign n28377 = n2876 ^ n2141 ^ n144 ;
  assign n28378 = ~n28376 & n28377 ;
  assign n28379 = ~n12409 & n28378 ;
  assign n28380 = n28379 ^ n24498 ^ 1'b0 ;
  assign n28381 = ( n3641 & n19062 ) | ( n3641 & n26931 ) | ( n19062 & n26931 ) ;
  assign n28382 = n8155 ^ n6973 ^ 1'b0 ;
  assign n28383 = n6467 & ~n28382 ;
  assign n28384 = ( n15161 & ~n22937 ) | ( n15161 & n28383 ) | ( ~n22937 & n28383 ) ;
  assign n28385 = ( ~n2920 & n14190 ) | ( ~n2920 & n23227 ) | ( n14190 & n23227 ) ;
  assign n28386 = ( n2286 & n3197 ) | ( n2286 & ~n17470 ) | ( n3197 & ~n17470 ) ;
  assign n28387 = n6381 ^ n4069 ^ n2706 ;
  assign n28388 = ( n5576 & n8658 ) | ( n5576 & n28387 ) | ( n8658 & n28387 ) ;
  assign n28389 = n28388 ^ n24367 ^ 1'b0 ;
  assign n28390 = ( n837 & n1697 ) | ( n837 & ~n4424 ) | ( n1697 & ~n4424 ) ;
  assign n28391 = ~n6107 & n28390 ;
  assign n28392 = n12461 | n15653 ;
  assign n28393 = n28392 ^ n14593 ^ 1'b0 ;
  assign n28394 = ( ~n2140 & n15237 ) | ( ~n2140 & n16808 ) | ( n15237 & n16808 ) ;
  assign n28395 = n1758 & n7928 ;
  assign n28396 = n23069 & n28395 ;
  assign n28397 = ( ~n14096 & n20517 ) | ( ~n14096 & n28396 ) | ( n20517 & n28396 ) ;
  assign n28398 = n16174 & ~n28397 ;
  assign n28399 = ( n6033 & n8718 ) | ( n6033 & n20413 ) | ( n8718 & n20413 ) ;
  assign n28400 = ( n137 & n7047 ) | ( n137 & n27896 ) | ( n7047 & n27896 ) ;
  assign n28401 = ( n2693 & n6895 ) | ( n2693 & n28400 ) | ( n6895 & n28400 ) ;
  assign n28402 = n27176 ^ n21223 ^ n17404 ;
  assign n28403 = n10750 ^ n9666 ^ n6678 ;
  assign n28404 = n20479 ^ n17930 ^ n9865 ;
  assign n28405 = n28404 ^ n23870 ^ n6215 ;
  assign n28406 = n3261 | n9786 ;
  assign n28407 = n8155 | n28406 ;
  assign n28408 = n14030 | n28407 ;
  assign n28409 = n5719 & n18549 ;
  assign n28410 = n16294 & n28409 ;
  assign n28411 = ~n20909 & n28410 ;
  assign n28413 = n23138 ^ n11270 ^ 1'b0 ;
  assign n28414 = n1375 | n28413 ;
  assign n28412 = ( n1143 & n1204 ) | ( n1143 & n7476 ) | ( n1204 & n7476 ) ;
  assign n28415 = n28414 ^ n28412 ^ n21667 ;
  assign n28416 = n434 | n15423 ;
  assign n28417 = n28416 ^ n6580 ^ 1'b0 ;
  assign n28418 = ( n3191 & n28415 ) | ( n3191 & ~n28417 ) | ( n28415 & ~n28417 ) ;
  assign n28419 = n16553 ^ n1395 ^ 1'b0 ;
  assign n28420 = n28419 ^ n7065 ^ n2941 ;
  assign n28421 = ( n7056 & n8935 ) | ( n7056 & n12885 ) | ( n8935 & n12885 ) ;
  assign n28422 = ~n9150 & n20754 ;
  assign n28423 = n8906 & n28422 ;
  assign n28424 = ( n384 & n18307 ) | ( n384 & n28423 ) | ( n18307 & n28423 ) ;
  assign n28425 = n21989 ^ n17529 ^ n7240 ;
  assign n28426 = n10518 & n21005 ;
  assign n28427 = ~n21005 & n28426 ;
  assign n28428 = n16567 | n18698 ;
  assign n28429 = ~n8283 & n27364 ;
  assign n28430 = n28429 ^ n17238 ^ n7351 ;
  assign n28431 = n28430 ^ n11761 ^ 1'b0 ;
  assign n28432 = ( n157 & n6805 ) | ( n157 & ~n25927 ) | ( n6805 & ~n25927 ) ;
  assign n28433 = n5341 ^ n1336 ^ 1'b0 ;
  assign n28434 = ( n26162 & n27428 ) | ( n26162 & n28433 ) | ( n27428 & n28433 ) ;
  assign n28435 = n9941 ^ n4035 ^ n3118 ;
  assign n28436 = ( n10533 & ~n19835 ) | ( n10533 & n28435 ) | ( ~n19835 & n28435 ) ;
  assign n28437 = ( n28432 & ~n28434 ) | ( n28432 & n28436 ) | ( ~n28434 & n28436 ) ;
  assign n28438 = ~n7824 & n20860 ;
  assign n28439 = ( n4730 & n9040 ) | ( n4730 & n15012 ) | ( n9040 & n15012 ) ;
  assign n28440 = ( n1833 & n3556 ) | ( n1833 & ~n26297 ) | ( n3556 & ~n26297 ) ;
  assign n28442 = n21053 ^ n9712 ^ 1'b0 ;
  assign n28443 = ~n25461 & n28442 ;
  assign n28441 = n18347 ^ n15322 ^ 1'b0 ;
  assign n28444 = n28443 ^ n28441 ^ n24518 ;
  assign n28445 = n2759 | n18618 ;
  assign n28446 = ( n3615 & n5293 ) | ( n3615 & ~n7531 ) | ( n5293 & ~n7531 ) ;
  assign n28447 = ( n1442 & ~n3186 ) | ( n1442 & n28446 ) | ( ~n3186 & n28446 ) ;
  assign n28449 = ( n4654 & n12896 ) | ( n4654 & n17156 ) | ( n12896 & n17156 ) ;
  assign n28450 = n28449 ^ n9216 ^ n1330 ;
  assign n28448 = n21165 & ~n22453 ;
  assign n28451 = n28450 ^ n28448 ^ 1'b0 ;
  assign n28452 = n13076 & n15006 ;
  assign n28453 = n3092 & ~n12393 ;
  assign n28454 = ( n1575 & n12483 ) | ( n1575 & ~n28453 ) | ( n12483 & ~n28453 ) ;
  assign n28455 = n28454 ^ n11501 ^ n8131 ;
  assign n28457 = n9854 ^ n4862 ^ n1217 ;
  assign n28456 = ( n4275 & ~n13867 ) | ( n4275 & n15778 ) | ( ~n13867 & n15778 ) ;
  assign n28458 = n28457 ^ n28456 ^ n19576 ;
  assign n28459 = n13973 & ~n15549 ;
  assign n28460 = ( n234 & n15962 ) | ( n234 & n16494 ) | ( n15962 & n16494 ) ;
  assign n28461 = n18720 ^ n11128 ^ n8284 ;
  assign n28462 = n13932 ^ n7564 ^ n1335 ;
  assign n28463 = ~n28461 & n28462 ;
  assign n28464 = n23449 ^ n14885 ^ 1'b0 ;
  assign n28467 = n1798 & ~n10826 ;
  assign n28466 = n12546 ^ n2988 ^ n2008 ;
  assign n28465 = ( x44 & n12314 ) | ( x44 & n23638 ) | ( n12314 & n23638 ) ;
  assign n28468 = n28467 ^ n28466 ^ n28465 ;
  assign n28469 = ( ~n17305 & n28464 ) | ( ~n17305 & n28468 ) | ( n28464 & n28468 ) ;
  assign n28470 = ( n7661 & n9162 ) | ( n7661 & ~n10524 ) | ( n9162 & ~n10524 ) ;
  assign n28471 = n10084 & n25789 ;
  assign n28472 = n3336 & n28471 ;
  assign n28473 = n8660 | n27177 ;
  assign n28474 = n28472 & ~n28473 ;
  assign n28475 = n13881 & ~n20131 ;
  assign n28476 = n2870 | n25272 ;
  assign n28477 = n698 | n28476 ;
  assign n28478 = n20120 & n28477 ;
  assign n28479 = n10572 | n28478 ;
  assign n28480 = n28479 ^ n13881 ^ 1'b0 ;
  assign n28481 = n1349 & n11525 ;
  assign n28482 = n2949 | n10711 ;
  assign n28483 = n4933 & ~n28482 ;
  assign n28484 = n6983 ^ n6057 ^ n1247 ;
  assign n28485 = n28484 ^ n12024 ^ n499 ;
  assign n28486 = ( n4687 & n12928 ) | ( n4687 & n28485 ) | ( n12928 & n28485 ) ;
  assign n28487 = ( ~n9565 & n28483 ) | ( ~n9565 & n28486 ) | ( n28483 & n28486 ) ;
  assign n28488 = ( n6327 & n7388 ) | ( n6327 & ~n15719 ) | ( n7388 & ~n15719 ) ;
  assign n28489 = ( n16415 & n20578 ) | ( n16415 & n28488 ) | ( n20578 & n28488 ) ;
  assign n28490 = ( n8488 & n17830 ) | ( n8488 & n26620 ) | ( n17830 & n26620 ) ;
  assign n28491 = ( n6020 & n8200 ) | ( n6020 & n9077 ) | ( n8200 & n9077 ) ;
  assign n28492 = n18015 & n19376 ;
  assign n28493 = n28492 ^ n16738 ^ n1017 ;
  assign n28494 = n6736 & ~n20360 ;
  assign n28495 = n28494 ^ n19551 ^ 1'b0 ;
  assign n28496 = ( ~n9908 & n16404 ) | ( ~n9908 & n28495 ) | ( n16404 & n28495 ) ;
  assign n28497 = n27556 ^ n3440 ^ 1'b0 ;
  assign n28498 = n4199 & n28497 ;
  assign n28499 = n21372 & n28498 ;
  assign n28500 = n28499 ^ n413 ^ 1'b0 ;
  assign n28501 = n3809 | n28500 ;
  assign n28502 = n25090 ^ n20750 ^ n7998 ;
  assign n28503 = n4524 & ~n5127 ;
  assign n28504 = n28502 & n28503 ;
  assign n28505 = ( n7638 & n10419 ) | ( n7638 & ~n20320 ) | ( n10419 & ~n20320 ) ;
  assign n28506 = ( n889 & n9813 ) | ( n889 & ~n21232 ) | ( n9813 & ~n21232 ) ;
  assign n28507 = n23420 ^ n14964 ^ n13371 ;
  assign n28508 = ( n1136 & ~n25266 ) | ( n1136 & n28507 ) | ( ~n25266 & n28507 ) ;
  assign n28509 = ( n7386 & n28506 ) | ( n7386 & ~n28508 ) | ( n28506 & ~n28508 ) ;
  assign n28510 = ~n16527 & n28509 ;
  assign n28512 = n15504 ^ n9370 ^ n2228 ;
  assign n28511 = ( ~n4062 & n11390 ) | ( ~n4062 & n12393 ) | ( n11390 & n12393 ) ;
  assign n28513 = n28512 ^ n28511 ^ 1'b0 ;
  assign n28514 = n28513 ^ n19357 ^ 1'b0 ;
  assign n28515 = n22638 ^ n18155 ^ n9178 ;
  assign n28516 = n25504 ^ n5114 ^ 1'b0 ;
  assign n28517 = ( ~n3511 & n5836 ) | ( ~n3511 & n28516 ) | ( n5836 & n28516 ) ;
  assign n28518 = n3732 ^ n1285 ^ n716 ;
  assign n28519 = n5697 & ~n18230 ;
  assign n28520 = ~n28518 & n28519 ;
  assign n28521 = n9693 & ~n14346 ;
  assign n28522 = n28521 ^ n21331 ^ n1151 ;
  assign n28523 = n9099 & n9972 ;
  assign n28524 = ( ~n4663 & n13073 ) | ( ~n4663 & n28523 ) | ( n13073 & n28523 ) ;
  assign n28525 = n28524 ^ n4655 ^ 1'b0 ;
  assign n28526 = ( n5412 & ~n15778 ) | ( n5412 & n28525 ) | ( ~n15778 & n28525 ) ;
  assign n28527 = n7685 & n13567 ;
  assign n28528 = n4862 & n28527 ;
  assign n28529 = n28528 ^ n7364 ^ n6302 ;
  assign n28530 = n3314 ^ n1503 ^ n1031 ;
  assign n28531 = ( n8216 & ~n8402 ) | ( n8216 & n28530 ) | ( ~n8402 & n28530 ) ;
  assign n28532 = n1282 | n28531 ;
  assign n28533 = n28529 & ~n28532 ;
  assign n28534 = n28533 ^ n25879 ^ n10066 ;
  assign n28535 = n10177 ^ n9046 ^ 1'b0 ;
  assign n28536 = ~n23504 & n28535 ;
  assign n28537 = ( n12644 & ~n16812 ) | ( n12644 & n28536 ) | ( ~n16812 & n28536 ) ;
  assign n28538 = ( ~n3935 & n21331 ) | ( ~n3935 & n28537 ) | ( n21331 & n28537 ) ;
  assign n28539 = ( ~n1601 & n5970 ) | ( ~n1601 & n14937 ) | ( n5970 & n14937 ) ;
  assign n28540 = n18756 ^ n8889 ^ n2575 ;
  assign n28541 = ( n2246 & ~n28539 ) | ( n2246 & n28540 ) | ( ~n28539 & n28540 ) ;
  assign n28542 = n14109 ^ n10777 ^ n7756 ;
  assign n28543 = n28542 ^ n21697 ^ 1'b0 ;
  assign n28544 = n14104 & ~n28543 ;
  assign n28545 = n6023 & ~n28544 ;
  assign n28546 = n28461 ^ n27835 ^ n6476 ;
  assign n28547 = n11602 & n26523 ;
  assign n28548 = n28546 & n28547 ;
  assign n28549 = n23725 ^ n23015 ^ n4919 ;
  assign n28550 = n28549 ^ n18522 ^ n17531 ;
  assign n28551 = ~n11402 & n13976 ;
  assign n28552 = n24918 & n28551 ;
  assign n28553 = ( n3559 & ~n10559 ) | ( n3559 & n28552 ) | ( ~n10559 & n28552 ) ;
  assign n28554 = n15766 ^ n14649 ^ 1'b0 ;
  assign n28555 = n3022 ^ n301 ^ 1'b0 ;
  assign n28556 = ( ~n2803 & n10131 ) | ( ~n2803 & n28555 ) | ( n10131 & n28555 ) ;
  assign n28557 = ( n7003 & ~n8731 ) | ( n7003 & n28556 ) | ( ~n8731 & n28556 ) ;
  assign n28558 = n9478 & ~n14584 ;
  assign n28559 = n28558 ^ n14435 ^ n933 ;
  assign n28561 = n6086 & n15170 ;
  assign n28560 = n19116 ^ n8939 ^ 1'b0 ;
  assign n28562 = n28561 ^ n28560 ^ n9218 ;
  assign n28563 = n21837 ^ n6845 ^ n5421 ;
  assign n28564 = ( n8861 & n16676 ) | ( n8861 & n28563 ) | ( n16676 & n28563 ) ;
  assign n28565 = n28564 ^ n14193 ^ n3424 ;
  assign n28566 = n27301 ^ n4911 ^ 1'b0 ;
  assign n28567 = ~n22097 & n22678 ;
  assign n28568 = ~n9651 & n28567 ;
  assign n28569 = n7582 ^ n300 ^ 1'b0 ;
  assign n28571 = n14068 | n21256 ;
  assign n28572 = n1174 & ~n28571 ;
  assign n28570 = ( n18394 & n22693 ) | ( n18394 & ~n27473 ) | ( n22693 & ~n27473 ) ;
  assign n28573 = n28572 ^ n28570 ^ 1'b0 ;
  assign n28574 = ~n11292 & n19969 ;
  assign n28575 = n28574 ^ n3707 ^ n524 ;
  assign n28576 = n8961 ^ n2237 ^ 1'b0 ;
  assign n28577 = ( n2328 & n8891 ) | ( n2328 & n28576 ) | ( n8891 & n28576 ) ;
  assign n28578 = ( n24724 & n28575 ) | ( n24724 & n28577 ) | ( n28575 & n28577 ) ;
  assign n28579 = n6485 & n11529 ;
  assign n28580 = ~n7460 & n8830 ;
  assign n28581 = n28580 ^ n7169 ^ 1'b0 ;
  assign n28582 = n6751 | n26044 ;
  assign n28583 = n18981 | n28582 ;
  assign n28584 = n28583 ^ n7859 ^ n931 ;
  assign n28585 = n28584 ^ n10259 ^ 1'b0 ;
  assign n28586 = ~n2015 & n28585 ;
  assign n28587 = n2412 ^ n495 ^ 1'b0 ;
  assign n28588 = n28587 ^ n16229 ^ n214 ;
  assign n28589 = ~n10122 & n28588 ;
  assign n28590 = n24697 ^ n18972 ^ n7420 ;
  assign n28591 = n4521 ^ n3581 ^ 1'b0 ;
  assign n28592 = n28591 ^ n16272 ^ n1810 ;
  assign n28593 = n28592 ^ n13227 ^ n5199 ;
  assign n28594 = n22750 & n28593 ;
  assign n28595 = n3099 ^ n154 ^ 1'b0 ;
  assign n28596 = n28595 ^ n12326 ^ n5975 ;
  assign n28597 = n7067 | n16502 ;
  assign n28598 = n28597 ^ n21665 ^ 1'b0 ;
  assign n28599 = n6467 | n28598 ;
  assign n28602 = ( n14755 & ~n16781 ) | ( n14755 & n18378 ) | ( ~n16781 & n18378 ) ;
  assign n28603 = n15809 ^ n261 ^ 1'b0 ;
  assign n28604 = ~n28602 & n28603 ;
  assign n28600 = n12050 ^ n7474 ^ 1'b0 ;
  assign n28601 = n5784 | n28600 ;
  assign n28605 = n28604 ^ n28601 ^ n24920 ;
  assign n28606 = n18095 & ~n19784 ;
  assign n28607 = n15865 ^ n11823 ^ 1'b0 ;
  assign n28608 = ~n7911 & n28607 ;
  assign n28609 = n26315 ^ n16463 ^ n7697 ;
  assign n28610 = n28609 ^ n24325 ^ n10565 ;
  assign n28611 = ( ~n14359 & n14661 ) | ( ~n14359 & n28610 ) | ( n14661 & n28610 ) ;
  assign n28612 = n13129 ^ n12713 ^ n12489 ;
  assign n28613 = n28612 ^ n25291 ^ n2219 ;
  assign n28614 = n18902 ^ n17860 ^ 1'b0 ;
  assign n28615 = n21946 ^ n19032 ^ n7006 ;
  assign n28616 = ( n3905 & n5746 ) | ( n3905 & n11588 ) | ( n5746 & n11588 ) ;
  assign n28617 = n28616 ^ n23564 ^ n3285 ;
  assign n28618 = n26690 & n28617 ;
  assign n28619 = n10689 ^ n5183 ^ 1'b0 ;
  assign n28620 = n26098 | n28619 ;
  assign n28621 = n8097 & ~n28620 ;
  assign n28622 = n28621 ^ n10532 ^ 1'b0 ;
  assign n28623 = n26959 ^ n18613 ^ n277 ;
  assign n28624 = n2561 & n4436 ;
  assign n28625 = n28624 ^ n2491 ^ 1'b0 ;
  assign n28626 = n4044 & n28625 ;
  assign n28627 = ( n16164 & n24610 ) | ( n16164 & ~n28626 ) | ( n24610 & ~n28626 ) ;
  assign n28628 = n28627 ^ n22602 ^ x116 ;
  assign n28629 = n861 | n12646 ;
  assign n28630 = n28629 ^ n28625 ^ 1'b0 ;
  assign n28631 = ( n10761 & n28628 ) | ( n10761 & ~n28630 ) | ( n28628 & ~n28630 ) ;
  assign n28632 = n20436 ^ n11178 ^ 1'b0 ;
  assign n28633 = n28632 ^ n5725 ^ 1'b0 ;
  assign n28634 = ( ~n2675 & n3175 ) | ( ~n2675 & n19335 ) | ( n3175 & n19335 ) ;
  assign n28635 = ( n3617 & ~n7545 ) | ( n3617 & n10494 ) | ( ~n7545 & n10494 ) ;
  assign n28637 = n12594 ^ n8722 ^ 1'b0 ;
  assign n28636 = ( n15489 & n18903 ) | ( n15489 & ~n20251 ) | ( n18903 & ~n20251 ) ;
  assign n28638 = n28637 ^ n28636 ^ n4365 ;
  assign n28639 = ( ~n1959 & n28635 ) | ( ~n1959 & n28638 ) | ( n28635 & n28638 ) ;
  assign n28640 = n2689 & n23571 ;
  assign n28641 = ~n28539 & n28640 ;
  assign n28642 = ~n728 & n18619 ;
  assign n28643 = n28642 ^ n5131 ^ 1'b0 ;
  assign n28644 = ~n3340 & n4137 ;
  assign n28645 = n28643 & n28644 ;
  assign n28646 = n2676 | n21160 ;
  assign n28647 = n28646 ^ n16242 ^ 1'b0 ;
  assign n28649 = ( n7282 & ~n16293 ) | ( n7282 & n18702 ) | ( ~n16293 & n18702 ) ;
  assign n28648 = n5546 & n17670 ;
  assign n28650 = n28649 ^ n28648 ^ 1'b0 ;
  assign n28651 = n12126 ^ n6146 ^ n3428 ;
  assign n28652 = n8035 | n28651 ;
  assign n28653 = ( x67 & ~n16096 ) | ( x67 & n28652 ) | ( ~n16096 & n28652 ) ;
  assign n28654 = ( n3688 & n5413 ) | ( n3688 & ~n15359 ) | ( n5413 & ~n15359 ) ;
  assign n28655 = n5514 ^ n4028 ^ n2741 ;
  assign n28656 = ( n2706 & n28654 ) | ( n2706 & ~n28655 ) | ( n28654 & ~n28655 ) ;
  assign n28657 = ( n4383 & n8374 ) | ( n4383 & ~n12654 ) | ( n8374 & ~n12654 ) ;
  assign n28658 = n25057 ^ n21790 ^ n4836 ;
  assign n28659 = ( n5862 & n10805 ) | ( n5862 & n28658 ) | ( n10805 & n28658 ) ;
  assign n28660 = n676 & n19109 ;
  assign n28661 = n28660 ^ n12464 ^ 1'b0 ;
  assign n28662 = ( n2785 & n3196 ) | ( n2785 & ~n26382 ) | ( n3196 & ~n26382 ) ;
  assign n28663 = n28662 ^ n17518 ^ n14849 ;
  assign n28664 = ( n9559 & ~n12467 ) | ( n9559 & n28663 ) | ( ~n12467 & n28663 ) ;
  assign n28665 = ~n2777 & n5453 ;
  assign n28666 = ~n28664 & n28665 ;
  assign n28667 = n998 | n11938 ;
  assign n28668 = n28667 ^ n7634 ^ 1'b0 ;
  assign n28669 = n9928 ^ n8806 ^ n5589 ;
  assign n28670 = n28669 ^ n21272 ^ n12335 ;
  assign n28671 = ( ~n6762 & n6772 ) | ( ~n6762 & n9805 ) | ( n6772 & n9805 ) ;
  assign n28672 = n8218 | n15579 ;
  assign n28676 = n2373 ^ n170 ^ 1'b0 ;
  assign n28675 = ( n4489 & n8222 ) | ( n4489 & ~n17699 ) | ( n8222 & ~n17699 ) ;
  assign n28673 = ( ~n2306 & n9725 ) | ( ~n2306 & n10904 ) | ( n9725 & n10904 ) ;
  assign n28674 = n28673 ^ n8101 ^ n4444 ;
  assign n28677 = n28676 ^ n28675 ^ n28674 ;
  assign n28678 = n28677 ^ n8192 ^ n6499 ;
  assign n28679 = ( n3809 & n28672 ) | ( n3809 & ~n28678 ) | ( n28672 & ~n28678 ) ;
  assign n28681 = n4326 | n6492 ;
  assign n28680 = n18642 ^ n15993 ^ n10675 ;
  assign n28682 = n28681 ^ n28680 ^ n14116 ;
  assign n28683 = ( n4967 & n15720 ) | ( n4967 & ~n24999 ) | ( n15720 & ~n24999 ) ;
  assign n28684 = n28683 ^ n12588 ^ n235 ;
  assign n28685 = n22025 | n22128 ;
  assign n28686 = n12481 & n18913 ;
  assign n28687 = ~n7490 & n28686 ;
  assign n28688 = n3592 & n28687 ;
  assign n28689 = n18153 ^ n6895 ^ n1607 ;
  assign n28690 = n28689 ^ n23854 ^ n8868 ;
  assign n28691 = n19181 ^ n12674 ^ 1'b0 ;
  assign n28692 = n9640 & ~n28691 ;
  assign n28693 = n28692 ^ n19904 ^ n17442 ;
  assign n28694 = n2886 & ~n16789 ;
  assign n28695 = n28694 ^ n20446 ^ 1'b0 ;
  assign n28696 = n28695 ^ n18342 ^ n8978 ;
  assign n28697 = n10652 ^ n7765 ^ n5412 ;
  assign n28698 = n16417 | n28697 ;
  assign n28699 = n22665 ^ n8530 ^ 1'b0 ;
  assign n28700 = n2493 | n28699 ;
  assign n28701 = n28700 ^ n20169 ^ 1'b0 ;
  assign n28702 = n28701 ^ n4205 ^ n3983 ;
  assign n28703 = n6614 & ~n13002 ;
  assign n28704 = n28703 ^ n25941 ^ 1'b0 ;
  assign n28705 = n7113 | n9628 ;
  assign n28706 = n28705 ^ n17021 ^ 1'b0 ;
  assign n28707 = ( n952 & n25743 ) | ( n952 & n28635 ) | ( n25743 & n28635 ) ;
  assign n28708 = ( n14416 & n27116 ) | ( n14416 & n28707 ) | ( n27116 & n28707 ) ;
  assign n28709 = ~n16440 & n28708 ;
  assign n28710 = ( n7675 & n8279 ) | ( n7675 & ~n11900 ) | ( n8279 & ~n11900 ) ;
  assign n28711 = n25588 ^ n3767 ^ n1488 ;
  assign n28712 = ( n2388 & n4285 ) | ( n2388 & ~n11811 ) | ( n4285 & ~n11811 ) ;
  assign n28713 = n20174 ^ n14212 ^ n12763 ;
  assign n28714 = ( ~n5978 & n12320 ) | ( ~n5978 & n17340 ) | ( n12320 & n17340 ) ;
  assign n28715 = n4931 & ~n28714 ;
  assign n28716 = n28713 & n28715 ;
  assign n28717 = n14479 ^ n12565 ^ 1'b0 ;
  assign n28722 = n19749 ^ n5194 ^ 1'b0 ;
  assign n28723 = n21592 | n28722 ;
  assign n28718 = n8527 ^ n5316 ^ n359 ;
  assign n28719 = ( n13956 & n23564 ) | ( n13956 & ~n28718 ) | ( n23564 & ~n28718 ) ;
  assign n28720 = n9581 & ~n28719 ;
  assign n28721 = n13004 & ~n28720 ;
  assign n28724 = n28723 ^ n28721 ^ 1'b0 ;
  assign n28725 = n19854 ^ n11033 ^ n4914 ;
  assign n28726 = n28725 ^ n12598 ^ 1'b0 ;
  assign n28727 = n2799 & n28726 ;
  assign n28728 = ~n7915 & n12181 ;
  assign n28729 = ~n10935 & n28728 ;
  assign n28730 = n5535 & ~n28701 ;
  assign n28731 = n20545 ^ n9584 ^ n3195 ;
  assign n28732 = n17336 ^ n4168 ^ n1490 ;
  assign n28733 = ~n1867 & n13575 ;
  assign n28734 = n28733 ^ n4148 ^ 1'b0 ;
  assign n28735 = n18337 ^ n6364 ^ 1'b0 ;
  assign n28736 = ~n6928 & n24232 ;
  assign n28737 = ~n21097 & n28736 ;
  assign n28738 = n11133 & n28737 ;
  assign n28739 = n20228 & n24574 ;
  assign n28740 = n28739 ^ n24680 ^ 1'b0 ;
  assign n28741 = n12531 ^ n3888 ^ n466 ;
  assign n28742 = n28741 ^ n7125 ^ 1'b0 ;
  assign n28743 = n25221 ^ n16581 ^ 1'b0 ;
  assign n28744 = ~n7443 & n28743 ;
  assign n28745 = ~n23810 & n28744 ;
  assign n28746 = ( n204 & n6424 ) | ( n204 & n16444 ) | ( n6424 & n16444 ) ;
  assign n28747 = ( n19105 & ~n20561 ) | ( n19105 & n27634 ) | ( ~n20561 & n27634 ) ;
  assign n28748 = ( n5504 & ~n16783 ) | ( n5504 & n26045 ) | ( ~n16783 & n26045 ) ;
  assign n28749 = ( ~n981 & n18679 ) | ( ~n981 & n28748 ) | ( n18679 & n28748 ) ;
  assign n28750 = n4015 & n6552 ;
  assign n28751 = n7244 & ~n18666 ;
  assign n28752 = ~n1914 & n14417 ;
  assign n28753 = n28752 ^ n10718 ^ n9115 ;
  assign n28754 = n9582 | n10873 ;
  assign n28755 = n1587 & ~n28754 ;
  assign n28756 = n9408 ^ n2798 ^ 1'b0 ;
  assign n28757 = n20314 | n28756 ;
  assign n28758 = ( n19067 & n28755 ) | ( n19067 & ~n28757 ) | ( n28755 & ~n28757 ) ;
  assign n28759 = ~n4292 & n14931 ;
  assign n28760 = n2613 | n21734 ;
  assign n28761 = n10675 | n25340 ;
  assign n28762 = n9215 ^ n2094 ^ 1'b0 ;
  assign n28763 = n28762 ^ n1252 ^ 1'b0 ;
  assign n28764 = n5805 | n16819 ;
  assign n28765 = n28764 ^ n10526 ^ 1'b0 ;
  assign n28766 = n5689 & n18110 ;
  assign n28767 = ~n8690 & n28766 ;
  assign n28768 = n21663 ^ n19191 ^ n7584 ;
  assign n28769 = n18794 & ~n22049 ;
  assign n28770 = n28768 & n28769 ;
  assign n28771 = n28770 ^ n19776 ^ n6711 ;
  assign n28772 = n1148 & n7185 ;
  assign n28773 = ( n5586 & ~n13439 ) | ( n5586 & n28772 ) | ( ~n13439 & n28772 ) ;
  assign n28774 = x125 & ~n26640 ;
  assign n28776 = n4646 ^ n3776 ^ 1'b0 ;
  assign n28777 = ~n14464 & n28776 ;
  assign n28775 = n7884 ^ n4177 ^ 1'b0 ;
  assign n28778 = n28777 ^ n28775 ^ n9471 ;
  assign n28779 = ( ~x1 & n6865 ) | ( ~x1 & n28778 ) | ( n6865 & n28778 ) ;
  assign n28780 = n5271 ^ n3915 ^ 1'b0 ;
  assign n28781 = n15496 | n28780 ;
  assign n28782 = n6580 | n28781 ;
  assign n28783 = ( ~n8451 & n20419 ) | ( ~n8451 & n28782 ) | ( n20419 & n28782 ) ;
  assign n28784 = ~n2927 & n23585 ;
  assign n28785 = n28784 ^ n22814 ^ 1'b0 ;
  assign n28786 = ( n1490 & ~n4447 ) | ( n1490 & n7748 ) | ( ~n4447 & n7748 ) ;
  assign n28787 = ( n866 & ~n28785 ) | ( n866 & n28786 ) | ( ~n28785 & n28786 ) ;
  assign n28788 = ( ~n2140 & n3689 ) | ( ~n2140 & n10318 ) | ( n3689 & n10318 ) ;
  assign n28789 = ~n18728 & n28788 ;
  assign n28790 = n4210 ^ n3006 ^ 1'b0 ;
  assign n28791 = n1306 & n16216 ;
  assign n28792 = n28655 ^ n22463 ^ n12734 ;
  assign n28793 = n28792 ^ n7462 ^ n1060 ;
  assign n28794 = n28793 ^ n10339 ^ n1579 ;
  assign n28795 = n12524 ^ n8018 ^ n6173 ;
  assign n28796 = n28795 ^ n16351 ^ n9308 ;
  assign n28797 = n13794 ^ n7931 ^ n3960 ;
  assign n28798 = ( n13036 & ~n17718 ) | ( n13036 & n23790 ) | ( ~n17718 & n23790 ) ;
  assign n28799 = n291 & n10424 ;
  assign n28800 = n28799 ^ n7337 ^ 1'b0 ;
  assign n28801 = ( n2324 & ~n17609 ) | ( n2324 & n26410 ) | ( ~n17609 & n26410 ) ;
  assign n28802 = n18882 ^ n10721 ^ 1'b0 ;
  assign n28803 = n28802 ^ n20105 ^ n4265 ;
  assign n28804 = ( n2668 & ~n19271 ) | ( n2668 & n22909 ) | ( ~n19271 & n22909 ) ;
  assign n28807 = ( n378 & n613 ) | ( n378 & ~n11221 ) | ( n613 & ~n11221 ) ;
  assign n28805 = n20099 ^ n2779 ^ n2599 ;
  assign n28806 = ( n12821 & ~n18739 ) | ( n12821 & n28805 ) | ( ~n18739 & n28805 ) ;
  assign n28808 = n28807 ^ n28806 ^ n21521 ;
  assign n28809 = n232 & n15761 ;
  assign n28811 = ( n5947 & ~n22767 ) | ( n5947 & n23004 ) | ( ~n22767 & n23004 ) ;
  assign n28812 = n28811 ^ n10181 ^ n4585 ;
  assign n28810 = n7322 & n10064 ;
  assign n28813 = n28812 ^ n28810 ^ 1'b0 ;
  assign n28814 = n3101 & ~n4377 ;
  assign n28815 = n28814 ^ n6626 ^ n5199 ;
  assign n28816 = n22857 ^ n10857 ^ 1'b0 ;
  assign n28817 = n28815 & ~n28816 ;
  assign n28818 = ( n1832 & ~n7205 ) | ( n1832 & n9751 ) | ( ~n7205 & n9751 ) ;
  assign n28819 = n28818 ^ n21451 ^ 1'b0 ;
  assign n28820 = ( n763 & n14313 ) | ( n763 & ~n15053 ) | ( n14313 & ~n15053 ) ;
  assign n28821 = ( n1921 & ~n14947 ) | ( n1921 & n28820 ) | ( ~n14947 & n28820 ) ;
  assign n28822 = n10534 ^ n10130 ^ n9844 ;
  assign n28823 = ~n21703 & n28822 ;
  assign n28824 = ( n6686 & ~n7842 ) | ( n6686 & n24920 ) | ( ~n7842 & n24920 ) ;
  assign n28825 = n18247 ^ n15005 ^ n10316 ;
  assign n28826 = n28825 ^ n3194 ^ 1'b0 ;
  assign n28827 = ~n10821 & n18759 ;
  assign n28828 = n15606 ^ n12805 ^ n5022 ;
  assign n28829 = n28828 ^ n11034 ^ n3188 ;
  assign n28830 = n28829 ^ n25354 ^ n919 ;
  assign n28831 = n907 | n22804 ;
  assign n28832 = ( ~n13126 & n17548 ) | ( ~n13126 & n28831 ) | ( n17548 & n28831 ) ;
  assign n28833 = ( ~n15378 & n22162 ) | ( ~n15378 & n24844 ) | ( n22162 & n24844 ) ;
  assign n28834 = n28833 ^ n15776 ^ n3556 ;
  assign n28835 = n2319 | n2348 ;
  assign n28836 = n28835 ^ n11721 ^ 1'b0 ;
  assign n28837 = n28836 ^ n1607 ^ 1'b0 ;
  assign n28838 = n4287 ^ n405 ^ 1'b0 ;
  assign n28839 = n28838 ^ n18557 ^ n16149 ;
  assign n28840 = n5302 & n5574 ;
  assign n28841 = n28840 ^ n8256 ^ 1'b0 ;
  assign n28842 = n9339 ^ n1264 ^ 1'b0 ;
  assign n28843 = n18868 & ~n28842 ;
  assign n28844 = ~n5891 & n19666 ;
  assign n28845 = ~n21467 & n28844 ;
  assign n28846 = n28845 ^ n5912 ^ n1553 ;
  assign n28847 = n4283 & ~n18813 ;
  assign n28848 = ~n25560 & n28847 ;
  assign n28849 = n28848 ^ n320 ^ 1'b0 ;
  assign n28850 = ~n28846 & n28849 ;
  assign n28851 = n5717 & ~n5928 ;
  assign n28852 = n28851 ^ n11420 ^ 1'b0 ;
  assign n28853 = n28852 ^ n6505 ^ 1'b0 ;
  assign n28854 = n24515 ^ n6874 ^ x44 ;
  assign n28855 = n14300 ^ n4831 ^ n2152 ;
  assign n28856 = ( ~n482 & n25244 ) | ( ~n482 & n28855 ) | ( n25244 & n28855 ) ;
  assign n28857 = ( n5477 & n10505 ) | ( n5477 & n19275 ) | ( n10505 & n19275 ) ;
  assign n28858 = n28637 ^ n17680 ^ n15847 ;
  assign n28859 = ( n3960 & n6380 ) | ( n3960 & ~n9801 ) | ( n6380 & ~n9801 ) ;
  assign n28860 = ~n380 & n20865 ;
  assign n28861 = ( n2558 & n22997 ) | ( n2558 & ~n28860 ) | ( n22997 & ~n28860 ) ;
  assign n28862 = n9060 ^ n8344 ^ 1'b0 ;
  assign n28863 = n28862 ^ n11609 ^ n5987 ;
  assign n28864 = n28273 ^ n14109 ^ 1'b0 ;
  assign n28865 = n1735 | n8644 ;
  assign n28866 = n2801 | n28865 ;
  assign n28867 = n28866 ^ n852 ^ 1'b0 ;
  assign n28868 = ~n28864 & n28867 ;
  assign n28870 = n14547 & n18698 ;
  assign n28871 = n28870 ^ n2613 ^ 1'b0 ;
  assign n28872 = ( ~n2729 & n21983 ) | ( ~n2729 & n28871 ) | ( n21983 & n28871 ) ;
  assign n28873 = n6737 ^ n3268 ^ 1'b0 ;
  assign n28874 = n28872 & ~n28873 ;
  assign n28875 = ( ~n805 & n8829 ) | ( ~n805 & n28874 ) | ( n8829 & n28874 ) ;
  assign n28869 = n222 & n14558 ;
  assign n28876 = n28875 ^ n28869 ^ 1'b0 ;
  assign n28877 = ( ~n2662 & n7233 ) | ( ~n2662 & n8376 ) | ( n7233 & n8376 ) ;
  assign n28879 = ~n1898 & n14780 ;
  assign n28880 = n28879 ^ n7661 ^ 1'b0 ;
  assign n28881 = n28880 ^ n753 ^ 1'b0 ;
  assign n28882 = ~n12429 & n28881 ;
  assign n28878 = ( n10266 & ~n18928 ) | ( n10266 & n24756 ) | ( ~n18928 & n24756 ) ;
  assign n28883 = n28882 ^ n28878 ^ n17470 ;
  assign n28884 = n26236 ^ n16691 ^ n5303 ;
  assign n28885 = ( n11563 & ~n19714 ) | ( n11563 & n28884 ) | ( ~n19714 & n28884 ) ;
  assign n28886 = n15003 ^ n6012 ^ n5574 ;
  assign n28887 = ( n7268 & ~n28885 ) | ( n7268 & n28886 ) | ( ~n28885 & n28886 ) ;
  assign n28888 = n20516 ^ n19340 ^ 1'b0 ;
  assign n28889 = n19489 ^ n9688 ^ 1'b0 ;
  assign n28890 = n13945 ^ n10750 ^ n5169 ;
  assign n28891 = ( ~n28620 & n28889 ) | ( ~n28620 & n28890 ) | ( n28889 & n28890 ) ;
  assign n28892 = n11807 ^ n3689 ^ 1'b0 ;
  assign n28893 = ~n22620 & n28892 ;
  assign n28897 = n6150 & n19047 ;
  assign n28894 = n1271 ^ n1258 ^ 1'b0 ;
  assign n28895 = n3075 & ~n28894 ;
  assign n28896 = n10935 & n28895 ;
  assign n28898 = n28897 ^ n28896 ^ 1'b0 ;
  assign n28899 = n22858 | n27958 ;
  assign n28900 = n28899 ^ n28308 ^ 1'b0 ;
  assign n28901 = n28900 ^ n1630 ^ n751 ;
  assign n28902 = n28901 ^ n25436 ^ 1'b0 ;
  assign n28903 = n20986 ^ n6134 ^ n2606 ;
  assign n28904 = n11208 & ~n28903 ;
  assign n28905 = ~n3339 & n8694 ;
  assign n28906 = n19013 & ~n28905 ;
  assign n28907 = ( n16288 & ~n19056 ) | ( n16288 & n28396 ) | ( ~n19056 & n28396 ) ;
  assign n28908 = n26601 ^ n13544 ^ n1396 ;
  assign n28910 = ( n3484 & ~n21532 ) | ( n3484 & n23480 ) | ( ~n21532 & n23480 ) ;
  assign n28909 = n6090 ^ n3475 ^ n2560 ;
  assign n28911 = n28910 ^ n28909 ^ n15460 ;
  assign n28912 = ( ~n11754 & n16262 ) | ( ~n11754 & n16595 ) | ( n16262 & n16595 ) ;
  assign n28913 = ( n3583 & n3591 ) | ( n3583 & ~n28912 ) | ( n3591 & ~n28912 ) ;
  assign n28914 = n234 & ~n11212 ;
  assign n28915 = ~n16677 & n28914 ;
  assign n28916 = n22120 ^ n14623 ^ 1'b0 ;
  assign n28917 = n7857 & ~n28916 ;
  assign n28918 = ~n230 & n13507 ;
  assign n28919 = ~n28917 & n28918 ;
  assign n28920 = ( n7612 & n14214 ) | ( n7612 & ~n26008 ) | ( n14214 & ~n26008 ) ;
  assign n28921 = ( x107 & ~n6724 ) | ( x107 & n26618 ) | ( ~n6724 & n26618 ) ;
  assign n28922 = n5238 & n28921 ;
  assign n28923 = n28920 & n28922 ;
  assign n28924 = n18235 ^ n13400 ^ n1731 ;
  assign n28925 = n28924 ^ n2246 ^ 1'b0 ;
  assign n28926 = n28925 ^ n7344 ^ 1'b0 ;
  assign n28927 = n14218 | n28926 ;
  assign n28928 = ~n9705 & n28927 ;
  assign n28929 = ( n7303 & n17597 ) | ( n7303 & n18878 ) | ( n17597 & n18878 ) ;
  assign n28930 = n27721 ^ n15917 ^ n9036 ;
  assign n28931 = x116 | n16780 ;
  assign n28932 = ( n20984 & ~n28930 ) | ( n20984 & n28931 ) | ( ~n28930 & n28931 ) ;
  assign n28933 = ~n2814 & n5464 ;
  assign n28934 = n24338 ^ n3912 ^ 1'b0 ;
  assign n28935 = ~n17129 & n28934 ;
  assign n28936 = ( ~x83 & n20221 ) | ( ~x83 & n28935 ) | ( n20221 & n28935 ) ;
  assign n28937 = n1901 & n20371 ;
  assign n28938 = ( n2741 & n3237 ) | ( n2741 & n12101 ) | ( n3237 & n12101 ) ;
  assign n28939 = ( ~n7690 & n12039 ) | ( ~n7690 & n28938 ) | ( n12039 & n28938 ) ;
  assign n28940 = n28381 ^ n3127 ^ 1'b0 ;
  assign n28941 = n1287 | n28940 ;
  assign n28942 = n12793 ^ n7712 ^ 1'b0 ;
  assign n28943 = n15726 & ~n28942 ;
  assign n28944 = n1382 & n7749 ;
  assign n28945 = n28944 ^ n7353 ^ 1'b0 ;
  assign n28946 = n28945 ^ n25039 ^ n1569 ;
  assign n28947 = n23632 ^ n20937 ^ n5609 ;
  assign n28948 = n9099 | n13668 ;
  assign n28949 = n465 | n28948 ;
  assign n28950 = n20535 ^ n13348 ^ n8097 ;
  assign n28951 = ( n13078 & n28949 ) | ( n13078 & n28950 ) | ( n28949 & n28950 ) ;
  assign n28952 = ( n409 & ~n13057 ) | ( n409 & n16915 ) | ( ~n13057 & n16915 ) ;
  assign n28953 = n7396 & n28952 ;
  assign n28954 = n28953 ^ n26244 ^ n7413 ;
  assign n28955 = ( n1932 & n10598 ) | ( n1932 & ~n22470 ) | ( n10598 & ~n22470 ) ;
  assign n28956 = n24255 ^ n11845 ^ n5168 ;
  assign n28957 = n9703 ^ n6467 ^ n3019 ;
  assign n28958 = n6473 | n12475 ;
  assign n28959 = n28958 ^ n5294 ^ 1'b0 ;
  assign n28960 = n7368 ^ n6443 ^ 1'b0 ;
  assign n28961 = ~n28959 & n28960 ;
  assign n28962 = n11510 ^ n434 ^ 1'b0 ;
  assign n28963 = n12111 | n28962 ;
  assign n28964 = n15026 | n15569 ;
  assign n28965 = n28964 ^ n1975 ^ 1'b0 ;
  assign n28966 = ( n24718 & ~n28963 ) | ( n24718 & n28965 ) | ( ~n28963 & n28965 ) ;
  assign n28967 = n4055 | n8318 ;
  assign n28968 = n28966 | n28967 ;
  assign n28969 = n24338 & ~n25130 ;
  assign n28970 = n28969 ^ n333 ^ 1'b0 ;
  assign n28971 = n13659 ^ n7110 ^ 1'b0 ;
  assign n28972 = ( x118 & ~n5796 ) | ( x118 & n15522 ) | ( ~n5796 & n15522 ) ;
  assign n28974 = n7314 & ~n24127 ;
  assign n28973 = ( ~n494 & n10766 ) | ( ~n494 & n19876 ) | ( n10766 & n19876 ) ;
  assign n28975 = n28974 ^ n28973 ^ n395 ;
  assign n28976 = ( n9089 & n28972 ) | ( n9089 & n28975 ) | ( n28972 & n28975 ) ;
  assign n28977 = n28976 ^ n13578 ^ n3452 ;
  assign n28978 = x98 & n1848 ;
  assign n28979 = n28978 ^ n2294 ^ 1'b0 ;
  assign n28980 = n28979 ^ n21608 ^ n245 ;
  assign n28981 = ( n8885 & ~n15455 ) | ( n8885 & n28980 ) | ( ~n15455 & n28980 ) ;
  assign n28982 = ( n3381 & n8693 ) | ( n3381 & n10359 ) | ( n8693 & n10359 ) ;
  assign n28983 = n22323 ^ n10745 ^ n2975 ;
  assign n28984 = n28182 | n28630 ;
  assign n28986 = ( n383 & n2364 ) | ( n383 & n5679 ) | ( n2364 & n5679 ) ;
  assign n28985 = ~n810 & n7924 ;
  assign n28987 = n28986 ^ n28985 ^ 1'b0 ;
  assign n28988 = n6492 | n28987 ;
  assign n28989 = n28988 ^ n21153 ^ 1'b0 ;
  assign n28990 = n8333 & n14360 ;
  assign n28991 = n28989 & n28990 ;
  assign n28992 = n28991 ^ n567 ^ 1'b0 ;
  assign n28993 = n16481 & n27052 ;
  assign n28994 = n2640 & n28993 ;
  assign n28995 = n3165 & n4141 ;
  assign n28996 = n5659 & n28995 ;
  assign n28997 = ( n4853 & n13556 ) | ( n4853 & ~n24040 ) | ( n13556 & ~n24040 ) ;
  assign n28998 = n24293 ^ n848 ^ 1'b0 ;
  assign n28999 = ~n9328 & n28998 ;
  assign n29000 = ( n7339 & n15128 ) | ( n7339 & ~n21731 ) | ( n15128 & ~n21731 ) ;
  assign n29001 = ( n4308 & ~n13580 ) | ( n4308 & n29000 ) | ( ~n13580 & n29000 ) ;
  assign n29002 = ( n23849 & n28999 ) | ( n23849 & n29001 ) | ( n28999 & n29001 ) ;
  assign n29003 = n28250 ^ n10708 ^ 1'b0 ;
  assign n29004 = n8871 & ~n19686 ;
  assign n29005 = ( n4624 & ~n11963 ) | ( n4624 & n15703 ) | ( ~n11963 & n15703 ) ;
  assign n29006 = n18453 ^ n13900 ^ 1'b0 ;
  assign n29007 = ~n9855 & n18565 ;
  assign n29008 = ( ~n2694 & n29006 ) | ( ~n2694 & n29007 ) | ( n29006 & n29007 ) ;
  assign n29009 = ~n1795 & n4458 ;
  assign n29010 = n29009 ^ n25055 ^ 1'b0 ;
  assign n29011 = n1122 | n21183 ;
  assign n29012 = n29010 & ~n29011 ;
  assign n29013 = n20169 ^ n13857 ^ n6498 ;
  assign n29014 = ( ~n15162 & n19069 ) | ( ~n15162 & n26734 ) | ( n19069 & n26734 ) ;
  assign n29015 = n2909 & ~n4202 ;
  assign n29016 = n12800 | n23250 ;
  assign n29017 = ( n18352 & ~n29015 ) | ( n18352 & n29016 ) | ( ~n29015 & n29016 ) ;
  assign n29018 = n29017 ^ n20133 ^ 1'b0 ;
  assign n29019 = n29014 & ~n29018 ;
  assign n29020 = ~n812 & n29019 ;
  assign n29021 = n12569 & n29020 ;
  assign n29022 = ( ~n6175 & n20160 ) | ( ~n6175 & n29021 ) | ( n20160 & n29021 ) ;
  assign n29023 = n1000 & ~n16052 ;
  assign n29024 = n29023 ^ n25561 ^ 1'b0 ;
  assign n29025 = ( ~n3422 & n20884 ) | ( ~n3422 & n29024 ) | ( n20884 & n29024 ) ;
  assign n29026 = n24895 ^ n22998 ^ n9528 ;
  assign n29027 = n12053 ^ n935 ^ 1'b0 ;
  assign n29028 = n28317 ^ n467 ^ 1'b0 ;
  assign n29029 = n11026 & n29028 ;
  assign n29030 = n140 & n29029 ;
  assign n29031 = n29030 ^ n24663 ^ 1'b0 ;
  assign n29032 = n27273 ^ n19980 ^ 1'b0 ;
  assign n29034 = n14668 ^ n14016 ^ n7912 ;
  assign n29033 = n7494 & n28480 ;
  assign n29035 = n29034 ^ n29033 ^ 1'b0 ;
  assign n29036 = n12524 & n14831 ;
  assign n29037 = n26207 & n29036 ;
  assign n29038 = n26299 ^ n3515 ^ 1'b0 ;
  assign n29039 = ( n14875 & n15805 ) | ( n14875 & n28604 ) | ( n15805 & n28604 ) ;
  assign n29040 = ~n5303 & n12555 ;
  assign n29041 = n29040 ^ n16241 ^ n927 ;
  assign n29042 = n14483 ^ n12044 ^ n1413 ;
  assign n29043 = n29042 ^ n23057 ^ n5525 ;
  assign n29045 = ( x1 & n1750 ) | ( x1 & n9423 ) | ( n1750 & n9423 ) ;
  assign n29044 = ~n15687 & n19357 ;
  assign n29046 = n29045 ^ n29044 ^ 1'b0 ;
  assign n29047 = n14892 ^ n9044 ^ n7885 ;
  assign n29048 = n29047 ^ n5819 ^ 1'b0 ;
  assign n29049 = n29046 & ~n29048 ;
  assign n29050 = n29049 ^ n23319 ^ n17582 ;
  assign n29051 = n10199 | n19482 ;
  assign n29052 = n29051 ^ n27689 ^ 1'b0 ;
  assign n29053 = n29052 ^ n13831 ^ n1973 ;
  assign n29054 = n29053 ^ n10445 ^ n3288 ;
  assign n29055 = n15319 | n27969 ;
  assign n29056 = n29055 ^ n8867 ^ 1'b0 ;
  assign n29057 = ( ~n201 & n1531 ) | ( ~n201 & n6960 ) | ( n1531 & n6960 ) ;
  assign n29058 = n29057 ^ n4356 ^ 1'b0 ;
  assign n29059 = n14471 | n29058 ;
  assign n29060 = n9996 & ~n14299 ;
  assign n29061 = n7492 | n24804 ;
  assign n29062 = n15152 | n29061 ;
  assign n29063 = n29062 ^ n19578 ^ n16060 ;
  assign n29064 = n23060 & ~n29063 ;
  assign n29065 = ( x115 & ~n22250 ) | ( x115 & n28022 ) | ( ~n22250 & n28022 ) ;
  assign n29066 = n20320 ^ n4438 ^ 1'b0 ;
  assign n29067 = n7824 ^ n2463 ^ 1'b0 ;
  assign n29068 = n29067 ^ n18202 ^ n13915 ;
  assign n29069 = n29068 ^ n484 ^ 1'b0 ;
  assign n29070 = n20266 ^ n5928 ^ 1'b0 ;
  assign n29071 = n29070 ^ n13361 ^ n6039 ;
  assign n29072 = ( n490 & n3481 ) | ( n490 & n27364 ) | ( n3481 & n27364 ) ;
  assign n29073 = n11737 & n22740 ;
  assign n29074 = n29072 & n29073 ;
  assign n29075 = x80 & ~n6226 ;
  assign n29076 = n12351 ^ n9508 ^ n8957 ;
  assign n29077 = n19207 & n29076 ;
  assign n29078 = ( ~n3703 & n5509 ) | ( ~n3703 & n21499 ) | ( n5509 & n21499 ) ;
  assign n29079 = ~n25052 & n29005 ;
  assign n29080 = n25461 ^ n3653 ^ 1'b0 ;
  assign n29081 = n14869 & n24397 ;
  assign n29084 = n24363 ^ n8684 ^ 1'b0 ;
  assign n29085 = ~n21127 & n29084 ;
  assign n29082 = n17808 ^ n8147 ^ n2334 ;
  assign n29083 = ~n27381 & n29082 ;
  assign n29086 = n29085 ^ n29083 ^ 1'b0 ;
  assign n29087 = ~n1313 & n8899 ;
  assign n29088 = n4525 | n7353 ;
  assign n29089 = n2112 & ~n29088 ;
  assign n29090 = n3679 | n22016 ;
  assign n29091 = n3241 ^ n1524 ^ 1'b0 ;
  assign n29092 = n29090 & n29091 ;
  assign n29093 = ( ~n9728 & n14761 ) | ( ~n9728 & n29038 ) | ( n14761 & n29038 ) ;
  assign n29094 = ( ~n4187 & n6813 ) | ( ~n4187 & n10505 ) | ( n6813 & n10505 ) ;
  assign n29095 = n29094 ^ n10721 ^ 1'b0 ;
  assign n29096 = n29095 ^ n9062 ^ n3385 ;
  assign n29097 = n26988 ^ n686 ^ 1'b0 ;
  assign n29098 = n29097 ^ n16757 ^ n295 ;
  assign n29099 = n11371 ^ n10094 ^ 1'b0 ;
  assign n29100 = ~n623 & n29099 ;
  assign n29101 = ( ~n5149 & n15060 ) | ( ~n5149 & n29100 ) | ( n15060 & n29100 ) ;
  assign n29102 = n29101 ^ n12306 ^ n8402 ;
  assign n29103 = n29102 ^ n13482 ^ 1'b0 ;
  assign n29104 = ~n29098 & n29103 ;
  assign n29105 = ( n6060 & ~n6090 ) | ( n6060 & n29104 ) | ( ~n6090 & n29104 ) ;
  assign n29106 = n9539 ^ x96 ^ 1'b0 ;
  assign n29107 = n29106 ^ n24167 ^ n12082 ;
  assign n29109 = ( n4354 & ~n15410 ) | ( n4354 & n16914 ) | ( ~n15410 & n16914 ) ;
  assign n29108 = n17047 ^ n15723 ^ n8576 ;
  assign n29110 = n29109 ^ n29108 ^ n20385 ;
  assign n29111 = ~n1118 & n10465 ;
  assign n29112 = n6388 & ~n15981 ;
  assign n29113 = n931 | n2526 ;
  assign n29114 = n29113 ^ n15248 ^ 1'b0 ;
  assign n29115 = n24832 ^ n7551 ^ 1'b0 ;
  assign n29116 = n3751 & n11134 ;
  assign n29117 = n29116 ^ n23006 ^ 1'b0 ;
  assign n29118 = n11080 & ~n29117 ;
  assign n29119 = n26410 ^ n22024 ^ n7244 ;
  assign n29120 = n13525 ^ n10151 ^ n8347 ;
  assign n29121 = ( n3684 & n15376 ) | ( n3684 & n29120 ) | ( n15376 & n29120 ) ;
  assign n29122 = n16309 ^ n6243 ^ n2360 ;
  assign n29123 = n14820 ^ n6740 ^ n4930 ;
  assign n29124 = n29123 ^ n14144 ^ 1'b0 ;
  assign n29125 = n21527 ^ n17347 ^ n1924 ;
  assign n29126 = ( n5565 & ~n23785 ) | ( n5565 & n24283 ) | ( ~n23785 & n24283 ) ;
  assign n29127 = ( n6870 & n11845 ) | ( n6870 & ~n22896 ) | ( n11845 & ~n22896 ) ;
  assign n29128 = n24255 ^ n9813 ^ 1'b0 ;
  assign n29129 = n29127 | n29128 ;
  assign n29134 = ( ~n6126 & n11653 ) | ( ~n6126 & n19524 ) | ( n11653 & n19524 ) ;
  assign n29135 = ( ~n258 & n10165 ) | ( ~n258 & n29134 ) | ( n10165 & n29134 ) ;
  assign n29130 = ( n8937 & n13317 ) | ( n8937 & n18843 ) | ( n13317 & n18843 ) ;
  assign n29131 = n29130 ^ n22339 ^ 1'b0 ;
  assign n29132 = n29131 ^ n27854 ^ 1'b0 ;
  assign n29133 = n21479 & n29132 ;
  assign n29136 = n29135 ^ n29133 ^ 1'b0 ;
  assign n29138 = ( n2558 & n3077 ) | ( n2558 & ~n5662 ) | ( n3077 & ~n5662 ) ;
  assign n29137 = n7058 & ~n18632 ;
  assign n29139 = n29138 ^ n29137 ^ 1'b0 ;
  assign n29140 = ( n5319 & n12421 ) | ( n5319 & ~n19725 ) | ( n12421 & ~n19725 ) ;
  assign n29141 = n10053 ^ n7091 ^ 1'b0 ;
  assign n29142 = ~n29140 & n29141 ;
  assign n29143 = ( n11112 & n12723 ) | ( n11112 & ~n20812 ) | ( n12723 & ~n20812 ) ;
  assign n29144 = n10368 & n29143 ;
  assign n29145 = ( x124 & n2483 ) | ( x124 & ~n24372 ) | ( n2483 & ~n24372 ) ;
  assign n29146 = n28649 ^ n26557 ^ n14862 ;
  assign n29147 = n29146 ^ x99 ^ 1'b0 ;
  assign n29148 = ( ~n27517 & n29145 ) | ( ~n27517 & n29147 ) | ( n29145 & n29147 ) ;
  assign n29149 = n25967 ^ n22347 ^ n9059 ;
  assign n29150 = n22257 ^ n4410 ^ 1'b0 ;
  assign n29151 = ( n1606 & ~n5675 ) | ( n1606 & n22087 ) | ( ~n5675 & n22087 ) ;
  assign n29152 = n15516 ^ n6264 ^ 1'b0 ;
  assign n29153 = n24230 | n29152 ;
  assign n29154 = n12040 ^ n7746 ^ 1'b0 ;
  assign n29155 = n6765 ^ n1492 ^ 1'b0 ;
  assign n29156 = ( n8235 & ~n23108 ) | ( n8235 & n29155 ) | ( ~n23108 & n29155 ) ;
  assign n29157 = n2339 & ~n13451 ;
  assign n29158 = ~n26745 & n29157 ;
  assign n29159 = n29158 ^ n9133 ^ n5818 ;
  assign n29160 = ( n4244 & ~n5447 ) | ( n4244 & n20623 ) | ( ~n5447 & n20623 ) ;
  assign n29161 = ( n553 & n8769 ) | ( n553 & n28317 ) | ( n8769 & n28317 ) ;
  assign n29162 = n29161 ^ n25721 ^ n14209 ;
  assign n29164 = ( n13181 & n15659 ) | ( n13181 & ~n27394 ) | ( n15659 & ~n27394 ) ;
  assign n29163 = n21736 ^ n8372 ^ n7187 ;
  assign n29165 = n29164 ^ n29163 ^ 1'b0 ;
  assign n29166 = n22414 ^ x49 ^ 1'b0 ;
  assign n29167 = n6271 | n12944 ;
  assign n29168 = n9814 & ~n29167 ;
  assign n29169 = ( n4497 & ~n29166 ) | ( n4497 & n29168 ) | ( ~n29166 & n29168 ) ;
  assign n29170 = n23560 ^ n21793 ^ n557 ;
  assign n29171 = n26552 ^ n9701 ^ 1'b0 ;
  assign n29172 = n29170 & n29171 ;
  assign n29173 = n28164 ^ n14940 ^ 1'b0 ;
  assign n29174 = n3202 & ~n29173 ;
  assign n29175 = n25157 ^ n22291 ^ n1927 ;
  assign n29176 = n24328 ^ n2015 ^ 1'b0 ;
  assign n29177 = ~n29175 & n29176 ;
  assign n29178 = ( n10002 & n15612 ) | ( n10002 & ~n19978 ) | ( n15612 & ~n19978 ) ;
  assign n29179 = n29178 ^ n25282 ^ n4964 ;
  assign n29180 = n13596 ^ n9382 ^ n5544 ;
  assign n29181 = n11250 ^ n2517 ^ 1'b0 ;
  assign n29182 = n12793 ^ n12221 ^ n795 ;
  assign n29183 = ( ~n1657 & n23108 ) | ( ~n1657 & n29182 ) | ( n23108 & n29182 ) ;
  assign n29184 = n7378 ^ n4795 ^ 1'b0 ;
  assign n29185 = ( n29181 & n29183 ) | ( n29181 & n29184 ) | ( n29183 & n29184 ) ;
  assign n29186 = n18864 ^ n1284 ^ 1'b0 ;
  assign n29187 = n29186 ^ n14096 ^ n1956 ;
  assign n29188 = n28689 ^ n1591 ^ 1'b0 ;
  assign n29189 = n29188 ^ n27762 ^ n13037 ;
  assign n29190 = ( ~n2668 & n14311 ) | ( ~n2668 & n22211 ) | ( n14311 & n22211 ) ;
  assign n29191 = n29190 ^ n9129 ^ n8303 ;
  assign n29192 = ( n4742 & n5704 ) | ( n4742 & ~n29191 ) | ( n5704 & ~n29191 ) ;
  assign n29193 = n2986 & n3168 ;
  assign n29194 = ~n6101 & n29193 ;
  assign n29195 = n826 | n29194 ;
  assign n29196 = n18306 ^ n10380 ^ 1'b0 ;
  assign n29197 = ~n1712 & n2218 ;
  assign n29199 = n10190 ^ n2061 ^ n835 ;
  assign n29198 = ( n6250 & ~n22082 ) | ( n6250 & n26078 ) | ( ~n22082 & n26078 ) ;
  assign n29200 = n29199 ^ n29198 ^ 1'b0 ;
  assign n29201 = n11059 | n29200 ;
  assign n29202 = n29201 ^ n10078 ^ n8255 ;
  assign n29204 = n11638 ^ n8516 ^ 1'b0 ;
  assign n29205 = ~n23060 & n29204 ;
  assign n29206 = ~n17309 & n29205 ;
  assign n29207 = n6872 & n29206 ;
  assign n29203 = n13875 ^ n13527 ^ n6997 ;
  assign n29208 = n29207 ^ n29203 ^ n3862 ;
  assign n29209 = n1325 ^ n183 ^ 1'b0 ;
  assign n29210 = n2218 & n23411 ;
  assign n29211 = ( ~n3075 & n14222 ) | ( ~n3075 & n28060 ) | ( n14222 & n28060 ) ;
  assign n29214 = n7919 | n12139 ;
  assign n29215 = n4115 & ~n29214 ;
  assign n29212 = ( n1257 & n7535 ) | ( n1257 & ~n9362 ) | ( n7535 & ~n9362 ) ;
  assign n29213 = n29212 ^ n9164 ^ n5267 ;
  assign n29216 = n29215 ^ n29213 ^ n21382 ;
  assign n29217 = n2249 ^ n1582 ^ 1'b0 ;
  assign n29218 = n466 | n29217 ;
  assign n29219 = n4758 ^ n4209 ^ n2994 ;
  assign n29220 = n29219 ^ n19971 ^ n17393 ;
  assign n29221 = ( ~n4903 & n5722 ) | ( ~n4903 & n10836 ) | ( n5722 & n10836 ) ;
  assign n29222 = n25434 | n29221 ;
  assign n29223 = n29220 & ~n29222 ;
  assign n29224 = n6991 ^ n4882 ^ 1'b0 ;
  assign n29225 = n17120 ^ n1409 ^ 1'b0 ;
  assign n29226 = n21728 ^ n14927 ^ 1'b0 ;
  assign n29227 = ( n255 & ~n10199 ) | ( n255 & n27641 ) | ( ~n10199 & n27641 ) ;
  assign n29228 = ( n11136 & ~n11596 ) | ( n11136 & n29227 ) | ( ~n11596 & n29227 ) ;
  assign n29229 = n14448 | n29228 ;
  assign n29230 = n29229 ^ n19532 ^ n6392 ;
  assign n29231 = n7759 ^ n3582 ^ n1840 ;
  assign n29232 = n29231 ^ n1680 ^ 1'b0 ;
  assign n29233 = ( n4884 & n26022 ) | ( n4884 & n29232 ) | ( n26022 & n29232 ) ;
  assign n29234 = n13479 ^ n11896 ^ n11484 ;
  assign n29235 = n1148 & n29234 ;
  assign n29236 = n2988 & n29235 ;
  assign n29237 = ( n11641 & n17014 ) | ( n11641 & ~n29236 ) | ( n17014 & ~n29236 ) ;
  assign n29238 = n21790 ^ n16435 ^ n5071 ;
  assign n29239 = ( n2024 & n4497 ) | ( n2024 & ~n29238 ) | ( n4497 & ~n29238 ) ;
  assign n29240 = n17582 ^ n11315 ^ 1'b0 ;
  assign n29241 = n12392 & n29240 ;
  assign n29242 = n27805 ^ n13941 ^ 1'b0 ;
  assign n29243 = n1004 & n29242 ;
  assign n29244 = ~n17336 & n19191 ;
  assign n29245 = n10197 & ~n15512 ;
  assign n29246 = n15309 ^ n14098 ^ n4732 ;
  assign n29247 = n2885 | n29246 ;
  assign n29248 = n8557 & ~n10774 ;
  assign n29249 = ( n511 & n6988 ) | ( n511 & n20575 ) | ( n6988 & n20575 ) ;
  assign n29250 = ( n15890 & n29248 ) | ( n15890 & n29249 ) | ( n29248 & n29249 ) ;
  assign n29251 = n29250 ^ n19515 ^ n19492 ;
  assign n29252 = ~n14490 & n29251 ;
  assign n29254 = n7412 ^ n3229 ^ n2645 ;
  assign n29253 = ( n9462 & n10840 ) | ( n9462 & n14422 ) | ( n10840 & n14422 ) ;
  assign n29255 = n29254 ^ n29253 ^ 1'b0 ;
  assign n29256 = n10684 ^ n9582 ^ n6514 ;
  assign n29257 = ( ~n13741 & n28260 ) | ( ~n13741 & n29256 ) | ( n28260 & n29256 ) ;
  assign n29258 = n29257 ^ n19419 ^ n3458 ;
  assign n29259 = n7395 ^ x82 ^ 1'b0 ;
  assign n29260 = n20402 ^ n12629 ^ n1101 ;
  assign n29263 = n7129 ^ n469 ^ 1'b0 ;
  assign n29264 = ~n6130 & n29263 ;
  assign n29261 = n8865 | n17792 ;
  assign n29262 = n18393 & ~n29261 ;
  assign n29265 = n29264 ^ n29262 ^ n8574 ;
  assign n29266 = ( n1295 & n29260 ) | ( n1295 & n29265 ) | ( n29260 & n29265 ) ;
  assign n29267 = n26910 ^ n25638 ^ 1'b0 ;
  assign n29268 = n21821 & ~n29267 ;
  assign n29269 = n29268 ^ n6370 ^ 1'b0 ;
  assign n29270 = n4159 ^ n2624 ^ 1'b0 ;
  assign n29271 = n15500 & ~n29270 ;
  assign n29272 = ~n5439 & n29271 ;
  assign n29273 = ( ~n16557 & n21534 ) | ( ~n16557 & n27424 ) | ( n21534 & n27424 ) ;
  assign n29274 = n716 & n13350 ;
  assign n29275 = n29274 ^ n24272 ^ 1'b0 ;
  assign n29276 = n12276 ^ n9076 ^ n3138 ;
  assign n29277 = n22978 & n29276 ;
  assign n29278 = ( n5107 & n29275 ) | ( n5107 & n29277 ) | ( n29275 & n29277 ) ;
  assign n29279 = n20786 ^ n13139 ^ 1'b0 ;
  assign n29280 = n860 & ~n29279 ;
  assign n29281 = ( ~n4520 & n24046 ) | ( ~n4520 & n29280 ) | ( n24046 & n29280 ) ;
  assign n29282 = n28028 ^ n8138 ^ 1'b0 ;
  assign n29283 = n13292 & n29282 ;
  assign n29284 = n10246 ^ n9344 ^ 1'b0 ;
  assign n29285 = ~n1557 & n29284 ;
  assign n29286 = n16627 | n24844 ;
  assign n29287 = n28449 ^ n7934 ^ n1184 ;
  assign n29288 = n1993 & ~n26942 ;
  assign n29289 = ~n188 & n29288 ;
  assign n29290 = n29289 ^ n21678 ^ n1793 ;
  assign n29291 = ( ~n17986 & n29287 ) | ( ~n17986 & n29290 ) | ( n29287 & n29290 ) ;
  assign n29292 = n17872 ^ n6238 ^ n5609 ;
  assign n29295 = ( n9765 & n18976 ) | ( n9765 & ~n19935 ) | ( n18976 & ~n19935 ) ;
  assign n29293 = n5930 & ~n7178 ;
  assign n29294 = n29293 ^ n6288 ^ 1'b0 ;
  assign n29296 = n29295 ^ n29294 ^ n26003 ;
  assign n29297 = n23458 ^ n197 ^ 1'b0 ;
  assign n29298 = n29297 ^ n10196 ^ n1330 ;
  assign n29299 = n28334 ^ n9019 ^ n4055 ;
  assign n29300 = n3820 | n9303 ;
  assign n29301 = n27992 | n29300 ;
  assign n29302 = n17801 ^ n2086 ^ 1'b0 ;
  assign n29303 = ( n715 & n3271 ) | ( n715 & ~n6168 ) | ( n3271 & ~n6168 ) ;
  assign n29304 = n1843 | n29303 ;
  assign n29305 = n19714 & ~n29304 ;
  assign n29306 = n3364 & n20961 ;
  assign n29307 = n29306 ^ n25015 ^ 1'b0 ;
  assign n29308 = ( n23030 & ~n28689 ) | ( n23030 & n29307 ) | ( ~n28689 & n29307 ) ;
  assign n29309 = ( ~n17176 & n19174 ) | ( ~n17176 & n21288 ) | ( n19174 & n21288 ) ;
  assign n29310 = ( n2906 & n4939 ) | ( n2906 & ~n6658 ) | ( n4939 & ~n6658 ) ;
  assign n29311 = ( n3127 & n13610 ) | ( n3127 & n15139 ) | ( n13610 & n15139 ) ;
  assign n29312 = n26257 ^ n19647 ^ n9207 ;
  assign n29314 = n5034 ^ n870 ^ 1'b0 ;
  assign n29313 = ( n1207 & n7718 ) | ( n1207 & n7878 ) | ( n7718 & n7878 ) ;
  assign n29315 = n29314 ^ n29313 ^ n3772 ;
  assign n29316 = n12550 & ~n26942 ;
  assign n29317 = ~n3243 & n29316 ;
  assign n29318 = n29317 ^ n13101 ^ 1'b0 ;
  assign n29319 = n21254 | n23874 ;
  assign n29320 = n7111 | n29319 ;
  assign n29321 = n1138 & ~n6961 ;
  assign n29322 = n29321 ^ n4223 ^ 1'b0 ;
  assign n29323 = n29322 ^ n22898 ^ n15270 ;
  assign n29324 = n12719 ^ n417 ^ 1'b0 ;
  assign n29325 = n787 & n16627 ;
  assign n29326 = ( n659 & ~n26995 ) | ( n659 & n29325 ) | ( ~n26995 & n29325 ) ;
  assign n29327 = n29326 ^ n8462 ^ n1851 ;
  assign n29328 = n5489 ^ n3963 ^ n1261 ;
  assign n29329 = n8487 & n18285 ;
  assign n29330 = ( n545 & n23501 ) | ( n545 & n29329 ) | ( n23501 & n29329 ) ;
  assign n29331 = ( ~n13641 & n20231 ) | ( ~n13641 & n23369 ) | ( n20231 & n23369 ) ;
  assign n29332 = n9133 ^ n5775 ^ 1'b0 ;
  assign n29333 = ( ~n4976 & n29331 ) | ( ~n4976 & n29332 ) | ( n29331 & n29332 ) ;
  assign n29334 = n18529 ^ n9048 ^ n1075 ;
  assign n29335 = n28485 ^ n22163 ^ 1'b0 ;
  assign n29336 = n5798 & ~n28303 ;
  assign n29337 = n29336 ^ n18683 ^ 1'b0 ;
  assign n29338 = n23181 & ~n23444 ;
  assign n29339 = n27228 | n29338 ;
  assign n29340 = n11131 | n29339 ;
  assign n29341 = n22190 ^ n3031 ^ 1'b0 ;
  assign n29342 = n5411 | n29341 ;
  assign n29343 = n7545 ^ n6346 ^ 1'b0 ;
  assign n29344 = n131 & ~n4683 ;
  assign n29345 = n29343 & n29344 ;
  assign n29346 = ( n4604 & n4813 ) | ( n4604 & n19809 ) | ( n4813 & n19809 ) ;
  assign n29347 = n29346 ^ n11838 ^ 1'b0 ;
  assign n29348 = ( n2998 & n29345 ) | ( n2998 & ~n29347 ) | ( n29345 & ~n29347 ) ;
  assign n29349 = n9206 | n10461 ;
  assign n29350 = n29349 ^ n27366 ^ n14537 ;
  assign n29353 = n12187 ^ n11745 ^ 1'b0 ;
  assign n29354 = n13362 & ~n29353 ;
  assign n29352 = n29182 ^ n8206 ^ 1'b0 ;
  assign n29351 = n8736 ^ n3910 ^ 1'b0 ;
  assign n29355 = n29354 ^ n29352 ^ n29351 ;
  assign n29356 = ( ~n4300 & n5709 ) | ( ~n4300 & n17644 ) | ( n5709 & n17644 ) ;
  assign n29357 = n17534 & ~n29356 ;
  assign n29358 = n17584 ^ n8781 ^ n5726 ;
  assign n29359 = n29358 ^ n25957 ^ n7652 ;
  assign n29360 = n3734 & ~n29359 ;
  assign n29361 = n29360 ^ n19059 ^ 1'b0 ;
  assign n29362 = n15356 ^ n14687 ^ n5414 ;
  assign n29363 = n4359 & n29362 ;
  assign n29364 = ( ~n8292 & n22962 ) | ( ~n8292 & n29363 ) | ( n22962 & n29363 ) ;
  assign n29365 = n2838 | n27043 ;
  assign n29366 = n26381 ^ n23118 ^ n2717 ;
  assign n29367 = n29366 ^ n9137 ^ n611 ;
  assign n29368 = n3916 | n4903 ;
  assign n29369 = n24054 ^ n14927 ^ n10827 ;
  assign n29370 = ( ~n2279 & n15395 ) | ( ~n2279 & n29369 ) | ( n15395 & n29369 ) ;
  assign n29371 = ( n14210 & ~n14724 ) | ( n14210 & n29370 ) | ( ~n14724 & n29370 ) ;
  assign n29372 = ( n7530 & ~n10404 ) | ( n7530 & n22255 ) | ( ~n10404 & n22255 ) ;
  assign n29373 = n29372 ^ n17556 ^ 1'b0 ;
  assign n29374 = n1913 & ~n5423 ;
  assign n29375 = n29374 ^ n27593 ^ n17222 ;
  assign n29376 = n29375 ^ n23120 ^ 1'b0 ;
  assign n29377 = n1540 ^ n1201 ^ 1'b0 ;
  assign n29378 = n22174 ^ n1996 ^ 1'b0 ;
  assign n29379 = n29377 & n29378 ;
  assign n29380 = n29379 ^ n11015 ^ n1543 ;
  assign n29381 = n21065 ^ n6572 ^ n3120 ;
  assign n29382 = n16673 & n27909 ;
  assign n29383 = n17431 ^ x46 ^ 1'b0 ;
  assign n29384 = n1129 & ~n10508 ;
  assign n29385 = n29384 ^ n3477 ^ n562 ;
  assign n29386 = n29383 | n29385 ;
  assign n29387 = n29386 ^ n17879 ^ n11262 ;
  assign n29388 = n23805 ^ n164 ^ 1'b0 ;
  assign n29389 = n28247 & ~n29388 ;
  assign n29390 = n15050 ^ n6916 ^ 1'b0 ;
  assign n29391 = n5263 ^ n3064 ^ 1'b0 ;
  assign n29392 = n29390 & n29391 ;
  assign n29393 = n5020 & n6451 ;
  assign n29394 = n29393 ^ n13512 ^ 1'b0 ;
  assign n29395 = n5661 | n9904 ;
  assign n29396 = n11651 & ~n29395 ;
  assign n29397 = ( n4053 & n8075 ) | ( n4053 & n23639 ) | ( n8075 & n23639 ) ;
  assign n29398 = ( n585 & n4234 ) | ( n585 & n29397 ) | ( n4234 & n29397 ) ;
  assign n29399 = n23951 ^ n4654 ^ n2818 ;
  assign n29401 = n3040 & n20244 ;
  assign n29402 = n6557 & n29401 ;
  assign n29400 = n3668 | n21066 ;
  assign n29403 = n29402 ^ n29400 ^ 1'b0 ;
  assign n29404 = n28855 ^ n10761 ^ 1'b0 ;
  assign n29405 = ~n29403 & n29404 ;
  assign n29406 = ( ~n3238 & n3790 ) | ( ~n3238 & n29405 ) | ( n3790 & n29405 ) ;
  assign n29407 = n26654 ^ n8949 ^ 1'b0 ;
  assign n29408 = n7328 & ~n29407 ;
  assign n29409 = n29408 ^ n10943 ^ 1'b0 ;
  assign n29410 = ( ~n2662 & n5730 ) | ( ~n2662 & n29409 ) | ( n5730 & n29409 ) ;
  assign n29411 = ~n1744 & n11997 ;
  assign n29412 = n20407 & n29411 ;
  assign n29413 = ( n7896 & ~n14471 ) | ( n7896 & n29412 ) | ( ~n14471 & n29412 ) ;
  assign n29414 = n17169 & ~n25954 ;
  assign n29417 = n16195 ^ n13971 ^ n10561 ;
  assign n29418 = n29417 ^ n17943 ^ n6984 ;
  assign n29419 = ( ~n15640 & n16494 ) | ( ~n15640 & n29418 ) | ( n16494 & n29418 ) ;
  assign n29420 = ~n2030 & n29419 ;
  assign n29421 = n29420 ^ n2727 ^ 1'b0 ;
  assign n29415 = n18386 ^ n16436 ^ n7858 ;
  assign n29416 = x0 & n29415 ;
  assign n29422 = n29421 ^ n29416 ^ 1'b0 ;
  assign n29423 = n7544 | n14200 ;
  assign n29424 = n24658 & ~n29423 ;
  assign n29425 = x37 & n9557 ;
  assign n29426 = ~n7287 & n29425 ;
  assign n29427 = ( n628 & ~n7175 ) | ( n628 & n7184 ) | ( ~n7175 & n7184 ) ;
  assign n29428 = ( ~n7218 & n13518 ) | ( ~n7218 & n29427 ) | ( n13518 & n29427 ) ;
  assign n29429 = n14824 ^ n3823 ^ n1990 ;
  assign n29430 = n20509 ^ n13186 ^ 1'b0 ;
  assign n29431 = ( n2296 & n29429 ) | ( n2296 & ~n29430 ) | ( n29429 & ~n29430 ) ;
  assign n29432 = ( n4456 & ~n16717 ) | ( n4456 & n28676 ) | ( ~n16717 & n28676 ) ;
  assign n29433 = n4843 | n26596 ;
  assign n29434 = n23770 ^ n14054 ^ n5409 ;
  assign n29435 = n27393 | n29434 ;
  assign n29436 = ~n10122 & n12817 ;
  assign n29437 = n29436 ^ n20850 ^ n7894 ;
  assign n29438 = n344 & n24404 ;
  assign n29439 = ~x79 & n29438 ;
  assign n29440 = n3561 & n19046 ;
  assign n29441 = n29440 ^ n4459 ^ 1'b0 ;
  assign n29442 = ( n9977 & n12138 ) | ( n9977 & n17881 ) | ( n12138 & n17881 ) ;
  assign n29443 = n13173 & n14604 ;
  assign n29444 = n29442 & n29443 ;
  assign n29448 = n1189 & ~n4798 ;
  assign n29449 = n3976 | n13596 ;
  assign n29450 = n29448 & n29449 ;
  assign n29445 = n8723 & ~n16510 ;
  assign n29446 = n29445 ^ n7912 ^ n5484 ;
  assign n29447 = ~n2209 & n29446 ;
  assign n29451 = n29450 ^ n29447 ^ 1'b0 ;
  assign n29452 = n29343 ^ n19540 ^ n15507 ;
  assign n29453 = n29452 ^ n27213 ^ n8192 ;
  assign n29454 = ( n334 & ~n16709 ) | ( n334 & n23419 ) | ( ~n16709 & n23419 ) ;
  assign n29455 = ( n17703 & n19263 ) | ( n17703 & ~n29454 ) | ( n19263 & ~n29454 ) ;
  assign n29456 = n2563 | n23051 ;
  assign n29457 = n29456 ^ n3425 ^ 1'b0 ;
  assign n29458 = n15017 & n29457 ;
  assign n29459 = n6158 ^ n4711 ^ n1696 ;
  assign n29460 = ~n8460 & n29459 ;
  assign n29461 = n29458 & n29460 ;
  assign n29462 = n29461 ^ n17350 ^ n16340 ;
  assign n29463 = n18265 & ~n25701 ;
  assign n29464 = n29463 ^ n16063 ^ 1'b0 ;
  assign n29465 = n29464 ^ n16071 ^ n5750 ;
  assign n29466 = n21706 ^ n4671 ^ 1'b0 ;
  assign n29467 = n12885 ^ n5448 ^ n1181 ;
  assign n29468 = n6148 & ~n29467 ;
  assign n29470 = ( n1312 & n7234 ) | ( n1312 & n18347 ) | ( n7234 & n18347 ) ;
  assign n29471 = ( n4011 & n5576 ) | ( n4011 & n29470 ) | ( n5576 & n29470 ) ;
  assign n29469 = n4664 & ~n8183 ;
  assign n29472 = n29471 ^ n29469 ^ 1'b0 ;
  assign n29473 = n2741 & ~n29472 ;
  assign n29474 = n29473 ^ n10177 ^ 1'b0 ;
  assign n29475 = n10129 ^ n7718 ^ n2070 ;
  assign n29476 = n6454 ^ n3061 ^ 1'b0 ;
  assign n29477 = ( n20175 & ~n29475 ) | ( n20175 & n29476 ) | ( ~n29475 & n29476 ) ;
  assign n29478 = n29477 ^ n17759 ^ n6525 ;
  assign n29479 = ( n4353 & ~n7599 ) | ( n4353 & n12024 ) | ( ~n7599 & n12024 ) ;
  assign n29480 = ( n8614 & n10106 ) | ( n8614 & ~n11605 ) | ( n10106 & ~n11605 ) ;
  assign n29481 = ( n4697 & n6648 ) | ( n4697 & n29480 ) | ( n6648 & n29480 ) ;
  assign n29482 = ( ~n2249 & n9283 ) | ( ~n2249 & n25372 ) | ( n9283 & n25372 ) ;
  assign n29483 = n29482 ^ n28049 ^ n24877 ;
  assign n29484 = ( n4567 & n7290 ) | ( n4567 & n29483 ) | ( n7290 & n29483 ) ;
  assign n29485 = n13183 ^ n7920 ^ n7111 ;
  assign n29486 = n18830 ^ n3352 ^ n1021 ;
  assign n29487 = n29486 ^ n19305 ^ 1'b0 ;
  assign n29488 = ( ~n2805 & n12576 ) | ( ~n2805 & n29487 ) | ( n12576 & n29487 ) ;
  assign n29489 = n27819 ^ n2660 ^ 1'b0 ;
  assign n29490 = n29489 ^ n16954 ^ n9872 ;
  assign n29491 = ~n11917 & n24299 ;
  assign n29492 = ~n19799 & n29491 ;
  assign n29493 = ~n9172 & n29492 ;
  assign n29494 = n29370 ^ n16660 ^ 1'b0 ;
  assign n29495 = n19529 & n29494 ;
  assign n29496 = n16873 & ~n20312 ;
  assign n29497 = n19147 ^ n141 ^ 1'b0 ;
  assign n29498 = ~n13956 & n29497 ;
  assign n29499 = ~n523 & n5679 ;
  assign n29500 = n28713 ^ n14841 ^ 1'b0 ;
  assign n29502 = n21753 ^ n2187 ^ 1'b0 ;
  assign n29501 = ( n3326 & ~n16420 ) | ( n3326 & n28488 ) | ( ~n16420 & n28488 ) ;
  assign n29503 = n29502 ^ n29501 ^ n16619 ;
  assign n29504 = n1927 & n19111 ;
  assign n29505 = n29504 ^ n7900 ^ n738 ;
  assign n29506 = n29505 ^ n27742 ^ 1'b0 ;
  assign n29507 = n13596 | n28781 ;
  assign n29508 = n6271 & ~n29507 ;
  assign n29509 = n23196 & n29508 ;
  assign n29510 = n29509 ^ n26638 ^ n10988 ;
  assign n29511 = n8785 | n12565 ;
  assign n29512 = n29511 ^ n3410 ^ 1'b0 ;
  assign n29513 = n29512 ^ n14603 ^ n1414 ;
  assign n29514 = ( n1046 & ~n6198 ) | ( n1046 & n17703 ) | ( ~n6198 & n17703 ) ;
  assign n29515 = n29514 ^ n22553 ^ n4750 ;
  assign n29516 = n27693 ^ n10483 ^ 1'b0 ;
  assign n29517 = n8597 & n29516 ;
  assign n29518 = ( n23991 & ~n29515 ) | ( n23991 & n29517 ) | ( ~n29515 & n29517 ) ;
  assign n29519 = n11998 ^ n9501 ^ 1'b0 ;
  assign n29520 = n27755 & ~n28864 ;
  assign n29521 = n29520 ^ n13367 ^ 1'b0 ;
  assign n29522 = n10231 ^ n3687 ^ 1'b0 ;
  assign n29523 = ~n12618 & n29522 ;
  assign n29524 = ( x2 & ~n9100 ) | ( x2 & n11086 ) | ( ~n9100 & n11086 ) ;
  assign n29525 = n29524 ^ n3792 ^ n3029 ;
  assign n29526 = ( n10256 & n14073 ) | ( n10256 & ~n24292 ) | ( n14073 & ~n24292 ) ;
  assign n29533 = ( n811 & ~n1628 ) | ( n811 & n2906 ) | ( ~n1628 & n2906 ) ;
  assign n29534 = ( n11432 & n12697 ) | ( n11432 & n29533 ) | ( n12697 & n29533 ) ;
  assign n29531 = n24996 ^ n10243 ^ 1'b0 ;
  assign n29528 = n12314 ^ n3389 ^ n3081 ;
  assign n29529 = n29528 ^ n12090 ^ n10996 ;
  assign n29527 = n3847 ^ n1736 ^ x65 ;
  assign n29530 = n29529 ^ n29527 ^ n15806 ;
  assign n29532 = n29531 ^ n29530 ^ n12730 ;
  assign n29535 = n29534 ^ n29532 ^ n29046 ;
  assign n29536 = ( ~n9676 & n17122 ) | ( ~n9676 & n29535 ) | ( n17122 & n29535 ) ;
  assign n29537 = n9741 | n18020 ;
  assign n29538 = ( ~n6783 & n10907 ) | ( ~n6783 & n13352 ) | ( n10907 & n13352 ) ;
  assign n29539 = n15691 | n29538 ;
  assign n29540 = n21673 ^ n13524 ^ 1'b0 ;
  assign n29541 = ( ~n5372 & n18506 ) | ( ~n5372 & n29540 ) | ( n18506 & n29540 ) ;
  assign n29542 = n17496 & n26638 ;
  assign n29543 = n19646 ^ n2016 ^ 1'b0 ;
  assign n29545 = n20168 ^ n3361 ^ n889 ;
  assign n29546 = n2502 | n29545 ;
  assign n29547 = n19773 & ~n29546 ;
  assign n29548 = ( ~n16438 & n26620 ) | ( ~n16438 & n29547 ) | ( n26620 & n29547 ) ;
  assign n29544 = n278 & n17786 ;
  assign n29549 = n29548 ^ n29544 ^ 1'b0 ;
  assign n29550 = ~n3214 & n29549 ;
  assign n29551 = ~n29543 & n29550 ;
  assign n29552 = n6814 ^ n374 ^ 1'b0 ;
  assign n29553 = n10521 ^ n5022 ^ 1'b0 ;
  assign n29554 = n16719 & ~n29553 ;
  assign n29555 = n12388 & n16352 ;
  assign n29556 = n6215 | n29555 ;
  assign n29557 = n3908 & ~n7627 ;
  assign n29558 = n6136 ^ n4040 ^ n2607 ;
  assign n29559 = ( n3842 & n17671 ) | ( n3842 & ~n19555 ) | ( n17671 & ~n19555 ) ;
  assign n29560 = n28729 ^ n20456 ^ n19404 ;
  assign n29561 = ( n2702 & n11278 ) | ( n2702 & n28030 ) | ( n11278 & n28030 ) ;
  assign n29562 = n26106 ^ n9354 ^ n1461 ;
  assign n29563 = ( n11147 & n22573 ) | ( n11147 & ~n29562 ) | ( n22573 & ~n29562 ) ;
  assign n29564 = n8087 ^ n4630 ^ n1765 ;
  assign n29565 = n16802 ^ n16281 ^ 1'b0 ;
  assign n29566 = ~n29564 & n29565 ;
  assign n29567 = n3033 | n18325 ;
  assign n29568 = n29567 ^ n19072 ^ 1'b0 ;
  assign n29569 = n14542 | n15768 ;
  assign n29570 = n29568 & ~n29569 ;
  assign n29571 = n16864 ^ n10568 ^ 1'b0 ;
  assign n29572 = n8246 & ~n29571 ;
  assign n29573 = n8546 & n28383 ;
  assign n29574 = n27692 ^ n26434 ^ n5037 ;
  assign n29575 = n29573 & n29574 ;
  assign n29576 = ( n8290 & ~n16612 ) | ( n8290 & n16857 ) | ( ~n16612 & n16857 ) ;
  assign n29577 = n16611 ^ n4006 ^ 1'b0 ;
  assign n29578 = ( n12520 & n22029 ) | ( n12520 & n25741 ) | ( n22029 & n25741 ) ;
  assign n29579 = ( n6227 & n29256 ) | ( n6227 & ~n29578 ) | ( n29256 & ~n29578 ) ;
  assign n29580 = n20742 ^ n7757 ^ 1'b0 ;
  assign n29581 = ~n1744 & n29580 ;
  assign n29582 = n29581 ^ n29164 ^ n4474 ;
  assign n29583 = n25988 ^ n12534 ^ n5177 ;
  assign n29584 = n2842 | n16123 ;
  assign n29585 = n19881 ^ n10840 ^ 1'b0 ;
  assign n29586 = n6289 | n29585 ;
  assign n29587 = ( n9600 & ~n29584 ) | ( n9600 & n29586 ) | ( ~n29584 & n29586 ) ;
  assign n29588 = ( ~n12606 & n29583 ) | ( ~n12606 & n29587 ) | ( n29583 & n29587 ) ;
  assign n29591 = n24756 ^ n15142 ^ 1'b0 ;
  assign n29589 = n10554 & ~n18336 ;
  assign n29590 = ( n1332 & ~n7323 ) | ( n1332 & n29589 ) | ( ~n7323 & n29589 ) ;
  assign n29592 = n29591 ^ n29590 ^ n17871 ;
  assign n29593 = n29592 ^ n21012 ^ n7818 ;
  assign n29594 = n755 & ~n15660 ;
  assign n29595 = ~n5043 & n19490 ;
  assign n29596 = n29594 & n29595 ;
  assign n29597 = n1747 | n29596 ;
  assign n29598 = n29597 ^ n22292 ^ 1'b0 ;
  assign n29599 = ( n1466 & n2501 ) | ( n1466 & ~n18149 ) | ( n2501 & ~n18149 ) ;
  assign n29600 = n29599 ^ n13596 ^ 1'b0 ;
  assign n29601 = n473 & ~n19022 ;
  assign n29602 = n5706 & ~n27404 ;
  assign n29603 = n23310 & n29602 ;
  assign n29604 = n20628 ^ n15211 ^ n1813 ;
  assign n29605 = ( n4964 & n9984 ) | ( n4964 & n28577 ) | ( n9984 & n28577 ) ;
  assign n29606 = ( n4486 & n7287 ) | ( n4486 & ~n14846 ) | ( n7287 & ~n14846 ) ;
  assign n29607 = ( ~n15522 & n16318 ) | ( ~n15522 & n29606 ) | ( n16318 & n29606 ) ;
  assign n29608 = ~n11004 & n26095 ;
  assign n29609 = ~n12464 & n29608 ;
  assign n29610 = n29609 ^ n19536 ^ n14669 ;
  assign n29611 = n7589 ^ n7204 ^ n6541 ;
  assign n29612 = ( n5222 & n5371 ) | ( n5222 & ~n10440 ) | ( n5371 & ~n10440 ) ;
  assign n29613 = ( n1744 & ~n20868 ) | ( n1744 & n29612 ) | ( ~n20868 & n29612 ) ;
  assign n29614 = ( n7171 & n16066 ) | ( n7171 & ~n18131 ) | ( n16066 & ~n18131 ) ;
  assign n29615 = n5429 ^ n4105 ^ n2946 ;
  assign n29616 = n29615 ^ n15729 ^ 1'b0 ;
  assign n29617 = n3970 & ~n24519 ;
  assign n29618 = ~n29616 & n29617 ;
  assign n29619 = n28513 ^ n26839 ^ n12034 ;
  assign n29620 = n29619 ^ n25998 ^ 1'b0 ;
  assign n29621 = n7220 & ~n29620 ;
  assign n29622 = n24731 ^ n11807 ^ n10664 ;
  assign n29623 = n4719 & ~n29622 ;
  assign n29624 = n16295 & n29623 ;
  assign n29625 = n6237 & ~n27179 ;
  assign n29626 = n29625 ^ n11838 ^ n5999 ;
  assign n29627 = n11197 ^ n2976 ^ 1'b0 ;
  assign n29628 = n13628 & n29627 ;
  assign n29629 = ( n9179 & n19507 ) | ( n9179 & n29628 ) | ( n19507 & n29628 ) ;
  assign n29630 = n9780 ^ n3643 ^ n2345 ;
  assign n29631 = ( n4899 & n8136 ) | ( n4899 & n29630 ) | ( n8136 & n29630 ) ;
  assign n29632 = n13881 ^ n3509 ^ n3139 ;
  assign n29633 = n29631 | n29632 ;
  assign n29634 = ( ~n7579 & n12681 ) | ( ~n7579 & n29633 ) | ( n12681 & n29633 ) ;
  assign n29635 = n29634 ^ n1341 ^ 1'b0 ;
  assign n29636 = ~n1780 & n29635 ;
  assign n29637 = n29636 ^ n28576 ^ n13392 ;
  assign n29638 = ( ~n2225 & n13215 ) | ( ~n2225 & n15936 ) | ( n13215 & n15936 ) ;
  assign n29639 = ( n1739 & n22812 ) | ( n1739 & n29638 ) | ( n22812 & n29638 ) ;
  assign n29647 = ( n6333 & n17247 ) | ( n6333 & ~n18516 ) | ( n17247 & ~n18516 ) ;
  assign n29648 = n29647 ^ n24589 ^ n7628 ;
  assign n29645 = n8175 & n8259 ;
  assign n29646 = ~n25349 & n29645 ;
  assign n29640 = n1738 & ~n10057 ;
  assign n29641 = n29640 ^ n6696 ^ 1'b0 ;
  assign n29642 = ( n4159 & n7759 ) | ( n4159 & n29641 ) | ( n7759 & n29641 ) ;
  assign n29643 = n29642 ^ n8669 ^ n7395 ;
  assign n29644 = n12396 | n29643 ;
  assign n29649 = n29648 ^ n29646 ^ n29644 ;
  assign n29650 = n15452 ^ n5324 ^ 1'b0 ;
  assign n29651 = n8491 & ~n29650 ;
  assign n29652 = n29651 ^ n19525 ^ n10026 ;
  assign n29653 = n4015 & n19191 ;
  assign n29654 = ( n8876 & n29652 ) | ( n8876 & ~n29653 ) | ( n29652 & ~n29653 ) ;
  assign n29655 = n21036 ^ n11855 ^ n11827 ;
  assign n29656 = n19028 ^ n3702 ^ 1'b0 ;
  assign n29657 = n29655 & ~n29656 ;
  assign n29658 = n29657 ^ n4671 ^ 1'b0 ;
  assign n29659 = n16507 ^ n4143 ^ n1965 ;
  assign n29660 = n3657 | n29659 ;
  assign n29661 = n3602 | n17253 ;
  assign n29662 = ( n1519 & n17624 ) | ( n1519 & n21677 ) | ( n17624 & n21677 ) ;
  assign n29663 = n3966 & ~n29662 ;
  assign n29664 = n29663 ^ n513 ^ 1'b0 ;
  assign n29665 = ( n5735 & ~n12140 ) | ( n5735 & n27350 ) | ( ~n12140 & n27350 ) ;
  assign n29666 = ( n19249 & n27381 ) | ( n19249 & ~n29665 ) | ( n27381 & ~n29665 ) ;
  assign n29667 = n8043 ^ n3438 ^ 1'b0 ;
  assign n29668 = ~n5993 & n29667 ;
  assign n29669 = n29668 ^ n16071 ^ n740 ;
  assign n29670 = ( n6703 & ~n10275 ) | ( n6703 & n29669 ) | ( ~n10275 & n29669 ) ;
  assign n29671 = n28884 ^ n12697 ^ n10201 ;
  assign n29672 = ( n1608 & n3453 ) | ( n1608 & ~n23826 ) | ( n3453 & ~n23826 ) ;
  assign n29673 = ( n2221 & n11934 ) | ( n2221 & n29672 ) | ( n11934 & n29672 ) ;
  assign n29674 = n5921 ^ n2485 ^ 1'b0 ;
  assign n29675 = n16231 & n23051 ;
  assign n29676 = n21849 & n29675 ;
  assign n29677 = n29676 ^ n20889 ^ n847 ;
  assign n29678 = ( ~n20522 & n29674 ) | ( ~n20522 & n29677 ) | ( n29674 & n29677 ) ;
  assign n29679 = ( n2234 & ~n2804 ) | ( n2234 & n3117 ) | ( ~n2804 & n3117 ) ;
  assign n29680 = n28467 ^ n21012 ^ n16768 ;
  assign n29681 = n20915 ^ n4986 ^ 1'b0 ;
  assign n29682 = n14682 ^ n12331 ^ n5117 ;
  assign n29683 = n29682 ^ n23802 ^ n2375 ;
  assign n29684 = n24457 ^ n3032 ^ 1'b0 ;
  assign n29685 = n29683 & n29684 ;
  assign n29686 = ~n1020 & n5180 ;
  assign n29687 = ~n29685 & n29686 ;
  assign n29688 = ( n14068 & n17729 ) | ( n14068 & n27188 ) | ( n17729 & n27188 ) ;
  assign n29689 = n28387 ^ n24295 ^ n22475 ;
  assign n29690 = n676 & n3415 ;
  assign n29691 = ~n8105 & n29690 ;
  assign n29692 = ( n12189 & n16063 ) | ( n12189 & n29691 ) | ( n16063 & n29691 ) ;
  assign n29693 = n3316 ^ n2622 ^ 1'b0 ;
  assign n29694 = n29693 ^ n3224 ^ n1982 ;
  assign n29695 = n451 & ~n8956 ;
  assign n29696 = n29695 ^ n3410 ^ 1'b0 ;
  assign n29697 = n29696 ^ n25579 ^ 1'b0 ;
  assign n29698 = n2155 ^ x45 ^ 1'b0 ;
  assign n29699 = ~n29697 & n29698 ;
  assign n29700 = ~n16796 & n19010 ;
  assign n29701 = n29700 ^ n5450 ^ 1'b0 ;
  assign n29702 = ( n8080 & ~n12040 ) | ( n8080 & n29701 ) | ( ~n12040 & n29701 ) ;
  assign n29703 = n29702 ^ n24244 ^ 1'b0 ;
  assign n29704 = n8897 & ~n16978 ;
  assign n29705 = n29704 ^ n21370 ^ n1059 ;
  assign n29706 = n23108 ^ n1186 ^ 1'b0 ;
  assign n29707 = n21144 & n23570 ;
  assign n29708 = n25039 ^ n1851 ^ 1'b0 ;
  assign n29709 = n29707 | n29708 ;
  assign n29710 = n29190 ^ n27388 ^ n24225 ;
  assign n29711 = ~n3574 & n29710 ;
  assign n29712 = ( n2295 & n29709 ) | ( n2295 & ~n29711 ) | ( n29709 & ~n29711 ) ;
  assign n29713 = n21230 ^ n15716 ^ 1'b0 ;
  assign n29714 = n8916 ^ n8240 ^ x50 ;
  assign n29715 = ( n2707 & n5295 ) | ( n2707 & ~n29714 ) | ( n5295 & ~n29714 ) ;
  assign n29716 = n11960 ^ n9137 ^ n8023 ;
  assign n29717 = ( n1140 & n13190 ) | ( n1140 & n29716 ) | ( n13190 & n29716 ) ;
  assign n29718 = ~n2458 & n13924 ;
  assign n29719 = ~n22774 & n29718 ;
  assign n29720 = n29719 ^ n7860 ^ 1'b0 ;
  assign n29721 = n18908 & ~n29720 ;
  assign n29722 = n21085 ^ n17881 ^ 1'b0 ;
  assign n29723 = n18466 & n29722 ;
  assign n29725 = n3173 ^ n2337 ^ 1'b0 ;
  assign n29726 = ~n2838 & n29725 ;
  assign n29724 = n8276 & ~n22951 ;
  assign n29727 = n29726 ^ n29724 ^ 1'b0 ;
  assign n29728 = ~n8984 & n26261 ;
  assign n29729 = ( ~n468 & n9055 ) | ( ~n468 & n29728 ) | ( n9055 & n29728 ) ;
  assign n29730 = ( n1271 & n14464 ) | ( n1271 & ~n29729 ) | ( n14464 & ~n29729 ) ;
  assign n29731 = n13477 ^ n374 ^ 1'b0 ;
  assign n29734 = n8059 ^ n4604 ^ 1'b0 ;
  assign n29735 = n22172 & ~n29734 ;
  assign n29736 = ~n20736 & n29735 ;
  assign n29737 = n3190 & n29736 ;
  assign n29732 = n25932 ^ n3991 ^ n1260 ;
  assign n29733 = n29732 ^ n13728 ^ n1778 ;
  assign n29738 = n29737 ^ n29733 ^ n18400 ;
  assign n29739 = ( n16196 & ~n29731 ) | ( n16196 & n29738 ) | ( ~n29731 & n29738 ) ;
  assign n29740 = ~n2685 & n12978 ;
  assign n29746 = n21656 ^ n10199 ^ 1'b0 ;
  assign n29741 = ~x108 & n3711 ;
  assign n29742 = n27745 & n29741 ;
  assign n29743 = n10386 & n29742 ;
  assign n29744 = n29743 ^ n24712 ^ n17160 ;
  assign n29745 = n10358 & n29744 ;
  assign n29747 = n29746 ^ n29745 ^ n22306 ;
  assign n29748 = n17837 ^ n16540 ^ 1'b0 ;
  assign n29749 = ~n16751 & n29748 ;
  assign n29750 = ( ~n20720 & n28348 ) | ( ~n20720 & n29749 ) | ( n28348 & n29749 ) ;
  assign n29751 = ( n6158 & ~n17965 ) | ( n6158 & n23970 ) | ( ~n17965 & n23970 ) ;
  assign n29752 = ( n360 & ~n12011 ) | ( n360 & n29751 ) | ( ~n12011 & n29751 ) ;
  assign n29753 = ( n6278 & n8105 ) | ( n6278 & ~n26953 ) | ( n8105 & ~n26953 ) ;
  assign n29754 = ( n3905 & ~n9317 ) | ( n3905 & n11044 ) | ( ~n9317 & n11044 ) ;
  assign n29755 = n5812 & ~n29754 ;
  assign n29756 = ( n17031 & ~n29753 ) | ( n17031 & n29755 ) | ( ~n29753 & n29755 ) ;
  assign n29757 = n20086 ^ n3937 ^ 1'b0 ;
  assign n29758 = n4869 & n29757 ;
  assign n29759 = n3782 | n7311 ;
  assign n29760 = n25496 & ~n29759 ;
  assign n29761 = ~n3039 & n11856 ;
  assign n29762 = n29761 ^ n13132 ^ 1'b0 ;
  assign n29763 = ( n3174 & n18615 ) | ( n3174 & ~n29762 ) | ( n18615 & ~n29762 ) ;
  assign n29764 = n17031 ^ n2075 ^ n1167 ;
  assign n29765 = n29764 ^ x92 ^ 1'b0 ;
  assign n29766 = ~n21600 & n29765 ;
  assign n29767 = n21849 & n29766 ;
  assign n29768 = n12004 ^ n5824 ^ n3610 ;
  assign n29769 = n16877 & n29768 ;
  assign n29770 = n20579 ^ n379 ^ 1'b0 ;
  assign n29771 = n139 & ~n29770 ;
  assign n29772 = n29771 ^ n19681 ^ 1'b0 ;
  assign n29773 = n27511 ^ n12562 ^ n9072 ;
  assign n29775 = n2498 & ~n9597 ;
  assign n29776 = n8702 ^ n5316 ^ n1994 ;
  assign n29777 = ~n13715 & n29776 ;
  assign n29778 = ( n4048 & n29775 ) | ( n4048 & n29777 ) | ( n29775 & n29777 ) ;
  assign n29774 = n472 & ~n3619 ;
  assign n29779 = n29778 ^ n29774 ^ n3179 ;
  assign n29780 = n1624 | n17798 ;
  assign n29781 = ~n3817 & n29780 ;
  assign n29782 = n21667 ^ n8038 ^ n2667 ;
  assign n29783 = n3140 & ~n29782 ;
  assign n29784 = n29783 ^ n19344 ^ 1'b0 ;
  assign n29785 = n6347 ^ n4740 ^ n858 ;
  assign n29786 = n3418 | n29785 ;
  assign n29787 = n1107 | n29786 ;
  assign n29788 = n8918 & n13690 ;
  assign n29789 = n29788 ^ n8855 ^ 1'b0 ;
  assign n29790 = ( n1483 & n10918 ) | ( n1483 & n24153 ) | ( n10918 & n24153 ) ;
  assign n29791 = n12862 & ~n19256 ;
  assign n29792 = n11351 ^ n8970 ^ n369 ;
  assign n29793 = n29792 ^ n26292 ^ n6471 ;
  assign n29794 = ( ~n1410 & n15934 ) | ( ~n1410 & n21121 ) | ( n15934 & n21121 ) ;
  assign n29798 = n4896 ^ n1201 ^ 1'b0 ;
  assign n29799 = ( n1293 & ~n27831 ) | ( n1293 & n29798 ) | ( ~n27831 & n29798 ) ;
  assign n29796 = n24067 ^ n14392 ^ n7896 ;
  assign n29795 = n25708 ^ n24283 ^ n7628 ;
  assign n29797 = n29796 ^ n29795 ^ n14704 ;
  assign n29800 = n29799 ^ n29797 ^ n10267 ;
  assign n29802 = n11383 ^ n2478 ^ 1'b0 ;
  assign n29801 = n6352 & ~n24636 ;
  assign n29803 = n29802 ^ n29801 ^ n23395 ;
  assign n29804 = ~n11739 & n15448 ;
  assign n29805 = n7476 & ~n8753 ;
  assign n29806 = ( n5106 & ~n16069 ) | ( n5106 & n16563 ) | ( ~n16069 & n16563 ) ;
  assign n29807 = ~n10840 & n29806 ;
  assign n29808 = n3227 ^ n1992 ^ 1'b0 ;
  assign n29809 = ~n13378 & n29808 ;
  assign n29811 = ( ~n7475 & n8811 ) | ( ~n7475 & n28979 ) | ( n8811 & n28979 ) ;
  assign n29810 = n11914 ^ n3395 ^ 1'b0 ;
  assign n29812 = n29811 ^ n29810 ^ n29254 ;
  assign n29813 = n29812 ^ n14446 ^ 1'b0 ;
  assign n29814 = n2145 & ~n15423 ;
  assign n29815 = n29000 ^ n19881 ^ n12699 ;
  assign n29816 = ( n8049 & n8097 ) | ( n8049 & ~n23967 ) | ( n8097 & ~n23967 ) ;
  assign n29817 = n16249 ^ n10023 ^ 1'b0 ;
  assign n29818 = ( n7698 & ~n11882 ) | ( n7698 & n29199 ) | ( ~n11882 & n29199 ) ;
  assign n29820 = n14335 ^ n13400 ^ 1'b0 ;
  assign n29821 = ~n16365 & n29820 ;
  assign n29819 = n20867 ^ n12326 ^ 1'b0 ;
  assign n29822 = n29821 ^ n29819 ^ n27436 ;
  assign n29823 = n460 | n26550 ;
  assign n29824 = n29823 ^ n12288 ^ 1'b0 ;
  assign n29825 = n12382 ^ n2977 ^ n2908 ;
  assign n29826 = n10497 & ~n11683 ;
  assign n29827 = ~n29825 & n29826 ;
  assign n29828 = n3347 | n29827 ;
  assign n29829 = n29828 ^ n10680 ^ n516 ;
  assign n29830 = ( ~n954 & n24996 ) | ( ~n954 & n29829 ) | ( n24996 & n29829 ) ;
  assign n29831 = n14556 & ~n29830 ;
  assign n29832 = n29831 ^ n15467 ^ 1'b0 ;
  assign n29833 = n4151 & ~n21747 ;
  assign n29834 = n18393 & n29833 ;
  assign n29835 = ( n2239 & ~n7806 ) | ( n2239 & n18358 ) | ( ~n7806 & n18358 ) ;
  assign n29836 = n29835 ^ n16087 ^ n5524 ;
  assign n29837 = n2457 & ~n2600 ;
  assign n29838 = ~n11218 & n29837 ;
  assign n29839 = n29838 ^ n14295 ^ n4537 ;
  assign n29840 = n29839 ^ n22792 ^ n15034 ;
  assign n29841 = n20451 ^ n7777 ^ n607 ;
  assign n29843 = n13712 ^ n240 ^ 1'b0 ;
  assign n29842 = n10481 & ~n11362 ;
  assign n29844 = n29843 ^ n29842 ^ n9534 ;
  assign n29845 = ~n1917 & n11371 ;
  assign n29846 = ( ~n2219 & n3995 ) | ( ~n2219 & n6797 ) | ( n3995 & n6797 ) ;
  assign n29847 = ( n6466 & n13215 ) | ( n6466 & n29846 ) | ( n13215 & n29846 ) ;
  assign n29848 = n3316 & ~n9118 ;
  assign n29849 = n29847 & n29848 ;
  assign n29850 = n2707 & ~n3899 ;
  assign n29851 = n29850 ^ n1727 ^ 1'b0 ;
  assign n29852 = ~n4536 & n12943 ;
  assign n29853 = n29852 ^ n28315 ^ 1'b0 ;
  assign n29854 = n16528 ^ n14429 ^ n3237 ;
  assign n29855 = n29854 ^ n8437 ^ n6492 ;
  assign n29856 = n11596 & ~n15121 ;
  assign n29857 = n19116 & n29856 ;
  assign n29858 = n29857 ^ n23817 ^ n9722 ;
  assign n29859 = n23195 ^ n9921 ^ n734 ;
  assign n29860 = ( n16071 & n20349 ) | ( n16071 & n29859 ) | ( n20349 & n29859 ) ;
  assign n29861 = ( n11002 & n13307 ) | ( n11002 & n29860 ) | ( n13307 & n29860 ) ;
  assign n29862 = ( ~n4129 & n11246 ) | ( ~n4129 & n20614 ) | ( n11246 & n20614 ) ;
  assign n29863 = n29862 ^ n8652 ^ 1'b0 ;
  assign n29864 = n16437 | n20706 ;
  assign n29865 = n29864 ^ n15537 ^ n7735 ;
  assign n29866 = n22406 ^ n14760 ^ n13875 ;
  assign n29867 = n11988 & ~n29866 ;
  assign n29868 = n23214 ^ n13328 ^ n11322 ;
  assign n29869 = n15520 ^ n746 ^ x2 ;
  assign n29870 = ~n9718 & n29869 ;
  assign n29871 = n29868 & n29870 ;
  assign n29872 = n10575 & n13073 ;
  assign n29873 = ~n11737 & n29872 ;
  assign n29874 = n21750 ^ n18820 ^ n6768 ;
  assign n29875 = n24523 ^ n19087 ^ n3347 ;
  assign n29876 = ( n616 & ~n3752 ) | ( n616 & n29369 ) | ( ~n3752 & n29369 ) ;
  assign n29877 = n22235 & ~n26247 ;
  assign n29878 = ( n2875 & n2995 ) | ( n2875 & ~n3232 ) | ( n2995 & ~n3232 ) ;
  assign n29879 = n29878 ^ n20812 ^ n3226 ;
  assign n29880 = n18832 ^ n4007 ^ x115 ;
  assign n29881 = n24462 | n29880 ;
  assign n29882 = n20349 ^ n12312 ^ n9072 ;
  assign n29883 = n7692 ^ n3000 ^ n362 ;
  assign n29884 = n6474 | n10640 ;
  assign n29885 = n29883 | n29884 ;
  assign n29886 = ( n8919 & n10579 ) | ( n8919 & n14228 ) | ( n10579 & n14228 ) ;
  assign n29887 = ( ~n1088 & n26942 ) | ( ~n1088 & n29886 ) | ( n26942 & n29886 ) ;
  assign n29888 = n29887 ^ n25066 ^ n8869 ;
  assign n29889 = n6268 | n14396 ;
  assign n29890 = n29888 & ~n29889 ;
  assign n29891 = n300 & n8696 ;
  assign n29892 = n29891 ^ n7312 ^ 1'b0 ;
  assign n29893 = ~n11763 & n14259 ;
  assign n29894 = n29893 ^ n16728 ^ 1'b0 ;
  assign n29895 = n7309 ^ n3543 ^ 1'b0 ;
  assign n29896 = n425 & ~n29895 ;
  assign n29897 = ( ~n4165 & n8413 ) | ( ~n4165 & n29896 ) | ( n8413 & n29896 ) ;
  assign n29898 = ( n11691 & ~n19246 ) | ( n11691 & n26344 ) | ( ~n19246 & n26344 ) ;
  assign n29899 = n234 & n29898 ;
  assign n29900 = ~n4570 & n6308 ;
  assign n29901 = ~n1989 & n29900 ;
  assign n29902 = n24798 ^ n2581 ^ 1'b0 ;
  assign n29903 = n28884 ^ n22110 ^ n15563 ;
  assign n29904 = ( ~n29901 & n29902 ) | ( ~n29901 & n29903 ) | ( n29902 & n29903 ) ;
  assign n29905 = n6684 & n7449 ;
  assign n29906 = n29905 ^ n12835 ^ n3272 ;
  assign n29907 = n5471 & ~n8041 ;
  assign n29908 = n29907 ^ n13198 ^ 1'b0 ;
  assign n29909 = n29908 ^ n5385 ^ x81 ;
  assign n29910 = n7641 & n16471 ;
  assign n29911 = n25583 | n29910 ;
  assign n29912 = n27689 ^ n19255 ^ 1'b0 ;
  assign n29913 = ~n1773 & n29912 ;
  assign n29914 = n27835 ^ n9943 ^ n5751 ;
  assign n29915 = ( n8286 & ~n8412 ) | ( n8286 & n29914 ) | ( ~n8412 & n29914 ) ;
  assign n29916 = n947 | n18243 ;
  assign n29917 = ( n7818 & n24327 ) | ( n7818 & n26345 ) | ( n24327 & n26345 ) ;
  assign n29918 = ( n9410 & n11585 ) | ( n9410 & n29917 ) | ( n11585 & n29917 ) ;
  assign n29919 = n19080 ^ n17922 ^ n6900 ;
  assign n29920 = n22632 ^ n15570 ^ 1'b0 ;
  assign n29921 = n29920 ^ n25596 ^ n2047 ;
  assign n29922 = n23735 ^ n14215 ^ n14186 ;
  assign n29923 = n29922 ^ n17644 ^ 1'b0 ;
  assign n29924 = ( n13584 & ~n18876 ) | ( n13584 & n22268 ) | ( ~n18876 & n22268 ) ;
  assign n29925 = ( n13707 & ~n29923 ) | ( n13707 & n29924 ) | ( ~n29923 & n29924 ) ;
  assign n29926 = n29925 ^ n12695 ^ 1'b0 ;
  assign n29927 = n29019 ^ n19799 ^ 1'b0 ;
  assign n29928 = n23881 & ~n29927 ;
  assign n29929 = n15564 ^ n9019 ^ n6591 ;
  assign n29930 = n29929 ^ n19979 ^ n5797 ;
  assign n29931 = n8015 ^ n5321 ^ n1394 ;
  assign n29932 = n29930 & ~n29931 ;
  assign n29933 = ( n7661 & ~n16147 ) | ( n7661 & n17408 ) | ( ~n16147 & n17408 ) ;
  assign n29934 = ( n5269 & ~n9079 ) | ( n5269 & n29933 ) | ( ~n9079 & n29933 ) ;
  assign n29936 = n984 & ~n20736 ;
  assign n29937 = n29936 ^ n4984 ^ 1'b0 ;
  assign n29935 = n21132 ^ n16587 ^ n9736 ;
  assign n29938 = n29937 ^ n29935 ^ n6209 ;
  assign n29939 = n25529 ^ n24987 ^ n6830 ;
  assign n29940 = n29939 ^ n11150 ^ n4130 ;
  assign n29941 = ( n3922 & n8809 ) | ( n3922 & ~n20274 ) | ( n8809 & ~n20274 ) ;
  assign n29942 = ( n4100 & n14047 ) | ( n4100 & n29941 ) | ( n14047 & n29941 ) ;
  assign n29943 = ( n15352 & n16242 ) | ( n15352 & n18355 ) | ( n16242 & n18355 ) ;
  assign n29944 = ( ~n3790 & n10200 ) | ( ~n3790 & n12351 ) | ( n10200 & n12351 ) ;
  assign n29945 = ( n4139 & n5434 ) | ( n4139 & ~n21479 ) | ( n5434 & ~n21479 ) ;
  assign n29946 = n29945 ^ n29189 ^ 1'b0 ;
  assign n29947 = n423 & ~n20678 ;
  assign n29948 = n20184 ^ n10699 ^ n633 ;
  assign n29949 = n17332 ^ n17264 ^ n14545 ;
  assign n29950 = ( n3916 & n10765 ) | ( n3916 & ~n11833 ) | ( n10765 & ~n11833 ) ;
  assign n29951 = ( n1705 & n29949 ) | ( n1705 & ~n29950 ) | ( n29949 & ~n29950 ) ;
  assign n29952 = n16253 | n29951 ;
  assign n29953 = n10421 ^ n217 ^ 1'b0 ;
  assign n29954 = n14476 ^ n7692 ^ n4581 ;
  assign n29955 = ( n25165 & n29953 ) | ( n25165 & n29954 ) | ( n29953 & n29954 ) ;
  assign n29956 = n14161 & ~n17891 ;
  assign n29957 = n21341 ^ n13975 ^ n1761 ;
  assign n29958 = n1416 | n5766 ;
  assign n29959 = n16576 | n29958 ;
  assign n29960 = ( n12475 & n29019 ) | ( n12475 & n29959 ) | ( n29019 & n29959 ) ;
  assign n29961 = n3600 & ~n19073 ;
  assign n29962 = ~n486 & n29961 ;
  assign n29963 = ~n10355 & n20501 ;
  assign n29964 = n3604 & n29963 ;
  assign n29965 = n14692 & ~n17645 ;
  assign n29966 = n21241 ^ n19842 ^ n16966 ;
  assign n29967 = ( n22509 & n29965 ) | ( n22509 & ~n29966 ) | ( n29965 & ~n29966 ) ;
  assign n29968 = n14792 ^ n8328 ^ n1874 ;
  assign n29969 = n29968 ^ n16189 ^ n12873 ;
  assign n29970 = n29969 ^ n20124 ^ n7446 ;
  assign n29971 = ( ~n810 & n9292 ) | ( ~n810 & n21028 ) | ( n9292 & n21028 ) ;
  assign n29972 = n29971 ^ n24351 ^ 1'b0 ;
  assign n29973 = ( n1238 & n5305 ) | ( n1238 & ~n15893 ) | ( n5305 & ~n15893 ) ;
  assign n29974 = ( ~n6221 & n11205 ) | ( ~n6221 & n29973 ) | ( n11205 & n29973 ) ;
  assign n29975 = n3623 | n5107 ;
  assign n29976 = n29975 ^ n5136 ^ 1'b0 ;
  assign n29977 = ( n722 & ~n5468 ) | ( n722 & n21651 ) | ( ~n5468 & n21651 ) ;
  assign n29978 = n29977 ^ n6619 ^ 1'b0 ;
  assign n29979 = n29976 & n29978 ;
  assign n29980 = n29979 ^ n21330 ^ n6589 ;
  assign n29981 = n1104 | n12498 ;
  assign n29982 = ( n5894 & n10090 ) | ( n5894 & n29716 ) | ( n10090 & n29716 ) ;
  assign n29983 = ( n4813 & ~n10233 ) | ( n4813 & n29982 ) | ( ~n10233 & n29982 ) ;
  assign n29984 = n24225 & ~n29983 ;
  assign n29985 = n19105 ^ n13819 ^ 1'b0 ;
  assign n29986 = ( n8399 & n13063 ) | ( n8399 & ~n29985 ) | ( n13063 & ~n29985 ) ;
  assign n29987 = n29986 ^ n1915 ^ 1'b0 ;
  assign n29988 = n26678 | n29987 ;
  assign n29989 = ~n15159 & n25122 ;
  assign n29990 = n26778 | n29989 ;
  assign n29991 = n20540 ^ n1948 ^ 1'b0 ;
  assign n29992 = n29990 & n29991 ;
  assign n29993 = n10006 & ~n19558 ;
  assign n29994 = n29993 ^ n14846 ^ 1'b0 ;
  assign n29995 = n16643 ^ n3373 ^ x60 ;
  assign n29996 = ( ~n5820 & n11346 ) | ( ~n5820 & n14392 ) | ( n11346 & n14392 ) ;
  assign n29997 = n4283 & ~n4465 ;
  assign n29998 = n29997 ^ n21323 ^ 1'b0 ;
  assign n29999 = ( ~n20725 & n29427 ) | ( ~n20725 & n29998 ) | ( n29427 & n29998 ) ;
  assign n30000 = n11218 ^ n10552 ^ x53 ;
  assign n30001 = ~n4676 & n30000 ;
  assign n30002 = n7453 & n14060 ;
  assign n30003 = ( n10907 & n12973 ) | ( n10907 & n30002 ) | ( n12973 & n30002 ) ;
  assign n30004 = ( n647 & n30001 ) | ( n647 & ~n30003 ) | ( n30001 & ~n30003 ) ;
  assign n30005 = n6630 & ~n14503 ;
  assign n30006 = n5715 & n30005 ;
  assign n30007 = n30006 ^ n20108 ^ n1537 ;
  assign n30008 = ( n1751 & n7254 ) | ( n1751 & n28632 ) | ( n7254 & n28632 ) ;
  assign n30009 = n30008 ^ n16993 ^ n11837 ;
  assign n30010 = n3111 | n17509 ;
  assign n30011 = n30010 ^ n5621 ^ 1'b0 ;
  assign n30012 = n7250 ^ n3156 ^ 1'b0 ;
  assign n30013 = ~n3798 & n30012 ;
  assign n30014 = n30013 ^ n16738 ^ 1'b0 ;
  assign n30015 = n30011 & ~n30014 ;
  assign n30016 = ( ~n1161 & n21528 ) | ( ~n1161 & n30015 ) | ( n21528 & n30015 ) ;
  assign n30017 = n8259 ^ n6225 ^ n472 ;
  assign n30018 = n30017 ^ n22656 ^ n6448 ;
  assign n30019 = ~n29773 & n30018 ;
  assign n30020 = n30019 ^ n13073 ^ 1'b0 ;
  assign n30021 = ~n3322 & n22810 ;
  assign n30022 = ~n4028 & n30021 ;
  assign n30023 = n2986 | n9556 ;
  assign n30024 = n19235 ^ n16667 ^ 1'b0 ;
  assign n30025 = n30023 | n30024 ;
  assign n30026 = n23480 ^ n15805 ^ n6336 ;
  assign n30027 = n4581 | n30026 ;
  assign n30028 = n10667 & ~n30027 ;
  assign n30029 = n1462 & n18242 ;
  assign n30030 = n4877 & ~n30029 ;
  assign n30031 = ~n26561 & n30030 ;
  assign n30032 = n30031 ^ n23072 ^ n10886 ;
  assign n30034 = n3308 | n6481 ;
  assign n30035 = n6159 | n30034 ;
  assign n30036 = n30035 ^ n8935 ^ n5841 ;
  assign n30033 = n2658 & ~n13905 ;
  assign n30037 = n30036 ^ n30033 ^ 1'b0 ;
  assign n30038 = ( ~n20577 & n21936 ) | ( ~n20577 & n30037 ) | ( n21936 & n30037 ) ;
  assign n30039 = n29524 ^ n13631 ^ n4097 ;
  assign n30040 = ( n5336 & ~n14056 ) | ( n5336 & n29583 ) | ( ~n14056 & n29583 ) ;
  assign n30041 = ~n3622 & n9110 ;
  assign n30042 = ( ~n8333 & n17212 ) | ( ~n8333 & n30041 ) | ( n17212 & n30041 ) ;
  assign n30043 = n8496 ^ n194 ^ 1'b0 ;
  assign n30044 = ~n10066 & n30043 ;
  assign n30045 = x119 & ~n18039 ;
  assign n30046 = n4369 & ~n8266 ;
  assign n30047 = n21919 ^ n13075 ^ 1'b0 ;
  assign n30048 = n10564 | n30047 ;
  assign n30049 = n14254 | n30048 ;
  assign n30050 = n30049 ^ n306 ^ 1'b0 ;
  assign n30051 = ( ~n14644 & n21943 ) | ( ~n14644 & n30050 ) | ( n21943 & n30050 ) ;
  assign n30052 = n8871 & n13234 ;
  assign n30053 = n1470 | n5849 ;
  assign n30054 = n11883 ^ n5854 ^ n1027 ;
  assign n30055 = ( n11321 & n23097 ) | ( n11321 & n30054 ) | ( n23097 & n30054 ) ;
  assign n30058 = n5035 ^ n4367 ^ n1098 ;
  assign n30059 = n30058 ^ n20827 ^ n6102 ;
  assign n30060 = ( n9259 & ~n9607 ) | ( n9259 & n30059 ) | ( ~n9607 & n30059 ) ;
  assign n30061 = n30060 ^ n3804 ^ x104 ;
  assign n30062 = n30061 ^ n28030 ^ n18538 ;
  assign n30056 = ~n487 & n2848 ;
  assign n30057 = n30056 ^ n12051 ^ 1'b0 ;
  assign n30063 = n30062 ^ n30057 ^ n1804 ;
  assign n30064 = n23052 ^ n5543 ^ n394 ;
  assign n30065 = n28852 ^ n1847 ^ 1'b0 ;
  assign n30066 = ~n24558 & n30065 ;
  assign n30067 = n12899 ^ n7127 ^ 1'b0 ;
  assign n30068 = n13866 & ~n30067 ;
  assign n30069 = n21533 ^ n4250 ^ 1'b0 ;
  assign n30070 = n13977 ^ n12388 ^ n9068 ;
  assign n30071 = ~n30069 & n30070 ;
  assign n30072 = ~n17238 & n28052 ;
  assign n30073 = n19127 ^ n7896 ^ n5910 ;
  assign n30074 = ( n6570 & n9229 ) | ( n6570 & ~n15752 ) | ( n9229 & ~n15752 ) ;
  assign n30075 = n30074 ^ n7401 ^ 1'b0 ;
  assign n30076 = n24938 ^ n2933 ^ n1250 ;
  assign n30077 = n14015 ^ n5078 ^ 1'b0 ;
  assign n30078 = n25967 ^ n365 ^ 1'b0 ;
  assign n30079 = ( n30076 & n30077 ) | ( n30076 & n30078 ) | ( n30077 & n30078 ) ;
  assign n30080 = n1017 & ~n2983 ;
  assign n30081 = n854 & ~n27822 ;
  assign n30082 = n30081 ^ n14044 ^ n7090 ;
  assign n30083 = ( ~n17032 & n17828 ) | ( ~n17032 & n28781 ) | ( n17828 & n28781 ) ;
  assign n30084 = n30083 ^ n18307 ^ n5058 ;
  assign n30085 = n8938 ^ n5863 ^ 1'b0 ;
  assign n30086 = n24158 & n30085 ;
  assign n30087 = n27594 & n30086 ;
  assign n30088 = n17566 & n18331 ;
  assign n30089 = n30088 ^ n11960 ^ 1'b0 ;
  assign n30090 = ~n2912 & n12354 ;
  assign n30091 = ~n2660 & n30090 ;
  assign n30092 = ( n1207 & n16911 ) | ( n1207 & n19815 ) | ( n16911 & n19815 ) ;
  assign n30093 = ( n6073 & ~n9261 ) | ( n6073 & n25109 ) | ( ~n9261 & n25109 ) ;
  assign n30094 = n30093 ^ n28001 ^ n13090 ;
  assign n30096 = n3377 ^ n1443 ^ 1'b0 ;
  assign n30095 = n2469 & ~n4626 ;
  assign n30097 = n30096 ^ n30095 ^ n12100 ;
  assign n30098 = ( ~n14319 & n17932 ) | ( ~n14319 & n30097 ) | ( n17932 & n30097 ) ;
  assign n30099 = ( ~n28059 & n29636 ) | ( ~n28059 & n30098 ) | ( n29636 & n30098 ) ;
  assign n30100 = ( n13014 & n13876 ) | ( n13014 & n28697 ) | ( n13876 & n28697 ) ;
  assign n30101 = n29268 ^ n16272 ^ n14063 ;
  assign n30102 = n5898 ^ n3290 ^ 1'b0 ;
  assign n30103 = ( n10346 & ~n13163 ) | ( n10346 & n30102 ) | ( ~n13163 & n30102 ) ;
  assign n30104 = ( n2593 & ~n19434 ) | ( n2593 & n30103 ) | ( ~n19434 & n30103 ) ;
  assign n30105 = n30104 ^ n23647 ^ n7688 ;
  assign n30106 = n7692 | n9540 ;
  assign n30107 = n3148 & ~n16689 ;
  assign n30108 = n30107 ^ n9362 ^ 1'b0 ;
  assign n30109 = n178 & ~n4153 ;
  assign n30110 = n30109 ^ n16244 ^ 1'b0 ;
  assign n30113 = ( n957 & ~n12539 ) | ( n957 & n24287 ) | ( ~n12539 & n24287 ) ;
  assign n30111 = n12613 & ~n19904 ;
  assign n30112 = n9198 & n30111 ;
  assign n30114 = n30113 ^ n30112 ^ 1'b0 ;
  assign n30116 = ( n6201 & n9217 ) | ( n6201 & ~n26811 ) | ( n9217 & ~n26811 ) ;
  assign n30115 = n2554 & ~n22149 ;
  assign n30117 = n30116 ^ n30115 ^ 1'b0 ;
  assign n30118 = n11087 ^ n10326 ^ n3732 ;
  assign n30119 = n5973 | n6953 ;
  assign n30120 = ( n13392 & ~n20623 ) | ( n13392 & n30119 ) | ( ~n20623 & n30119 ) ;
  assign n30121 = ( n424 & ~n11329 ) | ( n424 & n21626 ) | ( ~n11329 & n21626 ) ;
  assign n30122 = ( ~n4488 & n21680 ) | ( ~n4488 & n30121 ) | ( n21680 & n30121 ) ;
  assign n30123 = n8753 ^ n2213 ^ 1'b0 ;
  assign n30124 = ~n10549 & n30123 ;
  assign n30125 = ( ~n5916 & n24101 ) | ( ~n5916 & n30124 ) | ( n24101 & n30124 ) ;
  assign n30126 = n6928 | n24298 ;
  assign n30127 = n29638 | n30126 ;
  assign n30128 = ( ~n30122 & n30125 ) | ( ~n30122 & n30127 ) | ( n30125 & n30127 ) ;
  assign n30129 = n20827 ^ n6139 ^ 1'b0 ;
  assign n30130 = n12118 & ~n30129 ;
  assign n30131 = n30130 ^ n22587 ^ n20977 ;
  assign n30132 = n27114 ^ n19376 ^ n5970 ;
  assign n30133 = ~n1052 & n3529 ;
  assign n30134 = n23807 ^ n3007 ^ 1'b0 ;
  assign n30135 = n29049 & n30134 ;
  assign n30136 = n7844 ^ n7415 ^ 1'b0 ;
  assign n30137 = n10123 & n30136 ;
  assign n30138 = ~n1665 & n25437 ;
  assign n30139 = n9649 ^ n8054 ^ n2190 ;
  assign n30140 = n11719 ^ n7229 ^ 1'b0 ;
  assign n30141 = n30140 ^ n12973 ^ n7820 ;
  assign n30142 = n10492 ^ n6010 ^ n5710 ;
  assign n30143 = n30142 ^ n8676 ^ 1'b0 ;
  assign n30145 = n4040 | n26056 ;
  assign n30146 = n5149 | n30145 ;
  assign n30147 = n30146 ^ n12284 ^ 1'b0 ;
  assign n30148 = n30147 ^ n6746 ^ 1'b0 ;
  assign n30149 = n11516 & ~n30148 ;
  assign n30144 = n12809 ^ n5858 ^ 1'b0 ;
  assign n30150 = n30149 ^ n30144 ^ n19953 ;
  assign n30151 = n28523 ^ n16435 ^ 1'b0 ;
  assign n30152 = n27476 | n30151 ;
  assign n30154 = n20653 ^ n10777 ^ n8620 ;
  assign n30153 = n27485 & ~n27758 ;
  assign n30155 = n30154 ^ n30153 ^ 1'b0 ;
  assign n30156 = n9871 & n26522 ;
  assign n30157 = n30156 ^ n6746 ^ 1'b0 ;
  assign n30158 = n3118 & n30157 ;
  assign n30159 = ~n21428 & n30158 ;
  assign n30160 = n9844 ^ n386 ^ 1'b0 ;
  assign n30161 = n7399 & ~n30160 ;
  assign n30164 = n22634 ^ x95 ^ 1'b0 ;
  assign n30165 = n1541 | n30164 ;
  assign n30162 = n24443 ^ n2118 ^ n213 ;
  assign n30163 = n30162 ^ n25316 ^ n8931 ;
  assign n30166 = n30165 ^ n30163 ^ n22947 ;
  assign n30167 = n23894 ^ n18096 ^ n16943 ;
  assign n30169 = n5870 | n27657 ;
  assign n30170 = n29949 | n30169 ;
  assign n30168 = n25897 ^ n4721 ^ x80 ;
  assign n30171 = n30170 ^ n30168 ^ n24077 ;
  assign n30172 = ( n16457 & n17601 ) | ( n16457 & n19647 ) | ( n17601 & n19647 ) ;
  assign n30173 = n5360 ^ x10 ^ 1'b0 ;
  assign n30174 = ( n9599 & ~n14835 ) | ( n9599 & n30173 ) | ( ~n14835 & n30173 ) ;
  assign n30175 = n19327 ^ n3312 ^ n3153 ;
  assign n30176 = n8139 ^ n4761 ^ 1'b0 ;
  assign n30177 = n30176 ^ n28406 ^ n10795 ;
  assign n30179 = n25944 ^ n16228 ^ n12432 ;
  assign n30178 = n13733 | n28331 ;
  assign n30180 = n30179 ^ n30178 ^ 1'b0 ;
  assign n30181 = n10087 & ~n25646 ;
  assign n30182 = n30181 ^ n5837 ^ 1'b0 ;
  assign n30183 = ( ~n11038 & n28466 ) | ( ~n11038 & n28699 ) | ( n28466 & n28699 ) ;
  assign n30184 = ~n25910 & n30183 ;
  assign n30185 = n30184 ^ n7779 ^ 1'b0 ;
  assign n30186 = n18932 ^ n5193 ^ n3018 ;
  assign n30187 = ( ~n9031 & n12013 ) | ( ~n9031 & n22098 ) | ( n12013 & n22098 ) ;
  assign n30188 = n8454 ^ n7426 ^ n5973 ;
  assign n30189 = n17815 | n26599 ;
  assign n30190 = n13847 & ~n30189 ;
  assign n30191 = ( n7155 & n15067 ) | ( n7155 & ~n26200 ) | ( n15067 & ~n26200 ) ;
  assign n30192 = n13695 | n21554 ;
  assign n30193 = ( ~n9693 & n11907 ) | ( ~n9693 & n30192 ) | ( n11907 & n30192 ) ;
  assign n30194 = ( ~n2405 & n8226 ) | ( ~n2405 & n30193 ) | ( n8226 & n30193 ) ;
  assign n30195 = n30194 ^ n28923 ^ 1'b0 ;
  assign n30196 = n30191 & ~n30195 ;
  assign n30197 = n28675 ^ n25728 ^ n14785 ;
  assign n30198 = n25340 ^ n8086 ^ n1542 ;
  assign n30199 = n30198 ^ n21718 ^ n2142 ;
  assign n30200 = ( x40 & n1956 ) | ( x40 & n6240 ) | ( n1956 & n6240 ) ;
  assign n30201 = ~n8039 & n30200 ;
  assign n30202 = n30201 ^ n10012 ^ 1'b0 ;
  assign n30203 = ( ~n3200 & n17254 ) | ( ~n3200 & n30202 ) | ( n17254 & n30202 ) ;
  assign n30206 = n13697 & n29502 ;
  assign n30204 = n3033 | n28648 ;
  assign n30205 = n1172 | n30204 ;
  assign n30207 = n30206 ^ n30205 ^ n541 ;
  assign n30208 = n27697 ^ n19378 ^ n15270 ;
  assign n30209 = ( ~n3480 & n15324 ) | ( ~n3480 & n16438 ) | ( n15324 & n16438 ) ;
  assign n30210 = n30209 ^ n24459 ^ n11093 ;
  assign n30211 = n30208 | n30210 ;
  assign n30212 = ( ~n2849 & n6504 ) | ( ~n2849 & n24744 ) | ( n6504 & n24744 ) ;
  assign n30213 = n18335 ^ n11469 ^ 1'b0 ;
  assign n30214 = n19742 | n30213 ;
  assign n30215 = ~n13825 & n23210 ;
  assign n30216 = ~n23629 & n30215 ;
  assign n30217 = n27734 ^ n27241 ^ n9652 ;
  assign n30218 = n7674 & ~n25119 ;
  assign n30219 = n30218 ^ n4494 ^ 1'b0 ;
  assign n30220 = n30219 ^ n24896 ^ 1'b0 ;
  assign n30221 = ( ~n854 & n1506 ) | ( ~n854 & n19042 ) | ( n1506 & n19042 ) ;
  assign n30222 = ( n6042 & n25400 ) | ( n6042 & ~n30221 ) | ( n25400 & ~n30221 ) ;
  assign n30223 = n16914 ^ n10397 ^ n3687 ;
  assign n30224 = n30223 ^ n18193 ^ n13413 ;
  assign n30225 = ( ~n9303 & n12652 ) | ( ~n9303 & n30224 ) | ( n12652 & n30224 ) ;
  assign n30227 = n4467 & ~n21005 ;
  assign n30226 = n5444 ^ n2822 ^ n156 ;
  assign n30228 = n30227 ^ n30226 ^ n29697 ;
  assign n30229 = ( ~n6865 & n15674 ) | ( ~n6865 & n23660 ) | ( n15674 & n23660 ) ;
  assign n30230 = ( n5642 & ~n6534 ) | ( n5642 & n16277 ) | ( ~n6534 & n16277 ) ;
  assign n30231 = ( ~n2773 & n4920 ) | ( ~n2773 & n12464 ) | ( n4920 & n12464 ) ;
  assign n30232 = n30231 ^ n21699 ^ 1'b0 ;
  assign n30233 = n30230 & n30232 ;
  assign n30234 = n8719 & ~n15730 ;
  assign n30235 = n30234 ^ n29665 ^ 1'b0 ;
  assign n30236 = ~n7491 & n20950 ;
  assign n30237 = n14817 ^ n14726 ^ n12440 ;
  assign n30238 = n23721 & ~n30237 ;
  assign n30239 = n7551 & n30238 ;
  assign n30240 = n30239 ^ n29496 ^ 1'b0 ;
  assign n30241 = n16783 & ~n30240 ;
  assign n30242 = n18011 ^ n8135 ^ 1'b0 ;
  assign n30243 = ( n18944 & ~n22678 ) | ( n18944 & n26745 ) | ( ~n22678 & n26745 ) ;
  assign n30244 = ( n4221 & ~n6120 ) | ( n4221 & n7299 ) | ( ~n6120 & n7299 ) ;
  assign n30245 = n2261 | n16289 ;
  assign n30246 = n30244 | n30245 ;
  assign n30247 = n10838 | n13662 ;
  assign n30248 = ( ~n4179 & n30246 ) | ( ~n4179 & n30247 ) | ( n30246 & n30247 ) ;
  assign n30249 = n7085 | n10746 ;
  assign n30250 = n16102 ^ n12707 ^ n8695 ;
  assign n30251 = n30250 ^ n12328 ^ 1'b0 ;
  assign n30252 = n27822 ^ n10364 ^ n5965 ;
  assign n30254 = ~n2566 & n8658 ;
  assign n30255 = n30254 ^ n26516 ^ 1'b0 ;
  assign n30256 = ( n2872 & n24633 ) | ( n2872 & ~n30255 ) | ( n24633 & ~n30255 ) ;
  assign n30253 = n14010 | n14421 ;
  assign n30257 = n30256 ^ n30253 ^ 1'b0 ;
  assign n30258 = n16902 & ~n22468 ;
  assign n30259 = n7369 & n30258 ;
  assign n30260 = n16849 | n19605 ;
  assign n30261 = n30260 ^ n7841 ^ 1'b0 ;
  assign n30262 = n15785 ^ n15431 ^ 1'b0 ;
  assign n30263 = n926 & n30262 ;
  assign n30264 = ~n4257 & n7100 ;
  assign n30265 = n30264 ^ n18070 ^ n15151 ;
  assign n30266 = ( n2526 & ~n12456 ) | ( n2526 & n19575 ) | ( ~n12456 & n19575 ) ;
  assign n30267 = n18814 ^ n894 ^ 1'b0 ;
  assign n30268 = n7837 ^ n1694 ^ 1'b0 ;
  assign n30269 = ~n4033 & n20086 ;
  assign n30270 = n30269 ^ x52 ^ 1'b0 ;
  assign n30271 = n30270 ^ n17450 ^ n12825 ;
  assign n30272 = n1664 & ~n20674 ;
  assign n30273 = ~n10334 & n23001 ;
  assign n30274 = n30273 ^ n12425 ^ 1'b0 ;
  assign n30275 = n30274 ^ n7108 ^ n2858 ;
  assign n30276 = n30275 ^ n3646 ^ n2265 ;
  assign n30277 = ( ~n9149 & n30272 ) | ( ~n9149 & n30276 ) | ( n30272 & n30276 ) ;
  assign n30278 = n7143 ^ n2850 ^ 1'b0 ;
  assign n30279 = ( n2437 & ~n8433 ) | ( n2437 & n30278 ) | ( ~n8433 & n30278 ) ;
  assign n30280 = n4884 & ~n13733 ;
  assign n30281 = ~n22978 & n30280 ;
  assign n30282 = ~n2392 & n23794 ;
  assign n30283 = n30282 ^ n7909 ^ 1'b0 ;
  assign n30284 = ( n14706 & n17334 ) | ( n14706 & ~n19504 ) | ( n17334 & ~n19504 ) ;
  assign n30285 = n2580 & ~n30284 ;
  assign n30286 = ( n5241 & ~n6432 ) | ( n5241 & n7277 ) | ( ~n6432 & n7277 ) ;
  assign n30287 = n30286 ^ n24955 ^ n10552 ;
  assign n30288 = n23590 ^ n18360 ^ n11163 ;
  assign n30289 = n23874 ^ n22216 ^ n12619 ;
  assign n30290 = ~n16323 & n17872 ;
  assign n30291 = n28116 ^ n14748 ^ n3229 ;
  assign n30292 = n1291 | n30291 ;
  assign n30293 = n1992 & ~n28202 ;
  assign n30294 = n30293 ^ n1644 ^ 1'b0 ;
  assign n30295 = n28453 ^ n13219 ^ 1'b0 ;
  assign n30296 = ( n13468 & n15262 ) | ( n13468 & ~n30295 ) | ( n15262 & ~n30295 ) ;
  assign n30297 = n3265 | n12369 ;
  assign n30298 = n30297 ^ n7628 ^ 1'b0 ;
  assign n30299 = n4350 & ~n6157 ;
  assign n30300 = ~n10585 & n30299 ;
  assign n30301 = n30300 ^ n24627 ^ 1'b0 ;
  assign n30302 = n27939 | n30301 ;
  assign n30303 = ( n8923 & n17263 ) | ( n8923 & ~n29085 ) | ( n17263 & ~n29085 ) ;
  assign n30304 = ( n1761 & n6918 ) | ( n1761 & n12222 ) | ( n6918 & n12222 ) ;
  assign n30305 = ( n18161 & ~n25033 ) | ( n18161 & n30304 ) | ( ~n25033 & n30304 ) ;
  assign n30306 = n20194 ^ n17510 ^ n5638 ;
  assign n30307 = n26095 ^ n16614 ^ n3190 ;
  assign n30308 = n5335 ^ n4049 ^ 1'b0 ;
  assign n30309 = ( n5235 & n16693 ) | ( n5235 & n30308 ) | ( n16693 & n30308 ) ;
  assign n30310 = n1761 | n30309 ;
  assign n30312 = n17988 ^ n7518 ^ n3329 ;
  assign n30311 = n18635 ^ n2701 ^ 1'b0 ;
  assign n30313 = n30312 ^ n30311 ^ n2146 ;
  assign n30314 = n28725 ^ n7122 ^ 1'b0 ;
  assign n30315 = n20674 ^ n7202 ^ n7000 ;
  assign n30316 = ( n12606 & ~n22388 ) | ( n12606 & n30315 ) | ( ~n22388 & n30315 ) ;
  assign n30317 = n29038 & ~n30316 ;
  assign n30318 = n22712 & n30317 ;
  assign n30319 = n13572 | n24664 ;
  assign n30320 = n30319 ^ n9897 ^ 1'b0 ;
  assign n30321 = n28651 ^ n881 ^ 1'b0 ;
  assign n30322 = n10758 ^ n5978 ^ n1092 ;
  assign n30323 = n30322 ^ n12221 ^ 1'b0 ;
  assign n30324 = ~n30321 & n30323 ;
  assign n30325 = n6880 ^ n5012 ^ 1'b0 ;
  assign n30326 = n27947 ^ n14627 ^ n8891 ;
  assign n30327 = n30326 ^ n22672 ^ n773 ;
  assign n30328 = n30327 ^ n26764 ^ n1113 ;
  assign n30329 = n18742 ^ n17158 ^ n6108 ;
  assign n30330 = n19805 & n30329 ;
  assign n30331 = ( n17263 & ~n24798 ) | ( n17263 & n30330 ) | ( ~n24798 & n30330 ) ;
  assign n30332 = n2969 & n16466 ;
  assign n30333 = n23428 ^ n14523 ^ n13725 ;
  assign n30337 = n17515 ^ n15228 ^ n4161 ;
  assign n30334 = n3858 | n5281 ;
  assign n30335 = n23060 & ~n30334 ;
  assign n30336 = ( ~n9593 & n22386 ) | ( ~n9593 & n30335 ) | ( n22386 & n30335 ) ;
  assign n30338 = n30337 ^ n30336 ^ n18702 ;
  assign n30339 = n27822 ^ n27500 ^ n22316 ;
  assign n30340 = ( n3484 & n4678 ) | ( n3484 & ~n5276 ) | ( n4678 & ~n5276 ) ;
  assign n30341 = n30340 ^ n24191 ^ n11395 ;
  assign n30342 = ( ~n6914 & n15256 ) | ( ~n6914 & n26130 ) | ( n15256 & n26130 ) ;
  assign n30343 = n11578 & n30342 ;
  assign n30344 = ~n30341 & n30343 ;
  assign n30345 = n11594 ^ n4088 ^ 1'b0 ;
  assign n30346 = n13537 ^ n10091 ^ 1'b0 ;
  assign n30347 = n30345 & ~n30346 ;
  assign n30348 = n8391 ^ n7977 ^ n377 ;
  assign n30349 = n7157 & n30348 ;
  assign n30350 = n5816 & n30349 ;
  assign n30351 = x104 | n11797 ;
  assign n30352 = n7407 ^ n2716 ^ 1'b0 ;
  assign n30353 = ( n10568 & ~n30351 ) | ( n10568 & n30352 ) | ( ~n30351 & n30352 ) ;
  assign n30354 = n24957 ^ n10253 ^ n5782 ;
  assign n30355 = n28927 ^ n22467 ^ n13447 ;
  assign n30356 = n22472 ^ n22207 ^ n14396 ;
  assign n30357 = n30356 ^ n5056 ^ n2142 ;
  assign n30358 = ~n4464 & n11522 ;
  assign n30359 = n30357 & n30358 ;
  assign n30360 = n1114 & ~n30359 ;
  assign n30361 = n18511 ^ n14044 ^ n6271 ;
  assign n30362 = ( n9145 & n27716 ) | ( n9145 & n30275 ) | ( n27716 & n30275 ) ;
  assign n30363 = n6080 & ~n30362 ;
  assign n30364 = n967 & ~n7121 ;
  assign n30365 = n30364 ^ n2379 ^ 1'b0 ;
  assign n30366 = ( n13178 & n16636 ) | ( n13178 & n30365 ) | ( n16636 & n30365 ) ;
  assign n30367 = n25401 ^ n17860 ^ 1'b0 ;
  assign n30368 = n859 & ~n30367 ;
  assign n30369 = ~n11805 & n18349 ;
  assign n30370 = n30369 ^ n25694 ^ n23870 ;
  assign n30371 = n18322 ^ n16187 ^ n9121 ;
  assign n30372 = ( n2185 & ~n6783 ) | ( n2185 & n7524 ) | ( ~n6783 & n7524 ) ;
  assign n30373 = ( n5725 & n17991 ) | ( n5725 & n30372 ) | ( n17991 & n30372 ) ;
  assign n30374 = n19969 ^ n2011 ^ n1949 ;
  assign n30375 = n30374 ^ n11030 ^ 1'b0 ;
  assign n30376 = ~n5863 & n30375 ;
  assign n30377 = n30376 ^ n20754 ^ n1297 ;
  assign n30378 = ~n8421 & n23679 ;
  assign n30379 = n8509 & n30378 ;
  assign n30381 = n19939 ^ n12251 ^ n4444 ;
  assign n30380 = n464 | n6896 ;
  assign n30382 = n30381 ^ n30380 ^ 1'b0 ;
  assign n30383 = ( n12224 & n30379 ) | ( n12224 & ~n30382 ) | ( n30379 & ~n30382 ) ;
  assign n30384 = n4591 & n8829 ;
  assign n30385 = n30384 ^ n6850 ^ n3911 ;
  assign n30386 = n30154 ^ n28762 ^ n18591 ;
  assign n30387 = ( ~n12382 & n21045 ) | ( ~n12382 & n30386 ) | ( n21045 & n30386 ) ;
  assign n30388 = ( n16217 & ~n21712 ) | ( n16217 & n29810 ) | ( ~n21712 & n29810 ) ;
  assign n30389 = n30388 ^ n22024 ^ 1'b0 ;
  assign n30390 = ~n4823 & n23957 ;
  assign n30391 = n30390 ^ n15869 ^ 1'b0 ;
  assign n30392 = ( n1172 & n22126 ) | ( n1172 & ~n22207 ) | ( n22126 & ~n22207 ) ;
  assign n30393 = ~n12185 & n30392 ;
  assign n30394 = ( n20851 & ~n30391 ) | ( n20851 & n30393 ) | ( ~n30391 & n30393 ) ;
  assign n30395 = n21385 & ~n30394 ;
  assign n30396 = ~n21956 & n25275 ;
  assign n30397 = ( n1525 & n15789 ) | ( n1525 & ~n18409 ) | ( n15789 & ~n18409 ) ;
  assign n30398 = n30397 ^ n19760 ^ n2218 ;
  assign n30399 = ( n5099 & n20112 ) | ( n5099 & ~n22061 ) | ( n20112 & ~n22061 ) ;
  assign n30400 = n26110 ^ n22205 ^ n10945 ;
  assign n30402 = n16359 | n26647 ;
  assign n30401 = n7575 & ~n15572 ;
  assign n30403 = n30402 ^ n30401 ^ n8853 ;
  assign n30404 = ( n317 & n14041 ) | ( n317 & n14780 ) | ( n14041 & n14780 ) ;
  assign n30405 = n8259 & ~n10346 ;
  assign n30406 = n30405 ^ n17891 ^ 1'b0 ;
  assign n30407 = n19441 ^ n4381 ^ 1'b0 ;
  assign n30408 = n30406 & n30407 ;
  assign n30409 = ~n30404 & n30408 ;
  assign n30410 = n10950 ^ n10814 ^ n1688 ;
  assign n30411 = n713 | n7990 ;
  assign n30412 = ( n17934 & n30410 ) | ( n17934 & n30411 ) | ( n30410 & n30411 ) ;
  assign n30413 = ( n3635 & ~n28499 ) | ( n3635 & n30412 ) | ( ~n28499 & n30412 ) ;
  assign n30414 = ~n5967 & n10689 ;
  assign n30415 = ~n8323 & n30414 ;
  assign n30416 = ( ~n13437 & n17208 ) | ( ~n13437 & n30415 ) | ( n17208 & n30415 ) ;
  assign n30417 = n24795 ^ n13409 ^ 1'b0 ;
  assign n30418 = n13821 & n30417 ;
  assign n30419 = n268 & n9048 ;
  assign n30420 = n9645 & n30419 ;
  assign n30421 = n30420 ^ n23649 ^ 1'b0 ;
  assign n30423 = n27630 ^ n23069 ^ n12029 ;
  assign n30424 = ~n5909 & n30423 ;
  assign n30422 = n25773 & ~n27355 ;
  assign n30425 = n30424 ^ n30422 ^ 1'b0 ;
  assign n30426 = n20100 ^ n11115 ^ n5915 ;
  assign n30427 = ~n3922 & n15681 ;
  assign n30428 = n30427 ^ n8914 ^ 1'b0 ;
  assign n30429 = n30428 ^ n19368 ^ n16783 ;
  assign n30430 = ( n4936 & ~n6883 ) | ( n4936 & n26574 ) | ( ~n6883 & n26574 ) ;
  assign n30431 = n30430 ^ n13075 ^ 1'b0 ;
  assign n30432 = n2385 & n30431 ;
  assign n30433 = ( ~n2479 & n22054 ) | ( ~n2479 & n30432 ) | ( n22054 & n30432 ) ;
  assign n30435 = ~n12273 & n28164 ;
  assign n30434 = ( n5793 & n6198 ) | ( n5793 & ~n15424 ) | ( n6198 & ~n15424 ) ;
  assign n30436 = n30435 ^ n30434 ^ n7818 ;
  assign n30437 = ( n966 & ~n4850 ) | ( n966 & n20150 ) | ( ~n4850 & n20150 ) ;
  assign n30438 = n30437 ^ n12413 ^ n6954 ;
  assign n30439 = n30438 ^ n7936 ^ n2946 ;
  assign n30440 = n1660 | n30439 ;
  assign n30441 = ( x17 & n3397 ) | ( x17 & ~n10101 ) | ( n3397 & ~n10101 ) ;
  assign n30442 = ( n3999 & n26141 ) | ( n3999 & n30441 ) | ( n26141 & n30441 ) ;
  assign n30443 = ( n3984 & ~n12058 ) | ( n3984 & n30442 ) | ( ~n12058 & n30442 ) ;
  assign n30444 = n30443 ^ n15271 ^ n10974 ;
  assign n30445 = n9643 & ~n15144 ;
  assign n30446 = ~n27122 & n30445 ;
  assign n30447 = ( n2694 & ~n25134 ) | ( n2694 & n30446 ) | ( ~n25134 & n30446 ) ;
  assign n30448 = n16660 | n30447 ;
  assign n30449 = n13228 | n30448 ;
  assign n30450 = n3473 & ~n4418 ;
  assign n30451 = n5433 & n30450 ;
  assign n30454 = n7569 | n11348 ;
  assign n30455 = n29648 & ~n30454 ;
  assign n30452 = n10033 ^ n8167 ^ 1'b0 ;
  assign n30453 = n20302 | n30452 ;
  assign n30456 = n30455 ^ n30453 ^ 1'b0 ;
  assign n30459 = n4058 ^ n3592 ^ 1'b0 ;
  assign n30460 = n24213 & ~n30459 ;
  assign n30457 = ( n3139 & n4278 ) | ( n3139 & n4919 ) | ( n4278 & n4919 ) ;
  assign n30458 = ( x78 & ~n9336 ) | ( x78 & n30457 ) | ( ~n9336 & n30457 ) ;
  assign n30461 = n30460 ^ n30458 ^ n10142 ;
  assign n30462 = ~n12925 & n30461 ;
  assign n30463 = ~n17170 & n30462 ;
  assign n30464 = n18171 ^ n2644 ^ 1'b0 ;
  assign n30465 = ~n15901 & n29327 ;
  assign n30466 = ~n30464 & n30465 ;
  assign n30467 = n28279 ^ n8608 ^ n3603 ;
  assign n30468 = ( n6206 & n6790 ) | ( n6206 & ~n30467 ) | ( n6790 & ~n30467 ) ;
  assign n30469 = n13727 | n29937 ;
  assign n30474 = n12588 | n12896 ;
  assign n30475 = n30474 ^ n5333 ^ 1'b0 ;
  assign n30470 = n10998 ^ n10714 ^ n7839 ;
  assign n30471 = ( ~n966 & n6949 ) | ( ~n966 & n30470 ) | ( n6949 & n30470 ) ;
  assign n30472 = ~n6738 & n30471 ;
  assign n30473 = n3183 & n30472 ;
  assign n30476 = n30475 ^ n30473 ^ 1'b0 ;
  assign n30477 = n3097 & ~n25167 ;
  assign n30478 = n30477 ^ n13384 ^ 1'b0 ;
  assign n30479 = n30478 ^ n10225 ^ n3217 ;
  assign n30480 = ( n13687 & n20678 ) | ( n13687 & n30479 ) | ( n20678 & n30479 ) ;
  assign n30481 = n11916 ^ n3631 ^ 1'b0 ;
  assign n30482 = ~n13686 & n30481 ;
  assign n30483 = x62 & n30482 ;
  assign n30484 = ( ~n8047 & n11706 ) | ( ~n8047 & n30483 ) | ( n11706 & n30483 ) ;
  assign n30485 = n6413 | n12163 ;
  assign n30486 = n30485 ^ n9355 ^ 1'b0 ;
  assign n30487 = n30486 ^ n15311 ^ n5310 ;
  assign n30488 = ( ~n6503 & n11957 ) | ( ~n6503 & n24336 ) | ( n11957 & n24336 ) ;
  assign n30489 = ~n1462 & n13345 ;
  assign n30490 = ( n27137 & n30488 ) | ( n27137 & n30489 ) | ( n30488 & n30489 ) ;
  assign n30491 = n21081 | n30490 ;
  assign n30492 = ~n11546 & n18908 ;
  assign n30493 = n14227 | n20865 ;
  assign n30494 = n22900 & n30493 ;
  assign n30495 = ~n7473 & n8848 ;
  assign n30496 = ~n14984 & n30495 ;
  assign n30497 = n30496 ^ n9630 ^ 1'b0 ;
  assign n30498 = n12121 & n20873 ;
  assign n30499 = ~n7849 & n30498 ;
  assign n30500 = n28059 ^ n10920 ^ n7582 ;
  assign n30502 = ( n9163 & n12013 ) | ( n9163 & ~n12030 ) | ( n12013 & ~n12030 ) ;
  assign n30501 = n29524 ^ n5564 ^ 1'b0 ;
  assign n30503 = n30502 ^ n30501 ^ n19574 ;
  assign n30504 = ( n2210 & n9845 ) | ( n2210 & ~n14564 ) | ( n9845 & ~n14564 ) ;
  assign n30505 = n30504 ^ n28265 ^ n11701 ;
  assign n30506 = n30505 ^ n13664 ^ n681 ;
  assign n30507 = n13623 & ~n16213 ;
  assign n30508 = n30507 ^ n20804 ^ 1'b0 ;
  assign n30509 = ( ~n6578 & n11231 ) | ( ~n6578 & n30508 ) | ( n11231 & n30508 ) ;
  assign n30510 = n28219 ^ n14332 ^ 1'b0 ;
  assign n30511 = n25965 ^ n10369 ^ 1'b0 ;
  assign n30512 = ( ~n964 & n8513 ) | ( ~n964 & n13591 ) | ( n8513 & n13591 ) ;
  assign n30513 = n6207 | n18072 ;
  assign n30514 = n30512 | n30513 ;
  assign n30516 = n14780 ^ n3461 ^ 1'b0 ;
  assign n30515 = n6606 | n21520 ;
  assign n30517 = n30516 ^ n30515 ^ 1'b0 ;
  assign n30518 = ( ~n900 & n14639 ) | ( ~n900 & n18694 ) | ( n14639 & n18694 ) ;
  assign n30519 = ( n9553 & n10221 ) | ( n9553 & n29057 ) | ( n10221 & n29057 ) ;
  assign n30520 = n30519 ^ n16602 ^ 1'b0 ;
  assign n30521 = n30518 & ~n30520 ;
  assign n30522 = n7662 & n10303 ;
  assign n30523 = n30522 ^ n6580 ^ 1'b0 ;
  assign n30524 = n17138 & n22257 ;
  assign n30525 = n30524 ^ n4922 ^ 1'b0 ;
  assign n30526 = ( ~n8546 & n30523 ) | ( ~n8546 & n30525 ) | ( n30523 & n30525 ) ;
  assign n30532 = n22598 ^ n20960 ^ 1'b0 ;
  assign n30533 = n30532 ^ n11561 ^ n3525 ;
  assign n30531 = n20227 ^ n8539 ^ 1'b0 ;
  assign n30527 = n10431 ^ n3971 ^ 1'b0 ;
  assign n30528 = ~n8937 & n30527 ;
  assign n30529 = ( ~n5063 & n10288 ) | ( ~n5063 & n22052 ) | ( n10288 & n22052 ) ;
  assign n30530 = ( n9734 & ~n30528 ) | ( n9734 & n30529 ) | ( ~n30528 & n30529 ) ;
  assign n30534 = n30533 ^ n30531 ^ n30530 ;
  assign n30535 = ( n12044 & ~n22225 ) | ( n12044 & n29289 ) | ( ~n22225 & n29289 ) ;
  assign n30536 = ( n8876 & ~n23198 ) | ( n8876 & n30535 ) | ( ~n23198 & n30535 ) ;
  assign n30537 = n28917 ^ n25165 ^ n2777 ;
  assign n30538 = ( x51 & n751 ) | ( x51 & ~n3526 ) | ( n751 & ~n3526 ) ;
  assign n30539 = ( n2423 & ~n17607 ) | ( n2423 & n30112 ) | ( ~n17607 & n30112 ) ;
  assign n30540 = n3098 ^ n825 ^ 1'b0 ;
  assign n30541 = ~n4255 & n8958 ;
  assign n30542 = ~n21181 & n30541 ;
  assign n30543 = n13710 | n25413 ;
  assign n30544 = n30543 ^ n15876 ^ 1'b0 ;
  assign n30547 = n7175 ^ n1707 ^ 1'b0 ;
  assign n30548 = n13766 | n30547 ;
  assign n30546 = n10452 | n11870 ;
  assign n30545 = n24095 ^ n15600 ^ n5045 ;
  assign n30549 = n30548 ^ n30546 ^ n30545 ;
  assign n30550 = n5760 & ~n30549 ;
  assign n30551 = n3696 & n30550 ;
  assign n30552 = n24740 ^ n14182 ^ n5525 ;
  assign n30553 = n11509 ^ n9736 ^ n1958 ;
  assign n30554 = ( n3026 & ~n3935 ) | ( n3026 & n24443 ) | ( ~n3935 & n24443 ) ;
  assign n30555 = ( n4507 & n30553 ) | ( n4507 & ~n30554 ) | ( n30553 & ~n30554 ) ;
  assign n30556 = n6998 & ~n28187 ;
  assign n30557 = n30556 ^ n19549 ^ 1'b0 ;
  assign n30558 = ( ~n3740 & n12201 ) | ( ~n3740 & n30557 ) | ( n12201 & n30557 ) ;
  assign n30559 = n30558 ^ n16648 ^ 1'b0 ;
  assign n30560 = n19869 ^ n18842 ^ n7858 ;
  assign n30561 = n19746 | n30560 ;
  assign n30562 = n4093 & ~n27548 ;
  assign n30563 = n6149 | n6777 ;
  assign n30564 = n2351 & ~n30563 ;
  assign n30565 = n1206 | n5281 ;
  assign n30566 = n12472 & ~n30565 ;
  assign n30567 = n30566 ^ n5950 ^ n3259 ;
  assign n30568 = n5790 & n30567 ;
  assign n30569 = ( n9905 & ~n30564 ) | ( n9905 & n30568 ) | ( ~n30564 & n30568 ) ;
  assign n30570 = n22406 ^ n9306 ^ 1'b0 ;
  assign n30571 = n9716 ^ n7298 ^ n7146 ;
  assign n30572 = ( ~n22130 & n30570 ) | ( ~n22130 & n30571 ) | ( n30570 & n30571 ) ;
  assign n30573 = n30572 ^ n26761 ^ 1'b0 ;
  assign n30574 = n30573 ^ n22512 ^ n11948 ;
  assign n30575 = n15684 | n19413 ;
  assign n30576 = n28681 & ~n30575 ;
  assign n30577 = n19105 ^ n175 ^ 1'b0 ;
  assign n30578 = n30577 ^ n11784 ^ 1'b0 ;
  assign n30579 = n28584 ^ n11938 ^ n3167 ;
  assign n30580 = n4410 ^ n3526 ^ x77 ;
  assign n30581 = n30580 ^ n22890 ^ 1'b0 ;
  assign n30582 = ( ~n14867 & n23263 ) | ( ~n14867 & n29019 ) | ( n23263 & n29019 ) ;
  assign n30583 = n14817 | n27823 ;
  assign n30584 = n30583 ^ n6635 ^ 1'b0 ;
  assign n30585 = n30584 ^ n23333 ^ n1738 ;
  assign n30586 = ~n6233 & n9398 ;
  assign n30587 = n30554 ^ n20325 ^ 1'b0 ;
  assign n30588 = ( n11267 & n21643 ) | ( n11267 & ~n30587 ) | ( n21643 & ~n30587 ) ;
  assign n30589 = n4373 ^ n2759 ^ 1'b0 ;
  assign n30590 = ~n9777 & n21276 ;
  assign n30591 = n30590 ^ n19388 ^ 1'b0 ;
  assign n30592 = n8156 & ~n10450 ;
  assign n30593 = n30592 ^ n10033 ^ 1'b0 ;
  assign n30597 = ~n17391 & n22524 ;
  assign n30598 = ~n2053 & n30597 ;
  assign n30599 = n30598 ^ n22568 ^ n18237 ;
  assign n30600 = ( x83 & ~n27672 ) | ( x83 & n30599 ) | ( ~n27672 & n30599 ) ;
  assign n30594 = n28412 ^ n339 ^ 1'b0 ;
  assign n30595 = ~n15879 & n30594 ;
  assign n30596 = n30595 ^ n22114 ^ n13625 ;
  assign n30601 = n30600 ^ n30596 ^ n7266 ;
  assign n30602 = n20451 ^ n18534 ^ n12433 ;
  assign n30603 = n30602 ^ x7 ^ 1'b0 ;
  assign n30604 = n1900 & ~n18776 ;
  assign n30605 = n3113 & ~n24519 ;
  assign n30606 = n30604 & n30605 ;
  assign n30607 = ( ~n3503 & n25934 ) | ( ~n3503 & n30606 ) | ( n25934 & n30606 ) ;
  assign n30608 = n2734 & ~n30607 ;
  assign n30609 = n28949 ^ n25579 ^ n9291 ;
  assign n30610 = ( ~n2819 & n10654 ) | ( ~n2819 & n17888 ) | ( n10654 & n17888 ) ;
  assign n30611 = ( ~n1290 & n1965 ) | ( ~n1290 & n10600 ) | ( n1965 & n10600 ) ;
  assign n30612 = n30611 ^ n1051 ^ 1'b0 ;
  assign n30613 = ~n23965 & n30612 ;
  assign n30614 = ( n2003 & n18401 ) | ( n2003 & n30613 ) | ( n18401 & n30613 ) ;
  assign n30615 = n29080 ^ n10753 ^ n10232 ;
  assign n30616 = ( n24421 & n24874 ) | ( n24421 & n30615 ) | ( n24874 & n30615 ) ;
  assign n30617 = ( n11760 & ~n20184 ) | ( n11760 & n30616 ) | ( ~n20184 & n30616 ) ;
  assign n30618 = n22959 ^ n4442 ^ 1'b0 ;
  assign n30619 = ~n20317 & n30618 ;
  assign n30620 = n1348 & n5825 ;
  assign n30621 = ~n22171 & n30620 ;
  assign n30622 = ~n16346 & n29950 ;
  assign n30623 = n724 & n2307 ;
  assign n30624 = n30623 ^ n26680 ^ 1'b0 ;
  assign n30625 = n30624 ^ n10400 ^ 1'b0 ;
  assign n30626 = ~n30622 & n30625 ;
  assign n30631 = n2250 | n2995 ;
  assign n30627 = ~n505 & n2818 ;
  assign n30628 = ~n17759 & n30627 ;
  assign n30629 = ( ~n1842 & n23839 ) | ( ~n1842 & n30628 ) | ( n23839 & n30628 ) ;
  assign n30630 = ~n10827 & n30629 ;
  assign n30632 = n30631 ^ n30630 ^ 1'b0 ;
  assign n30633 = n29017 ^ n11350 ^ n628 ;
  assign n30634 = n22881 ^ n21719 ^ n8236 ;
  assign n30635 = n3887 & n26159 ;
  assign n30636 = ( ~n3571 & n4860 ) | ( ~n3571 & n27992 ) | ( n4860 & n27992 ) ;
  assign n30637 = n16890 ^ n7982 ^ 1'b0 ;
  assign n30638 = n20589 ^ n17094 ^ 1'b0 ;
  assign n30639 = ( n1528 & ~n2639 ) | ( n1528 & n30638 ) | ( ~n2639 & n30638 ) ;
  assign n30640 = n21544 | n22014 ;
  assign n30641 = n26768 | n30640 ;
  assign n30642 = n16411 & n25663 ;
  assign n30643 = n30642 ^ n13508 ^ 1'b0 ;
  assign n30644 = n20549 ^ n15489 ^ n1961 ;
  assign n30645 = ( n6125 & ~n16159 ) | ( n6125 & n30644 ) | ( ~n16159 & n30644 ) ;
  assign n30646 = n26879 ^ n26208 ^ n17005 ;
  assign n30647 = n30646 ^ n25598 ^ 1'b0 ;
  assign n30648 = n12224 ^ n4356 ^ n875 ;
  assign n30649 = n30648 ^ n13988 ^ 1'b0 ;
  assign n30650 = n24132 | n30649 ;
  assign n30652 = n7261 | n24996 ;
  assign n30651 = n5797 & ~n24293 ;
  assign n30653 = n30652 ^ n30651 ^ 1'b0 ;
  assign n30654 = ( n21360 & n30650 ) | ( n21360 & n30653 ) | ( n30650 & n30653 ) ;
  assign n30655 = ( ~n5124 & n18838 ) | ( ~n5124 & n30654 ) | ( n18838 & n30654 ) ;
  assign n30656 = n14835 ^ n3601 ^ 1'b0 ;
  assign n30657 = n23531 ^ n5194 ^ 1'b0 ;
  assign n30658 = x46 & ~n30657 ;
  assign n30659 = n27767 ^ n25977 ^ n20211 ;
  assign n30660 = ( n7765 & n17644 ) | ( n7765 & n30659 ) | ( n17644 & n30659 ) ;
  assign n30661 = ( n18637 & n30658 ) | ( n18637 & n30660 ) | ( n30658 & n30660 ) ;
  assign n30662 = n5909 | n7382 ;
  assign n30663 = n14168 & ~n30662 ;
  assign n30664 = n30663 ^ n28814 ^ n9389 ;
  assign n30665 = n5637 ^ n5300 ^ 1'b0 ;
  assign n30666 = n25968 ^ n6408 ^ n2896 ;
  assign n30667 = n1455 | n10674 ;
  assign n30668 = n30667 ^ n8958 ^ 1'b0 ;
  assign n30669 = n30666 & n30668 ;
  assign n30670 = n1832 & ~n5496 ;
  assign n30671 = n2642 & n30670 ;
  assign n30672 = n7439 | n16289 ;
  assign n30673 = n7056 | n30672 ;
  assign n30674 = n30673 ^ n20622 ^ n9065 ;
  assign n30675 = n2656 & ~n30674 ;
  assign n30676 = ( n4524 & ~n24223 ) | ( n4524 & n25993 ) | ( ~n24223 & n25993 ) ;
  assign n30677 = n16408 ^ n9722 ^ n4231 ;
  assign n30678 = n10157 ^ n5087 ^ 1'b0 ;
  assign n30679 = ( n814 & n12594 ) | ( n814 & n14505 ) | ( n12594 & n14505 ) ;
  assign n30680 = n4724 & ~n14373 ;
  assign n30681 = ( n3131 & n13796 ) | ( n3131 & n30680 ) | ( n13796 & n30680 ) ;
  assign n30682 = n13821 ^ n2011 ^ 1'b0 ;
  assign n30683 = n30682 ^ n27242 ^ n16639 ;
  assign n30684 = n10753 | n21572 ;
  assign n30685 = n30684 ^ n4178 ^ 1'b0 ;
  assign n30686 = n15325 & ~n18816 ;
  assign n30687 = n30686 ^ n28378 ^ 1'b0 ;
  assign n30688 = n18207 ^ n15813 ^ n10651 ;
  assign n30689 = n30688 ^ n8632 ^ 1'b0 ;
  assign n30690 = n1704 & n23872 ;
  assign n30691 = ( ~n14220 & n16761 ) | ( ~n14220 & n17575 ) | ( n16761 & n17575 ) ;
  assign n30692 = n11444 ^ n5269 ^ 1'b0 ;
  assign n30694 = n7108 | n9096 ;
  assign n30695 = n6172 & ~n30694 ;
  assign n30693 = x123 & ~n9242 ;
  assign n30696 = n30695 ^ n30693 ^ 1'b0 ;
  assign n30697 = ( n6890 & n8701 ) | ( n6890 & ~n30696 ) | ( n8701 & ~n30696 ) ;
  assign n30698 = n2132 | n14402 ;
  assign n30699 = n10822 | n30698 ;
  assign n30700 = n30699 ^ n11484 ^ 1'b0 ;
  assign n30701 = n16008 ^ n12910 ^ 1'b0 ;
  assign n30702 = n30701 ^ n4505 ^ n3713 ;
  assign n30703 = n4782 & ~n8098 ;
  assign n30704 = ( n1652 & n15244 ) | ( n1652 & ~n23196 ) | ( n15244 & ~n23196 ) ;
  assign n30705 = n11697 ^ n3334 ^ 1'b0 ;
  assign n30706 = n30704 & n30705 ;
  assign n30707 = n15557 & n30624 ;
  assign n30708 = n17420 ^ n16532 ^ 1'b0 ;
  assign n30709 = n30002 & n30708 ;
  assign n30710 = n30709 ^ n9475 ^ 1'b0 ;
  assign n30711 = n17323 ^ n1698 ^ 1'b0 ;
  assign n30712 = n25761 ^ n3723 ^ 1'b0 ;
  assign n30713 = n22452 & n30712 ;
  assign n30714 = ( ~n12912 & n30535 ) | ( ~n12912 & n30713 ) | ( n30535 & n30713 ) ;
  assign n30715 = n9096 & ~n14716 ;
  assign n30716 = ( n4990 & n18240 ) | ( n4990 & n24558 ) | ( n18240 & n24558 ) ;
  assign n30717 = n29047 ^ n23716 ^ 1'b0 ;
  assign n30718 = ~n8021 & n30717 ;
  assign n30719 = ~n10691 & n30667 ;
  assign n30720 = ~n16850 & n29198 ;
  assign n30721 = n2306 & ~n13549 ;
  assign n30722 = ~n253 & n7337 ;
  assign n30723 = ~n13292 & n30722 ;
  assign n30724 = ~n12298 & n15936 ;
  assign n30725 = n30724 ^ x26 ^ 1'b0 ;
  assign n30726 = n18020 ^ n17866 ^ n14940 ;
  assign n30727 = ( n3939 & ~n30725 ) | ( n3939 & n30726 ) | ( ~n30725 & n30726 ) ;
  assign n30728 = ( ~n3730 & n6911 ) | ( ~n3730 & n21816 ) | ( n6911 & n21816 ) ;
  assign n30729 = n30728 ^ n13224 ^ n10259 ;
  assign n30730 = n4246 ^ n491 ^ 1'b0 ;
  assign n30731 = n21179 & ~n30730 ;
  assign n30732 = n30731 ^ n9593 ^ 1'b0 ;
  assign n30733 = n4338 & ~n30732 ;
  assign n30734 = ( ~n6789 & n17100 ) | ( ~n6789 & n30733 ) | ( n17100 & n30733 ) ;
  assign n30735 = n9237 | n16441 ;
  assign n30736 = n5172 & ~n30735 ;
  assign n30737 = ( n15841 & n20120 ) | ( n15841 & ~n30736 ) | ( n20120 & ~n30736 ) ;
  assign n30738 = ~n4137 & n21425 ;
  assign n30739 = n30738 ^ n12356 ^ 1'b0 ;
  assign n30740 = ( n3816 & ~n6589 ) | ( n3816 & n30739 ) | ( ~n6589 & n30739 ) ;
  assign n30741 = ( n15461 & n15634 ) | ( n15461 & ~n28900 ) | ( n15634 & ~n28900 ) ;
  assign n30742 = n22301 | n30741 ;
  assign n30743 = n30742 ^ n30613 ^ n25039 ;
  assign n30744 = ( n5556 & n6281 ) | ( n5556 & n11102 ) | ( n6281 & n11102 ) ;
  assign n30745 = n30744 ^ n24891 ^ n6658 ;
  assign n30747 = ( n10584 & ~n15151 ) | ( n10584 & n20731 ) | ( ~n15151 & n20731 ) ;
  assign n30746 = n14092 ^ n6777 ^ n1211 ;
  assign n30748 = n30747 ^ n30746 ^ 1'b0 ;
  assign n30749 = n21807 | n30748 ;
  assign n30750 = ~n4936 & n5778 ;
  assign n30751 = n30750 ^ n9947 ^ n9715 ;
  assign n30752 = n30751 ^ n10407 ^ 1'b0 ;
  assign n30753 = n17704 & n30752 ;
  assign n30754 = n7670 ^ n4764 ^ 1'b0 ;
  assign n30755 = n4575 & n30754 ;
  assign n30756 = n270 & n19128 ;
  assign n30757 = n14501 ^ n11530 ^ n6381 ;
  assign n30758 = n30757 ^ n2839 ^ 1'b0 ;
  assign n30759 = n30756 & n30758 ;
  assign n30760 = ~n3038 & n6905 ;
  assign n30761 = ~n10893 & n21009 ;
  assign n30762 = ( n22778 & n30760 ) | ( n22778 & ~n30761 ) | ( n30760 & ~n30761 ) ;
  assign n30763 = ( ~n192 & n3949 ) | ( ~n192 & n12433 ) | ( n3949 & n12433 ) ;
  assign n30764 = n2876 & n16895 ;
  assign n30765 = n30763 & n30764 ;
  assign n30766 = n2813 & ~n30765 ;
  assign n30767 = n30766 ^ n10773 ^ n8387 ;
  assign n30768 = n8788 ^ n5948 ^ n3888 ;
  assign n30769 = n30768 ^ n10064 ^ n6532 ;
  assign n30771 = ( n591 & n14639 ) | ( n591 & n16549 ) | ( n14639 & n16549 ) ;
  assign n30772 = ( ~n5874 & n10997 ) | ( ~n5874 & n30771 ) | ( n10997 & n30771 ) ;
  assign n30773 = ( n23564 & n25157 ) | ( n23564 & ~n30772 ) | ( n25157 & ~n30772 ) ;
  assign n30770 = n1221 & n8404 ;
  assign n30774 = n30773 ^ n30770 ^ 1'b0 ;
  assign n30775 = n18329 & ~n29052 ;
  assign n30776 = ( n30769 & n30774 ) | ( n30769 & ~n30775 ) | ( n30774 & ~n30775 ) ;
  assign n30777 = n14038 ^ n12118 ^ 1'b0 ;
  assign n30778 = n28979 | n30777 ;
  assign n30779 = n23790 ^ n11751 ^ n1134 ;
  assign n30780 = ( n18104 & n30778 ) | ( n18104 & ~n30779 ) | ( n30778 & ~n30779 ) ;
  assign n30781 = n1242 ^ n706 ^ 1'b0 ;
  assign n30782 = n4920 | n5132 ;
  assign n30783 = ( n1958 & n13148 ) | ( n1958 & n30782 ) | ( n13148 & n30782 ) ;
  assign n30784 = ( ~n2360 & n9212 ) | ( ~n2360 & n17574 ) | ( n9212 & n17574 ) ;
  assign n30785 = n30784 ^ n24499 ^ 1'b0 ;
  assign n30786 = n21902 | n30785 ;
  assign n30787 = n5537 & n8370 ;
  assign n30788 = n30787 ^ n9164 ^ 1'b0 ;
  assign n30789 = n16096 ^ n6344 ^ 1'b0 ;
  assign n30790 = n30788 & ~n30789 ;
  assign n30791 = ( ~n21383 & n30786 ) | ( ~n21383 & n30790 ) | ( n30786 & n30790 ) ;
  assign n30792 = ( n5742 & ~n30783 ) | ( n5742 & n30791 ) | ( ~n30783 & n30791 ) ;
  assign n30793 = n14078 ^ n4664 ^ 1'b0 ;
  assign n30794 = n8285 & n16053 ;
  assign n30795 = n4930 & n30794 ;
  assign n30796 = n197 | n29175 ;
  assign n30797 = n7375 & ~n30796 ;
  assign n30798 = ( n3990 & ~n4452 ) | ( n3990 & n23692 ) | ( ~n4452 & n23692 ) ;
  assign n30799 = n8623 ^ n5556 ^ n2603 ;
  assign n30800 = ( n6000 & ~n22335 ) | ( n6000 & n26024 ) | ( ~n22335 & n26024 ) ;
  assign n30801 = ( n1480 & n4920 ) | ( n1480 & n19778 ) | ( n4920 & n19778 ) ;
  assign n30805 = n8145 & ~n25944 ;
  assign n30802 = n13589 ^ n2251 ^ 1'b0 ;
  assign n30803 = n30802 ^ n26072 ^ n7274 ;
  assign n30804 = n30803 ^ n16129 ^ 1'b0 ;
  assign n30806 = n30805 ^ n30804 ^ n26365 ;
  assign n30807 = n19310 ^ n14085 ^ 1'b0 ;
  assign n30808 = n8603 & ~n30807 ;
  assign n30809 = ( ~n17283 & n20940 ) | ( ~n17283 & n30808 ) | ( n20940 & n30808 ) ;
  assign n30810 = n21203 & ~n28256 ;
  assign n30811 = n30810 ^ x123 ^ 1'b0 ;
  assign n30812 = n10976 ^ n9534 ^ n9115 ;
  assign n30813 = n7240 & ~n30812 ;
  assign n30814 = n30813 ^ n6138 ^ 1'b0 ;
  assign n30815 = ( n852 & ~n1140 ) | ( n852 & n3666 ) | ( ~n1140 & n3666 ) ;
  assign n30816 = n30815 ^ n12934 ^ 1'b0 ;
  assign n30817 = n13746 | n30816 ;
  assign n30818 = n28556 ^ n24412 ^ n19698 ;
  assign n30819 = ( n10369 & n23350 ) | ( n10369 & ~n30818 ) | ( n23350 & ~n30818 ) ;
  assign n30820 = n18068 & n20862 ;
  assign n30821 = n17937 & n30820 ;
  assign n30822 = ( n1000 & ~n9001 ) | ( n1000 & n11170 ) | ( ~n9001 & n11170 ) ;
  assign n30823 = ( ~n11169 & n12523 ) | ( ~n11169 & n13524 ) | ( n12523 & n13524 ) ;
  assign n30824 = n30823 ^ n26905 ^ n2321 ;
  assign n30825 = ( n12331 & ~n30822 ) | ( n12331 & n30824 ) | ( ~n30822 & n30824 ) ;
  assign n30826 = n5889 | n11648 ;
  assign n30827 = n30826 ^ n9987 ^ 1'b0 ;
  assign n30828 = n30827 ^ n5080 ^ n3772 ;
  assign n30829 = n3188 & n16729 ;
  assign n30830 = ~n8998 & n30829 ;
  assign n30831 = n16042 | n30830 ;
  assign n30832 = n30831 ^ n11150 ^ 1'b0 ;
  assign n30833 = ( n12386 & n16719 ) | ( n12386 & ~n22523 ) | ( n16719 & ~n22523 ) ;
  assign n30834 = n26446 ^ n8530 ^ n1885 ;
  assign n30835 = n23087 | n30834 ;
  assign n30836 = n23209 ^ n21121 ^ 1'b0 ;
  assign n30837 = n30835 & ~n30836 ;
  assign n30838 = x6 & n15325 ;
  assign n30839 = ~n9016 & n30838 ;
  assign n30840 = n3179 & ~n5069 ;
  assign n30841 = n15156 & n30840 ;
  assign n30842 = ( n4724 & n14053 ) | ( n4724 & n25010 ) | ( n14053 & n25010 ) ;
  assign n30843 = ( n13066 & n14567 ) | ( n13066 & n28485 ) | ( n14567 & n28485 ) ;
  assign n30844 = n28598 | n30843 ;
  assign n30845 = ( n7576 & ~n30842 ) | ( n7576 & n30844 ) | ( ~n30842 & n30844 ) ;
  assign n30846 = ( n1089 & ~n3675 ) | ( n1089 & n30081 ) | ( ~n3675 & n30081 ) ;
  assign n30847 = n20238 ^ n17111 ^ n471 ;
  assign n30848 = ( ~n2421 & n13715 ) | ( ~n2421 & n23346 ) | ( n13715 & n23346 ) ;
  assign n30849 = ( ~n13722 & n30847 ) | ( ~n13722 & n30848 ) | ( n30847 & n30848 ) ;
  assign n30850 = n9834 ^ n2490 ^ n2101 ;
  assign n30851 = n30850 ^ n11900 ^ n9949 ;
  assign n30852 = n1402 | n6055 ;
  assign n30853 = n1989 | n30852 ;
  assign n30854 = ( ~n6165 & n16619 ) | ( ~n6165 & n30853 ) | ( n16619 & n30853 ) ;
  assign n30855 = ( n16654 & n17742 ) | ( n16654 & n30854 ) | ( n17742 & n30854 ) ;
  assign n30856 = n15791 ^ n3997 ^ 1'b0 ;
  assign n30857 = n9666 & ~n30856 ;
  assign n30858 = n30857 ^ n11051 ^ 1'b0 ;
  assign n30859 = n21017 ^ n14885 ^ 1'b0 ;
  assign n30860 = n14258 | n30859 ;
  assign n30861 = n7320 & n9620 ;
  assign n30862 = n30861 ^ n29631 ^ 1'b0 ;
  assign n30863 = ~n1120 & n30430 ;
  assign n30864 = ( n1630 & ~n3595 ) | ( n1630 & n30863 ) | ( ~n3595 & n30863 ) ;
  assign n30865 = n16576 & n17307 ;
  assign n30866 = n30865 ^ n12811 ^ n2648 ;
  assign n30867 = n30866 ^ n21952 ^ 1'b0 ;
  assign n30868 = ( ~n6481 & n10042 ) | ( ~n6481 & n14657 ) | ( n10042 & n14657 ) ;
  assign n30869 = n23920 ^ n8262 ^ n2275 ;
  assign n30870 = n30869 ^ n22834 ^ n20878 ;
  assign n30871 = n30870 ^ n11917 ^ n5748 ;
  assign n30872 = n9478 & n26879 ;
  assign n30873 = n30872 ^ n27301 ^ 1'b0 ;
  assign n30874 = ( n648 & n9544 ) | ( n648 & n11777 ) | ( n9544 & n11777 ) ;
  assign n30875 = n30874 ^ n21133 ^ n11042 ;
  assign n30876 = ( n2769 & ~n13125 ) | ( n2769 & n29352 ) | ( ~n13125 & n29352 ) ;
  assign n30877 = n2389 | n30876 ;
  assign n30878 = n30875 | n30877 ;
  assign n30879 = ( n7944 & ~n13831 ) | ( n7944 & n22392 ) | ( ~n13831 & n22392 ) ;
  assign n30880 = ( n13500 & n21176 ) | ( n13500 & ~n24584 ) | ( n21176 & ~n24584 ) ;
  assign n30884 = ( ~n1359 & n24328 ) | ( ~n1359 & n29709 ) | ( n24328 & n29709 ) ;
  assign n30881 = n21518 ^ n12053 ^ 1'b0 ;
  assign n30882 = n214 & n30881 ;
  assign n30883 = n3837 & n30882 ;
  assign n30885 = n30884 ^ n30883 ^ n20333 ;
  assign n30886 = ( n4893 & n16988 ) | ( n4893 & ~n28465 ) | ( n16988 & ~n28465 ) ;
  assign n30887 = ~n22850 & n26499 ;
  assign n30888 = n12979 & n30887 ;
  assign n30889 = ( ~n467 & n18522 ) | ( ~n467 & n30888 ) | ( n18522 & n30888 ) ;
  assign n30890 = ( x52 & n10587 ) | ( x52 & n16354 ) | ( n10587 & n16354 ) ;
  assign n30891 = ( x5 & n19595 ) | ( x5 & n22814 ) | ( n19595 & n22814 ) ;
  assign n30892 = n30891 ^ n24000 ^ n10374 ;
  assign n30893 = n3651 & n10129 ;
  assign n30894 = ~n8400 & n30893 ;
  assign n30895 = n2260 ^ n716 ^ 1'b0 ;
  assign n30896 = ( n1936 & ~n9115 ) | ( n1936 & n13995 ) | ( ~n9115 & n13995 ) ;
  assign n30897 = n30896 ^ n2940 ^ 1'b0 ;
  assign n30898 = n9813 | n30897 ;
  assign n30899 = ( ~n4079 & n4429 ) | ( ~n4079 & n10353 ) | ( n4429 & n10353 ) ;
  assign n30900 = n18240 ^ n2897 ^ 1'b0 ;
  assign n30901 = ~n2957 & n30900 ;
  assign n30902 = ( n11540 & n19397 ) | ( n11540 & n22276 ) | ( n19397 & n22276 ) ;
  assign n30903 = n30901 & n30902 ;
  assign n30906 = n17211 ^ n3799 ^ 1'b0 ;
  assign n30904 = n6096 ^ n3752 ^ 1'b0 ;
  assign n30905 = ~n14614 & n30904 ;
  assign n30907 = n30906 ^ n30905 ^ n5711 ;
  assign n30908 = n24182 ^ n13894 ^ 1'b0 ;
  assign n30909 = n15217 & ~n30908 ;
  assign n30910 = n30909 ^ n30315 ^ n4191 ;
  assign n30911 = n4681 | n16884 ;
  assign n30912 = n13073 & n19356 ;
  assign n30913 = ( ~n11986 & n13489 ) | ( ~n11986 & n18706 ) | ( n13489 & n18706 ) ;
  assign n30914 = ( ~n2375 & n13999 ) | ( ~n2375 & n30913 ) | ( n13999 & n30913 ) ;
  assign n30915 = n21051 ^ n10922 ^ n9586 ;
  assign n30916 = ( ~n4589 & n19704 ) | ( ~n4589 & n30915 ) | ( n19704 & n30915 ) ;
  assign n30917 = n8320 | n13556 ;
  assign n30918 = n30916 | n30917 ;
  assign n30919 = n11354 & ~n13540 ;
  assign n30920 = n2047 & n30919 ;
  assign n30921 = ( n7046 & n19983 ) | ( n7046 & n27548 ) | ( n19983 & n27548 ) ;
  assign n30922 = n7571 & ~n11577 ;
  assign n30923 = n30922 ^ n24735 ^ n245 ;
  assign n30925 = n7563 ^ n5156 ^ 1'b0 ;
  assign n30926 = ~n9475 & n30925 ;
  assign n30927 = n1551 & n30926 ;
  assign n30924 = ( ~n923 & n2670 ) | ( ~n923 & n5896 ) | ( n2670 & n5896 ) ;
  assign n30928 = n30927 ^ n30924 ^ n7012 ;
  assign n30929 = n24244 ^ n8844 ^ n5269 ;
  assign n30930 = ( n5928 & n17777 ) | ( n5928 & ~n30929 ) | ( n17777 & ~n30929 ) ;
  assign n30931 = ( n11133 & ~n13907 ) | ( n11133 & n14451 ) | ( ~n13907 & n14451 ) ;
  assign n30932 = n21989 ^ n9869 ^ n8625 ;
  assign n30933 = n1260 & n2412 ;
  assign n30934 = n28148 ^ n7115 ^ 1'b0 ;
  assign n30935 = ~n20810 & n30934 ;
  assign n30936 = n8335 & ~n29525 ;
  assign n30937 = n30936 ^ n2860 ^ 1'b0 ;
  assign n30938 = ( n478 & n3495 ) | ( n478 & ~n4405 ) | ( n3495 & ~n4405 ) ;
  assign n30939 = n30938 ^ n30112 ^ n6167 ;
  assign n30940 = n24185 ^ n9501 ^ n3395 ;
  assign n30941 = ( n3979 & n6976 ) | ( n3979 & n23006 ) | ( n6976 & n23006 ) ;
  assign n30942 = ( n838 & ~n16298 ) | ( n838 & n16761 ) | ( ~n16298 & n16761 ) ;
  assign n30943 = n14194 ^ n9657 ^ n8343 ;
  assign n30944 = n29838 ^ n13881 ^ 1'b0 ;
  assign n30945 = n869 | n5259 ;
  assign n30946 = n30945 ^ n12215 ^ 1'b0 ;
  assign n30947 = n30946 ^ n20468 ^ n2262 ;
  assign n30948 = n17930 | n20399 ;
  assign n30949 = ~n6189 & n6766 ;
  assign n30950 = n16252 ^ n7476 ^ n330 ;
  assign n30951 = n30950 ^ n25022 ^ 1'b0 ;
  assign n30952 = n20120 | n30951 ;
  assign n30953 = n30952 ^ n11862 ^ n7816 ;
  assign n30954 = n8037 & ~n15697 ;
  assign n30955 = ~n10333 & n30954 ;
  assign n30956 = ( n14761 & n25967 ) | ( n14761 & ~n30955 ) | ( n25967 & ~n30955 ) ;
  assign n30957 = ( ~n5106 & n10386 ) | ( ~n5106 & n30956 ) | ( n10386 & n30956 ) ;
  assign n30958 = ( x67 & n18876 ) | ( x67 & ~n24230 ) | ( n18876 & ~n24230 ) ;
  assign n30959 = n23844 ^ n23746 ^ n3321 ;
  assign n30960 = n4179 & n15664 ;
  assign n30961 = n30960 ^ n11633 ^ n6146 ;
  assign n30962 = n5412 & ~n11716 ;
  assign n30963 = n6371 | n8359 ;
  assign n30964 = n16421 & ~n30963 ;
  assign n30965 = n6014 & n9458 ;
  assign n30966 = n30965 ^ n4061 ^ 1'b0 ;
  assign n30967 = n17535 ^ n12189 ^ 1'b0 ;
  assign n30968 = n1934 & n30967 ;
  assign n30969 = n30968 ^ n20946 ^ n17506 ;
  assign n30970 = n30969 ^ n1957 ^ n173 ;
  assign n30971 = n16819 ^ n6773 ^ n6222 ;
  assign n30972 = n30971 ^ n28601 ^ n9643 ;
  assign n30973 = n30972 ^ n22858 ^ n21043 ;
  assign n30974 = n17514 ^ n5390 ^ 1'b0 ;
  assign n30975 = n5024 & ~n30974 ;
  assign n30976 = n2888 & ~n3196 ;
  assign n30977 = n30976 ^ n1607 ^ 1'b0 ;
  assign n30978 = n30977 ^ n15345 ^ n4325 ;
  assign n30979 = n30978 ^ n30017 ^ 1'b0 ;
  assign n30980 = n7177 & n30979 ;
  assign n30981 = n19229 ^ n8201 ^ n3219 ;
  assign n30982 = ( n30975 & ~n30980 ) | ( n30975 & n30981 ) | ( ~n30980 & n30981 ) ;
  assign n30983 = n29854 ^ n24287 ^ n13414 ;
  assign n30984 = n10992 ^ n10573 ^ 1'b0 ;
  assign n30985 = n30984 ^ n14734 ^ n12375 ;
  assign n30986 = n17704 ^ n10374 ^ n5883 ;
  assign n30987 = n22276 ^ n21173 ^ n1745 ;
  assign n30988 = n30987 ^ n22626 ^ n898 ;
  assign n30989 = n24596 | n30988 ;
  assign n30991 = n22280 ^ n12943 ^ 1'b0 ;
  assign n30992 = n12816 | n30991 ;
  assign n30993 = n30992 ^ n12817 ^ n10062 ;
  assign n30990 = n1450 | n16874 ;
  assign n30994 = n30993 ^ n30990 ^ 1'b0 ;
  assign n30995 = ( n4513 & ~n6016 ) | ( n4513 & n11078 ) | ( ~n6016 & n11078 ) ;
  assign n30996 = n8370 & n30995 ;
  assign n30997 = n30996 ^ n25375 ^ 1'b0 ;
  assign n30998 = n24180 ^ n3465 ^ 1'b0 ;
  assign n30999 = n12469 & n30998 ;
  assign n31001 = ( ~n2033 & n21047 ) | ( ~n2033 & n23940 ) | ( n21047 & n23940 ) ;
  assign n31002 = ( ~n13135 & n29475 ) | ( ~n13135 & n31001 ) | ( n29475 & n31001 ) ;
  assign n31000 = n3965 & n12889 ;
  assign n31003 = n31002 ^ n31000 ^ 1'b0 ;
  assign n31004 = n15453 ^ n11277 ^ 1'b0 ;
  assign n31005 = n27350 ^ n7844 ^ n2888 ;
  assign n31008 = ~n5070 & n26580 ;
  assign n31009 = ~n5684 & n31008 ;
  assign n31006 = ~n1890 & n12927 ;
  assign n31007 = n31006 ^ n4797 ^ 1'b0 ;
  assign n31010 = n31009 ^ n31007 ^ n15228 ;
  assign n31011 = n27011 ^ n4650 ^ 1'b0 ;
  assign n31012 = ( n13547 & n29375 ) | ( n13547 & ~n31011 ) | ( n29375 & ~n31011 ) ;
  assign n31013 = n11735 & n25204 ;
  assign n31014 = ( ~n3952 & n7641 ) | ( ~n3952 & n31013 ) | ( n7641 & n31013 ) ;
  assign n31015 = ( n7173 & ~n7346 ) | ( n7173 & n8899 ) | ( ~n7346 & n8899 ) ;
  assign n31016 = n31015 ^ n22919 ^ n6785 ;
  assign n31017 = ( ~n23546 & n30827 ) | ( ~n23546 & n31016 ) | ( n30827 & n31016 ) ;
  assign n31018 = n26358 ^ n22913 ^ 1'b0 ;
  assign n31019 = ~n9167 & n31018 ;
  assign n31020 = n12909 ^ n8545 ^ 1'b0 ;
  assign n31021 = ~n2049 & n31020 ;
  assign n31022 = n5219 & n31021 ;
  assign n31023 = n12528 & ~n12529 ;
  assign n31024 = ~n7427 & n31023 ;
  assign n31025 = ( n7875 & n22065 ) | ( n7875 & ~n24437 ) | ( n22065 & ~n24437 ) ;
  assign n31026 = n27871 ^ n8728 ^ n6129 ;
  assign n31028 = n13825 ^ n5176 ^ n371 ;
  assign n31027 = ~n5291 & n27356 ;
  assign n31029 = n31028 ^ n31027 ^ 1'b0 ;
  assign n31030 = n31029 ^ n25654 ^ n10460 ;
  assign n31031 = n31030 ^ n20454 ^ 1'b0 ;
  assign n31032 = ( n2256 & n4150 ) | ( n2256 & ~n10532 ) | ( n4150 & ~n10532 ) ;
  assign n31033 = n14782 & ~n31032 ;
  assign n31034 = n31033 ^ n6431 ^ 1'b0 ;
  assign n31035 = ( n13492 & ~n22525 ) | ( n13492 & n31034 ) | ( ~n22525 & n31034 ) ;
  assign n31036 = ( ~n2041 & n16260 ) | ( ~n2041 & n22425 ) | ( n16260 & n22425 ) ;
  assign n31037 = n23351 ^ n8252 ^ 1'b0 ;
  assign n31038 = n23290 ^ n7467 ^ n1242 ;
  assign n31039 = ( n11159 & ~n17843 ) | ( n11159 & n31038 ) | ( ~n17843 & n31038 ) ;
  assign n31040 = n5686 ^ n4129 ^ 1'b0 ;
  assign n31041 = n7399 & n31040 ;
  assign n31042 = n31041 ^ n3200 ^ 1'b0 ;
  assign n31043 = n22931 & ~n29713 ;
  assign n31044 = n31043 ^ n29868 ^ 1'b0 ;
  assign n31045 = n29829 ^ n29524 ^ n2729 ;
  assign n31046 = n8759 ^ n7961 ^ n3049 ;
  assign n31047 = ( n395 & n14007 ) | ( n395 & n31046 ) | ( n14007 & n31046 ) ;
  assign n31048 = n7269 ^ n6910 ^ n1618 ;
  assign n31049 = ( n7992 & ~n15221 ) | ( n7992 & n19492 ) | ( ~n15221 & n19492 ) ;
  assign n31050 = n822 & ~n15671 ;
  assign n31051 = ~n7208 & n31050 ;
  assign n31052 = ( n31048 & n31049 ) | ( n31048 & ~n31051 ) | ( n31049 & ~n31051 ) ;
  assign n31053 = n7301 ^ n5659 ^ n2876 ;
  assign n31054 = n22729 ^ n4845 ^ n2157 ;
  assign n31055 = ( n14368 & ~n29728 ) | ( n14368 & n31054 ) | ( ~n29728 & n31054 ) ;
  assign n31056 = n8096 ^ n588 ^ n541 ;
  assign n31057 = ( n866 & n1434 ) | ( n866 & n15115 ) | ( n1434 & n15115 ) ;
  assign n31058 = n31057 ^ n15397 ^ 1'b0 ;
  assign n31059 = n3174 & ~n3187 ;
  assign n31060 = n25241 & n31059 ;
  assign n31061 = ~n7206 & n16060 ;
  assign n31062 = ~n22510 & n31061 ;
  assign n31063 = ( n9682 & ~n16336 ) | ( n9682 & n23802 ) | ( ~n16336 & n23802 ) ;
  assign n31064 = n31063 ^ n22279 ^ 1'b0 ;
  assign n31066 = n24070 ^ n2664 ^ 1'b0 ;
  assign n31065 = ( n6552 & n16599 ) | ( n6552 & ~n16966 ) | ( n16599 & ~n16966 ) ;
  assign n31067 = n31066 ^ n31065 ^ n15110 ;
  assign n31068 = n31067 ^ n22692 ^ n16508 ;
  assign n31069 = n7657 ^ n4437 ^ n2772 ;
  assign n31070 = ( ~n3532 & n7332 ) | ( ~n3532 & n31069 ) | ( n7332 & n31069 ) ;
  assign n31071 = n14824 ^ n3022 ^ n1507 ;
  assign n31072 = n31071 ^ n21476 ^ 1'b0 ;
  assign n31073 = n31072 ^ n21567 ^ n12029 ;
  assign n31075 = n5139 & n9625 ;
  assign n31076 = n31075 ^ n4111 ^ 1'b0 ;
  assign n31077 = n11370 ^ n8809 ^ 1'b0 ;
  assign n31078 = n31076 | n31077 ;
  assign n31079 = n14727 & ~n31078 ;
  assign n31074 = n5373 & ~n6020 ;
  assign n31080 = n31079 ^ n31074 ^ 1'b0 ;
  assign n31081 = n4092 & n8802 ;
  assign n31082 = ( ~n3466 & n31080 ) | ( ~n3466 & n31081 ) | ( n31080 & n31081 ) ;
  assign n31086 = n21617 ^ n11414 ^ n4416 ;
  assign n31083 = n15993 ^ n10002 ^ n1999 ;
  assign n31084 = ( n8570 & n9026 ) | ( n8570 & ~n31083 ) | ( n9026 & ~n31083 ) ;
  assign n31085 = n31084 ^ n28368 ^ n9194 ;
  assign n31087 = n31086 ^ n31085 ^ n25858 ;
  assign n31088 = n4549 ^ n502 ^ 1'b0 ;
  assign n31089 = n31088 ^ n30898 ^ 1'b0 ;
  assign n31090 = n22287 & n31089 ;
  assign n31091 = n6714 ^ n3588 ^ 1'b0 ;
  assign n31092 = n28433 & ~n31091 ;
  assign n31093 = ~n4906 & n7047 ;
  assign n31094 = ~n31092 & n31093 ;
  assign n31095 = ~n1093 & n28401 ;
  assign n31096 = n31095 ^ n7683 ^ 1'b0 ;
  assign n31097 = ( ~n1620 & n5609 ) | ( ~n1620 & n8203 ) | ( n5609 & n8203 ) ;
  assign n31098 = n31097 ^ n16045 ^ n13508 ;
  assign n31099 = n18880 ^ n18601 ^ n8277 ;
  assign n31100 = n31099 ^ n30058 ^ n15985 ;
  assign n31109 = n14786 ^ n9254 ^ n4048 ;
  assign n31102 = ( n620 & ~n3511 ) | ( n620 & n15159 ) | ( ~n3511 & n15159 ) ;
  assign n31103 = ( n8116 & n10777 ) | ( n8116 & n31102 ) | ( n10777 & n31102 ) ;
  assign n31104 = n31103 ^ n27945 ^ 1'b0 ;
  assign n31105 = n8725 & ~n31104 ;
  assign n31106 = n31105 ^ n19495 ^ 1'b0 ;
  assign n31107 = n8356 & n31106 ;
  assign n31101 = ( n2070 & ~n20593 ) | ( n2070 & n28092 ) | ( ~n20593 & n28092 ) ;
  assign n31108 = n31107 ^ n31101 ^ 1'b0 ;
  assign n31110 = n31109 ^ n31108 ^ n13453 ;
  assign n31111 = ( n5566 & n23524 ) | ( n5566 & n25558 ) | ( n23524 & n25558 ) ;
  assign n31112 = ( n5131 & n10493 ) | ( n5131 & n19889 ) | ( n10493 & n19889 ) ;
  assign n31113 = ~n10197 & n10942 ;
  assign n31114 = n27030 ^ n8164 ^ n5554 ;
  assign n31115 = n31114 ^ n3421 ^ 1'b0 ;
  assign n31116 = ~n14063 & n31115 ;
  assign n31117 = n1381 & n13295 ;
  assign n31118 = n31117 ^ n21408 ^ n14474 ;
  assign n31119 = ( n5780 & n31116 ) | ( n5780 & ~n31118 ) | ( n31116 & ~n31118 ) ;
  assign n31120 = n2910 & n17379 ;
  assign n31121 = ~n21576 & n31120 ;
  assign n31122 = n22398 ^ n21595 ^ n21470 ;
  assign n31123 = ~n25706 & n31122 ;
  assign n31124 = n20159 ^ x34 ^ 1'b0 ;
  assign n31125 = n23008 ^ n8615 ^ n3460 ;
  assign n31126 = ( ~n605 & n12360 ) | ( ~n605 & n17199 ) | ( n12360 & n17199 ) ;
  assign n31127 = ( n17788 & ~n28031 ) | ( n17788 & n31126 ) | ( ~n28031 & n31126 ) ;
  assign n31128 = ( ~n3790 & n16314 ) | ( ~n3790 & n26681 ) | ( n16314 & n26681 ) ;
  assign n31129 = ( n3065 & ~n5586 ) | ( n3065 & n8539 ) | ( ~n5586 & n8539 ) ;
  assign n31130 = n31129 ^ n5683 ^ 1'b0 ;
  assign n31131 = n9233 & ~n16980 ;
  assign n31132 = n5979 & n20689 ;
  assign n31133 = n2683 ^ n1971 ^ 1'b0 ;
  assign n31134 = ~n384 & n31133 ;
  assign n31135 = n14065 ^ n3881 ^ 1'b0 ;
  assign n31136 = ( n2860 & ~n7788 ) | ( n2860 & n16516 ) | ( ~n7788 & n16516 ) ;
  assign n31137 = n31136 ^ n21667 ^ n1107 ;
  assign n31138 = ( ~n1581 & n9600 ) | ( ~n1581 & n10739 ) | ( n9600 & n10739 ) ;
  assign n31139 = n14069 ^ n635 ^ 1'b0 ;
  assign n31140 = ( n3529 & ~n18928 ) | ( n3529 & n31139 ) | ( ~n18928 & n31139 ) ;
  assign n31141 = n31140 ^ n12878 ^ n3203 ;
  assign n31142 = n12183 ^ n7371 ^ n7323 ;
  assign n31143 = n24119 ^ n8746 ^ n3657 ;
  assign n31144 = n31143 ^ n21175 ^ n4015 ;
  assign n31145 = ( n1016 & n7443 ) | ( n1016 & ~n13865 ) | ( n7443 & ~n13865 ) ;
  assign n31146 = ~n11732 & n31145 ;
  assign n31147 = n31146 ^ n22291 ^ 1'b0 ;
  assign n31148 = n9432 & ~n9579 ;
  assign n31149 = n31148 ^ n17853 ^ 1'b0 ;
  assign n31151 = ( ~n10691 & n21879 ) | ( ~n10691 & n30309 ) | ( n21879 & n30309 ) ;
  assign n31150 = n15692 & ~n21556 ;
  assign n31152 = n31151 ^ n31150 ^ n6360 ;
  assign n31155 = n3161 & n12793 ;
  assign n31156 = n31155 ^ n13704 ^ 1'b0 ;
  assign n31154 = n4143 | n9883 ;
  assign n31153 = n13628 ^ n13547 ^ n7652 ;
  assign n31157 = n31156 ^ n31154 ^ n31153 ;
  assign n31158 = n21821 ^ n17093 ^ n14464 ;
  assign n31159 = ( n15768 & n23743 ) | ( n15768 & n30376 ) | ( n23743 & n30376 ) ;
  assign n31160 = ~n3966 & n11600 ;
  assign n31161 = n31160 ^ n7822 ^ 1'b0 ;
  assign n31162 = ( n3906 & ~n15241 ) | ( n3906 & n31161 ) | ( ~n15241 & n31161 ) ;
  assign n31163 = ( n1982 & ~n8690 ) | ( n1982 & n9738 ) | ( ~n8690 & n9738 ) ;
  assign n31166 = ( n950 & n4330 ) | ( n950 & n10732 ) | ( n4330 & n10732 ) ;
  assign n31164 = n14946 ^ n4768 ^ n2376 ;
  assign n31165 = n6647 & n31164 ;
  assign n31167 = n31166 ^ n31165 ^ 1'b0 ;
  assign n31168 = ~n22693 & n31167 ;
  assign n31169 = n8350 & ~n20069 ;
  assign n31170 = n27558 ^ n3747 ^ 1'b0 ;
  assign n31171 = n28855 ^ n13886 ^ 1'b0 ;
  assign n31172 = n8029 ^ n5300 ^ 1'b0 ;
  assign n31173 = n22634 | n31172 ;
  assign n31174 = n31173 ^ n2373 ^ 1'b0 ;
  assign n31175 = n31174 ^ n21232 ^ n19371 ;
  assign n31176 = ( n8241 & n17994 ) | ( n8241 & n29508 ) | ( n17994 & n29508 ) ;
  assign n31177 = n7959 & ~n22943 ;
  assign n31178 = n19933 ^ n7126 ^ 1'b0 ;
  assign n31179 = n6399 | n31178 ;
  assign n31180 = n31179 ^ n27861 ^ 1'b0 ;
  assign n31182 = n13936 ^ n12602 ^ n7275 ;
  assign n31181 = n12555 | n20812 ;
  assign n31183 = n31182 ^ n31181 ^ n20566 ;
  assign n31184 = ~n5715 & n10179 ;
  assign n31185 = ~n25437 & n31184 ;
  assign n31186 = n18028 ^ n15957 ^ n770 ;
  assign n31187 = n31186 ^ n7051 ^ 1'b0 ;
  assign n31188 = n24809 | n31187 ;
  assign n31189 = n2375 & n19060 ;
  assign n31190 = n31189 ^ n1989 ^ 1'b0 ;
  assign n31191 = ~n230 & n10605 ;
  assign n31192 = n31191 ^ n9651 ^ 1'b0 ;
  assign n31193 = n31192 ^ n14423 ^ n10449 ;
  assign n31194 = n23345 ^ n17315 ^ n572 ;
  assign n31195 = ( n1851 & ~n8498 ) | ( n1851 & n31194 ) | ( ~n8498 & n31194 ) ;
  assign n31196 = n27699 ^ n11828 ^ n10092 ;
  assign n31197 = n31196 ^ n15917 ^ n12416 ;
  assign n31198 = n16281 ^ n14272 ^ 1'b0 ;
  assign n31199 = n6078 & ~n28266 ;
  assign n31200 = n30006 ^ n21731 ^ 1'b0 ;
  assign n31202 = ( ~n7173 & n18375 ) | ( ~n7173 & n19837 ) | ( n18375 & n19837 ) ;
  assign n31201 = n27989 & ~n28568 ;
  assign n31203 = n31202 ^ n31201 ^ 1'b0 ;
  assign n31204 = x67 & n24487 ;
  assign n31205 = n16856 & n31204 ;
  assign n31206 = n19077 & ~n21594 ;
  assign n31207 = n31206 ^ n20065 ^ 1'b0 ;
  assign n31208 = n10609 | n28787 ;
  assign n31209 = n29905 | n31208 ;
  assign n31210 = n16052 ^ n14887 ^ 1'b0 ;
  assign n31211 = n4520 & n31210 ;
  assign n31212 = n31211 ^ n21045 ^ n10383 ;
  assign n31213 = ( n7448 & ~n24654 ) | ( n7448 & n31212 ) | ( ~n24654 & n31212 ) ;
  assign n31214 = n12755 ^ n3904 ^ n1753 ;
  assign n31215 = ~n8135 & n10461 ;
  assign n31216 = n31214 & n31215 ;
  assign n31217 = n15248 | n31216 ;
  assign n31218 = n31217 ^ n29140 ^ n21712 ;
  assign n31219 = ( n7066 & n10926 ) | ( n7066 & ~n31218 ) | ( n10926 & ~n31218 ) ;
  assign n31220 = n10440 ^ n10344 ^ n1185 ;
  assign n31221 = n28897 ^ n21331 ^ 1'b0 ;
  assign n31222 = n5434 | n31221 ;
  assign n31223 = ( n20135 & n31220 ) | ( n20135 & ~n31222 ) | ( n31220 & ~n31222 ) ;
  assign n31225 = n2986 & ~n12586 ;
  assign n31224 = n175 & ~n22547 ;
  assign n31226 = n31225 ^ n31224 ^ 1'b0 ;
  assign n31227 = n14085 ^ n7569 ^ n7176 ;
  assign n31228 = ( n4721 & n11086 ) | ( n4721 & ~n31227 ) | ( n11086 & ~n31227 ) ;
  assign n31229 = n14423 ^ n7254 ^ n3340 ;
  assign n31230 = n31229 ^ n10535 ^ 1'b0 ;
  assign n31231 = n27712 ^ n8340 ^ n6354 ;
  assign n31233 = n16693 ^ n11528 ^ n5905 ;
  assign n31234 = n31233 ^ n26679 ^ n4758 ;
  assign n31235 = ~n1158 & n31234 ;
  assign n31232 = n8136 & n19974 ;
  assign n31236 = n31235 ^ n31232 ^ 1'b0 ;
  assign n31237 = n7417 & ~n10413 ;
  assign n31238 = n31237 ^ n4770 ^ 1'b0 ;
  assign n31239 = ( n2721 & ~n21823 ) | ( n2721 & n31238 ) | ( ~n21823 & n31238 ) ;
  assign n31240 = n31239 ^ n18883 ^ 1'b0 ;
  assign n31242 = n27945 ^ n8552 ^ n1653 ;
  assign n31241 = n24315 ^ n23822 ^ n981 ;
  assign n31243 = n31242 ^ n31241 ^ n30560 ;
  assign n31244 = n2138 & n19375 ;
  assign n31245 = n8630 & n31244 ;
  assign n31246 = ( n676 & ~n3998 ) | ( n676 & n31245 ) | ( ~n3998 & n31245 ) ;
  assign n31247 = n31246 ^ n7862 ^ 1'b0 ;
  assign n31248 = ( ~n4311 & n7080 ) | ( ~n4311 & n22475 ) | ( n7080 & n22475 ) ;
  assign n31251 = n5924 & ~n8433 ;
  assign n31249 = n28529 ^ n4431 ^ 1'b0 ;
  assign n31250 = n11998 & n31249 ;
  assign n31252 = n31251 ^ n31250 ^ n8412 ;
  assign n31253 = n31252 ^ n22636 ^ n6790 ;
  assign n31254 = ( n16400 & n23770 ) | ( n16400 & ~n25961 ) | ( n23770 & ~n25961 ) ;
  assign n31255 = ( n3293 & n4878 ) | ( n3293 & ~n6094 ) | ( n4878 & ~n6094 ) ;
  assign n31256 = n4014 | n16567 ;
  assign n31257 = n31256 ^ n3495 ^ 1'b0 ;
  assign n31258 = n31255 & n31257 ;
  assign n31259 = ( ~n3831 & n10343 ) | ( ~n3831 & n31258 ) | ( n10343 & n31258 ) ;
  assign n31260 = n29586 ^ n2526 ^ 1'b0 ;
  assign n31261 = ~n6813 & n31260 ;
  assign n31262 = n18826 ^ n9517 ^ 1'b0 ;
  assign n31263 = n10585 & ~n31262 ;
  assign n31264 = ~n10931 & n29776 ;
  assign n31265 = n31264 ^ n20418 ^ 1'b0 ;
  assign n31266 = ~n19802 & n31265 ;
  assign n31268 = ~n7031 & n17528 ;
  assign n31269 = n31268 ^ n11450 ^ 1'b0 ;
  assign n31267 = n2000 & n20071 ;
  assign n31270 = n31269 ^ n31267 ^ 1'b0 ;
  assign n31271 = n27729 ^ n11182 ^ n1808 ;
  assign n31272 = n6845 & n28275 ;
  assign n31273 = n31272 ^ n29227 ^ 1'b0 ;
  assign n31274 = ( n3518 & n23822 ) | ( n3518 & n31273 ) | ( n23822 & n31273 ) ;
  assign n31275 = n27191 ^ n10452 ^ n2648 ;
  assign n31276 = ( n3179 & n10805 ) | ( n3179 & n31275 ) | ( n10805 & n31275 ) ;
  assign n31277 = n31276 ^ n20933 ^ 1'b0 ;
  assign n31278 = n31277 ^ n14357 ^ 1'b0 ;
  assign n31279 = n758 & ~n11738 ;
  assign n31280 = n16450 ^ n2367 ^ 1'b0 ;
  assign n31281 = ( ~n13466 & n25872 ) | ( ~n13466 & n31280 ) | ( n25872 & n31280 ) ;
  assign n31284 = n7661 ^ n3380 ^ n1430 ;
  assign n31285 = ( n6419 & ~n15900 ) | ( n6419 & n31284 ) | ( ~n15900 & n31284 ) ;
  assign n31286 = ( n12852 & n30977 ) | ( n12852 & ~n31285 ) | ( n30977 & ~n31285 ) ;
  assign n31282 = n27894 ^ n22016 ^ n9330 ;
  assign n31283 = n31282 ^ n18855 ^ 1'b0 ;
  assign n31287 = n31286 ^ n31283 ^ n8867 ;
  assign n31288 = ~n27043 & n31287 ;
  assign n31289 = ~n7404 & n31288 ;
  assign n31290 = n31289 ^ n21663 ^ 1'b0 ;
  assign n31291 = n11401 & n15395 ;
  assign n31292 = ~n16675 & n31291 ;
  assign n31293 = n22414 ^ n18298 ^ 1'b0 ;
  assign n31294 = n5790 & ~n5800 ;
  assign n31295 = ~n28181 & n31294 ;
  assign n31296 = n30470 & ~n31295 ;
  assign n31297 = n3308 | n23817 ;
  assign n31298 = n31296 | n31297 ;
  assign n31299 = n3413 | n29410 ;
  assign n31300 = n31298 | n31299 ;
  assign n31301 = ( n3316 & n5535 ) | ( n3316 & ~n12682 ) | ( n5535 & ~n12682 ) ;
  assign n31302 = n31301 ^ n17881 ^ n16187 ;
  assign n31303 = n31302 ^ n17854 ^ n5254 ;
  assign n31304 = ( n5201 & n15434 ) | ( n5201 & ~n22485 ) | ( n15434 & ~n22485 ) ;
  assign n31305 = ( n18961 & n26577 ) | ( n18961 & ~n31304 ) | ( n26577 & ~n31304 ) ;
  assign n31306 = n31305 ^ n16270 ^ n3261 ;
  assign n31307 = n3382 & n25280 ;
  assign n31309 = n6067 & ~n16134 ;
  assign n31310 = n6724 & n31309 ;
  assign n31308 = ( n7537 & n8443 ) | ( n7537 & n18095 ) | ( n8443 & n18095 ) ;
  assign n31311 = n31310 ^ n31308 ^ n5491 ;
  assign n31312 = n25448 ^ n13815 ^ n3798 ;
  assign n31313 = ( n10133 & ~n16676 ) | ( n10133 & n24061 ) | ( ~n16676 & n24061 ) ;
  assign n31314 = ( n2646 & n4389 ) | ( n2646 & ~n24367 ) | ( n4389 & ~n24367 ) ;
  assign n31315 = n184 | n31314 ;
  assign n31316 = n31315 ^ n12288 ^ 1'b0 ;
  assign n31317 = n31316 ^ n29527 ^ n25607 ;
  assign n31318 = ( n16339 & ~n28950 ) | ( n16339 & n31317 ) | ( ~n28950 & n31317 ) ;
  assign n31319 = ( n2052 & ~n4425 ) | ( n2052 & n5397 ) | ( ~n4425 & n5397 ) ;
  assign n31320 = n24334 ^ n16984 ^ n4032 ;
  assign n31321 = ( n18514 & ~n31319 ) | ( n18514 & n31320 ) | ( ~n31319 & n31320 ) ;
  assign n31322 = n31321 ^ n15880 ^ n3310 ;
  assign n31323 = ~n9801 & n31322 ;
  assign n31324 = n31323 ^ n807 ^ 1'b0 ;
  assign n31325 = n5960 ^ n209 ^ 1'b0 ;
  assign n31326 = ~n26341 & n31325 ;
  assign n31327 = n6726 ^ n704 ^ 1'b0 ;
  assign n31328 = n919 & ~n31327 ;
  assign n31329 = n15736 ^ n8205 ^ n6992 ;
  assign n31330 = n31329 ^ n28920 ^ n10140 ;
  assign n31331 = n18662 ^ n6346 ^ 1'b0 ;
  assign n31332 = ( n15449 & n16157 ) | ( n15449 & n31331 ) | ( n16157 & n31331 ) ;
  assign n31335 = n31143 ^ n15958 ^ n9925 ;
  assign n31333 = ~n17671 & n28111 ;
  assign n31334 = n6074 & n31333 ;
  assign n31336 = n31335 ^ n31334 ^ n10256 ;
  assign n31337 = ( n3005 & n4739 ) | ( n3005 & ~n5287 ) | ( n4739 & ~n5287 ) ;
  assign n31338 = ( n5639 & ~n11339 ) | ( n5639 & n31337 ) | ( ~n11339 & n31337 ) ;
  assign n31339 = n31338 ^ n27531 ^ 1'b0 ;
  assign n31340 = n31339 ^ n5912 ^ n1713 ;
  assign n31341 = n26303 ^ n9727 ^ n2823 ;
  assign n31342 = n10535 ^ n10102 ^ 1'b0 ;
  assign n31343 = n31342 ^ n12156 ^ n8146 ;
  assign n31344 = n10060 & n11657 ;
  assign n31345 = n31344 ^ n4101 ^ 1'b0 ;
  assign n31346 = ( n25718 & ~n26993 ) | ( n25718 & n31345 ) | ( ~n26993 & n31345 ) ;
  assign n31347 = n5307 ^ n4879 ^ n789 ;
  assign n31348 = n31347 ^ n378 ^ 1'b0 ;
  assign n31349 = ~n27011 & n31348 ;
  assign n31350 = n5524 & n9327 ;
  assign n31351 = n31350 ^ n12969 ^ 1'b0 ;
  assign n31352 = n22712 ^ n5276 ^ n4761 ;
  assign n31353 = n4492 ^ n2923 ^ n1451 ;
  assign n31354 = ( n1474 & ~n27467 ) | ( n1474 & n31353 ) | ( ~n27467 & n31353 ) ;
  assign n31355 = ( n3515 & n10554 ) | ( n3515 & n31354 ) | ( n10554 & n31354 ) ;
  assign n31358 = ( n2302 & n3593 ) | ( n2302 & n7710 ) | ( n3593 & n7710 ) ;
  assign n31356 = ( n3396 & n9907 ) | ( n3396 & ~n20091 ) | ( n9907 & ~n20091 ) ;
  assign n31357 = n31356 ^ n23874 ^ n1961 ;
  assign n31359 = n31358 ^ n31357 ^ n3511 ;
  assign n31360 = n11737 & n15324 ;
  assign n31361 = n31359 & n31360 ;
  assign n31362 = ( n4538 & n16962 ) | ( n4538 & ~n31361 ) | ( n16962 & ~n31361 ) ;
  assign n31363 = ( n2043 & n18097 ) | ( n2043 & n22624 ) | ( n18097 & n22624 ) ;
  assign n31364 = n6550 ^ n349 ^ 1'b0 ;
  assign n31365 = ( n370 & n6380 ) | ( n370 & n14547 ) | ( n6380 & n14547 ) ;
  assign n31366 = n31365 ^ n24683 ^ n10856 ;
  assign n31367 = ( n1682 & n4543 ) | ( n1682 & ~n6711 ) | ( n4543 & ~n6711 ) ;
  assign n31371 = n10588 | n15377 ;
  assign n31372 = n13219 & ~n31371 ;
  assign n31368 = n20233 ^ n3947 ^ 1'b0 ;
  assign n31369 = n17026 & n31368 ;
  assign n31370 = ( n14226 & n31150 ) | ( n14226 & n31369 ) | ( n31150 & n31369 ) ;
  assign n31373 = n31372 ^ n31370 ^ 1'b0 ;
  assign n31374 = n11947 ^ n9665 ^ n8574 ;
  assign n31375 = ( ~n1887 & n25867 ) | ( ~n1887 & n31374 ) | ( n25867 & n31374 ) ;
  assign n31376 = n4518 & n31375 ;
  assign n31377 = n31376 ^ n957 ^ 1'b0 ;
  assign n31378 = n8690 & ~n25583 ;
  assign n31379 = n9237 & n31378 ;
  assign n31380 = ~n5433 & n19041 ;
  assign n31382 = ( n3950 & n5275 ) | ( n3950 & ~n22194 ) | ( n5275 & ~n22194 ) ;
  assign n31381 = ~n2519 & n19181 ;
  assign n31383 = n31382 ^ n31381 ^ 1'b0 ;
  assign n31384 = n5115 ^ n3129 ^ n341 ;
  assign n31385 = ( n1972 & n31383 ) | ( n1972 & ~n31384 ) | ( n31383 & ~n31384 ) ;
  assign n31386 = x11 | n4108 ;
  assign n31387 = ( n587 & n29205 ) | ( n587 & ~n31386 ) | ( n29205 & ~n31386 ) ;
  assign n31388 = n17134 ^ n12306 ^ n10318 ;
  assign n31389 = ( n2069 & ~n5285 ) | ( n2069 & n5367 ) | ( ~n5285 & n5367 ) ;
  assign n31390 = n29070 ^ n17309 ^ n14601 ;
  assign n31391 = n306 & ~n5566 ;
  assign n31392 = ( n6823 & n14997 ) | ( n6823 & ~n31391 ) | ( n14997 & ~n31391 ) ;
  assign n31393 = n14874 ^ n2360 ^ 1'b0 ;
  assign n31394 = n31393 ^ n12102 ^ n10590 ;
  assign n31395 = n12521 & ~n31394 ;
  assign n31396 = n30029 & n31395 ;
  assign n31397 = ~n7909 & n28358 ;
  assign n31399 = ( n7746 & ~n12619 ) | ( n7746 & n13804 ) | ( ~n12619 & n13804 ) ;
  assign n31398 = n8096 & n16617 ;
  assign n31400 = n31399 ^ n31398 ^ 1'b0 ;
  assign n31401 = n29476 ^ n26193 ^ n14957 ;
  assign n31402 = n31401 ^ n25910 ^ n11899 ;
  assign n31403 = ( n1498 & n6280 ) | ( n1498 & n22954 ) | ( n6280 & n22954 ) ;
  assign n31404 = n15401 ^ n6528 ^ 1'b0 ;
  assign n31405 = n31404 ^ n17900 ^ n5996 ;
  assign n31406 = n1050 | n16495 ;
  assign n31407 = n31406 ^ n17238 ^ 1'b0 ;
  assign n31408 = n29464 ^ n21651 ^ n4650 ;
  assign n31409 = n20172 | n26479 ;
  assign n31410 = n31409 ^ n4012 ^ 1'b0 ;
  assign n31411 = n31410 ^ n23989 ^ n12419 ;
  assign n31412 = n19795 ^ n12190 ^ n909 ;
  assign n31413 = ~n1699 & n3053 ;
  assign n31414 = ~n30257 & n31413 ;
  assign n31415 = n5306 & n10799 ;
  assign n31416 = n31415 ^ n8140 ^ 1'b0 ;
  assign n31417 = ( n5987 & ~n7072 ) | ( n5987 & n21335 ) | ( ~n7072 & n21335 ) ;
  assign n31418 = n4868 | n12727 ;
  assign n31419 = n31417 & ~n31418 ;
  assign n31422 = ( n6308 & n16873 ) | ( n6308 & n18632 ) | ( n16873 & n18632 ) ;
  assign n31420 = n5863 | n6433 ;
  assign n31421 = n7780 | n31420 ;
  assign n31423 = n31422 ^ n31421 ^ n24631 ;
  assign n31424 = n6164 & n31423 ;
  assign n31425 = n5523 | n19705 ;
  assign n31426 = n17535 | n31425 ;
  assign n31427 = n12621 & ~n13425 ;
  assign n31428 = ~n16954 & n31427 ;
  assign n31429 = n31428 ^ n19617 ^ 1'b0 ;
  assign n31430 = ( n379 & n31426 ) | ( n379 & ~n31429 ) | ( n31426 & ~n31429 ) ;
  assign n31431 = n20032 ^ n11618 ^ 1'b0 ;
  assign n31432 = n13769 ^ n4444 ^ n1769 ;
  assign n31433 = n31432 ^ n26247 ^ n13740 ;
  assign n31434 = n4287 ^ n3711 ^ 1'b0 ;
  assign n31435 = ( ~n2785 & n9062 ) | ( ~n2785 & n23133 ) | ( n9062 & n23133 ) ;
  assign n31439 = n18938 ^ n8738 ^ 1'b0 ;
  assign n31440 = ~n15444 & n31439 ;
  assign n31441 = n31440 ^ n14296 ^ n13315 ;
  assign n31442 = n23866 & ~n31441 ;
  assign n31436 = ( n8981 & ~n10400 ) | ( n8981 & n20114 ) | ( ~n10400 & n20114 ) ;
  assign n31437 = ( n14150 & n27518 ) | ( n14150 & ~n31436 ) | ( n27518 & ~n31436 ) ;
  assign n31438 = n31437 ^ n10916 ^ 1'b0 ;
  assign n31443 = n31442 ^ n31438 ^ 1'b0 ;
  assign n31444 = n9641 | n29165 ;
  assign n31445 = ~n1203 & n7974 ;
  assign n31446 = ~n313 & n31445 ;
  assign n31447 = n3083 | n31446 ;
  assign n31448 = n22780 ^ n21597 ^ n5419 ;
  assign n31449 = n13725 ^ n407 ^ 1'b0 ;
  assign n31450 = n31448 & ~n31449 ;
  assign n31451 = n20426 ^ n5409 ^ 1'b0 ;
  assign n31452 = n21353 & ~n31451 ;
  assign n31453 = n27169 ^ n15255 ^ n538 ;
  assign n31454 = n21519 ^ n3352 ^ n2457 ;
  assign n31455 = ~n18591 & n24100 ;
  assign n31457 = n28434 ^ n7346 ^ 1'b0 ;
  assign n31458 = n24306 & n31457 ;
  assign n31456 = n15300 ^ n10025 ^ n7384 ;
  assign n31459 = n31458 ^ n31456 ^ n11219 ;
  assign n31460 = n28006 ^ n20990 ^ n552 ;
  assign n31461 = n2575 | n3839 ;
  assign n31462 = n31227 ^ n10656 ^ 1'b0 ;
  assign n31463 = n31462 ^ n7819 ^ n7638 ;
  assign n31464 = ( ~n31460 & n31461 ) | ( ~n31460 & n31463 ) | ( n31461 & n31463 ) ;
  assign n31465 = n31464 ^ n27762 ^ n22162 ;
  assign n31466 = n10341 ^ n6132 ^ 1'b0 ;
  assign n31467 = n31466 ^ n14545 ^ n666 ;
  assign n31468 = n3486 | n29693 ;
  assign n31469 = n31468 ^ n6602 ^ 1'b0 ;
  assign n31470 = ( n7083 & n10498 ) | ( n7083 & n31469 ) | ( n10498 & n31469 ) ;
  assign n31471 = ~n18113 & n19977 ;
  assign n31472 = ~n12800 & n31471 ;
  assign n31475 = ( ~n10898 & n12694 ) | ( ~n10898 & n21793 ) | ( n12694 & n21793 ) ;
  assign n31473 = ( ~n135 & n4719 ) | ( ~n135 & n22678 ) | ( n4719 & n22678 ) ;
  assign n31474 = ~n11104 & n31473 ;
  assign n31476 = n31475 ^ n31474 ^ 1'b0 ;
  assign n31477 = n26965 ^ n17082 ^ n16149 ;
  assign n31478 = ~n23970 & n31477 ;
  assign n31479 = n26601 ^ n5998 ^ n4111 ;
  assign n31480 = n31479 ^ n25324 ^ n14254 ;
  assign n31482 = n21441 ^ n2805 ^ 1'b0 ;
  assign n31483 = n27092 & ~n31482 ;
  assign n31481 = n7523 ^ n6207 ^ n3322 ;
  assign n31484 = n31483 ^ n31481 ^ n26797 ;
  assign n31485 = n31105 ^ n20474 ^ n18182 ;
  assign n31486 = n31485 ^ n19362 ^ n3045 ;
  assign n31487 = n14024 ^ n5848 ^ 1'b0 ;
  assign n31488 = n15949 & ~n31487 ;
  assign n31489 = ( n6655 & ~n16521 ) | ( n6655 & n31488 ) | ( ~n16521 & n31488 ) ;
  assign n31490 = n25077 ^ n20110 ^ n1644 ;
  assign n31491 = n14706 | n15752 ;
  assign n31492 = n2747 ^ n1794 ^ x22 ;
  assign n31493 = n14191 ^ n9856 ^ n7992 ;
  assign n31494 = n6509 ^ n4779 ^ n619 ;
  assign n31495 = ( ~n23897 & n31493 ) | ( ~n23897 & n31494 ) | ( n31493 & n31494 ) ;
  assign n31496 = ( n7595 & n31492 ) | ( n7595 & ~n31495 ) | ( n31492 & ~n31495 ) ;
  assign n31497 = ( n10888 & n11899 ) | ( n10888 & ~n24191 ) | ( n11899 & ~n24191 ) ;
  assign n31498 = n31497 ^ n13818 ^ 1'b0 ;
  assign n31499 = ( n3409 & n5423 ) | ( n3409 & n9524 ) | ( n5423 & n9524 ) ;
  assign n31500 = n31499 ^ n2507 ^ 1'b0 ;
  assign n31501 = n1828 & n5079 ;
  assign n31502 = n12750 & n31501 ;
  assign n31503 = ( n25833 & n28673 ) | ( n25833 & ~n31502 ) | ( n28673 & ~n31502 ) ;
  assign n31504 = n10309 ^ n9886 ^ n2058 ;
  assign n31505 = n14847 ^ n7360 ^ n4899 ;
  assign n31506 = ( n5487 & n11110 ) | ( n5487 & n31505 ) | ( n11110 & n31505 ) ;
  assign n31507 = n15062 ^ n11850 ^ 1'b0 ;
  assign n31508 = n8777 & ~n11322 ;
  assign n31509 = ~n2514 & n8728 ;
  assign n31510 = n31509 ^ n25771 ^ 1'b0 ;
  assign n31511 = n1725 | n15786 ;
  assign n31512 = n31511 ^ n7029 ^ 1'b0 ;
  assign n31513 = n10456 ^ n8293 ^ 1'b0 ;
  assign n31514 = n16308 | n31513 ;
  assign n31515 = ~n12409 & n31514 ;
  assign n31518 = n26661 ^ n7779 ^ n3084 ;
  assign n31519 = ( n6916 & n9289 ) | ( n6916 & n31518 ) | ( n9289 & n31518 ) ;
  assign n31516 = ( n799 & n6299 ) | ( n799 & n8530 ) | ( n6299 & n8530 ) ;
  assign n31517 = n31516 ^ n22120 ^ 1'b0 ;
  assign n31520 = n31519 ^ n31517 ^ n18242 ;
  assign n31521 = ( n25679 & n29599 ) | ( n25679 & n31520 ) | ( n29599 & n31520 ) ;
  assign n31522 = n26330 | n31521 ;
  assign n31523 = n31515 & ~n31522 ;
  assign n31524 = ( ~x11 & x32 ) | ( ~x11 & n291 ) | ( x32 & n291 ) ;
  assign n31525 = ~n255 & n555 ;
  assign n31526 = n31525 ^ n11355 ^ 1'b0 ;
  assign n31527 = n14841 ^ n4945 ^ 1'b0 ;
  assign n31528 = ~n542 & n31527 ;
  assign n31529 = ~n10716 & n31528 ;
  assign n31530 = n31526 & n31529 ;
  assign n31531 = ( ~n23704 & n29356 ) | ( ~n23704 & n31530 ) | ( n29356 & n31530 ) ;
  assign n31532 = n29475 ^ n27052 ^ n19653 ;
  assign n31533 = n26075 ^ n25599 ^ n4728 ;
  assign n31534 = n21116 ^ n19976 ^ n4227 ;
  assign n31535 = n11222 ^ n3267 ^ 1'b0 ;
  assign n31536 = n13773 & n26408 ;
  assign n31537 = ( ~n1545 & n5452 ) | ( ~n1545 & n16905 ) | ( n5452 & n16905 ) ;
  assign n31538 = n31537 ^ n20195 ^ 1'b0 ;
  assign n31539 = n15707 & ~n31538 ;
  assign n31540 = n6015 ^ n2192 ^ 1'b0 ;
  assign n31541 = n4132 & ~n31540 ;
  assign n31546 = n1253 & n5312 ;
  assign n31547 = n31546 ^ n23826 ^ 1'b0 ;
  assign n31542 = n1557 | n6214 ;
  assign n31543 = n31542 ^ n23713 ^ 1'b0 ;
  assign n31544 = n31543 ^ n13344 ^ n5680 ;
  assign n31545 = n31544 ^ n13478 ^ n8702 ;
  assign n31548 = n31547 ^ n31545 ^ 1'b0 ;
  assign n31549 = n31548 ^ n5351 ^ 1'b0 ;
  assign n31550 = n31541 & ~n31549 ;
  assign n31551 = n5016 ^ n1744 ^ 1'b0 ;
  assign n31552 = n2388 | n12551 ;
  assign n31553 = ~n6541 & n31552 ;
  assign n31554 = n31551 & n31553 ;
  assign n31556 = n1880 & ~n8828 ;
  assign n31555 = n3224 & ~n15625 ;
  assign n31557 = n31556 ^ n31555 ^ 1'b0 ;
  assign n31558 = ( n4378 & n25713 ) | ( n4378 & ~n31557 ) | ( n25713 & ~n31557 ) ;
  assign n31559 = ( ~n2600 & n15893 ) | ( ~n2600 & n27609 ) | ( n15893 & n27609 ) ;
  assign n31560 = n25242 & n31559 ;
  assign n31561 = n27600 ^ n14388 ^ n5717 ;
  assign n31562 = n21478 ^ n8177 ^ n6257 ;
  assign n31563 = n11815 ^ n5750 ^ n4083 ;
  assign n31564 = n31563 ^ n15664 ^ n5433 ;
  assign n31565 = n10899 ^ n6639 ^ n4598 ;
  assign n31566 = n31565 ^ n30766 ^ n6143 ;
  assign n31567 = n14389 ^ n3615 ^ 1'b0 ;
  assign n31568 = n7874 & ~n7975 ;
  assign n31569 = n31568 ^ n27665 ^ 1'b0 ;
  assign n31570 = ~n966 & n3501 ;
  assign n31574 = n7716 & ~n17527 ;
  assign n31575 = ~n11433 & n31574 ;
  assign n31576 = n16467 | n31575 ;
  assign n31571 = n702 & n2379 ;
  assign n31572 = n11280 & n31571 ;
  assign n31573 = n1669 & ~n31572 ;
  assign n31577 = n31576 ^ n31573 ^ 1'b0 ;
  assign n31578 = n21528 | n26087 ;
  assign n31579 = n31578 ^ n686 ^ 1'b0 ;
  assign n31580 = n23353 ^ n11764 ^ 1'b0 ;
  assign n31581 = ( n7988 & n12566 ) | ( n7988 & ~n23592 ) | ( n12566 & ~n23592 ) ;
  assign n31582 = n18599 ^ n2970 ^ 1'b0 ;
  assign n31583 = n19881 ^ n12878 ^ n2921 ;
  assign n31584 = ( n31581 & n31582 ) | ( n31581 & ~n31583 ) | ( n31582 & ~n31583 ) ;
  assign n31585 = ~n31580 & n31584 ;
  assign n31586 = n3805 & n27377 ;
  assign n31589 = n19258 ^ n8655 ^ n3187 ;
  assign n31587 = n22778 | n23947 ;
  assign n31588 = n31587 ^ n25860 ^ 1'b0 ;
  assign n31590 = n31589 ^ n31588 ^ n8253 ;
  assign n31591 = ( n2228 & n2372 ) | ( n2228 & ~n5306 ) | ( n2372 & ~n5306 ) ;
  assign n31592 = n31591 ^ n18934 ^ n10390 ;
  assign n31593 = n10460 ^ n10136 ^ n8509 ;
  assign n31594 = n31593 ^ n22888 ^ n493 ;
  assign n31595 = n18511 ^ n5123 ^ n2712 ;
  assign n31596 = ( n8913 & n23011 ) | ( n8913 & ~n29354 ) | ( n23011 & ~n29354 ) ;
  assign n31597 = ( n14927 & ~n28331 ) | ( n14927 & n31596 ) | ( ~n28331 & n31596 ) ;
  assign n31598 = n846 | n28396 ;
  assign n31599 = n31598 ^ n13759 ^ 1'b0 ;
  assign n31605 = ( n4980 & n13190 ) | ( n4980 & n18251 ) | ( n13190 & n18251 ) ;
  assign n31600 = n5639 | n7425 ;
  assign n31601 = n3461 & ~n31600 ;
  assign n31602 = n13982 ^ n11041 ^ n3849 ;
  assign n31603 = ( n21437 & n31601 ) | ( n21437 & n31602 ) | ( n31601 & n31602 ) ;
  assign n31604 = ~n7932 & n31603 ;
  assign n31606 = n31605 ^ n31604 ^ 1'b0 ;
  assign n31607 = n27223 ^ n21349 ^ n3080 ;
  assign n31608 = n2725 & n26284 ;
  assign n31609 = n31607 & n31608 ;
  assign n31610 = n18176 & ~n23544 ;
  assign n31611 = n31610 ^ n293 ^ 1'b0 ;
  assign n31612 = n12298 ^ n4417 ^ 1'b0 ;
  assign n31613 = ( n3533 & n25146 ) | ( n3533 & n25540 ) | ( n25146 & n25540 ) ;
  assign n31614 = n23522 ^ n2410 ^ 1'b0 ;
  assign n31615 = n20499 ^ n10769 ^ 1'b0 ;
  assign n31616 = n31615 ^ n23475 ^ n13371 ;
  assign n31617 = ( n1584 & n16654 ) | ( n1584 & ~n23419 ) | ( n16654 & ~n23419 ) ;
  assign n31618 = n31518 ^ n9471 ^ n7582 ;
  assign n31619 = n19523 ^ n17868 ^ n17651 ;
  assign n31620 = ( n14220 & n31618 ) | ( n14220 & n31619 ) | ( n31618 & n31619 ) ;
  assign n31621 = n14540 | n24812 ;
  assign n31622 = ( n582 & ~n8139 ) | ( n582 & n13168 ) | ( ~n8139 & n13168 ) ;
  assign n31623 = n17998 & ~n31622 ;
  assign n31624 = n31623 ^ n10329 ^ 1'b0 ;
  assign n31625 = n4129 | n24918 ;
  assign n31626 = n31625 ^ n4708 ^ 1'b0 ;
  assign n31627 = ( n10816 & n11473 ) | ( n10816 & n13585 ) | ( n11473 & n13585 ) ;
  assign n31629 = n1630 ^ n1480 ^ 1'b0 ;
  assign n31630 = ~n4725 & n31629 ;
  assign n31628 = ( n1212 & ~n6352 ) | ( n1212 & n24474 ) | ( ~n6352 & n24474 ) ;
  assign n31631 = n31630 ^ n31628 ^ n11708 ;
  assign n31632 = n4966 | n15623 ;
  assign n31633 = n31632 ^ n14049 ^ n11815 ;
  assign n31634 = n15914 & ~n18063 ;
  assign n31635 = n17767 ^ n3752 ^ 1'b0 ;
  assign n31636 = ~n5918 & n31635 ;
  assign n31637 = n31636 ^ n7891 ^ 1'b0 ;
  assign n31638 = ( ~x101 & n15077 ) | ( ~x101 & n31637 ) | ( n15077 & n31637 ) ;
  assign n31639 = ( n4888 & ~n12990 ) | ( n4888 & n26725 ) | ( ~n12990 & n26725 ) ;
  assign n31640 = ( n2164 & n14227 ) | ( n2164 & ~n20617 ) | ( n14227 & ~n20617 ) ;
  assign n31641 = ( ~n12010 & n31639 ) | ( ~n12010 & n31640 ) | ( n31639 & n31640 ) ;
  assign n31642 = ~n6846 & n7839 ;
  assign n31643 = ( n20015 & ~n23185 ) | ( n20015 & n31642 ) | ( ~n23185 & n31642 ) ;
  assign n31644 = n31643 ^ n20117 ^ n15094 ;
  assign n31645 = ( ~n919 & n13094 ) | ( ~n919 & n31644 ) | ( n13094 & n31644 ) ;
  assign n31647 = n6730 & ~n12831 ;
  assign n31646 = n2953 | n7022 ;
  assign n31648 = n31647 ^ n31646 ^ 1'b0 ;
  assign n31649 = n183 & ~n8216 ;
  assign n31650 = ~n19241 & n31649 ;
  assign n31651 = n8327 | n14263 ;
  assign n31652 = n31651 ^ n12219 ^ 1'b0 ;
  assign n31653 = ~n3552 & n15378 ;
  assign n31654 = n31653 ^ n21718 ^ 1'b0 ;
  assign n31655 = ~n26909 & n31654 ;
  assign n31656 = ( n2136 & n6893 ) | ( n2136 & n10002 ) | ( n6893 & n10002 ) ;
  assign n31657 = n29303 ^ n3900 ^ 1'b0 ;
  assign n31658 = n15191 & n31657 ;
  assign n31659 = n10861 ^ n289 ^ 1'b0 ;
  assign n31660 = n31658 & n31659 ;
  assign n31661 = ( n222 & ~n8663 ) | ( n222 & n31660 ) | ( ~n8663 & n31660 ) ;
  assign n31662 = n28483 ^ n19179 ^ n19005 ;
  assign n31663 = n31662 ^ n16757 ^ 1'b0 ;
  assign n31664 = n31663 ^ n27044 ^ n17316 ;
  assign n31665 = n25798 ^ n9758 ^ n2694 ;
  assign n31666 = n20078 ^ n17142 ^ n4965 ;
  assign n31667 = ~n1059 & n19945 ;
  assign n31668 = ( n4685 & n5894 ) | ( n4685 & ~n17063 ) | ( n5894 & ~n17063 ) ;
  assign n31669 = ( n7136 & n15663 ) | ( n7136 & ~n31668 ) | ( n15663 & ~n31668 ) ;
  assign n31670 = n8474 & ~n27639 ;
  assign n31671 = n31670 ^ n9012 ^ 1'b0 ;
  assign n31672 = ~n6263 & n18669 ;
  assign n31673 = n6128 ^ n733 ^ 1'b0 ;
  assign n31674 = ~n13276 & n31673 ;
  assign n31675 = n23677 ^ n14329 ^ n7788 ;
  assign n31676 = n18484 ^ n16917 ^ n1340 ;
  assign n31677 = n31676 ^ n14966 ^ 1'b0 ;
  assign n31678 = n23378 ^ n19386 ^ n6572 ;
  assign n31679 = n31370 ^ n30017 ^ n3944 ;
  assign n31681 = ( n1645 & n21621 ) | ( n1645 & n22656 ) | ( n21621 & n22656 ) ;
  assign n31680 = n1745 | n11406 ;
  assign n31682 = n31681 ^ n31680 ^ 1'b0 ;
  assign n31683 = n23006 & ~n31682 ;
  assign n31684 = n26482 ^ n19459 ^ n14588 ;
  assign n31685 = ~n2733 & n21755 ;
  assign n31686 = n18862 & n18923 ;
  assign n31687 = ( n26216 & ~n31685 ) | ( n26216 & n31686 ) | ( ~n31685 & n31686 ) ;
  assign n31688 = n30747 ^ n4989 ^ 1'b0 ;
  assign n31690 = n13244 ^ n11756 ^ n9212 ;
  assign n31689 = n12922 & n29517 ;
  assign n31691 = n31690 ^ n31689 ^ 1'b0 ;
  assign n31692 = n2204 & n7664 ;
  assign n31693 = ~n19240 & n31692 ;
  assign n31696 = n15896 ^ n439 ^ 1'b0 ;
  assign n31697 = n8479 & ~n31696 ;
  assign n31694 = ( ~n5083 & n7510 ) | ( ~n5083 & n8362 ) | ( n7510 & n8362 ) ;
  assign n31695 = n31694 ^ n21554 ^ n14184 ;
  assign n31698 = n31697 ^ n31695 ^ n19938 ;
  assign n31699 = ( n4499 & n11235 ) | ( n4499 & n21893 ) | ( n11235 & n21893 ) ;
  assign n31700 = ( n5394 & n12343 ) | ( n5394 & ~n31699 ) | ( n12343 & ~n31699 ) ;
  assign n31701 = ( x121 & ~n7867 ) | ( x121 & n8972 ) | ( ~n7867 & n8972 ) ;
  assign n31702 = ( ~n7171 & n7404 ) | ( ~n7171 & n31701 ) | ( n7404 & n31701 ) ;
  assign n31703 = ~n11530 & n16136 ;
  assign n31704 = n7097 & ~n28187 ;
  assign n31705 = n11714 & n31704 ;
  assign n31706 = ~n3843 & n4116 ;
  assign n31707 = n7767 & n31706 ;
  assign n31708 = ( n4285 & ~n31705 ) | ( n4285 & n31707 ) | ( ~n31705 & n31707 ) ;
  assign n31709 = n14699 & n23808 ;
  assign n31710 = ( n3192 & n3685 ) | ( n3192 & ~n14450 ) | ( n3685 & ~n14450 ) ;
  assign n31711 = n31710 ^ n23993 ^ n23761 ;
  assign n31712 = n27470 ^ n23409 ^ n12138 ;
  assign n31713 = n5313 & n17170 ;
  assign n31714 = n31713 ^ n16033 ^ 1'b0 ;
  assign n31715 = n16527 ^ n8451 ^ 1'b0 ;
  assign n31716 = ( n4797 & n6321 ) | ( n4797 & n19074 ) | ( n6321 & n19074 ) ;
  assign n31717 = n31716 ^ n23771 ^ 1'b0 ;
  assign n31718 = n23181 ^ n11028 ^ n2168 ;
  assign n31720 = ( n3692 & n24423 ) | ( n3692 & ~n28372 ) | ( n24423 & ~n28372 ) ;
  assign n31721 = ( ~n18337 & n23310 ) | ( ~n18337 & n31720 ) | ( n23310 & n31720 ) ;
  assign n31719 = n3653 & ~n29383 ;
  assign n31722 = n31721 ^ n31719 ^ 1'b0 ;
  assign n31723 = ( n15568 & n31718 ) | ( n15568 & ~n31722 ) | ( n31718 & ~n31722 ) ;
  assign n31724 = n7408 ^ n2230 ^ n457 ;
  assign n31725 = ( n3321 & ~n24122 ) | ( n3321 & n31724 ) | ( ~n24122 & n31724 ) ;
  assign n31726 = n5758 ^ n666 ^ 1'b0 ;
  assign n31727 = ~n5369 & n31726 ;
  assign n31728 = n15532 ^ n7860 ^ 1'b0 ;
  assign n31729 = n31727 & n31728 ;
  assign n31730 = n31729 ^ n25244 ^ n9354 ;
  assign n31731 = ( ~n971 & n2436 ) | ( ~n971 & n3335 ) | ( n2436 & n3335 ) ;
  assign n31732 = n31731 ^ n27989 ^ n16189 ;
  assign n31733 = n31732 ^ n19522 ^ n3573 ;
  assign n31736 = n18449 ^ n4570 ^ 1'b0 ;
  assign n31737 = n31736 ^ n8260 ^ n5060 ;
  assign n31734 = ~n8923 & n26910 ;
  assign n31735 = ~n21271 & n31734 ;
  assign n31738 = n31737 ^ n31735 ^ n2292 ;
  assign n31739 = n27594 ^ n21301 ^ x25 ;
  assign n31742 = ( n14656 & n25775 ) | ( n14656 & ~n29954 ) | ( n25775 & ~n29954 ) ;
  assign n31740 = n3537 & n27446 ;
  assign n31741 = ~n6811 & n31740 ;
  assign n31743 = n31742 ^ n31741 ^ 1'b0 ;
  assign n31744 = n5480 | n27242 ;
  assign n31745 = n31744 ^ n17340 ^ 1'b0 ;
  assign n31748 = n10702 ^ n4433 ^ n2117 ;
  assign n31746 = n11111 ^ n4428 ^ 1'b0 ;
  assign n31747 = n9233 & ~n31746 ;
  assign n31749 = n31748 ^ n31747 ^ n20294 ;
  assign n31750 = ( n12324 & ~n29792 ) | ( n12324 & n31749 ) | ( ~n29792 & n31749 ) ;
  assign n31751 = ( ~n1576 & n16880 ) | ( ~n1576 & n18054 ) | ( n16880 & n18054 ) ;
  assign n31752 = n14340 | n28243 ;
  assign n31753 = n17045 & ~n31752 ;
  assign n31754 = n29234 & ~n31753 ;
  assign n31755 = n13243 & n31754 ;
  assign n31756 = ( n11100 & ~n26964 ) | ( n11100 & n31755 ) | ( ~n26964 & n31755 ) ;
  assign n31757 = ~n15947 & n25845 ;
  assign n31758 = n14754 ^ n9053 ^ n5611 ;
  assign n31759 = ~n931 & n6963 ;
  assign n31760 = n31759 ^ n12015 ^ 1'b0 ;
  assign n31761 = ( ~n6497 & n24135 ) | ( ~n6497 & n31760 ) | ( n24135 & n31760 ) ;
  assign n31762 = n830 & ~n12618 ;
  assign n31763 = n21282 ^ n13954 ^ 1'b0 ;
  assign n31764 = ~n18398 & n31763 ;
  assign n31765 = n13660 & n29118 ;
  assign n31766 = n6912 & ~n8338 ;
  assign n31767 = n18745 ^ n12675 ^ n1606 ;
  assign n31769 = n7199 ^ n4302 ^ x70 ;
  assign n31768 = ( n1361 & ~n8591 ) | ( n1361 & n22239 ) | ( ~n8591 & n22239 ) ;
  assign n31770 = n31769 ^ n31768 ^ n10231 ;
  assign n31771 = ( n12490 & n13929 ) | ( n12490 & ~n31770 ) | ( n13929 & ~n31770 ) ;
  assign n31772 = ( n12144 & n17238 ) | ( n12144 & ~n27393 ) | ( n17238 & ~n27393 ) ;
  assign n31773 = n9229 & n31772 ;
  assign n31774 = ~n5434 & n14812 ;
  assign n31775 = ~n1606 & n31774 ;
  assign n31776 = ( n4786 & n31773 ) | ( n4786 & ~n31775 ) | ( n31773 & ~n31775 ) ;
  assign n31777 = n825 | n25486 ;
  assign n31778 = n1652 | n31777 ;
  assign n31779 = n31778 ^ n20520 ^ 1'b0 ;
  assign n31780 = n12360 & ~n31779 ;
  assign n31781 = ( n4742 & n11777 ) | ( n4742 & n31780 ) | ( n11777 & n31780 ) ;
  assign n31782 = ( n6928 & ~n15633 ) | ( n6928 & n26754 ) | ( ~n15633 & n26754 ) ;
  assign n31783 = n14697 ^ n13497 ^ 1'b0 ;
  assign n31784 = n31782 & n31783 ;
  assign n31785 = n31784 ^ n25950 ^ 1'b0 ;
  assign n31786 = ( n2948 & n6309 ) | ( n2948 & n20434 ) | ( n6309 & n20434 ) ;
  assign n31787 = n8898 ^ n6078 ^ n591 ;
  assign n31788 = n10424 | n31787 ;
  assign n31789 = n31788 ^ n16780 ^ n8445 ;
  assign n31790 = n31789 ^ n9057 ^ n7563 ;
  assign n31791 = n8136 ^ n7064 ^ 1'b0 ;
  assign n31792 = ~n9633 & n14581 ;
  assign n31793 = ~n29651 & n31792 ;
  assign n31794 = n7376 & n15663 ;
  assign n31795 = n8233 & n31794 ;
  assign n31796 = ( n8815 & n17962 ) | ( n8815 & ~n23332 ) | ( n17962 & ~n23332 ) ;
  assign n31797 = ( ~n19672 & n26011 ) | ( ~n19672 & n31796 ) | ( n26011 & n31796 ) ;
  assign n31798 = n11574 ^ n1630 ^ n1326 ;
  assign n31799 = n31798 ^ n26942 ^ n3651 ;
  assign n31802 = n12011 ^ n10412 ^ n1232 ;
  assign n31801 = n22039 ^ n14973 ^ n12323 ;
  assign n31800 = n2111 ^ n333 ^ 1'b0 ;
  assign n31803 = n31802 ^ n31801 ^ n31800 ;
  assign n31804 = n4600 ^ x62 ^ 1'b0 ;
  assign n31805 = ( n11378 & ~n13358 ) | ( n11378 & n31804 ) | ( ~n13358 & n31804 ) ;
  assign n31806 = n10183 & ~n13144 ;
  assign n31807 = ( n4090 & n8363 ) | ( n4090 & n17618 ) | ( n8363 & n17618 ) ;
  assign n31808 = ( ~x91 & n31806 ) | ( ~x91 & n31807 ) | ( n31806 & n31807 ) ;
  assign n31809 = n5658 ^ n3951 ^ 1'b0 ;
  assign n31811 = n760 & n7612 ;
  assign n31812 = n31811 ^ n6885 ^ n3296 ;
  assign n31813 = n31812 ^ n13012 ^ n5683 ;
  assign n31814 = n17334 & n31813 ;
  assign n31810 = n16908 & ~n23097 ;
  assign n31815 = n31814 ^ n31810 ^ 1'b0 ;
  assign n31816 = ( ~x82 & n17547 ) | ( ~x82 & n23074 ) | ( n17547 & n23074 ) ;
  assign n31817 = n31816 ^ n2992 ^ 1'b0 ;
  assign n31818 = n30595 & ~n31817 ;
  assign n31819 = ~n3946 & n16535 ;
  assign n31820 = n19702 ^ n16053 ^ 1'b0 ;
  assign n31821 = n31819 | n31820 ;
  assign n31822 = ( n5052 & ~n28035 ) | ( n5052 & n30600 ) | ( ~n28035 & n30600 ) ;
  assign n31823 = n9925 ^ n7515 ^ n378 ;
  assign n31824 = ( n7894 & n21556 ) | ( n7894 & ~n31823 ) | ( n21556 & ~n31823 ) ;
  assign n31825 = n31824 ^ n21788 ^ n1459 ;
  assign n31826 = n21946 ^ n20882 ^ 1'b0 ;
  assign n31827 = n14059 & n21048 ;
  assign n31828 = n18022 ^ n15145 ^ n2497 ;
  assign n31829 = n20269 & n23570 ;
  assign n31830 = ( ~n1060 & n8350 ) | ( ~n1060 & n29903 ) | ( n8350 & n29903 ) ;
  assign n31831 = x74 & n6329 ;
  assign n31832 = n31831 ^ n12428 ^ 1'b0 ;
  assign n31833 = ( n15549 & n17548 ) | ( n15549 & ~n23336 ) | ( n17548 & ~n23336 ) ;
  assign n31834 = n31833 ^ n3482 ^ 1'b0 ;
  assign n31835 = n22638 | n26882 ;
  assign n31836 = n31835 ^ n6167 ^ 1'b0 ;
  assign n31837 = n29517 ^ n7911 ^ 1'b0 ;
  assign n31838 = ~n6228 & n23500 ;
  assign n31839 = n31838 ^ n24248 ^ 1'b0 ;
  assign n31840 = n31839 ^ n4366 ^ n499 ;
  assign n31841 = n31807 ^ n5730 ^ n1573 ;
  assign n31842 = n26392 ^ n23301 ^ n2624 ;
  assign n31847 = n20838 ^ n18121 ^ 1'b0 ;
  assign n31843 = n16719 ^ n5740 ^ 1'b0 ;
  assign n31844 = n9672 | n31843 ;
  assign n31845 = n25584 & ~n31844 ;
  assign n31846 = n31845 ^ n25954 ^ n14290 ;
  assign n31848 = n31847 ^ n31846 ^ n8416 ;
  assign n31849 = ( ~n24840 & n31842 ) | ( ~n24840 & n31848 ) | ( n31842 & n31848 ) ;
  assign n31850 = ~n811 & n18603 ;
  assign n31851 = n31850 ^ n2158 ^ n2065 ;
  assign n31852 = n13002 | n31591 ;
  assign n31853 = n31852 ^ n13927 ^ 1'b0 ;
  assign n31854 = n31853 ^ n18289 ^ n2389 ;
  assign n31855 = n5462 | n31854 ;
  assign n31856 = ~n5351 & n24158 ;
  assign n31857 = n8061 & ~n28350 ;
  assign n31858 = n24153 & n31857 ;
  assign n31859 = n4848 ^ n4757 ^ n1772 ;
  assign n31860 = n23164 ^ n7728 ^ 1'b0 ;
  assign n31861 = ~n31859 & n31860 ;
  assign n31862 = n2339 & n6951 ;
  assign n31863 = ~n31861 & n31862 ;
  assign n31864 = n19798 ^ n15959 ^ 1'b0 ;
  assign n31865 = ~n28447 & n31864 ;
  assign n31866 = ~n28576 & n31865 ;
  assign n31867 = n12023 & ~n12393 ;
  assign n31868 = ( n8556 & n11270 ) | ( n8556 & ~n30001 ) | ( n11270 & ~n30001 ) ;
  assign n31869 = n22997 ^ n17930 ^ n14266 ;
  assign n31870 = n31869 ^ n20589 ^ n12602 ;
  assign n31871 = ( n3202 & n9649 ) | ( n3202 & ~n31870 ) | ( n9649 & ~n31870 ) ;
  assign n31872 = ( ~n2247 & n4468 ) | ( ~n2247 & n12792 ) | ( n4468 & n12792 ) ;
  assign n31873 = n31872 ^ n22817 ^ n16059 ;
  assign n31874 = ( n5652 & n12238 ) | ( n5652 & n19342 ) | ( n12238 & n19342 ) ;
  assign n31875 = ( n8366 & n10784 ) | ( n8366 & ~n25695 ) | ( n10784 & ~n25695 ) ;
  assign n31876 = ~n10201 & n22474 ;
  assign n31877 = n31876 ^ n17156 ^ 1'b0 ;
  assign n31878 = ( n1971 & ~n31875 ) | ( n1971 & n31877 ) | ( ~n31875 & n31877 ) ;
  assign n31879 = n31878 ^ n22493 ^ n13908 ;
  assign n31880 = n14936 ^ n13797 ^ n8888 ;
  assign n31881 = n13366 ^ n7820 ^ 1'b0 ;
  assign n31882 = n21249 & ~n31881 ;
  assign n31883 = n27841 ^ n13074 ^ 1'b0 ;
  assign n31884 = n14859 & ~n31883 ;
  assign n31885 = n23317 ^ n7419 ^ 1'b0 ;
  assign n31886 = n3062 & n31885 ;
  assign n31887 = n9191 & n26639 ;
  assign n31888 = n21627 & ~n31887 ;
  assign n31889 = ( n20125 & n22113 ) | ( n20125 & n31888 ) | ( n22113 & n31888 ) ;
  assign n31890 = n8996 ^ n6507 ^ 1'b0 ;
  assign n31891 = ~n31889 & n31890 ;
  assign n31892 = n4284 & n8763 ;
  assign n31893 = ( n583 & n14991 ) | ( n583 & n16714 ) | ( n14991 & n16714 ) ;
  assign n31894 = n15368 & ~n26344 ;
  assign n31895 = ( n7304 & ~n31893 ) | ( n7304 & n31894 ) | ( ~n31893 & n31894 ) ;
  assign n31896 = ( n1671 & n15300 ) | ( n1671 & n30882 ) | ( n15300 & n30882 ) ;
  assign n31897 = ~n6739 & n7342 ;
  assign n31898 = ( n2509 & n7190 ) | ( n2509 & n17161 ) | ( n7190 & n17161 ) ;
  assign n31899 = ( n8466 & n31897 ) | ( n8466 & ~n31898 ) | ( n31897 & ~n31898 ) ;
  assign n31900 = n12101 ^ n6865 ^ n2803 ;
  assign n31901 = n31900 ^ n9392 ^ 1'b0 ;
  assign n31902 = ( ~n3883 & n8330 ) | ( ~n3883 & n31901 ) | ( n8330 & n31901 ) ;
  assign n31903 = ( n7911 & ~n18850 ) | ( n7911 & n31902 ) | ( ~n18850 & n31902 ) ;
  assign n31904 = n25337 ^ n24768 ^ n10441 ;
  assign n31905 = n23735 ^ n13317 ^ n473 ;
  assign n31906 = n11587 | n14849 ;
  assign n31907 = n31906 ^ n28281 ^ 1'b0 ;
  assign n31908 = ( n4259 & n4610 ) | ( n4259 & ~n24554 ) | ( n4610 & ~n24554 ) ;
  assign n31909 = n16359 ^ n661 ^ 1'b0 ;
  assign n31910 = n8105 & n31909 ;
  assign n31911 = n31910 ^ n16939 ^ n9067 ;
  assign n31912 = n22893 ^ n8082 ^ n5638 ;
  assign n31913 = n5553 & n24059 ;
  assign n31914 = ~n12323 & n18590 ;
  assign n31915 = ( ~n31662 & n31913 ) | ( ~n31662 & n31914 ) | ( n31913 & n31914 ) ;
  assign n31916 = ( n2390 & n12238 ) | ( n2390 & n14794 ) | ( n12238 & n14794 ) ;
  assign n31917 = n31916 ^ n29369 ^ 1'b0 ;
  assign n31918 = n5124 & ~n6657 ;
  assign n31919 = n31918 ^ n10178 ^ 1'b0 ;
  assign n31920 = n31919 ^ n14912 ^ n14752 ;
  assign n31921 = n31920 ^ n28234 ^ n20589 ;
  assign n31922 = n4008 ^ n477 ^ 1'b0 ;
  assign n31923 = n6452 | n6681 ;
  assign n31924 = n8065 | n31923 ;
  assign n31925 = ~n2257 & n24798 ;
  assign n31926 = ~n7998 & n31925 ;
  assign n31927 = n31926 ^ n1019 ^ 1'b0 ;
  assign n31928 = ( ~n2488 & n9339 ) | ( ~n2488 & n18677 ) | ( n9339 & n18677 ) ;
  assign n31929 = n31928 ^ n511 ^ 1'b0 ;
  assign n31930 = n31927 & n31929 ;
  assign n31931 = n2306 & n7584 ;
  assign n31932 = n31931 ^ n3954 ^ 1'b0 ;
  assign n31933 = ( n24415 & n25846 ) | ( n24415 & ~n31932 ) | ( n25846 & ~n31932 ) ;
  assign n31934 = ( ~n931 & n7594 ) | ( ~n931 & n23286 ) | ( n7594 & n23286 ) ;
  assign n31935 = ( n31930 & n31933 ) | ( n31930 & ~n31934 ) | ( n31933 & ~n31934 ) ;
  assign n31936 = n19066 ^ n15784 ^ 1'b0 ;
  assign n31937 = n12520 & n31936 ;
  assign n31938 = ( ~n1983 & n14258 ) | ( ~n1983 & n31937 ) | ( n14258 & n31937 ) ;
  assign n31940 = ( n5522 & n7468 ) | ( n5522 & ~n10002 ) | ( n7468 & ~n10002 ) ;
  assign n31939 = n7903 ^ n698 ^ 1'b0 ;
  assign n31941 = n31940 ^ n31939 ^ 1'b0 ;
  assign n31942 = n13035 | n13986 ;
  assign n31943 = n13233 & ~n31942 ;
  assign n31944 = ( n1713 & n8727 ) | ( n1713 & n31943 ) | ( n8727 & n31943 ) ;
  assign n31945 = n6257 ^ n1448 ^ 1'b0 ;
  assign n31946 = ( n4544 & n17007 ) | ( n4544 & ~n31945 ) | ( n17007 & ~n31945 ) ;
  assign n31947 = n15264 ^ n7517 ^ 1'b0 ;
  assign n31948 = n31947 ^ n16775 ^ n3018 ;
  assign n31949 = ( ~n28336 & n31946 ) | ( ~n28336 & n31948 ) | ( n31946 & n31948 ) ;
  assign n31950 = ( n17690 & n30731 ) | ( n17690 & n31949 ) | ( n30731 & n31949 ) ;
  assign n31951 = n25968 ^ n22272 ^ n3947 ;
  assign n31952 = ( n20165 & ~n20864 ) | ( n20165 & n31951 ) | ( ~n20864 & n31951 ) ;
  assign n31953 = n31607 ^ n22287 ^ n19874 ;
  assign n31958 = n1424 & ~n18626 ;
  assign n31959 = ~n23095 & n31958 ;
  assign n31960 = n31959 ^ n20854 ^ n11239 ;
  assign n31961 = n23012 ^ n19939 ^ 1'b0 ;
  assign n31962 = n31960 | n31961 ;
  assign n31954 = ( n8454 & ~n16399 ) | ( n8454 & n17733 ) | ( ~n16399 & n17733 ) ;
  assign n31955 = n31954 ^ n16470 ^ n10858 ;
  assign n31956 = ( n5670 & n30775 ) | ( n5670 & n31955 ) | ( n30775 & n31955 ) ;
  assign n31957 = n4537 | n31956 ;
  assign n31963 = n31962 ^ n31957 ^ 1'b0 ;
  assign n31964 = ( n2935 & ~n3531 ) | ( n2935 & n12380 ) | ( ~n3531 & n12380 ) ;
  assign n31965 = n8199 & n29160 ;
  assign n31966 = ~n31964 & n31965 ;
  assign n31967 = n29911 ^ n18612 ^ 1'b0 ;
  assign n31968 = n9343 & ~n31967 ;
  assign n31969 = n28561 ^ n24599 ^ n3630 ;
  assign n31970 = ( n8755 & n27291 ) | ( n8755 & ~n31969 ) | ( n27291 & ~n31969 ) ;
  assign n31971 = n18025 & n24696 ;
  assign n31972 = n31971 ^ n12763 ^ x93 ;
  assign n31973 = n31972 ^ n26530 ^ n16200 ;
  assign n31974 = n21039 ^ n2773 ^ 1'b0 ;
  assign n31975 = n31974 ^ n28980 ^ n5668 ;
  assign n31976 = ( ~n2785 & n8430 ) | ( ~n2785 & n18415 ) | ( n8430 & n18415 ) ;
  assign n31977 = n31976 ^ n10707 ^ n7296 ;
  assign n31978 = n8821 ^ n3699 ^ 1'b0 ;
  assign n31979 = n22662 | n31978 ;
  assign n31980 = ( ~n4232 & n12377 ) | ( ~n4232 & n31979 ) | ( n12377 & n31979 ) ;
  assign n31981 = n9853 & n31980 ;
  assign n31982 = n31981 ^ n24323 ^ n16098 ;
  assign n31983 = ( n7138 & n9677 ) | ( n7138 & ~n29675 ) | ( n9677 & ~n29675 ) ;
  assign n31984 = n8929 ^ n666 ^ 1'b0 ;
  assign n31985 = n3680 & n31984 ;
  assign n31986 = ( n8679 & n31983 ) | ( n8679 & ~n31985 ) | ( n31983 & ~n31985 ) ;
  assign n31987 = ( x18 & ~n8215 ) | ( x18 & n31986 ) | ( ~n8215 & n31986 ) ;
  assign n31988 = n27620 ^ n14710 ^ 1'b0 ;
  assign n31989 = n20078 | n31988 ;
  assign n31990 = n10555 ^ n9934 ^ n3773 ;
  assign n31991 = n31990 ^ n10395 ^ 1'b0 ;
  assign n31992 = n16936 & n31991 ;
  assign n31993 = n29652 ^ n6445 ^ 1'b0 ;
  assign n31994 = ~n1090 & n1853 ;
  assign n31995 = n31994 ^ n16904 ^ n1236 ;
  assign n31996 = n20253 ^ n14080 ^ 1'b0 ;
  assign n31997 = ~n2173 & n31996 ;
  assign n31998 = ( n6568 & n31372 ) | ( n6568 & ~n31997 ) | ( n31372 & ~n31997 ) ;
  assign n31999 = ( n15919 & n22194 ) | ( n15919 & n31998 ) | ( n22194 & n31998 ) ;
  assign n32000 = ~n19436 & n20118 ;
  assign n32001 = n32000 ^ n21490 ^ 1'b0 ;
  assign n32002 = n15426 ^ n6887 ^ n4476 ;
  assign n32004 = ( x64 & n9722 ) | ( x64 & n25907 ) | ( n9722 & n25907 ) ;
  assign n32003 = n22066 ^ n13627 ^ n8695 ;
  assign n32005 = n32004 ^ n32003 ^ 1'b0 ;
  assign n32006 = ( ~n9993 & n32002 ) | ( ~n9993 & n32005 ) | ( n32002 & n32005 ) ;
  assign n32007 = n28895 ^ n259 ^ 1'b0 ;
  assign n32008 = ( ~n15250 & n15735 ) | ( ~n15250 & n22466 ) | ( n15735 & n22466 ) ;
  assign n32009 = ( n5106 & n5805 ) | ( n5106 & ~n24453 ) | ( n5805 & ~n24453 ) ;
  assign n32010 = n32009 ^ n25032 ^ n12829 ;
  assign n32011 = n12101 ^ n9001 ^ n3126 ;
  assign n32012 = n32011 ^ n11193 ^ 1'b0 ;
  assign n32013 = ~n32010 & n32012 ;
  assign n32014 = n1667 & n32013 ;
  assign n32015 = ~n20072 & n32014 ;
  assign n32016 = n7238 & ~n17704 ;
  assign n32017 = ( n9797 & n19758 ) | ( n9797 & ~n32016 ) | ( n19758 & ~n32016 ) ;
  assign n32018 = ( n11739 & n12627 ) | ( n11739 & ~n13870 ) | ( n12627 & ~n13870 ) ;
  assign n32019 = ( n27906 & n32017 ) | ( n27906 & n32018 ) | ( n32017 & n32018 ) ;
  assign n32020 = n4015 | n32019 ;
  assign n32021 = n32020 ^ n14584 ^ 1'b0 ;
  assign n32022 = ~n13328 & n13756 ;
  assign n32023 = n32022 ^ n25244 ^ 1'b0 ;
  assign n32024 = n14294 ^ n11856 ^ 1'b0 ;
  assign n32025 = n30789 ^ n19483 ^ 1'b0 ;
  assign n32026 = ( x51 & n14885 ) | ( x51 & ~n22716 ) | ( n14885 & ~n22716 ) ;
  assign n32027 = ( n12010 & n18493 ) | ( n12010 & n32026 ) | ( n18493 & n32026 ) ;
  assign n32028 = n28672 ^ n20735 ^ 1'b0 ;
  assign n32029 = n31565 ^ n18594 ^ 1'b0 ;
  assign n32030 = ( ~n841 & n21460 ) | ( ~n841 & n32029 ) | ( n21460 & n32029 ) ;
  assign n32031 = n32030 ^ n30119 ^ n24239 ;
  assign n32032 = n21722 ^ n6521 ^ 1'b0 ;
  assign n32033 = n14640 ^ n13878 ^ 1'b0 ;
  assign n32034 = ~n19098 & n23416 ;
  assign n32035 = ~n32033 & n32034 ;
  assign n32036 = n7949 & n23081 ;
  assign n32037 = n32036 ^ n8746 ^ 1'b0 ;
  assign n32038 = n4922 & n31620 ;
  assign n32039 = n1919 & n32038 ;
  assign n32040 = ~n3667 & n10792 ;
  assign n32041 = ~x89 & n32040 ;
  assign n32042 = ( n5068 & ~n22902 ) | ( n5068 & n27358 ) | ( ~n22902 & n27358 ) ;
  assign n32043 = n14209 ^ n13217 ^ n9449 ;
  assign n32044 = n32043 ^ n26849 ^ n9302 ;
  assign n32045 = n30437 ^ n29950 ^ n7551 ;
  assign n32046 = ( n310 & ~n9246 ) | ( n310 & n32045 ) | ( ~n9246 & n32045 ) ;
  assign n32047 = n15293 ^ n9380 ^ n2882 ;
  assign n32048 = n32046 | n32047 ;
  assign n32049 = n30256 ^ n29726 ^ n7751 ;
  assign n32050 = n7622 | n11762 ;
  assign n32051 = ~n12366 & n32050 ;
  assign n32052 = n32051 ^ n15316 ^ n5153 ;
  assign n32053 = n20314 ^ n16188 ^ n7803 ;
  assign n32054 = ~n5169 & n11359 ;
  assign n32055 = n8345 & n32054 ;
  assign n32056 = ( ~n5472 & n20867 ) | ( ~n5472 & n32055 ) | ( n20867 & n32055 ) ;
  assign n32057 = ( n11140 & n32053 ) | ( n11140 & ~n32056 ) | ( n32053 & ~n32056 ) ;
  assign n32058 = n27487 ^ n20692 ^ 1'b0 ;
  assign n32059 = n7524 & n30784 ;
  assign n32060 = ~n3883 & n32059 ;
  assign n32061 = n6030 & ~n6105 ;
  assign n32062 = ~n16281 & n32061 ;
  assign n32063 = n27145 ^ n4195 ^ 1'b0 ;
  assign n32064 = n8282 & n32063 ;
  assign n32065 = n32064 ^ n28464 ^ n6118 ;
  assign n32066 = n13667 ^ n11313 ^ n4856 ;
  assign n32067 = n30365 | n32066 ;
  assign n32068 = n5374 ^ n1455 ^ 1'b0 ;
  assign n32069 = n1953 | n5108 ;
  assign n32070 = n32069 ^ n13868 ^ n6238 ;
  assign n32073 = ( ~n18119 & n23633 ) | ( ~n18119 & n27968 ) | ( n23633 & n27968 ) ;
  assign n32074 = n32073 ^ n26711 ^ n17529 ;
  assign n32071 = n21798 ^ n15200 ^ n14170 ;
  assign n32072 = n32071 ^ n13580 ^ 1'b0 ;
  assign n32075 = n32074 ^ n32072 ^ n15653 ;
  assign n32076 = n24050 ^ n16022 ^ n13651 ;
  assign n32077 = n3135 & n30041 ;
  assign n32078 = ~n6664 & n32077 ;
  assign n32079 = ( n15368 & ~n32076 ) | ( n15368 & n32078 ) | ( ~n32076 & n32078 ) ;
  assign n32080 = n21138 ^ n11949 ^ n8280 ;
  assign n32081 = n32080 ^ n5862 ^ n348 ;
  assign n32082 = n3461 | n20973 ;
  assign n32083 = n8493 | n32082 ;
  assign n32084 = n15272 & ~n19158 ;
  assign n32085 = n1862 & n7084 ;
  assign n32086 = n32085 ^ n20418 ^ 1'b0 ;
  assign n32087 = n32086 ^ n13930 ^ 1'b0 ;
  assign n32088 = n3257 & n32087 ;
  assign y0 = x0 ;
  assign y1 = x3 ;
  assign y2 = x4 ;
  assign y3 = x6 ;
  assign y4 = x13 ;
  assign y5 = x16 ;
  assign y6 = x24 ;
  assign y7 = x30 ;
  assign y8 = x42 ;
  assign y9 = x58 ;
  assign y10 = x78 ;
  assign y11 = x85 ;
  assign y12 = x110 ;
  assign y13 = n129 ;
  assign y14 = n130 ;
  assign y15 = n131 ;
  assign y16 = ~n133 ;
  assign y17 = ~1'b0 ;
  assign y18 = ~n136 ;
  assign y19 = n137 ;
  assign y20 = n140 ;
  assign y21 = n144 ;
  assign y22 = n145 ;
  assign y23 = n148 ;
  assign y24 = ~n153 ;
  assign y25 = ~n159 ;
  assign y26 = n161 ;
  assign y27 = ~n163 ;
  assign y28 = ~n164 ;
  assign y29 = ~n167 ;
  assign y30 = n172 ;
  assign y31 = n178 ;
  assign y32 = n179 ;
  assign y33 = ~1'b0 ;
  assign y34 = ~n190 ;
  assign y35 = n192 ;
  assign y36 = ~n194 ;
  assign y37 = ~1'b0 ;
  assign y38 = ~n197 ;
  assign y39 = n200 ;
  assign y40 = ~n209 ;
  assign y41 = ~n220 ;
  assign y42 = ~n230 ;
  assign y43 = n233 ;
  assign y44 = ~n236 ;
  assign y45 = n238 ;
  assign y46 = ~n242 ;
  assign y47 = n251 ;
  assign y48 = ~n253 ;
  assign y49 = n266 ;
  assign y50 = n271 ;
  assign y51 = n272 ;
  assign y52 = ~1'b0 ;
  assign y53 = n273 ;
  assign y54 = ~n285 ;
  assign y55 = n289 ;
  assign y56 = n292 ;
  assign y57 = n296 ;
  assign y58 = n300 ;
  assign y59 = ~n303 ;
  assign y60 = n305 ;
  assign y61 = ~n312 ;
  assign y62 = n314 ;
  assign y63 = ~1'b0 ;
  assign y64 = ~n320 ;
  assign y65 = ~1'b0 ;
  assign y66 = n325 ;
  assign y67 = ~n339 ;
  assign y68 = n344 ;
  assign y69 = n345 ;
  assign y70 = n350 ;
  assign y71 = ~n357 ;
  assign y72 = ~1'b0 ;
  assign y73 = n367 ;
  assign y74 = n374 ;
  assign y75 = n378 ;
  assign y76 = ~n386 ;
  assign y77 = n389 ;
  assign y78 = ~n405 ;
  assign y79 = ~n407 ;
  assign y80 = ~1'b0 ;
  assign y81 = ~n415 ;
  assign y82 = n420 ;
  assign y83 = ~n426 ;
  assign y84 = n429 ;
  assign y85 = ~n434 ;
  assign y86 = ~1'b0 ;
  assign y87 = ~n436 ;
  assign y88 = ~1'b0 ;
  assign y89 = ~n442 ;
  assign y90 = ~1'b0 ;
  assign y91 = ~n445 ;
  assign y92 = n458 ;
  assign y93 = ~n460 ;
  assign y94 = ~n462 ;
  assign y95 = ~n464 ;
  assign y96 = n476 ;
  assign y97 = n201 ;
  assign y98 = ~n477 ;
  assign y99 = n480 ;
  assign y100 = n489 ;
  assign y101 = n491 ;
  assign y102 = ~1'b0 ;
  assign y103 = n494 ;
  assign y104 = ~1'b0 ;
  assign y105 = ~n508 ;
  assign y106 = ~1'b0 ;
  assign y107 = n511 ;
  assign y108 = n528 ;
  assign y109 = n547 ;
  assign y110 = ~n553 ;
  assign y111 = n555 ;
  assign y112 = n559 ;
  assign y113 = n561 ;
  assign y114 = n563 ;
  assign y115 = ~n578 ;
  assign y116 = n594 ;
  assign y117 = ~n602 ;
  assign y118 = n605 ;
  assign y119 = ~n614 ;
  assign y120 = ~n630 ;
  assign y121 = n634 ;
  assign y122 = ~n637 ;
  assign y123 = ~n645 ;
  assign y124 = n648 ;
  assign y125 = ~n650 ;
  assign y126 = n651 ;
  assign y127 = ~n653 ;
  assign y128 = ~n657 ;
  assign y129 = ~n668 ;
  assign y130 = ~n673 ;
  assign y131 = ~n680 ;
  assign y132 = n689 ;
  assign y133 = ~n690 ;
  assign y134 = n695 ;
  assign y135 = ~1'b0 ;
  assign y136 = ~n704 ;
  assign y137 = n709 ;
  assign y138 = n711 ;
  assign y139 = ~n718 ;
  assign y140 = n724 ;
  assign y141 = n459 ;
  assign y142 = n725 ;
  assign y143 = n731 ;
  assign y144 = n733 ;
  assign y145 = ~n735 ;
  assign y146 = ~n737 ;
  assign y147 = n744 ;
  assign y148 = n754 ;
  assign y149 = ~n759 ;
  assign y150 = n767 ;
  assign y151 = ~n771 ;
  assign y152 = ~n774 ;
  assign y153 = n778 ;
  assign y154 = ~n779 ;
  assign y155 = ~n782 ;
  assign y156 = ~n784 ;
  assign y157 = ~n785 ;
  assign y158 = ~n789 ;
  assign y159 = n794 ;
  assign y160 = ~1'b0 ;
  assign y161 = n796 ;
  assign y162 = n798 ;
  assign y163 = ~n809 ;
  assign y164 = n810 ;
  assign y165 = n822 ;
  assign y166 = ~n826 ;
  assign y167 = n827 ;
  assign y168 = n829 ;
  assign y169 = ~n835 ;
  assign y170 = ~1'b0 ;
  assign y171 = ~n837 ;
  assign y172 = ~n838 ;
  assign y173 = ~n839 ;
  assign y174 = n845 ;
  assign y175 = ~n846 ;
  assign y176 = ~n848 ;
  assign y177 = n852 ;
  assign y178 = n853 ;
  assign y179 = ~n855 ;
  assign y180 = ~n858 ;
  assign y181 = n860 ;
  assign y182 = ~n861 ;
  assign y183 = ~n393 ;
  assign y184 = n865 ;
  assign y185 = ~1'b0 ;
  assign y186 = ~n867 ;
  assign y187 = ~n869 ;
  assign y188 = ~n878 ;
  assign y189 = ~n887 ;
  assign y190 = ~n896 ;
  assign y191 = ~n901 ;
  assign y192 = ~n904 ;
  assign y193 = ~n908 ;
  assign y194 = n921 ;
  assign y195 = ~n923 ;
  assign y196 = n927 ;
  assign y197 = ~n928 ;
  assign y198 = ~n931 ;
  assign y199 = n945 ;
  assign y200 = ~n953 ;
  assign y201 = n963 ;
  assign y202 = ~n964 ;
  assign y203 = n971 ;
  assign y204 = ~1'b0 ;
  assign y205 = n973 ;
  assign y206 = n976 ;
  assign y207 = ~n977 ;
  assign y208 = ~n990 ;
  assign y209 = n993 ;
  assign y210 = n996 ;
  assign y211 = ~n998 ;
  assign y212 = ~n1009 ;
  assign y213 = ~n1013 ;
  assign y214 = n1019 ;
  assign y215 = ~n1020 ;
  assign y216 = ~n1023 ;
  assign y217 = ~n1028 ;
  assign y218 = n1036 ;
  assign y219 = ~n1039 ;
  assign y220 = ~n1045 ;
  assign y221 = ~n1051 ;
  assign y222 = n1055 ;
  assign y223 = ~n1056 ;
  assign y224 = n1058 ;
  assign y225 = n1061 ;
  assign y226 = ~1'b0 ;
  assign y227 = ~n1062 ;
  assign y228 = n1064 ;
  assign y229 = n1068 ;
  assign y230 = n1086 ;
  assign y231 = n1095 ;
  assign y232 = ~n1106 ;
  assign y233 = ~n1109 ;
  assign y234 = n1118 ;
  assign y235 = ~n1123 ;
  assign y236 = ~n1127 ;
  assign y237 = n1139 ;
  assign y238 = ~n1141 ;
  assign y239 = n1148 ;
  assign y240 = ~1'b0 ;
  assign y241 = ~1'b0 ;
  assign y242 = ~n1153 ;
  assign y243 = n1162 ;
  assign y244 = ~n1183 ;
  assign y245 = n1187 ;
  assign y246 = n1219 ;
  assign y247 = n1221 ;
  assign y248 = ~n1223 ;
  assign y249 = ~1'b0 ;
  assign y250 = ~1'b0 ;
  assign y251 = n1231 ;
  assign y252 = ~n1234 ;
  assign y253 = n1247 ;
  assign y254 = ~n1255 ;
  assign y255 = n1257 ;
  assign y256 = ~1'b0 ;
  assign y257 = ~n1258 ;
  assign y258 = ~n1259 ;
  assign y259 = n1263 ;
  assign y260 = ~n1264 ;
  assign y261 = ~n1266 ;
  assign y262 = n1274 ;
  assign y263 = ~n1277 ;
  assign y264 = ~1'b0 ;
  assign y265 = ~1'b0 ;
  assign y266 = n1278 ;
  assign y267 = ~n1282 ;
  assign y268 = ~n1283 ;
  assign y269 = ~n1284 ;
  assign y270 = ~n1288 ;
  assign y271 = ~n1289 ;
  assign y272 = ~n1301 ;
  assign y273 = n1306 ;
  assign y274 = ~n1308 ;
  assign y275 = ~1'b0 ;
  assign y276 = n1313 ;
  assign y277 = ~n1315 ;
  assign y278 = ~n1322 ;
  assign y279 = ~n1333 ;
  assign y280 = ~n1334 ;
  assign y281 = ~n1341 ;
  assign y282 = n214 ;
  assign y283 = n1352 ;
  assign y284 = ~n1353 ;
  assign y285 = ~n1354 ;
  assign y286 = ~n1357 ;
  assign y287 = ~n1369 ;
  assign y288 = n1371 ;
  assign y289 = n1380 ;
  assign y290 = ~n1386 ;
  assign y291 = n1399 ;
  assign y292 = ~n1402 ;
  assign y293 = n1407 ;
  assign y294 = ~n1408 ;
  assign y295 = ~n1413 ;
  assign y296 = ~n1414 ;
  assign y297 = n1418 ;
  assign y298 = ~n1420 ;
  assign y299 = n1431 ;
  assign y300 = ~n1433 ;
  assign y301 = n1434 ;
  assign y302 = ~n1450 ;
  assign y303 = n1453 ;
  assign y304 = n1463 ;
  assign y305 = n1466 ;
  assign y306 = ~n1467 ;
  assign y307 = ~n1475 ;
  assign y308 = n1476 ;
  assign y309 = ~n1484 ;
  assign y310 = ~1'b0 ;
  assign y311 = ~1'b0 ;
  assign y312 = ~n1489 ;
  assign y313 = n1492 ;
  assign y314 = ~n1495 ;
  assign y315 = ~n1504 ;
  assign y316 = ~n1507 ;
  assign y317 = ~n1516 ;
  assign y318 = n1521 ;
  assign y319 = ~n1524 ;
  assign y320 = n1532 ;
  assign y321 = n1534 ;
  assign y322 = ~n1535 ;
  assign y323 = n1538 ;
  assign y324 = n1545 ;
  assign y325 = ~n1571 ;
  assign y326 = ~n1578 ;
  assign y327 = ~n1583 ;
  assign y328 = ~n1589 ;
  assign y329 = ~n1595 ;
  assign y330 = ~n1605 ;
  assign y331 = ~n1610 ;
  assign y332 = ~n1619 ;
  assign y333 = n1621 ;
  assign y334 = ~n1628 ;
  assign y335 = ~n1638 ;
  assign y336 = ~1'b0 ;
  assign y337 = ~1'b0 ;
  assign y338 = ~n1645 ;
  assign y339 = n1646 ;
  assign y340 = ~n1648 ;
  assign y341 = ~n1653 ;
  assign y342 = ~n1659 ;
  assign y343 = n1662 ;
  assign y344 = ~n1666 ;
  assign y345 = n1667 ;
  assign y346 = ~1'b0 ;
  assign y347 = ~1'b0 ;
  assign y348 = n1669 ;
  assign y349 = ~n1670 ;
  assign y350 = ~n1672 ;
  assign y351 = n1679 ;
  assign y352 = n1688 ;
  assign y353 = ~n1695 ;
  assign y354 = ~n1709 ;
  assign y355 = n1716 ;
  assign y356 = ~n1718 ;
  assign y357 = ~n1719 ;
  assign y358 = ~n1722 ;
  assign y359 = ~n1725 ;
  assign y360 = ~1'b0 ;
  assign y361 = n1728 ;
  assign y362 = ~n1731 ;
  assign y363 = ~1'b0 ;
  assign y364 = ~n1735 ;
  assign y365 = ~n1740 ;
  assign y366 = n1743 ;
  assign y367 = ~n1745 ;
  assign y368 = ~n1746 ;
  assign y369 = ~n1747 ;
  assign y370 = n1758 ;
  assign y371 = n1762 ;
  assign y372 = ~1'b0 ;
  assign y373 = n1769 ;
  assign y374 = ~n1773 ;
  assign y375 = n1779 ;
  assign y376 = n1781 ;
  assign y377 = n1788 ;
  assign y378 = ~n1793 ;
  assign y379 = n1797 ;
  assign y380 = n1800 ;
  assign y381 = ~n1801 ;
  assign y382 = n1806 ;
  assign y383 = n1819 ;
  assign y384 = n1832 ;
  assign y385 = n1833 ;
  assign y386 = n1834 ;
  assign y387 = ~n1843 ;
  assign y388 = ~1'b0 ;
  assign y389 = n1847 ;
  assign y390 = ~n1858 ;
  assign y391 = ~1'b0 ;
  assign y392 = ~1'b0 ;
  assign y393 = ~n1859 ;
  assign y394 = n1860 ;
  assign y395 = ~1'b0 ;
  assign y396 = ~1'b0 ;
  assign y397 = ~n1863 ;
  assign y398 = ~n1870 ;
  assign y399 = n1873 ;
  assign y400 = n1882 ;
  assign y401 = n1888 ;
  assign y402 = ~n1890 ;
  assign y403 = ~n1899 ;
  assign y404 = ~n1905 ;
  assign y405 = ~n1906 ;
  assign y406 = n1908 ;
  assign y407 = n1911 ;
  assign y408 = ~n1912 ;
  assign y409 = n1915 ;
  assign y410 = n1929 ;
  assign y411 = ~n1939 ;
  assign y412 = n1941 ;
  assign y413 = ~n1944 ;
  assign y414 = n1948 ;
  assign y415 = ~n1950 ;
  assign y416 = ~1'b0 ;
  assign y417 = ~1'b0 ;
  assign y418 = n1952 ;
  assign y419 = ~n1962 ;
  assign y420 = n1964 ;
  assign y421 = n1967 ;
  assign y422 = ~n1969 ;
  assign y423 = ~n1977 ;
  assign y424 = ~n1986 ;
  assign y425 = ~n1987 ;
  assign y426 = n1992 ;
  assign y427 = ~n2005 ;
  assign y428 = ~n2007 ;
  assign y429 = ~n2008 ;
  assign y430 = ~n2015 ;
  assign y431 = ~n2017 ;
  assign y432 = n2025 ;
  assign y433 = ~1'b0 ;
  assign y434 = ~n2030 ;
  assign y435 = ~n2032 ;
  assign y436 = n2053 ;
  assign y437 = n2059 ;
  assign y438 = ~n810 ;
  assign y439 = ~n2068 ;
  assign y440 = ~1'b0 ;
  assign y441 = n2071 ;
  assign y442 = n2079 ;
  assign y443 = ~n2086 ;
  assign y444 = ~n2089 ;
  assign y445 = ~n2099 ;
  assign y446 = ~n2102 ;
  assign y447 = n2103 ;
  assign y448 = n2114 ;
  assign y449 = ~n2115 ;
  assign y450 = ~n2120 ;
  assign y451 = ~n2132 ;
  assign y452 = n2143 ;
  assign y453 = n2155 ;
  assign y454 = n2159 ;
  assign y455 = ~n2162 ;
  assign y456 = n2170 ;
  assign y457 = ~1'b0 ;
  assign y458 = n2174 ;
  assign y459 = ~n2179 ;
  assign y460 = n2192 ;
  assign y461 = ~n2196 ;
  assign y462 = ~n2201 ;
  assign y463 = ~n2202 ;
  assign y464 = n2204 ;
  assign y465 = ~n2205 ;
  assign y466 = ~n2209 ;
  assign y467 = ~n2213 ;
  assign y468 = n2220 ;
  assign y469 = ~n2226 ;
  assign y470 = ~1'b0 ;
  assign y471 = n2232 ;
  assign y472 = n2235 ;
  assign y473 = n2238 ;
  assign y474 = ~n2244 ;
  assign y475 = n2249 ;
  assign y476 = ~n2250 ;
  assign y477 = n2251 ;
  assign y478 = n2253 ;
  assign y479 = n2260 ;
  assign y480 = ~n2261 ;
  assign y481 = n2270 ;
  assign y482 = ~n2271 ;
  assign y483 = n2278 ;
  assign y484 = ~n2280 ;
  assign y485 = ~1'b0 ;
  assign y486 = ~n2303 ;
  assign y487 = n2308 ;
  assign y488 = ~n2319 ;
  assign y489 = ~n2326 ;
  assign y490 = ~n2327 ;
  assign y491 = n2339 ;
  assign y492 = ~1'b0 ;
  assign y493 = ~n2341 ;
  assign y494 = n2346 ;
  assign y495 = n2364 ;
  assign y496 = n2368 ;
  assign y497 = ~n2371 ;
  assign y498 = n2376 ;
  assign y499 = n2379 ;
  assign y500 = ~n2387 ;
  assign y501 = ~n2389 ;
  assign y502 = ~n2390 ;
  assign y503 = ~n2396 ;
  assign y504 = n2398 ;
  assign y505 = n2412 ;
  assign y506 = ~n2420 ;
  assign y507 = ~n2425 ;
  assign y508 = ~n2427 ;
  assign y509 = ~n2433 ;
  assign y510 = ~n2447 ;
  assign y511 = n2455 ;
  assign y512 = ~n2458 ;
  assign y513 = n2460 ;
  assign y514 = ~n2471 ;
  assign y515 = n2473 ;
  assign y516 = 1'b0 ;
  assign y517 = ~n2476 ;
  assign y518 = n2484 ;
  assign y519 = ~1'b0 ;
  assign y520 = ~n2486 ;
  assign y521 = n2489 ;
  assign y522 = ~n2491 ;
  assign y523 = ~n2502 ;
  assign y524 = ~n2510 ;
  assign y525 = ~n2516 ;
  assign y526 = n2518 ;
  assign y527 = ~n2526 ;
  assign y528 = ~n2535 ;
  assign y529 = ~n2538 ;
  assign y530 = ~n2548 ;
  assign y531 = ~n2549 ;
  assign y532 = n2550 ;
  assign y533 = n2554 ;
  assign y534 = n2555 ;
  assign y535 = ~1'b0 ;
  assign y536 = ~n2559 ;
  assign y537 = n2562 ;
  assign y538 = ~n2566 ;
  assign y539 = n2580 ;
  assign y540 = n2582 ;
  assign y541 = n2583 ;
  assign y542 = ~n2587 ;
  assign y543 = ~1'b0 ;
  assign y544 = ~1'b0 ;
  assign y545 = ~1'b0 ;
  assign y546 = n2590 ;
  assign y547 = ~n2592 ;
  assign y548 = ~n2594 ;
  assign y549 = n2601 ;
  assign y550 = ~n2606 ;
  assign y551 = ~n2609 ;
  assign y552 = n2615 ;
  assign y553 = ~1'b0 ;
  assign y554 = ~n2617 ;
  assign y555 = ~1'b0 ;
  assign y556 = n2618 ;
  assign y557 = n2622 ;
  assign y558 = n2629 ;
  assign y559 = ~n2632 ;
  assign y560 = n2635 ;
  assign y561 = n2650 ;
  assign y562 = ~n2652 ;
  assign y563 = n2656 ;
  assign y564 = n2658 ;
  assign y565 = n2664 ;
  assign y566 = ~n2668 ;
  assign y567 = ~n2676 ;
  assign y568 = ~n2679 ;
  assign y569 = n2681 ;
  assign y570 = ~1'b0 ;
  assign y571 = n2689 ;
  assign y572 = ~n2690 ;
  assign y573 = ~n2696 ;
  assign y574 = n2707 ;
  assign y575 = ~n2710 ;
  assign y576 = ~n2714 ;
  assign y577 = n2716 ;
  assign y578 = n2725 ;
  assign y579 = n2732 ;
  assign y580 = n2741 ;
  assign y581 = ~n2744 ;
  assign y582 = ~n2745 ;
  assign y583 = n2752 ;
  assign y584 = ~n2757 ;
  assign y585 = ~n2768 ;
  assign y586 = ~n2772 ;
  assign y587 = ~n2789 ;
  assign y588 = n2798 ;
  assign y589 = n2802 ;
  assign y590 = n2803 ;
  assign y591 = n2804 ;
  assign y592 = ~n2812 ;
  assign y593 = n2813 ;
  assign y594 = ~n2820 ;
  assign y595 = ~n2821 ;
  assign y596 = n2822 ;
  assign y597 = ~n2830 ;
  assign y598 = ~1'b0 ;
  assign y599 = ~n2835 ;
  assign y600 = n2839 ;
  assign y601 = n2846 ;
  assign y602 = n2848 ;
  assign y603 = n2853 ;
  assign y604 = ~n2854 ;
  assign y605 = ~n2861 ;
  assign y606 = n2866 ;
  assign y607 = ~n2868 ;
  assign y608 = ~n2869 ;
  assign y609 = n2876 ;
  assign y610 = ~n2877 ;
  assign y611 = n2886 ;
  assign y612 = ~n2898 ;
  assign y613 = n2901 ;
  assign y614 = n2910 ;
  assign y615 = ~n2917 ;
  assign y616 = ~n2923 ;
  assign y617 = ~n2927 ;
  assign y618 = n2937 ;
  assign y619 = ~n2940 ;
  assign y620 = ~1'b0 ;
  assign y621 = ~n2953 ;
  assign y622 = ~n2954 ;
  assign y623 = ~n2957 ;
  assign y624 = n2962 ;
  assign y625 = n2964 ;
  assign y626 = ~1'b0 ;
  assign y627 = ~n2965 ;
  assign y628 = ~n2971 ;
  assign y629 = ~n2976 ;
  assign y630 = n2980 ;
  assign y631 = n2990 ;
  assign y632 = n2992 ;
  assign y633 = n3003 ;
  assign y634 = n3005 ;
  assign y635 = n3008 ;
  assign y636 = n3012 ;
  assign y637 = ~n3016 ;
  assign y638 = ~n3017 ;
  assign y639 = ~n3021 ;
  assign y640 = n3032 ;
  assign y641 = ~n3033 ;
  assign y642 = n3035 ;
  assign y643 = n3037 ;
  assign y644 = n3041 ;
  assign y645 = ~n3050 ;
  assign y646 = n3054 ;
  assign y647 = n3057 ;
  assign y648 = n3058 ;
  assign y649 = ~n3063 ;
  assign y650 = ~n3067 ;
  assign y651 = n3076 ;
  assign y652 = ~n3083 ;
  assign y653 = ~1'b0 ;
  assign y654 = ~n3087 ;
  assign y655 = ~n3089 ;
  assign y656 = ~1'b0 ;
  assign y657 = ~n3090 ;
  assign y658 = ~n3095 ;
  assign y659 = ~n3100 ;
  assign y660 = ~1'b0 ;
  assign y661 = ~n3101 ;
  assign y662 = n3106 ;
  assign y663 = ~n3111 ;
  assign y664 = n3118 ;
  assign y665 = n3121 ;
  assign y666 = n3134 ;
  assign y667 = ~1'b0 ;
  assign y668 = n3135 ;
  assign y669 = n3140 ;
  assign y670 = n3144 ;
  assign y671 = n3148 ;
  assign y672 = ~n3151 ;
  assign y673 = ~n3156 ;
  assign y674 = ~1'b0 ;
  assign y675 = ~1'b0 ;
  assign y676 = ~1'b0 ;
  assign y677 = ~1'b0 ;
  assign y678 = ~n3159 ;
  assign y679 = n3161 ;
  assign y680 = n3162 ;
  assign y681 = ~n3170 ;
  assign y682 = n3179 ;
  assign y683 = ~n3185 ;
  assign y684 = ~n3187 ;
  assign y685 = ~1'b0 ;
  assign y686 = ~n3194 ;
  assign y687 = ~n3206 ;
  assign y688 = ~n3212 ;
  assign y689 = ~n3214 ;
  assign y690 = ~n3229 ;
  assign y691 = ~n3230 ;
  assign y692 = n3234 ;
  assign y693 = n3244 ;
  assign y694 = ~1'b0 ;
  assign y695 = n3248 ;
  assign y696 = n3264 ;
  assign y697 = ~1'b0 ;
  assign y698 = ~n3266 ;
  assign y699 = n3268 ;
  assign y700 = ~n3281 ;
  assign y701 = ~n3286 ;
  assign y702 = ~1'b0 ;
  assign y703 = ~n3290 ;
  assign y704 = n3297 ;
  assign y705 = ~n3300 ;
  assign y706 = n3301 ;
  assign y707 = ~1'b0 ;
  assign y708 = ~n3308 ;
  assign y709 = ~n3314 ;
  assign y710 = ~n3317 ;
  assign y711 = ~n3322 ;
  assign y712 = n3328 ;
  assign y713 = n3334 ;
  assign y714 = ~1'b0 ;
  assign y715 = ~n3339 ;
  assign y716 = ~n3342 ;
  assign y717 = n3344 ;
  assign y718 = ~n3351 ;
  assign y719 = ~n3360 ;
  assign y720 = ~1'b0 ;
  assign y721 = ~n3377 ;
  assign y722 = ~n3389 ;
  assign y723 = ~1'b0 ;
  assign y724 = ~1'b0 ;
  assign y725 = ~n3390 ;
  assign y726 = n3391 ;
  assign y727 = ~n3402 ;
  assign y728 = ~n3407 ;
  assign y729 = ~n3408 ;
  assign y730 = ~n3411 ;
  assign y731 = ~n3418 ;
  assign y732 = ~1'b0 ;
  assign y733 = n3425 ;
  assign y734 = n3442 ;
  assign y735 = ~n3449 ;
  assign y736 = ~1'b0 ;
  assign y737 = ~1'b0 ;
  assign y738 = ~n3461 ;
  assign y739 = ~1'b0 ;
  assign y740 = ~n3465 ;
  assign y741 = n3467 ;
  assign y742 = ~n3477 ;
  assign y743 = n3482 ;
  assign y744 = ~n3484 ;
  assign y745 = n3500 ;
  assign y746 = ~n3501 ;
  assign y747 = ~n3506 ;
  assign y748 = n3507 ;
  assign y749 = ~n3508 ;
  assign y750 = ~n3514 ;
  assign y751 = n3522 ;
  assign y752 = ~n3527 ;
  assign y753 = ~1'b0 ;
  assign y754 = n3534 ;
  assign y755 = ~n3535 ;
  assign y756 = n3538 ;
  assign y757 = n3550 ;
  assign y758 = n3551 ;
  assign y759 = ~n3552 ;
  assign y760 = n3561 ;
  assign y761 = n3563 ;
  assign y762 = ~1'b0 ;
  assign y763 = ~n3566 ;
  assign y764 = n3577 ;
  assign y765 = ~n3586 ;
  assign y766 = n3594 ;
  assign y767 = n3600 ;
  assign y768 = ~n3602 ;
  assign y769 = n3609 ;
  assign y770 = n3612 ;
  assign y771 = ~n3620 ;
  assign y772 = n3624 ;
  assign y773 = ~n3630 ;
  assign y774 = ~1'b0 ;
  assign y775 = n3631 ;
  assign y776 = ~n3632 ;
  assign y777 = ~n3633 ;
  assign y778 = ~n3638 ;
  assign y779 = ~n3640 ;
  assign y780 = n3644 ;
  assign y781 = ~n3656 ;
  assign y782 = n3657 ;
  assign y783 = ~n3662 ;
  assign y784 = n3665 ;
  assign y785 = ~n3668 ;
  assign y786 = n3674 ;
  assign y787 = ~n3679 ;
  assign y788 = ~n3681 ;
  assign y789 = ~n3689 ;
  assign y790 = n3695 ;
  assign y791 = ~n3697 ;
  assign y792 = n3705 ;
  assign y793 = n3706 ;
  assign y794 = n3734 ;
  assign y795 = ~n3739 ;
  assign y796 = n3741 ;
  assign y797 = n3744 ;
  assign y798 = n3751 ;
  assign y799 = ~n3760 ;
  assign y800 = n3769 ;
  assign y801 = n3780 ;
  assign y802 = ~n3781 ;
  assign y803 = ~n3782 ;
  assign y804 = n3787 ;
  assign y805 = n3795 ;
  assign y806 = ~n3796 ;
  assign y807 = ~n3803 ;
  assign y808 = ~n3807 ;
  assign y809 = ~n3819 ;
  assign y810 = ~n3820 ;
  assign y811 = ~n3822 ;
  assign y812 = n3823 ;
  assign y813 = ~n3830 ;
  assign y814 = n3838 ;
  assign y815 = ~1'b0 ;
  assign y816 = ~n3839 ;
  assign y817 = ~1'b0 ;
  assign y818 = ~n3843 ;
  assign y819 = n3848 ;
  assign y820 = n3853 ;
  assign y821 = ~n3855 ;
  assign y822 = ~n3858 ;
  assign y823 = ~n3861 ;
  assign y824 = n3870 ;
  assign y825 = n3875 ;
  assign y826 = ~n3878 ;
  assign y827 = ~n3882 ;
  assign y828 = n3886 ;
  assign y829 = ~n3889 ;
  assign y830 = ~1'b0 ;
  assign y831 = ~n3892 ;
  assign y832 = n3895 ;
  assign y833 = ~n3905 ;
  assign y834 = ~n3924 ;
  assign y835 = n3932 ;
  assign y836 = n3937 ;
  assign y837 = ~n3938 ;
  assign y838 = n3945 ;
  assign y839 = ~1'b0 ;
  assign y840 = n3948 ;
  assign y841 = ~n3950 ;
  assign y842 = ~n3964 ;
  assign y843 = n3965 ;
  assign y844 = ~1'b0 ;
  assign y845 = n3970 ;
  assign y846 = n3973 ;
  assign y847 = n3983 ;
  assign y848 = ~1'b0 ;
  assign y849 = n3989 ;
  assign y850 = n3997 ;
  assign y851 = ~n3999 ;
  assign y852 = ~n4001 ;
  assign y853 = ~n4013 ;
  assign y854 = ~n4015 ;
  assign y855 = n4017 ;
  assign y856 = ~n4020 ;
  assign y857 = n4021 ;
  assign y858 = ~n4023 ;
  assign y859 = ~n4033 ;
  assign y860 = ~n4035 ;
  assign y861 = ~n4038 ;
  assign y862 = ~n4039 ;
  assign y863 = ~n4048 ;
  assign y864 = n4076 ;
  assign y865 = ~1'b0 ;
  assign y866 = n4082 ;
  assign y867 = ~n4087 ;
  assign y868 = ~n4108 ;
  assign y869 = ~n4109 ;
  assign y870 = ~n4110 ;
  assign y871 = ~n4114 ;
  assign y872 = ~n4121 ;
  assign y873 = ~n4122 ;
  assign y874 = n4125 ;
  assign y875 = ~1'b0 ;
  assign y876 = ~1'b0 ;
  assign y877 = ~n4126 ;
  assign y878 = ~n4128 ;
  assign y879 = ~n4129 ;
  assign y880 = ~n4134 ;
  assign y881 = n4136 ;
  assign y882 = n4137 ;
  assign y883 = n4138 ;
  assign y884 = n4141 ;
  assign y885 = n4149 ;
  assign y886 = ~n4162 ;
  assign y887 = n1971 ;
  assign y888 = ~n4169 ;
  assign y889 = ~n4172 ;
  assign y890 = ~n4181 ;
  assign y891 = ~n4187 ;
  assign y892 = n4192 ;
  assign y893 = ~n4193 ;
  assign y894 = n4201 ;
  assign y895 = ~n4210 ;
  assign y896 = n4219 ;
  assign y897 = n4222 ;
  assign y898 = ~n4225 ;
  assign y899 = ~n4229 ;
  assign y900 = n4233 ;
  assign y901 = ~n4255 ;
  assign y902 = ~1'b0 ;
  assign y903 = n4257 ;
  assign y904 = ~n4261 ;
  assign y905 = ~n4263 ;
  assign y906 = ~n4267 ;
  assign y907 = n4268 ;
  assign y908 = ~n4270 ;
  assign y909 = ~n4276 ;
  assign y910 = n4280 ;
  assign y911 = n4283 ;
  assign y912 = n4296 ;
  assign y913 = n4298 ;
  assign y914 = ~n4306 ;
  assign y915 = n4308 ;
  assign y916 = n4313 ;
  assign y917 = ~n4319 ;
  assign y918 = ~1'b0 ;
  assign y919 = ~n4322 ;
  assign y920 = ~n4327 ;
  assign y921 = n4332 ;
  assign y922 = ~n4335 ;
  assign y923 = n4339 ;
  assign y924 = n4340 ;
  assign y925 = ~n4345 ;
  assign y926 = ~n4356 ;
  assign y927 = n4359 ;
  assign y928 = ~n4360 ;
  assign y929 = ~n4363 ;
  assign y930 = n4369 ;
  assign y931 = ~n4381 ;
  assign y932 = ~n4385 ;
  assign y933 = n4387 ;
  assign y934 = ~n4390 ;
  assign y935 = n4394 ;
  assign y936 = n4398 ;
  assign y937 = n4404 ;
  assign y938 = ~n4408 ;
  assign y939 = ~n4418 ;
  assign y940 = ~n4422 ;
  assign y941 = ~n4427 ;
  assign y942 = ~1'b0 ;
  assign y943 = ~n4430 ;
  assign y944 = ~n4431 ;
  assign y945 = n4435 ;
  assign y946 = n4436 ;
  assign y947 = n4440 ;
  assign y948 = n4449 ;
  assign y949 = n4458 ;
  assign y950 = n4466 ;
  assign y951 = ~n4468 ;
  assign y952 = ~n4477 ;
  assign y953 = ~1'b0 ;
  assign y954 = n4482 ;
  assign y955 = n4487 ;
  assign y956 = n4493 ;
  assign y957 = n4500 ;
  assign y958 = ~n4513 ;
  assign y959 = ~1'b0 ;
  assign y960 = ~n4515 ;
  assign y961 = n4517 ;
  assign y962 = n4518 ;
  assign y963 = ~1'b0 ;
  assign y964 = ~n4525 ;
  assign y965 = ~n4537 ;
  assign y966 = ~n1826 ;
  assign y967 = n4539 ;
  assign y968 = ~1'b0 ;
  assign y969 = n4548 ;
  assign y970 = n4569 ;
  assign y971 = n4571 ;
  assign y972 = n4573 ;
  assign y973 = ~n4576 ;
  assign y974 = n4586 ;
  assign y975 = n4601 ;
  assign y976 = ~n4609 ;
  assign y977 = ~n4614 ;
  assign y978 = ~n4615 ;
  assign y979 = ~n4625 ;
  assign y980 = ~n4641 ;
  assign y981 = n4642 ;
  assign y982 = ~n4644 ;
  assign y983 = ~n4647 ;
  assign y984 = n4655 ;
  assign y985 = n4657 ;
  assign y986 = ~1'b0 ;
  assign y987 = ~n4660 ;
  assign y988 = n4664 ;
  assign y989 = n4666 ;
  assign y990 = ~1'b0 ;
  assign y991 = ~n4679 ;
  assign y992 = ~n4680 ;
  assign y993 = ~n4683 ;
  assign y994 = ~n4694 ;
  assign y995 = n4697 ;
  assign y996 = ~n4707 ;
  assign y997 = ~n4710 ;
  assign y998 = n4712 ;
  assign y999 = ~n4715 ;
  assign y1000 = n4719 ;
  assign y1001 = ~n4720 ;
  assign y1002 = ~n4723 ;
  assign y1003 = n4726 ;
  assign y1004 = ~n4727 ;
  assign y1005 = ~n4729 ;
  assign y1006 = ~1'b0 ;
  assign y1007 = n4744 ;
  assign y1008 = ~n4757 ;
  assign y1009 = n4758 ;
  assign y1010 = n4760 ;
  assign y1011 = n4765 ;
  assign y1012 = ~n4783 ;
  assign y1013 = ~n4788 ;
  assign y1014 = n4799 ;
  assign y1015 = n4802 ;
  assign y1016 = ~1'b0 ;
  assign y1017 = ~n4811 ;
  assign y1018 = ~n4814 ;
  assign y1019 = ~n4818 ;
  assign y1020 = ~1'b0 ;
  assign y1021 = ~n4823 ;
  assign y1022 = n4829 ;
  assign y1023 = ~n4835 ;
  assign y1024 = ~n4839 ;
  assign y1025 = ~n4851 ;
  assign y1026 = n4857 ;
  assign y1027 = ~n4868 ;
  assign y1028 = ~1'b0 ;
  assign y1029 = n4872 ;
  assign y1030 = n4877 ;
  assign y1031 = ~1'b0 ;
  assign y1032 = n4879 ;
  assign y1033 = n4880 ;
  assign y1034 = ~1'b0 ;
  assign y1035 = ~n4881 ;
  assign y1036 = ~n4883 ;
  assign y1037 = ~1'b0 ;
  assign y1038 = ~n4888 ;
  assign y1039 = n4896 ;
  assign y1040 = ~n4897 ;
  assign y1041 = ~1'b0 ;
  assign y1042 = ~1'b0 ;
  assign y1043 = ~n4908 ;
  assign y1044 = ~n4909 ;
  assign y1045 = n4912 ;
  assign y1046 = ~n4923 ;
  assign y1047 = ~n4933 ;
  assign y1048 = n4937 ;
  assign y1049 = n4945 ;
  assign y1050 = n4958 ;
  assign y1051 = ~n4960 ;
  assign y1052 = ~1'b0 ;
  assign y1053 = ~n4963 ;
  assign y1054 = n4970 ;
  assign y1055 = n4982 ;
  assign y1056 = n4989 ;
  assign y1057 = ~n4992 ;
  assign y1058 = ~n4997 ;
  assign y1059 = n5000 ;
  assign y1060 = ~n5001 ;
  assign y1061 = ~n5002 ;
  assign y1062 = ~n5007 ;
  assign y1063 = ~n5009 ;
  assign y1064 = n5011 ;
  assign y1065 = ~n5022 ;
  assign y1066 = n5030 ;
  assign y1067 = ~n5035 ;
  assign y1068 = n5037 ;
  assign y1069 = ~n5039 ;
  assign y1070 = ~1'b0 ;
  assign y1071 = ~n5040 ;
  assign y1072 = ~n5043 ;
  assign y1073 = ~n5053 ;
  assign y1074 = n5057 ;
  assign y1075 = ~n5059 ;
  assign y1076 = ~n5061 ;
  assign y1077 = 1'b0 ;
  assign y1078 = ~n5063 ;
  assign y1079 = ~n5065 ;
  assign y1080 = ~n5067 ;
  assign y1081 = ~n5073 ;
  assign y1082 = ~n5082 ;
  assign y1083 = ~1'b0 ;
  assign y1084 = n5093 ;
  assign y1085 = ~n5097 ;
  assign y1086 = n5098 ;
  assign y1087 = ~n5113 ;
  assign y1088 = ~1'b0 ;
  assign y1089 = ~1'b0 ;
  assign y1090 = n5117 ;
  assign y1091 = ~n5120 ;
  assign y1092 = n5122 ;
  assign y1093 = ~n5127 ;
  assign y1094 = n5129 ;
  assign y1095 = ~n5138 ;
  assign y1096 = n5139 ;
  assign y1097 = n5141 ;
  assign y1098 = ~n5148 ;
  assign y1099 = n5151 ;
  assign y1100 = n5159 ;
  assign y1101 = ~n5160 ;
  assign y1102 = ~n5167 ;
  assign y1103 = ~n5176 ;
  assign y1104 = ~n5177 ;
  assign y1105 = ~n5183 ;
  assign y1106 = n5184 ;
  assign y1107 = ~1'b0 ;
  assign y1108 = ~n5194 ;
  assign y1109 = ~n5197 ;
  assign y1110 = n5204 ;
  assign y1111 = n5207 ;
  assign y1112 = ~1'b0 ;
  assign y1113 = n5210 ;
  assign y1114 = ~n5219 ;
  assign y1115 = ~n5223 ;
  assign y1116 = ~1'b0 ;
  assign y1117 = n5234 ;
  assign y1118 = n5238 ;
  assign y1119 = n5246 ;
  assign y1120 = ~n5250 ;
  assign y1121 = n5253 ;
  assign y1122 = n5256 ;
  assign y1123 = n5263 ;
  assign y1124 = ~n5268 ;
  assign y1125 = n5270 ;
  assign y1126 = ~1'b0 ;
  assign y1127 = ~1'b0 ;
  assign y1128 = n5271 ;
  assign y1129 = ~1'b0 ;
  assign y1130 = n5273 ;
  assign y1131 = n5297 ;
  assign y1132 = n5298 ;
  assign y1133 = ~n5320 ;
  assign y1134 = ~n5328 ;
  assign y1135 = ~n5331 ;
  assign y1136 = n5362 ;
  assign y1137 = n2517 ;
  assign y1138 = ~n5365 ;
  assign y1139 = ~n5368 ;
  assign y1140 = ~n5369 ;
  assign y1141 = n5379 ;
  assign y1142 = n5383 ;
  assign y1143 = ~n5386 ;
  assign y1144 = ~n5392 ;
  assign y1145 = ~n1877 ;
  assign y1146 = n5393 ;
  assign y1147 = ~n5397 ;
  assign y1148 = ~1'b0 ;
  assign y1149 = n5409 ;
  assign y1150 = n5413 ;
  assign y1151 = ~n5418 ;
  assign y1152 = n5422 ;
  assign y1153 = ~n5423 ;
  assign y1154 = n5432 ;
  assign y1155 = ~n5437 ;
  assign y1156 = n5450 ;
  assign y1157 = n5453 ;
  assign y1158 = n5457 ;
  assign y1159 = ~n5458 ;
  assign y1160 = ~1'b0 ;
  assign y1161 = ~n5459 ;
  assign y1162 = ~n5460 ;
  assign y1163 = n5471 ;
  assign y1164 = n5479 ;
  assign y1165 = ~n5480 ;
  assign y1166 = ~n5481 ;
  assign y1167 = ~1'b0 ;
  assign y1168 = n5500 ;
  assign y1169 = ~n5501 ;
  assign y1170 = ~n5502 ;
  assign y1171 = ~n5503 ;
  assign y1172 = ~n5508 ;
  assign y1173 = n5510 ;
  assign y1174 = ~n5513 ;
  assign y1175 = n5518 ;
  assign y1176 = ~1'b0 ;
  assign y1177 = n5524 ;
  assign y1178 = ~n5525 ;
  assign y1179 = n5529 ;
  assign y1180 = ~n5531 ;
  assign y1181 = n5536 ;
  assign y1182 = n5548 ;
  assign y1183 = ~n5558 ;
  assign y1184 = ~n5564 ;
  assign y1185 = n5570 ;
  assign y1186 = n5574 ;
  assign y1187 = n5580 ;
  assign y1188 = n5581 ;
  assign y1189 = n5583 ;
  assign y1190 = n5585 ;
  assign y1191 = ~n5590 ;
  assign y1192 = n5603 ;
  assign y1193 = n5621 ;
  assign y1194 = ~n5627 ;
  assign y1195 = n5629 ;
  assign y1196 = n5641 ;
  assign y1197 = ~1'b0 ;
  assign y1198 = ~n5647 ;
  assign y1199 = ~n5660 ;
  assign y1200 = ~1'b0 ;
  assign y1201 = ~n5664 ;
  assign y1202 = n5665 ;
  assign y1203 = n5674 ;
  assign y1204 = n5681 ;
  assign y1205 = n5684 ;
  assign y1206 = ~n5688 ;
  assign y1207 = n5696 ;
  assign y1208 = n3935 ;
  assign y1209 = n5697 ;
  assign y1210 = n5703 ;
  assign y1211 = n5706 ;
  assign y1212 = ~1'b0 ;
  assign y1213 = ~n5715 ;
  assign y1214 = ~n5721 ;
  assign y1215 = n5728 ;
  assign y1216 = ~n5729 ;
  assign y1217 = ~1'b0 ;
  assign y1218 = ~n5733 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~n5739 ;
  assign y1221 = ~n5756 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = n5759 ;
  assign y1224 = n5760 ;
  assign y1225 = ~n5762 ;
  assign y1226 = ~1'b0 ;
  assign y1227 = ~n5763 ;
  assign y1228 = ~n5766 ;
  assign y1229 = n5771 ;
  assign y1230 = n5773 ;
  assign y1231 = ~1'b0 ;
  assign y1232 = n5774 ;
  assign y1233 = n5776 ;
  assign y1234 = ~n5786 ;
  assign y1235 = ~n5788 ;
  assign y1236 = ~1'b0 ;
  assign y1237 = ~n5789 ;
  assign y1238 = ~n5792 ;
  assign y1239 = n5794 ;
  assign y1240 = ~n5805 ;
  assign y1241 = n336 ;
  assign y1242 = ~n5812 ;
  assign y1243 = n5825 ;
  assign y1244 = ~n5826 ;
  assign y1245 = ~n5830 ;
  assign y1246 = ~n5832 ;
  assign y1247 = n5834 ;
  assign y1248 = ~n5838 ;
  assign y1249 = ~1'b0 ;
  assign y1250 = ~1'b0 ;
  assign y1251 = n5844 ;
  assign y1252 = n5845 ;
  assign y1253 = n5859 ;
  assign y1254 = ~n5860 ;
  assign y1255 = n5861 ;
  assign y1256 = ~n5870 ;
  assign y1257 = ~n5872 ;
  assign y1258 = ~1'b0 ;
  assign y1259 = ~n5873 ;
  assign y1260 = n5880 ;
  assign y1261 = ~n5886 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = ~n5891 ;
  assign y1264 = n5898 ;
  assign y1265 = ~n5899 ;
  assign y1266 = ~n5902 ;
  assign y1267 = n5904 ;
  assign y1268 = ~n5905 ;
  assign y1269 = n5917 ;
  assign y1270 = ~n5918 ;
  assign y1271 = n5922 ;
  assign y1272 = ~1'b0 ;
  assign y1273 = ~n5925 ;
  assign y1274 = ~n5927 ;
  assign y1275 = ~n5929 ;
  assign y1276 = n5930 ;
  assign y1277 = ~n5933 ;
  assign y1278 = ~n5937 ;
  assign y1279 = ~n5940 ;
  assign y1280 = ~n5946 ;
  assign y1281 = n5952 ;
  assign y1282 = n5959 ;
  assign y1283 = ~1'b0 ;
  assign y1284 = ~n5971 ;
  assign y1285 = ~n5974 ;
  assign y1286 = n5980 ;
  assign y1287 = n5988 ;
  assign y1288 = ~n5991 ;
  assign y1289 = n5994 ;
  assign y1290 = ~n5995 ;
  assign y1291 = ~n6006 ;
  assign y1292 = n6014 ;
  assign y1293 = ~n6015 ;
  assign y1294 = ~n6021 ;
  assign y1295 = n6030 ;
  assign y1296 = ~n6031 ;
  assign y1297 = ~n6038 ;
  assign y1298 = ~n6040 ;
  assign y1299 = ~n6041 ;
  assign y1300 = n4424 ;
  assign y1301 = ~n6048 ;
  assign y1302 = ~1'b0 ;
  assign y1303 = n6054 ;
  assign y1304 = n6056 ;
  assign y1305 = ~n6058 ;
  assign y1306 = n6062 ;
  assign y1307 = ~n6066 ;
  assign y1308 = ~1'b0 ;
  assign y1309 = ~n6067 ;
  assign y1310 = n6068 ;
  assign y1311 = ~n6075 ;
  assign y1312 = n6079 ;
  assign y1313 = ~n6085 ;
  assign y1314 = n6086 ;
  assign y1315 = ~n6096 ;
  assign y1316 = n6100 ;
  assign y1317 = n6111 ;
  assign y1318 = ~n6115 ;
  assign y1319 = ~n6121 ;
  assign y1320 = ~n6122 ;
  assign y1321 = ~n6124 ;
  assign y1322 = n6126 ;
  assign y1323 = ~n6140 ;
  assign y1324 = n6148 ;
  assign y1325 = n6152 ;
  assign y1326 = n6154 ;
  assign y1327 = ~n6157 ;
  assign y1328 = n6159 ;
  assign y1329 = ~n6170 ;
  assign y1330 = ~1'b0 ;
  assign y1331 = ~n6174 ;
  assign y1332 = n6177 ;
  assign y1333 = ~n6179 ;
  assign y1334 = ~1'b0 ;
  assign y1335 = ~1'b0 ;
  assign y1336 = ~n6180 ;
  assign y1337 = ~1'b0 ;
  assign y1338 = ~n6207 ;
  assign y1339 = n6208 ;
  assign y1340 = ~n6214 ;
  assign y1341 = ~n6216 ;
  assign y1342 = ~n6223 ;
  assign y1343 = ~n6228 ;
  assign y1344 = n6244 ;
  assign y1345 = ~n6252 ;
  assign y1346 = ~n6253 ;
  assign y1347 = ~n6254 ;
  assign y1348 = ~1'b0 ;
  assign y1349 = n6264 ;
  assign y1350 = n6269 ;
  assign y1351 = n6270 ;
  assign y1352 = ~n6272 ;
  assign y1353 = n6273 ;
  assign y1354 = ~n6274 ;
  assign y1355 = n6276 ;
  assign y1356 = n6277 ;
  assign y1357 = ~n6282 ;
  assign y1358 = n6293 ;
  assign y1359 = n6295 ;
  assign y1360 = ~n6299 ;
  assign y1361 = ~n6300 ;
  assign y1362 = n6304 ;
  assign y1363 = ~1'b0 ;
  assign y1364 = ~n6307 ;
  assign y1365 = n6308 ;
  assign y1366 = ~1'b0 ;
  assign y1367 = ~n6310 ;
  assign y1368 = ~1'b0 ;
  assign y1369 = ~1'b0 ;
  assign y1370 = ~n6312 ;
  assign y1371 = n6322 ;
  assign y1372 = n6329 ;
  assign y1373 = ~n6332 ;
  assign y1374 = ~n6334 ;
  assign y1375 = ~n6336 ;
  assign y1376 = ~1'b0 ;
  assign y1377 = n6342 ;
  assign y1378 = ~n6356 ;
  assign y1379 = n6358 ;
  assign y1380 = n6365 ;
  assign y1381 = ~n6367 ;
  assign y1382 = ~n6371 ;
  assign y1383 = ~n6373 ;
  assign y1384 = n6375 ;
  assign y1385 = n6376 ;
  assign y1386 = ~n6379 ;
  assign y1387 = ~n6392 ;
  assign y1388 = ~n6397 ;
  assign y1389 = n6418 ;
  assign y1390 = ~n6419 ;
  assign y1391 = ~n6423 ;
  assign y1392 = n6428 ;
  assign y1393 = ~n6433 ;
  assign y1394 = ~n6434 ;
  assign y1395 = n6436 ;
  assign y1396 = n6441 ;
  assign y1397 = ~n6444 ;
  assign y1398 = n6445 ;
  assign y1399 = ~n6449 ;
  assign y1400 = n6451 ;
  assign y1401 = ~n6452 ;
  assign y1402 = ~n6465 ;
  assign y1403 = n6469 ;
  assign y1404 = ~n6474 ;
  assign y1405 = ~1'b0 ;
  assign y1406 = n6475 ;
  assign y1407 = n6484 ;
  assign y1408 = ~n6502 ;
  assign y1409 = ~1'b0 ;
  assign y1410 = n6504 ;
  assign y1411 = n6507 ;
  assign y1412 = n6513 ;
  assign y1413 = ~1'b0 ;
  assign y1414 = ~n6528 ;
  assign y1415 = n6531 ;
  assign y1416 = ~n6534 ;
  assign y1417 = n6535 ;
  assign y1418 = n6540 ;
  assign y1419 = ~1'b0 ;
  assign y1420 = ~n6541 ;
  assign y1421 = ~1'b0 ;
  assign y1422 = ~n6543 ;
  assign y1423 = ~n6551 ;
  assign y1424 = n6552 ;
  assign y1425 = ~n6554 ;
  assign y1426 = n6559 ;
  assign y1427 = n6569 ;
  assign y1428 = ~n6570 ;
  assign y1429 = ~n6573 ;
  assign y1430 = n6577 ;
  assign y1431 = ~n6594 ;
  assign y1432 = ~n6600 ;
  assign y1433 = n6605 ;
  assign y1434 = n6608 ;
  assign y1435 = ~n6619 ;
  assign y1436 = ~n6623 ;
  assign y1437 = n6627 ;
  assign y1438 = n6630 ;
  assign y1439 = n6631 ;
  assign y1440 = ~n6634 ;
  assign y1441 = ~n6638 ;
  assign y1442 = n6644 ;
  assign y1443 = n6647 ;
  assign y1444 = ~n6657 ;
  assign y1445 = n6668 ;
  assign y1446 = n6673 ;
  assign y1447 = ~n6675 ;
  assign y1448 = n6676 ;
  assign y1449 = ~n6679 ;
  assign y1450 = n6681 ;
  assign y1451 = ~n6683 ;
  assign y1452 = ~n6685 ;
  assign y1453 = ~n6690 ;
  assign y1454 = ~n6697 ;
  assign y1455 = n6699 ;
  assign y1456 = ~n6715 ;
  assign y1457 = n6718 ;
  assign y1458 = ~n6723 ;
  assign y1459 = ~n6729 ;
  assign y1460 = n6733 ;
  assign y1461 = ~n6738 ;
  assign y1462 = ~n6745 ;
  assign y1463 = ~n6751 ;
  assign y1464 = n6758 ;
  assign y1465 = ~n6763 ;
  assign y1466 = n6764 ;
  assign y1467 = ~n6765 ;
  assign y1468 = n6775 ;
  assign y1469 = ~n6777 ;
  assign y1470 = ~n6782 ;
  assign y1471 = ~1'b0 ;
  assign y1472 = ~n6787 ;
  assign y1473 = n6788 ;
  assign y1474 = n6797 ;
  assign y1475 = n6799 ;
  assign y1476 = n6800 ;
  assign y1477 = n6806 ;
  assign y1478 = ~n6811 ;
  assign y1479 = ~n6819 ;
  assign y1480 = ~n6822 ;
  assign y1481 = n6825 ;
  assign y1482 = n6831 ;
  assign y1483 = n6833 ;
  assign y1484 = ~1'b0 ;
  assign y1485 = ~n6835 ;
  assign y1486 = n6840 ;
  assign y1487 = ~n6842 ;
  assign y1488 = n6845 ;
  assign y1489 = ~n6849 ;
  assign y1490 = ~n6852 ;
  assign y1491 = n6875 ;
  assign y1492 = ~n6878 ;
  assign y1493 = ~n6884 ;
  assign y1494 = n6891 ;
  assign y1495 = ~n6892 ;
  assign y1496 = n6903 ;
  assign y1497 = ~n6906 ;
  assign y1498 = ~1'b0 ;
  assign y1499 = n6912 ;
  assign y1500 = n6913 ;
  assign y1501 = ~1'b0 ;
  assign y1502 = n6920 ;
  assign y1503 = n6921 ;
  assign y1504 = ~n6924 ;
  assign y1505 = n6925 ;
  assign y1506 = ~n6928 ;
  assign y1507 = n6929 ;
  assign y1508 = ~n6935 ;
  assign y1509 = ~n6941 ;
  assign y1510 = n6945 ;
  assign y1511 = n6948 ;
  assign y1512 = ~n6949 ;
  assign y1513 = ~n6952 ;
  assign y1514 = n6958 ;
  assign y1515 = ~1'b0 ;
  assign y1516 = ~n6959 ;
  assign y1517 = n6966 ;
  assign y1518 = n6978 ;
  assign y1519 = ~n6980 ;
  assign y1520 = n6984 ;
  assign y1521 = ~n6993 ;
  assign y1522 = n6998 ;
  assign y1523 = ~n7008 ;
  assign y1524 = ~1'b0 ;
  assign y1525 = n7010 ;
  assign y1526 = ~n7016 ;
  assign y1527 = ~n7017 ;
  assign y1528 = n7018 ;
  assign y1529 = ~1'b0 ;
  assign y1530 = n7023 ;
  assign y1531 = ~n7025 ;
  assign y1532 = n7027 ;
  assign y1533 = ~n7039 ;
  assign y1534 = ~n7042 ;
  assign y1535 = n7047 ;
  assign y1536 = n7049 ;
  assign y1537 = ~1'b0 ;
  assign y1538 = n7051 ;
  assign y1539 = ~n7055 ;
  assign y1540 = ~1'b0 ;
  assign y1541 = n7058 ;
  assign y1542 = ~n7067 ;
  assign y1543 = ~n7070 ;
  assign y1544 = ~1'b0 ;
  assign y1545 = n7081 ;
  assign y1546 = n7085 ;
  assign y1547 = ~n7087 ;
  assign y1548 = n7089 ;
  assign y1549 = n7092 ;
  assign y1550 = ~n7093 ;
  assign y1551 = n7097 ;
  assign y1552 = n7100 ;
  assign y1553 = n7102 ;
  assign y1554 = ~n7105 ;
  assign y1555 = n7107 ;
  assign y1556 = n7109 ;
  assign y1557 = ~n7115 ;
  assign y1558 = ~n7118 ;
  assign y1559 = ~n7123 ;
  assign y1560 = ~n7126 ;
  assign y1561 = n7127 ;
  assign y1562 = ~n7137 ;
  assign y1563 = n6485 ;
  assign y1564 = ~n3900 ;
  assign y1565 = n7143 ;
  assign y1566 = ~n7144 ;
  assign y1567 = n7153 ;
  assign y1568 = ~1'b0 ;
  assign y1569 = n7157 ;
  assign y1570 = n7166 ;
  assign y1571 = ~1'b0 ;
  assign y1572 = ~1'b0 ;
  assign y1573 = n7175 ;
  assign y1574 = ~n7178 ;
  assign y1575 = ~n7184 ;
  assign y1576 = ~n7191 ;
  assign y1577 = ~n7196 ;
  assign y1578 = n7197 ;
  assign y1579 = ~n7206 ;
  assign y1580 = ~n7212 ;
  assign y1581 = n7223 ;
  assign y1582 = n7226 ;
  assign y1583 = n7230 ;
  assign y1584 = ~n7237 ;
  assign y1585 = ~1'b0 ;
  assign y1586 = n7240 ;
  assign y1587 = ~1'b0 ;
  assign y1588 = ~n7241 ;
  assign y1589 = n7247 ;
  assign y1590 = n7252 ;
  assign y1591 = n7261 ;
  assign y1592 = ~n7267 ;
  assign y1593 = ~n7269 ;
  assign y1594 = ~n7276 ;
  assign y1595 = ~1'b0 ;
  assign y1596 = n7279 ;
  assign y1597 = ~n7285 ;
  assign y1598 = n7286 ;
  assign y1599 = n7288 ;
  assign y1600 = ~n7298 ;
  assign y1601 = ~n7308 ;
  assign y1602 = ~n7313 ;
  assign y1603 = ~n7315 ;
  assign y1604 = n7320 ;
  assign y1605 = n7322 ;
  assign y1606 = n7324 ;
  assign y1607 = n7328 ;
  assign y1608 = ~n7335 ;
  assign y1609 = n7344 ;
  assign y1610 = ~n7346 ;
  assign y1611 = n7348 ;
  assign y1612 = ~n7349 ;
  assign y1613 = n7358 ;
  assign y1614 = n7361 ;
  assign y1615 = ~n7362 ;
  assign y1616 = ~n7368 ;
  assign y1617 = ~n7378 ;
  assign y1618 = n7380 ;
  assign y1619 = n7381 ;
  assign y1620 = ~1'b0 ;
  assign y1621 = ~n7390 ;
  assign y1622 = n7399 ;
  assign y1623 = n7402 ;
  assign y1624 = n7403 ;
  assign y1625 = n7405 ;
  assign y1626 = ~n7410 ;
  assign y1627 = ~1'b0 ;
  assign y1628 = ~n7411 ;
  assign y1629 = ~n7413 ;
  assign y1630 = n7414 ;
  assign y1631 = n7417 ;
  assign y1632 = ~n7424 ;
  assign y1633 = ~n7425 ;
  assign y1634 = n7447 ;
  assign y1635 = ~n7451 ;
  assign y1636 = ~n7455 ;
  assign y1637 = ~n7473 ;
  assign y1638 = n7477 ;
  assign y1639 = ~n7480 ;
  assign y1640 = ~n7481 ;
  assign y1641 = n7482 ;
  assign y1642 = ~n7487 ;
  assign y1643 = ~n7490 ;
  assign y1644 = ~1'b0 ;
  assign y1645 = ~n7491 ;
  assign y1646 = ~n7492 ;
  assign y1647 = ~n7503 ;
  assign y1648 = ~n7506 ;
  assign y1649 = n7524 ;
  assign y1650 = ~n7526 ;
  assign y1651 = ~n7528 ;
  assign y1652 = n7537 ;
  assign y1653 = ~n7540 ;
  assign y1654 = ~n7551 ;
  assign y1655 = n7564 ;
  assign y1656 = ~n7565 ;
  assign y1657 = ~1'b0 ;
  assign y1658 = ~1'b0 ;
  assign y1659 = ~1'b0 ;
  assign y1660 = ~n7569 ;
  assign y1661 = ~n7571 ;
  assign y1662 = ~n7573 ;
  assign y1663 = ~n7578 ;
  assign y1664 = ~1'b0 ;
  assign y1665 = ~n7586 ;
  assign y1666 = ~n7598 ;
  assign y1667 = n7600 ;
  assign y1668 = ~1'b0 ;
  assign y1669 = ~n7605 ;
  assign y1670 = n7606 ;
  assign y1671 = ~n7611 ;
  assign y1672 = ~n7612 ;
  assign y1673 = n7618 ;
  assign y1674 = ~n7622 ;
  assign y1675 = ~n7624 ;
  assign y1676 = n7636 ;
  assign y1677 = n7639 ;
  assign y1678 = n4888 ;
  assign y1679 = ~n7642 ;
  assign y1680 = ~1'b0 ;
  assign y1681 = ~n7643 ;
  assign y1682 = n7647 ;
  assign y1683 = n7648 ;
  assign y1684 = ~n7649 ;
  assign y1685 = n7656 ;
  assign y1686 = ~n7659 ;
  assign y1687 = ~1'b0 ;
  assign y1688 = n7663 ;
  assign y1689 = ~n7665 ;
  assign y1690 = ~n7670 ;
  assign y1691 = n7672 ;
  assign y1692 = n7674 ;
  assign y1693 = n7681 ;
  assign y1694 = ~n7694 ;
  assign y1695 = n7707 ;
  assign y1696 = ~n7708 ;
  assign y1697 = ~1'b0 ;
  assign y1698 = ~n7712 ;
  assign y1699 = n7713 ;
  assign y1700 = n7716 ;
  assign y1701 = n7718 ;
  assign y1702 = ~1'b0 ;
  assign y1703 = ~n7720 ;
  assign y1704 = ~n7722 ;
  assign y1705 = ~n7729 ;
  assign y1706 = ~1'b0 ;
  assign y1707 = ~1'b0 ;
  assign y1708 = ~n7730 ;
  assign y1709 = ~n7732 ;
  assign y1710 = n7750 ;
  assign y1711 = n7768 ;
  assign y1712 = ~1'b0 ;
  assign y1713 = ~n7770 ;
  assign y1714 = n7774 ;
  assign y1715 = ~n7776 ;
  assign y1716 = ~n7781 ;
  assign y1717 = n7786 ;
  assign y1718 = ~n7790 ;
  assign y1719 = ~n7796 ;
  assign y1720 = ~n7817 ;
  assign y1721 = n7820 ;
  assign y1722 = n7823 ;
  assign y1723 = n7832 ;
  assign y1724 = n7843 ;
  assign y1725 = ~n7850 ;
  assign y1726 = n7860 ;
  assign y1727 = n7865 ;
  assign y1728 = n7870 ;
  assign y1729 = ~n7871 ;
  assign y1730 = ~n7879 ;
  assign y1731 = ~n7881 ;
  assign y1732 = n7884 ;
  assign y1733 = n7885 ;
  assign y1734 = ~n7887 ;
  assign y1735 = ~n7897 ;
  assign y1736 = n7898 ;
  assign y1737 = ~n7909 ;
  assign y1738 = ~n7915 ;
  assign y1739 = n7918 ;
  assign y1740 = ~n7919 ;
  assign y1741 = n7924 ;
  assign y1742 = ~n7926 ;
  assign y1743 = ~1'b0 ;
  assign y1744 = n7930 ;
  assign y1745 = n7931 ;
  assign y1746 = ~n7932 ;
  assign y1747 = n7939 ;
  assign y1748 = ~n7946 ;
  assign y1749 = n7949 ;
  assign y1750 = ~n7960 ;
  assign y1751 = n7965 ;
  assign y1752 = ~n7973 ;
  assign y1753 = n7974 ;
  assign y1754 = ~n7975 ;
  assign y1755 = n7976 ;
  assign y1756 = n7978 ;
  assign y1757 = n7980 ;
  assign y1758 = ~n7985 ;
  assign y1759 = n7999 ;
  assign y1760 = ~n8001 ;
  assign y1761 = n8003 ;
  assign y1762 = n8008 ;
  assign y1763 = n8014 ;
  assign y1764 = ~n8026 ;
  assign y1765 = n6495 ;
  assign y1766 = ~n8027 ;
  assign y1767 = ~n8039 ;
  assign y1768 = ~n8041 ;
  assign y1769 = n8043 ;
  assign y1770 = ~1'b0 ;
  assign y1771 = ~n8046 ;
  assign y1772 = n8053 ;
  assign y1773 = n8056 ;
  assign y1774 = ~n8059 ;
  assign y1775 = ~n8063 ;
  assign y1776 = ~n8065 ;
  assign y1777 = n8069 ;
  assign y1778 = n8089 ;
  assign y1779 = ~n8098 ;
  assign y1780 = n8100 ;
  assign y1781 = n8103 ;
  assign y1782 = ~n8107 ;
  assign y1783 = n8108 ;
  assign y1784 = ~n8113 ;
  assign y1785 = ~n8114 ;
  assign y1786 = ~n8117 ;
  assign y1787 = ~1'b0 ;
  assign y1788 = ~n8118 ;
  assign y1789 = ~n8128 ;
  assign y1790 = n8129 ;
  assign y1791 = n8130 ;
  assign y1792 = n8136 ;
  assign y1793 = ~n8138 ;
  assign y1794 = ~n8145 ;
  assign y1795 = n8148 ;
  assign y1796 = ~n8155 ;
  assign y1797 = n8157 ;
  assign y1798 = n8158 ;
  assign y1799 = n8169 ;
  assign y1800 = ~1'b0 ;
  assign y1801 = ~n8172 ;
  assign y1802 = n8175 ;
  assign y1803 = n8179 ;
  assign y1804 = ~n8180 ;
  assign y1805 = n8185 ;
  assign y1806 = ~n8189 ;
  assign y1807 = n8202 ;
  assign y1808 = ~n8216 ;
  assign y1809 = ~n8217 ;
  assign y1810 = n8220 ;
  assign y1811 = ~n8224 ;
  assign y1812 = ~1'b0 ;
  assign y1813 = n8227 ;
  assign y1814 = ~n8238 ;
  assign y1815 = n8248 ;
  assign y1816 = ~n8254 ;
  assign y1817 = ~n8262 ;
  assign y1818 = n8265 ;
  assign y1819 = ~n8274 ;
  assign y1820 = ~1'b0 ;
  assign y1821 = ~n8275 ;
  assign y1822 = n8276 ;
  assign y1823 = n8279 ;
  assign y1824 = n8285 ;
  assign y1825 = n8287 ;
  assign y1826 = ~n8293 ;
  assign y1827 = n8297 ;
  assign y1828 = n8304 ;
  assign y1829 = n8306 ;
  assign y1830 = ~n8320 ;
  assign y1831 = ~n8321 ;
  assign y1832 = ~1'b0 ;
  assign y1833 = n8326 ;
  assign y1834 = n8327 ;
  assign y1835 = ~n8328 ;
  assign y1836 = ~n8332 ;
  assign y1837 = ~n8334 ;
  assign y1838 = n8349 ;
  assign y1839 = n8351 ;
  assign y1840 = n8356 ;
  assign y1841 = 1'b0 ;
  assign y1842 = ~1'b0 ;
  assign y1843 = ~n8357 ;
  assign y1844 = ~n8361 ;
  assign y1845 = n8364 ;
  assign y1846 = ~n8368 ;
  assign y1847 = n8370 ;
  assign y1848 = ~n8373 ;
  assign y1849 = ~n8377 ;
  assign y1850 = n8378 ;
  assign y1851 = n8380 ;
  assign y1852 = ~1'b0 ;
  assign y1853 = n8389 ;
  assign y1854 = n8396 ;
  assign y1855 = ~n8403 ;
  assign y1856 = ~n8405 ;
  assign y1857 = n8406 ;
  assign y1858 = n8415 ;
  assign y1859 = ~n8417 ;
  assign y1860 = ~n8418 ;
  assign y1861 = n8419 ;
  assign y1862 = n8424 ;
  assign y1863 = n8435 ;
  assign y1864 = n8451 ;
  assign y1865 = ~n8452 ;
  assign y1866 = n8457 ;
  assign y1867 = n8459 ;
  assign y1868 = ~n8460 ;
  assign y1869 = ~n8464 ;
  assign y1870 = n8467 ;
  assign y1871 = n8474 ;
  assign y1872 = ~n8477 ;
  assign y1873 = n8479 ;
  assign y1874 = n8486 ;
  assign y1875 = ~n8489 ;
  assign y1876 = ~n8499 ;
  assign y1877 = n8502 ;
  assign y1878 = ~n8505 ;
  assign y1879 = ~n8510 ;
  assign y1880 = ~n8515 ;
  assign y1881 = ~n8518 ;
  assign y1882 = ~n8523 ;
  assign y1883 = ~n8525 ;
  assign y1884 = n8526 ;
  assign y1885 = n8528 ;
  assign y1886 = ~n8537 ;
  assign y1887 = n8545 ;
  assign y1888 = ~n8548 ;
  assign y1889 = ~n8550 ;
  assign y1890 = ~n8553 ;
  assign y1891 = n8557 ;
  assign y1892 = ~1'b0 ;
  assign y1893 = n8563 ;
  assign y1894 = n8578 ;
  assign y1895 = ~n8582 ;
  assign y1896 = ~n8587 ;
  assign y1897 = ~n8598 ;
  assign y1898 = ~n8601 ;
  assign y1899 = n8610 ;
  assign y1900 = n8613 ;
  assign y1901 = n8616 ;
  assign y1902 = n8617 ;
  assign y1903 = n8626 ;
  assign y1904 = ~n8636 ;
  assign y1905 = ~1'b0 ;
  assign y1906 = ~n8637 ;
  assign y1907 = n8640 ;
  assign y1908 = ~n8642 ;
  assign y1909 = n8645 ;
  assign y1910 = n8646 ;
  assign y1911 = n8647 ;
  assign y1912 = n8648 ;
  assign y1913 = ~n8653 ;
  assign y1914 = n8657 ;
  assign y1915 = n8661 ;
  assign y1916 = n8664 ;
  assign y1917 = ~n8667 ;
  assign y1918 = n8674 ;
  assign y1919 = n8675 ;
  assign y1920 = ~1'b0 ;
  assign y1921 = ~n8678 ;
  assign y1922 = ~n8682 ;
  assign y1923 = n8683 ;
  assign y1924 = n8684 ;
  assign y1925 = n8685 ;
  assign y1926 = ~n8687 ;
  assign y1927 = n8690 ;
  assign y1928 = n8700 ;
  assign y1929 = n8706 ;
  assign y1930 = ~1'b0 ;
  assign y1931 = ~1'b0 ;
  assign y1932 = n8707 ;
  assign y1933 = ~n8708 ;
  assign y1934 = n8712 ;
  assign y1935 = ~1'b0 ;
  assign y1936 = ~n8714 ;
  assign y1937 = ~1'b0 ;
  assign y1938 = n8719 ;
  assign y1939 = n8723 ;
  assign y1940 = n8725 ;
  assign y1941 = ~1'b0 ;
  assign y1942 = n8726 ;
  assign y1943 = n8728 ;
  assign y1944 = n8732 ;
  assign y1945 = ~n8735 ;
  assign y1946 = ~n8743 ;
  assign y1947 = n8757 ;
  assign y1948 = ~1'b0 ;
  assign y1949 = ~n8762 ;
  assign y1950 = n8767 ;
  assign y1951 = n8772 ;
  assign y1952 = ~n8773 ;
  assign y1953 = ~n8778 ;
  assign y1954 = ~n8782 ;
  assign y1955 = ~1'b0 ;
  assign y1956 = n8783 ;
  assign y1957 = ~n8787 ;
  assign y1958 = n8795 ;
  assign y1959 = ~n8798 ;
  assign y1960 = ~n8799 ;
  assign y1961 = n8800 ;
  assign y1962 = ~1'b0 ;
  assign y1963 = ~n8805 ;
  assign y1964 = n8809 ;
  assign y1965 = ~n8814 ;
  assign y1966 = n8818 ;
  assign y1967 = n8830 ;
  assign y1968 = n8832 ;
  assign y1969 = ~n8836 ;
  assign y1970 = ~n8841 ;
  assign y1971 = ~n8847 ;
  assign y1972 = ~n8850 ;
  assign y1973 = ~n8852 ;
  assign y1974 = n8857 ;
  assign y1975 = n8859 ;
  assign y1976 = ~n8863 ;
  assign y1977 = ~n8870 ;
  assign y1978 = ~n8873 ;
  assign y1979 = n8875 ;
  assign y1980 = n8880 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = n8882 ;
  assign y1983 = n8897 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = n8901 ;
  assign y1986 = ~n8902 ;
  assign y1987 = n8904 ;
  assign y1988 = ~n8907 ;
  assign y1989 = n8910 ;
  assign y1990 = ~n8911 ;
  assign y1991 = n8916 ;
  assign y1992 = ~n8922 ;
  assign y1993 = ~n8925 ;
  assign y1994 = ~1'b0 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = n8929 ;
  assign y1997 = n8933 ;
  assign y1998 = ~n8940 ;
  assign y1999 = ~n8942 ;
  assign y2000 = ~n8948 ;
  assign y2001 = n8954 ;
  assign y2002 = n8958 ;
  assign y2003 = ~n8959 ;
  assign y2004 = n8960 ;
  assign y2005 = n8961 ;
  assign y2006 = n8963 ;
  assign y2007 = ~1'b0 ;
  assign y2008 = n8964 ;
  assign y2009 = ~n8965 ;
  assign y2010 = n8968 ;
  assign y2011 = ~n8979 ;
  assign y2012 = n8980 ;
  assign y2013 = n8981 ;
  assign y2014 = n8985 ;
  assign y2015 = ~n8987 ;
  assign y2016 = ~n8991 ;
  assign y2017 = n8993 ;
  assign y2018 = n9000 ;
  assign y2019 = ~1'b0 ;
  assign y2020 = n9002 ;
  assign y2021 = ~n9004 ;
  assign y2022 = ~n9008 ;
  assign y2023 = n9013 ;
  assign y2024 = n9017 ;
  assign y2025 = ~n9022 ;
  assign y2026 = ~n9024 ;
  assign y2027 = ~1'b0 ;
  assign y2028 = ~n9027 ;
  assign y2029 = ~1'b0 ;
  assign y2030 = n9033 ;
  assign y2031 = n9038 ;
  assign y2032 = n9041 ;
  assign y2033 = ~1'b0 ;
  assign y2034 = n9046 ;
  assign y2035 = n9051 ;
  assign y2036 = ~n9069 ;
  assign y2037 = n9073 ;
  assign y2038 = ~1'b0 ;
  assign y2039 = ~n9082 ;
  assign y2040 = ~1'b0 ;
  assign y2041 = ~1'b0 ;
  assign y2042 = ~1'b0 ;
  assign y2043 = n9085 ;
  assign y2044 = n9087 ;
  assign y2045 = n9090 ;
  assign y2046 = ~n9091 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = ~n9099 ;
  assign y2049 = ~n9103 ;
  assign y2050 = ~n9110 ;
  assign y2051 = ~n9114 ;
  assign y2052 = ~1'b0 ;
  assign y2053 = ~n9118 ;
  assign y2054 = ~n9122 ;
  assign y2055 = ~1'b0 ;
  assign y2056 = ~n9127 ;
  assign y2057 = ~n9134 ;
  assign y2058 = n9136 ;
  assign y2059 = n9141 ;
  assign y2060 = ~n9142 ;
  assign y2061 = ~n9148 ;
  assign y2062 = ~n6584 ;
  assign y2063 = n9155 ;
  assign y2064 = ~n9160 ;
  assign y2065 = n9166 ;
  assign y2066 = ~n9169 ;
  assign y2067 = n9180 ;
  assign y2068 = ~n9182 ;
  assign y2069 = ~n9183 ;
  assign y2070 = n9189 ;
  assign y2071 = ~n9196 ;
  assign y2072 = n9204 ;
  assign y2073 = ~n9209 ;
  assign y2074 = n9210 ;
  assign y2075 = ~n9213 ;
  assign y2076 = ~n9218 ;
  assign y2077 = ~n9226 ;
  assign y2078 = n9234 ;
  assign y2079 = n9235 ;
  assign y2080 = n9236 ;
  assign y2081 = n9252 ;
  assign y2082 = ~n9264 ;
  assign y2083 = ~1'b0 ;
  assign y2084 = ~n9266 ;
  assign y2085 = ~1'b0 ;
  assign y2086 = n9281 ;
  assign y2087 = ~n9282 ;
  assign y2088 = n9292 ;
  assign y2089 = ~1'b0 ;
  assign y2090 = ~1'b0 ;
  assign y2091 = ~n9297 ;
  assign y2092 = n9299 ;
  assign y2093 = n9304 ;
  assign y2094 = ~n9305 ;
  assign y2095 = ~n9307 ;
  assign y2096 = ~n9311 ;
  assign y2097 = ~n9313 ;
  assign y2098 = ~n9324 ;
  assign y2099 = ~n9325 ;
  assign y2100 = ~n9332 ;
  assign y2101 = ~n9333 ;
  assign y2102 = ~n9334 ;
  assign y2103 = n9339 ;
  assign y2104 = ~n9340 ;
  assign y2105 = ~n9344 ;
  assign y2106 = ~1'b0 ;
  assign y2107 = ~n9345 ;
  assign y2108 = ~n9347 ;
  assign y2109 = n9348 ;
  assign y2110 = n9350 ;
  assign y2111 = n9353 ;
  assign y2112 = ~n9357 ;
  assign y2113 = n9358 ;
  assign y2114 = n9366 ;
  assign y2115 = ~n9372 ;
  assign y2116 = ~n9375 ;
  assign y2117 = ~n9377 ;
  assign y2118 = n9378 ;
  assign y2119 = ~1'b0 ;
  assign y2120 = ~1'b0 ;
  assign y2121 = n9379 ;
  assign y2122 = n9381 ;
  assign y2123 = ~1'b0 ;
  assign y2124 = ~n9384 ;
  assign y2125 = ~n9385 ;
  assign y2126 = ~n9394 ;
  assign y2127 = ~n9397 ;
  assign y2128 = ~n9399 ;
  assign y2129 = ~n9411 ;
  assign y2130 = ~n9414 ;
  assign y2131 = ~n9417 ;
  assign y2132 = ~1'b0 ;
  assign y2133 = ~1'b0 ;
  assign y2134 = ~n9418 ;
  assign y2135 = ~n9428 ;
  assign y2136 = n9432 ;
  assign y2137 = ~n9438 ;
  assign y2138 = n9442 ;
  assign y2139 = ~n9453 ;
  assign y2140 = n9455 ;
  assign y2141 = ~n9465 ;
  assign y2142 = n9485 ;
  assign y2143 = ~n9491 ;
  assign y2144 = ~n9495 ;
  assign y2145 = n9500 ;
  assign y2146 = n9509 ;
  assign y2147 = ~n9515 ;
  assign y2148 = ~n9518 ;
  assign y2149 = n9520 ;
  assign y2150 = ~n9527 ;
  assign y2151 = ~n9529 ;
  assign y2152 = ~n9541 ;
  assign y2153 = n9547 ;
  assign y2154 = n9552 ;
  assign y2155 = ~n9554 ;
  assign y2156 = n9557 ;
  assign y2157 = ~n9564 ;
  assign y2158 = n9570 ;
  assign y2159 = ~n9575 ;
  assign y2160 = ~n9576 ;
  assign y2161 = n9580 ;
  assign y2162 = n9589 ;
  assign y2163 = n9596 ;
  assign y2164 = n9603 ;
  assign y2165 = n9606 ;
  assign y2166 = n9610 ;
  assign y2167 = n9616 ;
  assign y2168 = ~n9628 ;
  assign y2169 = ~n9639 ;
  assign y2170 = ~n9644 ;
  assign y2171 = n9645 ;
  assign y2172 = ~n9650 ;
  assign y2173 = ~n9655 ;
  assign y2174 = n9656 ;
  assign y2175 = ~n9663 ;
  assign y2176 = ~1'b0 ;
  assign y2177 = ~n9667 ;
  assign y2178 = n9668 ;
  assign y2179 = ~n9669 ;
  assign y2180 = n9675 ;
  assign y2181 = ~n9679 ;
  assign y2182 = ~n9681 ;
  assign y2183 = ~1'b0 ;
  assign y2184 = n9692 ;
  assign y2185 = n9695 ;
  assign y2186 = n9698 ;
  assign y2187 = ~n9700 ;
  assign y2188 = n9712 ;
  assign y2189 = ~n9718 ;
  assign y2190 = n9721 ;
  assign y2191 = ~1'b0 ;
  assign y2192 = n9733 ;
  assign y2193 = ~n9735 ;
  assign y2194 = n9740 ;
  assign y2195 = ~n9743 ;
  assign y2196 = ~1'b0 ;
  assign y2197 = n9747 ;
  assign y2198 = n9754 ;
  assign y2199 = ~n9759 ;
  assign y2200 = ~n9761 ;
  assign y2201 = n9763 ;
  assign y2202 = ~n9772 ;
  assign y2203 = ~n9774 ;
  assign y2204 = ~n9777 ;
  assign y2205 = n9784 ;
  assign y2206 = ~1'b0 ;
  assign y2207 = ~n9789 ;
  assign y2208 = ~n9795 ;
  assign y2209 = ~n9796 ;
  assign y2210 = ~1'b0 ;
  assign y2211 = n9798 ;
  assign y2212 = n9799 ;
  assign y2213 = ~n9801 ;
  assign y2214 = ~1'b0 ;
  assign y2215 = n9804 ;
  assign y2216 = n9810 ;
  assign y2217 = n9816 ;
  assign y2218 = n9818 ;
  assign y2219 = n9820 ;
  assign y2220 = ~n9822 ;
  assign y2221 = ~n9823 ;
  assign y2222 = ~n9825 ;
  assign y2223 = ~n9828 ;
  assign y2224 = ~n9837 ;
  assign y2225 = ~n9843 ;
  assign y2226 = ~n9846 ;
  assign y2227 = ~n9847 ;
  assign y2228 = ~1'b0 ;
  assign y2229 = ~n9852 ;
  assign y2230 = ~n9858 ;
  assign y2231 = ~1'b0 ;
  assign y2232 = n9861 ;
  assign y2233 = n9864 ;
  assign y2234 = ~n9875 ;
  assign y2235 = n9878 ;
  assign y2236 = ~n9881 ;
  assign y2237 = ~n9882 ;
  assign y2238 = ~n9888 ;
  assign y2239 = n9893 ;
  assign y2240 = ~1'b0 ;
  assign y2241 = ~n9895 ;
  assign y2242 = ~n9904 ;
  assign y2243 = ~n9910 ;
  assign y2244 = n9914 ;
  assign y2245 = n9916 ;
  assign y2246 = ~1'b0 ;
  assign y2247 = ~1'b0 ;
  assign y2248 = n9923 ;
  assign y2249 = n9924 ;
  assign y2250 = ~n9927 ;
  assign y2251 = n9935 ;
  assign y2252 = ~n9940 ;
  assign y2253 = ~n9944 ;
  assign y2254 = ~n9959 ;
  assign y2255 = ~n9963 ;
  assign y2256 = n4435 ;
  assign y2257 = ~n9966 ;
  assign y2258 = ~n9968 ;
  assign y2259 = n9970 ;
  assign y2260 = ~1'b0 ;
  assign y2261 = n9977 ;
  assign y2262 = n9980 ;
  assign y2263 = ~n9983 ;
  assign y2264 = ~1'b0 ;
  assign y2265 = ~n9986 ;
  assign y2266 = n9989 ;
  assign y2267 = n9990 ;
  assign y2268 = ~n9991 ;
  assign y2269 = n9996 ;
  assign y2270 = n10005 ;
  assign y2271 = ~n10009 ;
  assign y2272 = n10011 ;
  assign y2273 = n10018 ;
  assign y2274 = ~n10022 ;
  assign y2275 = ~n10025 ;
  assign y2276 = ~n10027 ;
  assign y2277 = n10032 ;
  assign y2278 = ~n10034 ;
  assign y2279 = n10036 ;
  assign y2280 = n10045 ;
  assign y2281 = ~1'b0 ;
  assign y2282 = n10046 ;
  assign y2283 = n10051 ;
  assign y2284 = ~n10053 ;
  assign y2285 = n10056 ;
  assign y2286 = ~n10061 ;
  assign y2287 = n10068 ;
  assign y2288 = ~n10076 ;
  assign y2289 = n10082 ;
  assign y2290 = n10084 ;
  assign y2291 = n10089 ;
  assign y2292 = ~n10097 ;
  assign y2293 = n10099 ;
  assign y2294 = ~1'b0 ;
  assign y2295 = n10105 ;
  assign y2296 = n10107 ;
  assign y2297 = ~n10113 ;
  assign y2298 = ~1'b0 ;
  assign y2299 = ~n10126 ;
  assign y2300 = ~n1856 ;
  assign y2301 = ~n10130 ;
  assign y2302 = n10137 ;
  assign y2303 = ~n10139 ;
  assign y2304 = n10143 ;
  assign y2305 = n10144 ;
  assign y2306 = n10148 ;
  assign y2307 = ~n10156 ;
  assign y2308 = n10159 ;
  assign y2309 = n10164 ;
  assign y2310 = n10167 ;
  assign y2311 = ~n10169 ;
  assign y2312 = ~1'b0 ;
  assign y2313 = ~n10170 ;
  assign y2314 = ~n10172 ;
  assign y2315 = n10180 ;
  assign y2316 = n10186 ;
  assign y2317 = n10187 ;
  assign y2318 = n10209 ;
  assign y2319 = ~n10216 ;
  assign y2320 = ~n10218 ;
  assign y2321 = ~n10220 ;
  assign y2322 = n10227 ;
  assign y2323 = ~n2479 ;
  assign y2324 = ~n10230 ;
  assign y2325 = n10231 ;
  assign y2326 = ~1'b0 ;
  assign y2327 = n10233 ;
  assign y2328 = ~n10234 ;
  assign y2329 = ~n10236 ;
  assign y2330 = ~n10249 ;
  assign y2331 = ~n10250 ;
  assign y2332 = n10264 ;
  assign y2333 = ~n10268 ;
  assign y2334 = n10272 ;
  assign y2335 = n10279 ;
  assign y2336 = ~n10286 ;
  assign y2337 = n10287 ;
  assign y2338 = ~n10289 ;
  assign y2339 = n10292 ;
  assign y2340 = n10295 ;
  assign y2341 = n10297 ;
  assign y2342 = n10300 ;
  assign y2343 = ~n10302 ;
  assign y2344 = n10305 ;
  assign y2345 = n10308 ;
  assign y2346 = ~n10310 ;
  assign y2347 = n10321 ;
  assign y2348 = n10323 ;
  assign y2349 = n10327 ;
  assign y2350 = n10330 ;
  assign y2351 = ~n10334 ;
  assign y2352 = n10338 ;
  assign y2353 = ~n10340 ;
  assign y2354 = n10356 ;
  assign y2355 = ~n10360 ;
  assign y2356 = n10362 ;
  assign y2357 = ~n10366 ;
  assign y2358 = ~n10371 ;
  assign y2359 = ~n10375 ;
  assign y2360 = ~n10385 ;
  assign y2361 = n10388 ;
  assign y2362 = n10393 ;
  assign y2363 = n10395 ;
  assign y2364 = n10396 ;
  assign y2365 = n10400 ;
  assign y2366 = n10407 ;
  assign y2367 = ~n10408 ;
  assign y2368 = n10409 ;
  assign y2369 = n10414 ;
  assign y2370 = ~n10415 ;
  assign y2371 = n10417 ;
  assign y2372 = n10424 ;
  assign y2373 = n10426 ;
  assign y2374 = ~n10427 ;
  assign y2375 = ~n10431 ;
  assign y2376 = n10433 ;
  assign y2377 = ~n10435 ;
  assign y2378 = ~n10438 ;
  assign y2379 = ~1'b0 ;
  assign y2380 = ~n10439 ;
  assign y2381 = ~n10442 ;
  assign y2382 = ~n10450 ;
  assign y2383 = n10453 ;
  assign y2384 = n10457 ;
  assign y2385 = ~n10458 ;
  assign y2386 = ~1'b0 ;
  assign y2387 = n10462 ;
  assign y2388 = ~n10463 ;
  assign y2389 = ~n10464 ;
  assign y2390 = ~n10467 ;
  assign y2391 = n10472 ;
  assign y2392 = ~n10473 ;
  assign y2393 = ~n10476 ;
  assign y2394 = n10481 ;
  assign y2395 = ~n10483 ;
  assign y2396 = ~n10490 ;
  assign y2397 = n10491 ;
  assign y2398 = ~n10495 ;
  assign y2399 = ~n10496 ;
  assign y2400 = ~n10499 ;
  assign y2401 = n10503 ;
  assign y2402 = ~n10507 ;
  assign y2403 = ~n10516 ;
  assign y2404 = n10518 ;
  assign y2405 = n10519 ;
  assign y2406 = ~n10527 ;
  assign y2407 = n10529 ;
  assign y2408 = n10530 ;
  assign y2409 = n10534 ;
  assign y2410 = n10536 ;
  assign y2411 = n10539 ;
  assign y2412 = ~1'b0 ;
  assign y2413 = ~n10540 ;
  assign y2414 = ~n10544 ;
  assign y2415 = n10550 ;
  assign y2416 = n10552 ;
  assign y2417 = ~n10556 ;
  assign y2418 = ~n10558 ;
  assign y2419 = ~n10564 ;
  assign y2420 = n10565 ;
  assign y2421 = ~n10569 ;
  assign y2422 = ~1'b0 ;
  assign y2423 = n10570 ;
  assign y2424 = ~n10572 ;
  assign y2425 = ~1'b0 ;
  assign y2426 = n10576 ;
  assign y2427 = n10580 ;
  assign y2428 = ~n10588 ;
  assign y2429 = n10606 ;
  assign y2430 = ~n10611 ;
  assign y2431 = n10614 ;
  assign y2432 = n10621 ;
  assign y2433 = n10628 ;
  assign y2434 = ~n10631 ;
  assign y2435 = ~n10633 ;
  assign y2436 = ~n10637 ;
  assign y2437 = ~n10638 ;
  assign y2438 = n10643 ;
  assign y2439 = ~n10644 ;
  assign y2440 = ~n10648 ;
  assign y2441 = n10650 ;
  assign y2442 = ~1'b0 ;
  assign y2443 = n10658 ;
  assign y2444 = n10660 ;
  assign y2445 = ~n10661 ;
  assign y2446 = ~1'b0 ;
  assign y2447 = n10663 ;
  assign y2448 = ~n10668 ;
  assign y2449 = ~n10677 ;
  assign y2450 = ~n10679 ;
  assign y2451 = ~n10683 ;
  assign y2452 = ~n10685 ;
  assign y2453 = n10686 ;
  assign y2454 = n10692 ;
  assign y2455 = n10694 ;
  assign y2456 = ~n10704 ;
  assign y2457 = ~n10709 ;
  assign y2458 = ~n10713 ;
  assign y2459 = ~n10716 ;
  assign y2460 = ~n10722 ;
  assign y2461 = ~n10737 ;
  assign y2462 = ~n10738 ;
  assign y2463 = ~n10740 ;
  assign y2464 = ~1'b0 ;
  assign y2465 = ~n10742 ;
  assign y2466 = ~n10743 ;
  assign y2467 = ~n10749 ;
  assign y2468 = ~n10751 ;
  assign y2469 = ~n10753 ;
  assign y2470 = ~n10757 ;
  assign y2471 = ~1'b0 ;
  assign y2472 = n10759 ;
  assign y2473 = n10762 ;
  assign y2474 = ~1'b0 ;
  assign y2475 = ~n10763 ;
  assign y2476 = ~1'b0 ;
  assign y2477 = ~n10770 ;
  assign y2478 = ~n10775 ;
  assign y2479 = ~n10780 ;
  assign y2480 = n10783 ;
  assign y2481 = ~n10787 ;
  assign y2482 = n10790 ;
  assign y2483 = n10792 ;
  assign y2484 = n10794 ;
  assign y2485 = n10797 ;
  assign y2486 = ~n10798 ;
  assign y2487 = n10799 ;
  assign y2488 = ~n10800 ;
  assign y2489 = n10802 ;
  assign y2490 = n10804 ;
  assign y2491 = ~n10811 ;
  assign y2492 = ~n10813 ;
  assign y2493 = n10822 ;
  assign y2494 = ~n10827 ;
  assign y2495 = n10833 ;
  assign y2496 = ~n10834 ;
  assign y2497 = ~n10837 ;
  assign y2498 = ~1'b0 ;
  assign y2499 = ~n10840 ;
  assign y2500 = ~n10841 ;
  assign y2501 = n10847 ;
  assign y2502 = n10850 ;
  assign y2503 = n10853 ;
  assign y2504 = ~n10862 ;
  assign y2505 = n10869 ;
  assign y2506 = ~n10871 ;
  assign y2507 = ~n10873 ;
  assign y2508 = n10874 ;
  assign y2509 = ~n10881 ;
  assign y2510 = ~n10885 ;
  assign y2511 = ~n10895 ;
  assign y2512 = ~n10896 ;
  assign y2513 = n10898 ;
  assign y2514 = ~1'b0 ;
  assign y2515 = ~n588 ;
  assign y2516 = ~1'b0 ;
  assign y2517 = ~n10905 ;
  assign y2518 = ~n10908 ;
  assign y2519 = n10911 ;
  assign y2520 = n10914 ;
  assign y2521 = n10922 ;
  assign y2522 = ~n10927 ;
  assign y2523 = ~n10931 ;
  assign y2524 = n10935 ;
  assign y2525 = n10944 ;
  assign y2526 = ~1'b0 ;
  assign y2527 = ~1'b0 ;
  assign y2528 = n10947 ;
  assign y2529 = n10951 ;
  assign y2530 = n10958 ;
  assign y2531 = n10964 ;
  assign y2532 = n10967 ;
  assign y2533 = ~n10968 ;
  assign y2534 = ~n10970 ;
  assign y2535 = ~n10971 ;
  assign y2536 = ~1'b0 ;
  assign y2537 = n10982 ;
  assign y2538 = ~n10992 ;
  assign y2539 = ~n10994 ;
  assign y2540 = ~n10999 ;
  assign y2541 = n11000 ;
  assign y2542 = ~n11004 ;
  assign y2543 = ~1'b0 ;
  assign y2544 = n11005 ;
  assign y2545 = ~n11008 ;
  assign y2546 = ~n11011 ;
  assign y2547 = ~n11014 ;
  assign y2548 = n11018 ;
  assign y2549 = ~n11021 ;
  assign y2550 = ~n11027 ;
  assign y2551 = ~1'b0 ;
  assign y2552 = ~n11031 ;
  assign y2553 = ~1'b0 ;
  assign y2554 = ~n11036 ;
  assign y2555 = n11043 ;
  assign y2556 = ~n11044 ;
  assign y2557 = ~n11048 ;
  assign y2558 = ~1'b0 ;
  assign y2559 = n11049 ;
  assign y2560 = n11053 ;
  assign y2561 = n11056 ;
  assign y2562 = ~n11057 ;
  assign y2563 = n11060 ;
  assign y2564 = ~n11070 ;
  assign y2565 = n11071 ;
  assign y2566 = n11073 ;
  assign y2567 = n11081 ;
  assign y2568 = n11084 ;
  assign y2569 = ~n11088 ;
  assign y2570 = n11097 ;
  assign y2571 = ~n11098 ;
  assign y2572 = n11099 ;
  assign y2573 = n11101 ;
  assign y2574 = ~n11104 ;
  assign y2575 = n5170 ;
  assign y2576 = n11114 ;
  assign y2577 = ~n11117 ;
  assign y2578 = ~n11123 ;
  assign y2579 = n11124 ;
  assign y2580 = n11130 ;
  assign y2581 = n11137 ;
  assign y2582 = ~n11141 ;
  assign y2583 = ~n11145 ;
  assign y2584 = ~n11149 ;
  assign y2585 = ~n11154 ;
  assign y2586 = n11175 ;
  assign y2587 = ~n11176 ;
  assign y2588 = ~n11183 ;
  assign y2589 = ~n11184 ;
  assign y2590 = ~n11186 ;
  assign y2591 = ~n11188 ;
  assign y2592 = n11192 ;
  assign y2593 = ~n11193 ;
  assign y2594 = ~n11195 ;
  assign y2595 = n11196 ;
  assign y2596 = ~n11201 ;
  assign y2597 = ~n11209 ;
  assign y2598 = n11214 ;
  assign y2599 = n11217 ;
  assign y2600 = n11221 ;
  assign y2601 = ~1'b0 ;
  assign y2602 = n11224 ;
  assign y2603 = ~n11233 ;
  assign y2604 = ~n11237 ;
  assign y2605 = n11238 ;
  assign y2606 = ~n11240 ;
  assign y2607 = ~n11242 ;
  assign y2608 = n11244 ;
  assign y2609 = ~n11248 ;
  assign y2610 = ~n11256 ;
  assign y2611 = ~n11261 ;
  assign y2612 = ~n11265 ;
  assign y2613 = ~n11269 ;
  assign y2614 = ~n11279 ;
  assign y2615 = ~n11281 ;
  assign y2616 = ~n11288 ;
  assign y2617 = n11290 ;
  assign y2618 = ~n11293 ;
  assign y2619 = n11294 ;
  assign y2620 = n11298 ;
  assign y2621 = n11299 ;
  assign y2622 = ~n11301 ;
  assign y2623 = n11302 ;
  assign y2624 = ~n11307 ;
  assign y2625 = ~n11309 ;
  assign y2626 = n11315 ;
  assign y2627 = ~n11324 ;
  assign y2628 = n11332 ;
  assign y2629 = ~1'b0 ;
  assign y2630 = ~n11333 ;
  assign y2631 = ~n11335 ;
  assign y2632 = n11344 ;
  assign y2633 = n11347 ;
  assign y2634 = ~n7596 ;
  assign y2635 = n11358 ;
  assign y2636 = n11367 ;
  assign y2637 = ~n11371 ;
  assign y2638 = n11379 ;
  assign y2639 = n11384 ;
  assign y2640 = n11386 ;
  assign y2641 = n11393 ;
  assign y2642 = n11396 ;
  assign y2643 = n11399 ;
  assign y2644 = ~n11400 ;
  assign y2645 = n11401 ;
  assign y2646 = ~n11402 ;
  assign y2647 = ~n11403 ;
  assign y2648 = ~n11408 ;
  assign y2649 = n11412 ;
  assign y2650 = ~1'b0 ;
  assign y2651 = n11416 ;
  assign y2652 = ~n11417 ;
  assign y2653 = ~n11421 ;
  assign y2654 = ~n997 ;
  assign y2655 = ~n11423 ;
  assign y2656 = ~n11425 ;
  assign y2657 = ~n11434 ;
  assign y2658 = ~n11436 ;
  assign y2659 = ~1'b0 ;
  assign y2660 = ~n11439 ;
  assign y2661 = ~n11443 ;
  assign y2662 = ~n11446 ;
  assign y2663 = ~1'b0 ;
  assign y2664 = n11451 ;
  assign y2665 = n11455 ;
  assign y2666 = ~n11456 ;
  assign y2667 = ~n11461 ;
  assign y2668 = ~n11466 ;
  assign y2669 = ~n11471 ;
  assign y2670 = ~n11475 ;
  assign y2671 = n11479 ;
  assign y2672 = ~n11482 ;
  assign y2673 = n11491 ;
  assign y2674 = n11493 ;
  assign y2675 = n11497 ;
  assign y2676 = ~n11502 ;
  assign y2677 = n11510 ;
  assign y2678 = ~n11513 ;
  assign y2679 = ~1'b0 ;
  assign y2680 = n11520 ;
  assign y2681 = n11522 ;
  assign y2682 = n11523 ;
  assign y2683 = ~n11532 ;
  assign y2684 = n11534 ;
  assign y2685 = ~n11539 ;
  assign y2686 = ~n11547 ;
  assign y2687 = n11549 ;
  assign y2688 = ~n11552 ;
  assign y2689 = ~n11554 ;
  assign y2690 = ~1'b0 ;
  assign y2691 = n11556 ;
  assign y2692 = ~n11559 ;
  assign y2693 = ~n11562 ;
  assign y2694 = n11566 ;
  assign y2695 = ~n11572 ;
  assign y2696 = n11573 ;
  assign y2697 = n11578 ;
  assign y2698 = ~n4893 ;
  assign y2699 = n11582 ;
  assign y2700 = ~n11587 ;
  assign y2701 = ~1'b0 ;
  assign y2702 = n11595 ;
  assign y2703 = ~n11603 ;
  assign y2704 = ~n11606 ;
  assign y2705 = n11610 ;
  assign y2706 = ~n11614 ;
  assign y2707 = ~n11615 ;
  assign y2708 = n11619 ;
  assign y2709 = n11622 ;
  assign y2710 = n11624 ;
  assign y2711 = ~n11628 ;
  assign y2712 = n11640 ;
  assign y2713 = ~n11643 ;
  assign y2714 = ~n11644 ;
  assign y2715 = ~n11648 ;
  assign y2716 = n11652 ;
  assign y2717 = n11661 ;
  assign y2718 = n11663 ;
  assign y2719 = n11666 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = n11668 ;
  assign y2722 = ~n11670 ;
  assign y2723 = ~n11672 ;
  assign y2724 = ~n11673 ;
  assign y2725 = n10900 ;
  assign y2726 = n11678 ;
  assign y2727 = ~n11682 ;
  assign y2728 = n11684 ;
  assign y2729 = n11686 ;
  assign y2730 = ~n11690 ;
  assign y2731 = n11692 ;
  assign y2732 = n11703 ;
  assign y2733 = n11709 ;
  assign y2734 = n11710 ;
  assign y2735 = n11712 ;
  assign y2736 = ~1'b0 ;
  assign y2737 = ~n11719 ;
  assign y2738 = n11724 ;
  assign y2739 = n11726 ;
  assign y2740 = ~n11730 ;
  assign y2741 = ~n11732 ;
  assign y2742 = ~n11736 ;
  assign y2743 = n11737 ;
  assign y2744 = n11740 ;
  assign y2745 = ~n11744 ;
  assign y2746 = n11748 ;
  assign y2747 = n11750 ;
  assign y2748 = ~n11755 ;
  assign y2749 = n11759 ;
  assign y2750 = ~1'b0 ;
  assign y2751 = ~n11761 ;
  assign y2752 = ~n11766 ;
  assign y2753 = n11768 ;
  assign y2754 = n11778 ;
  assign y2755 = ~n11784 ;
  assign y2756 = ~n11787 ;
  assign y2757 = n11790 ;
  assign y2758 = ~n11793 ;
  assign y2759 = ~1'b0 ;
  assign y2760 = ~n11801 ;
  assign y2761 = ~n11804 ;
  assign y2762 = n11808 ;
  assign y2763 = ~n11812 ;
  assign y2764 = n11816 ;
  assign y2765 = ~n11822 ;
  assign y2766 = n11826 ;
  assign y2767 = n11835 ;
  assign y2768 = ~n11842 ;
  assign y2769 = ~1'b0 ;
  assign y2770 = ~n11843 ;
  assign y2771 = ~n11851 ;
  assign y2772 = ~1'b0 ;
  assign y2773 = ~n11854 ;
  assign y2774 = n11860 ;
  assign y2775 = n11865 ;
  assign y2776 = ~1'b0 ;
  assign y2777 = n11869 ;
  assign y2778 = ~n11874 ;
  assign y2779 = ~n11877 ;
  assign y2780 = ~1'b0 ;
  assign y2781 = n11879 ;
  assign y2782 = n11887 ;
  assign y2783 = ~1'b0 ;
  assign y2784 = ~n11890 ;
  assign y2785 = ~n11891 ;
  assign y2786 = n11893 ;
  assign y2787 = ~1'b0 ;
  assign y2788 = ~n11905 ;
  assign y2789 = n11911 ;
  assign y2790 = ~n11912 ;
  assign y2791 = n11913 ;
  assign y2792 = n11923 ;
  assign y2793 = ~n11928 ;
  assign y2794 = n11932 ;
  assign y2795 = ~n11943 ;
  assign y2796 = ~n11944 ;
  assign y2797 = ~1'b0 ;
  assign y2798 = ~n11950 ;
  assign y2799 = ~n11952 ;
  assign y2800 = n11953 ;
  assign y2801 = ~1'b0 ;
  assign y2802 = n11955 ;
  assign y2803 = ~n11962 ;
  assign y2804 = n11967 ;
  assign y2805 = ~n11968 ;
  assign y2806 = n11971 ;
  assign y2807 = ~n11972 ;
  assign y2808 = ~1'b0 ;
  assign y2809 = ~1'b0 ;
  assign y2810 = n11973 ;
  assign y2811 = n11975 ;
  assign y2812 = n11977 ;
  assign y2813 = ~n11980 ;
  assign y2814 = n11983 ;
  assign y2815 = ~n11987 ;
  assign y2816 = n11997 ;
  assign y2817 = n11999 ;
  assign y2818 = n12001 ;
  assign y2819 = n12007 ;
  assign y2820 = n12009 ;
  assign y2821 = ~n12017 ;
  assign y2822 = ~n12019 ;
  assign y2823 = ~n12021 ;
  assign y2824 = ~n12026 ;
  assign y2825 = n12031 ;
  assign y2826 = ~1'b0 ;
  assign y2827 = n12036 ;
  assign y2828 = ~n12037 ;
  assign y2829 = n12045 ;
  assign y2830 = n12052 ;
  assign y2831 = n12059 ;
  assign y2832 = n12061 ;
  assign y2833 = ~1'b0 ;
  assign y2834 = ~n12064 ;
  assign y2835 = n12066 ;
  assign y2836 = ~n12067 ;
  assign y2837 = n12080 ;
  assign y2838 = n12083 ;
  assign y2839 = ~n12086 ;
  assign y2840 = n12087 ;
  assign y2841 = n12088 ;
  assign y2842 = ~1'b0 ;
  assign y2843 = ~n12092 ;
  assign y2844 = n12102 ;
  assign y2845 = n12107 ;
  assign y2846 = ~1'b0 ;
  assign y2847 = ~n12112 ;
  assign y2848 = ~n12115 ;
  assign y2849 = ~n12116 ;
  assign y2850 = ~n12117 ;
  assign y2851 = n12120 ;
  assign y2852 = n12121 ;
  assign y2853 = n12123 ;
  assign y2854 = ~n12135 ;
  assign y2855 = ~n12136 ;
  assign y2856 = ~n12137 ;
  assign y2857 = ~n12138 ;
  assign y2858 = ~1'b0 ;
  assign y2859 = ~n3658 ;
  assign y2860 = n12145 ;
  assign y2861 = n12147 ;
  assign y2862 = n12153 ;
  assign y2863 = n12155 ;
  assign y2864 = n12159 ;
  assign y2865 = ~n12164 ;
  assign y2866 = ~n12167 ;
  assign y2867 = n12169 ;
  assign y2868 = ~1'b0 ;
  assign y2869 = ~1'b0 ;
  assign y2870 = ~n12170 ;
  assign y2871 = n12175 ;
  assign y2872 = ~n12178 ;
  assign y2873 = ~n12180 ;
  assign y2874 = n12184 ;
  assign y2875 = n12194 ;
  assign y2876 = ~n12210 ;
  assign y2877 = ~1'b0 ;
  assign y2878 = n12212 ;
  assign y2879 = ~n12214 ;
  assign y2880 = ~n12216 ;
  assign y2881 = ~n12221 ;
  assign y2882 = ~n12232 ;
  assign y2883 = n12236 ;
  assign y2884 = ~n12241 ;
  assign y2885 = n12246 ;
  assign y2886 = n12253 ;
  assign y2887 = ~n12254 ;
  assign y2888 = n12255 ;
  assign y2889 = ~n12268 ;
  assign y2890 = n12269 ;
  assign y2891 = ~n12274 ;
  assign y2892 = ~n12276 ;
  assign y2893 = ~n6505 ;
  assign y2894 = n12280 ;
  assign y2895 = n12282 ;
  assign y2896 = n12284 ;
  assign y2897 = n12285 ;
  assign y2898 = n12292 ;
  assign y2899 = ~1'b0 ;
  assign y2900 = ~n12294 ;
  assign y2901 = ~n12299 ;
  assign y2902 = ~n12301 ;
  assign y2903 = n12302 ;
  assign y2904 = n12304 ;
  assign y2905 = n12309 ;
  assign y2906 = ~n12319 ;
  assign y2907 = n12321 ;
  assign y2908 = n12323 ;
  assign y2909 = ~n12330 ;
  assign y2910 = ~n12340 ;
  assign y2911 = n12345 ;
  assign y2912 = ~1'b0 ;
  assign y2913 = ~n12355 ;
  assign y2914 = ~n12366 ;
  assign y2915 = n12368 ;
  assign y2916 = ~n12369 ;
  assign y2917 = ~n12371 ;
  assign y2918 = ~n12378 ;
  assign y2919 = ~n12383 ;
  assign y2920 = ~n3460 ;
  assign y2921 = ~n12388 ;
  assign y2922 = n12389 ;
  assign y2923 = ~1'b0 ;
  assign y2924 = n12390 ;
  assign y2925 = ~n12391 ;
  assign y2926 = n12395 ;
  assign y2927 = ~n12402 ;
  assign y2928 = ~1'b0 ;
  assign y2929 = n12406 ;
  assign y2930 = ~n12410 ;
  assign y2931 = ~n12411 ;
  assign y2932 = n12415 ;
  assign y2933 = ~n12417 ;
  assign y2934 = ~n12431 ;
  assign y2935 = n12436 ;
  assign y2936 = n12438 ;
  assign y2937 = ~1'b0 ;
  assign y2938 = ~n12441 ;
  assign y2939 = ~n12443 ;
  assign y2940 = n12445 ;
  assign y2941 = ~n12446 ;
  assign y2942 = n12453 ;
  assign y2943 = ~1'b0 ;
  assign y2944 = n12454 ;
  assign y2945 = ~n12460 ;
  assign y2946 = ~n12461 ;
  assign y2947 = ~1'b0 ;
  assign y2948 = ~1'b0 ;
  assign y2949 = n12466 ;
  assign y2950 = ~n12468 ;
  assign y2951 = n12470 ;
  assign y2952 = n12473 ;
  assign y2953 = n12485 ;
  assign y2954 = ~n12488 ;
  assign y2955 = ~n12491 ;
  assign y2956 = ~n12494 ;
  assign y2957 = n12495 ;
  assign y2958 = ~n12503 ;
  assign y2959 = ~n12507 ;
  assign y2960 = ~n12508 ;
  assign y2961 = n12511 ;
  assign y2962 = n12519 ;
  assign y2963 = n12521 ;
  assign y2964 = ~1'b0 ;
  assign y2965 = n12524 ;
  assign y2966 = ~n12527 ;
  assign y2967 = ~n12529 ;
  assign y2968 = ~n12535 ;
  assign y2969 = ~n12537 ;
  assign y2970 = n12543 ;
  assign y2971 = ~n12549 ;
  assign y2972 = n12550 ;
  assign y2973 = ~n12557 ;
  assign y2974 = n12561 ;
  assign y2975 = n12563 ;
  assign y2976 = ~1'b0 ;
  assign y2977 = n12568 ;
  assign y2978 = ~n12572 ;
  assign y2979 = n12580 ;
  assign y2980 = ~n12581 ;
  assign y2981 = n12582 ;
  assign y2982 = n12589 ;
  assign y2983 = n12591 ;
  assign y2984 = n12592 ;
  assign y2985 = ~n12597 ;
  assign y2986 = n12599 ;
  assign y2987 = n12600 ;
  assign y2988 = ~n12603 ;
  assign y2989 = ~1'b0 ;
  assign y2990 = ~1'b0 ;
  assign y2991 = n12607 ;
  assign y2992 = n12609 ;
  assign y2993 = ~n12610 ;
  assign y2994 = n12624 ;
  assign y2995 = n12625 ;
  assign y2996 = ~n12631 ;
  assign y2997 = ~n12637 ;
  assign y2998 = ~n12638 ;
  assign y2999 = ~n12641 ;
  assign y3000 = ~n12645 ;
  assign y3001 = n12651 ;
  assign y3002 = n12661 ;
  assign y3003 = ~1'b0 ;
  assign y3004 = n12665 ;
  assign y3005 = n12668 ;
  assign y3006 = ~n12669 ;
  assign y3007 = ~n12671 ;
  assign y3008 = ~n12672 ;
  assign y3009 = ~n12673 ;
  assign y3010 = ~n12680 ;
  assign y3011 = ~n12681 ;
  assign y3012 = ~n12684 ;
  assign y3013 = ~n12685 ;
  assign y3014 = ~1'b0 ;
  assign y3015 = ~n12688 ;
  assign y3016 = ~n12689 ;
  assign y3017 = ~1'b0 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = ~n12695 ;
  assign y3020 = n12696 ;
  assign y3021 = ~n12715 ;
  assign y3022 = n12716 ;
  assign y3023 = ~n12736 ;
  assign y3024 = ~n12747 ;
  assign y3025 = n12749 ;
  assign y3026 = ~n12751 ;
  assign y3027 = n12758 ;
  assign y3028 = n12761 ;
  assign y3029 = ~n12765 ;
  assign y3030 = n12767 ;
  assign y3031 = ~n12773 ;
  assign y3032 = n12775 ;
  assign y3033 = ~n12776 ;
  assign y3034 = ~n12779 ;
  assign y3035 = n12782 ;
  assign y3036 = ~n12789 ;
  assign y3037 = ~n12790 ;
  assign y3038 = ~n12804 ;
  assign y3039 = n12807 ;
  assign y3040 = ~1'b0 ;
  assign y3041 = ~n12813 ;
  assign y3042 = n12814 ;
  assign y3043 = ~1'b0 ;
  assign y3044 = n12822 ;
  assign y3045 = n12823 ;
  assign y3046 = ~n12824 ;
  assign y3047 = ~n12831 ;
  assign y3048 = ~1'b0 ;
  assign y3049 = ~n12832 ;
  assign y3050 = ~n12833 ;
  assign y3051 = n12836 ;
  assign y3052 = n12838 ;
  assign y3053 = n12846 ;
  assign y3054 = ~n12847 ;
  assign y3055 = n12848 ;
  assign y3056 = n12850 ;
  assign y3057 = n12858 ;
  assign y3058 = ~n12863 ;
  assign y3059 = ~1'b0 ;
  assign y3060 = ~n12865 ;
  assign y3061 = ~1'b0 ;
  assign y3062 = ~1'b0 ;
  assign y3063 = n12866 ;
  assign y3064 = n12871 ;
  assign y3065 = ~n12874 ;
  assign y3066 = ~n12875 ;
  assign y3067 = n12879 ;
  assign y3068 = ~n12886 ;
  assign y3069 = ~n12888 ;
  assign y3070 = n12890 ;
  assign y3071 = n12891 ;
  assign y3072 = ~n12897 ;
  assign y3073 = ~1'b0 ;
  assign y3074 = n12902 ;
  assign y3075 = n12907 ;
  assign y3076 = ~n12915 ;
  assign y3077 = n12917 ;
  assign y3078 = ~n12919 ;
  assign y3079 = ~n1663 ;
  assign y3080 = ~n12925 ;
  assign y3081 = n12930 ;
  assign y3082 = ~n12934 ;
  assign y3083 = ~n12939 ;
  assign y3084 = n12941 ;
  assign y3085 = n12943 ;
  assign y3086 = n12946 ;
  assign y3087 = ~n12947 ;
  assign y3088 = n12354 ;
  assign y3089 = ~n12951 ;
  assign y3090 = ~n12952 ;
  assign y3091 = n12953 ;
  assign y3092 = n12956 ;
  assign y3093 = ~n12962 ;
  assign y3094 = ~n12964 ;
  assign y3095 = n12965 ;
  assign y3096 = ~n12972 ;
  assign y3097 = ~n12977 ;
  assign y3098 = ~n12982 ;
  assign y3099 = ~n12983 ;
  assign y3100 = ~1'b0 ;
  assign y3101 = ~n12984 ;
  assign y3102 = ~n12985 ;
  assign y3103 = n12986 ;
  assign y3104 = ~n12987 ;
  assign y3105 = ~n12988 ;
  assign y3106 = ~1'b0 ;
  assign y3107 = n12992 ;
  assign y3108 = ~n13002 ;
  assign y3109 = ~n13003 ;
  assign y3110 = n13004 ;
  assign y3111 = n13010 ;
  assign y3112 = n13017 ;
  assign y3113 = n13020 ;
  assign y3114 = ~n13025 ;
  assign y3115 = ~n13029 ;
  assign y3116 = ~n13033 ;
  assign y3117 = n13048 ;
  assign y3118 = n13065 ;
  assign y3119 = ~n13070 ;
  assign y3120 = ~1'b0 ;
  assign y3121 = ~n13071 ;
  assign y3122 = n13074 ;
  assign y3123 = n13075 ;
  assign y3124 = ~n13082 ;
  assign y3125 = ~n13083 ;
  assign y3126 = ~n13085 ;
  assign y3127 = ~n13086 ;
  assign y3128 = ~n13095 ;
  assign y3129 = ~n13096 ;
  assign y3130 = n13101 ;
  assign y3131 = n13104 ;
  assign y3132 = ~n13105 ;
  assign y3133 = n13107 ;
  assign y3134 = ~n13113 ;
  assign y3135 = n13115 ;
  assign y3136 = ~1'b0 ;
  assign y3137 = ~n13117 ;
  assign y3138 = ~n13120 ;
  assign y3139 = n13137 ;
  assign y3140 = ~n13139 ;
  assign y3141 = n13140 ;
  assign y3142 = ~1'b0 ;
  assign y3143 = n13144 ;
  assign y3144 = ~n13149 ;
  assign y3145 = n13155 ;
  assign y3146 = ~n13156 ;
  assign y3147 = ~n13161 ;
  assign y3148 = n13165 ;
  assign y3149 = n13170 ;
  assign y3150 = n13185 ;
  assign y3151 = n13188 ;
  assign y3152 = ~n13191 ;
  assign y3153 = n13195 ;
  assign y3154 = ~n13200 ;
  assign y3155 = n13202 ;
  assign y3156 = n13207 ;
  assign y3157 = ~n13210 ;
  assign y3158 = n13212 ;
  assign y3159 = ~1'b0 ;
  assign y3160 = n13216 ;
  assign y3161 = ~n13221 ;
  assign y3162 = n13223 ;
  assign y3163 = ~1'b0 ;
  assign y3164 = n13227 ;
  assign y3165 = ~n13229 ;
  assign y3166 = ~n13230 ;
  assign y3167 = ~n13233 ;
  assign y3168 = n13237 ;
  assign y3169 = ~1'b0 ;
  assign y3170 = n13241 ;
  assign y3171 = ~n13245 ;
  assign y3172 = ~n13250 ;
  assign y3173 = ~n13252 ;
  assign y3174 = n13253 ;
  assign y3175 = ~n13265 ;
  assign y3176 = n13267 ;
  assign y3177 = ~n13268 ;
  assign y3178 = n13274 ;
  assign y3179 = n13277 ;
  assign y3180 = ~n13280 ;
  assign y3181 = ~n13281 ;
  assign y3182 = ~n13283 ;
  assign y3183 = n13288 ;
  assign y3184 = n13302 ;
  assign y3185 = ~1'b0 ;
  assign y3186 = n13304 ;
  assign y3187 = ~n13310 ;
  assign y3188 = ~n13314 ;
  assign y3189 = n13320 ;
  assign y3190 = n13327 ;
  assign y3191 = ~n13328 ;
  assign y3192 = ~n13329 ;
  assign y3193 = ~1'b0 ;
  assign y3194 = n13332 ;
  assign y3195 = ~n13336 ;
  assign y3196 = ~n13339 ;
  assign y3197 = n13341 ;
  assign y3198 = ~n13343 ;
  assign y3199 = ~1'b0 ;
  assign y3200 = n13346 ;
  assign y3201 = ~n13349 ;
  assign y3202 = n13351 ;
  assign y3203 = ~n13356 ;
  assign y3204 = n13364 ;
  assign y3205 = ~n13365 ;
  assign y3206 = n13369 ;
  assign y3207 = ~n1051 ;
  assign y3208 = ~1'b0 ;
  assign y3209 = ~n13370 ;
  assign y3210 = n13376 ;
  assign y3211 = ~n13378 ;
  assign y3212 = ~n13380 ;
  assign y3213 = n13386 ;
  assign y3214 = ~1'b0 ;
  assign y3215 = ~1'b0 ;
  assign y3216 = n13387 ;
  assign y3217 = n13394 ;
  assign y3218 = ~n13398 ;
  assign y3219 = n13401 ;
  assign y3220 = ~n13403 ;
  assign y3221 = n13405 ;
  assign y3222 = ~n13409 ;
  assign y3223 = ~n2251 ;
  assign y3224 = ~n13411 ;
  assign y3225 = ~n13412 ;
  assign y3226 = n13417 ;
  assign y3227 = ~n13424 ;
  assign y3228 = ~n13425 ;
  assign y3229 = ~n13426 ;
  assign y3230 = ~n13427 ;
  assign y3231 = ~1'b0 ;
  assign y3232 = n13434 ;
  assign y3233 = ~n13442 ;
  assign y3234 = n13446 ;
  assign y3235 = ~n13469 ;
  assign y3236 = ~n13470 ;
  assign y3237 = n13471 ;
  assign y3238 = n13474 ;
  assign y3239 = ~n13479 ;
  assign y3240 = ~1'b0 ;
  assign y3241 = ~n13482 ;
  assign y3242 = n13494 ;
  assign y3243 = ~1'b0 ;
  assign y3244 = ~n13497 ;
  assign y3245 = n13498 ;
  assign y3246 = ~1'b0 ;
  assign y3247 = n13501 ;
  assign y3248 = ~n13503 ;
  assign y3249 = n13505 ;
  assign y3250 = ~n13511 ;
  assign y3251 = ~n13514 ;
  assign y3252 = n13520 ;
  assign y3253 = ~n13522 ;
  assign y3254 = ~n13533 ;
  assign y3255 = ~1'b0 ;
  assign y3256 = n13536 ;
  assign y3257 = ~n13537 ;
  assign y3258 = n13539 ;
  assign y3259 = ~n13540 ;
  assign y3260 = ~n13543 ;
  assign y3261 = ~n13549 ;
  assign y3262 = n13555 ;
  assign y3263 = ~n13557 ;
  assign y3264 = n13558 ;
  assign y3265 = ~n13561 ;
  assign y3266 = ~n13563 ;
  assign y3267 = n13574 ;
  assign y3268 = ~n13576 ;
  assign y3269 = ~n13577 ;
  assign y3270 = n13581 ;
  assign y3271 = n13588 ;
  assign y3272 = n13590 ;
  assign y3273 = ~n13595 ;
  assign y3274 = ~n13596 ;
  assign y3275 = n13602 ;
  assign y3276 = n13604 ;
  assign y3277 = ~n13606 ;
  assign y3278 = ~n13607 ;
  assign y3279 = n13611 ;
  assign y3280 = ~1'b0 ;
  assign y3281 = ~n13612 ;
  assign y3282 = ~n13617 ;
  assign y3283 = n13618 ;
  assign y3284 = n13623 ;
  assign y3285 = n13632 ;
  assign y3286 = n13637 ;
  assign y3287 = ~n13647 ;
  assign y3288 = n13649 ;
  assign y3289 = n13655 ;
  assign y3290 = ~n13658 ;
  assign y3291 = ~n13661 ;
  assign y3292 = n13663 ;
  assign y3293 = n13671 ;
  assign y3294 = n13672 ;
  assign y3295 = ~n13677 ;
  assign y3296 = n13678 ;
  assign y3297 = n13681 ;
  assign y3298 = ~n13683 ;
  assign y3299 = n13685 ;
  assign y3300 = n13690 ;
  assign y3301 = ~n13693 ;
  assign y3302 = n13696 ;
  assign y3303 = n13698 ;
  assign y3304 = ~1'b0 ;
  assign y3305 = ~n13702 ;
  assign y3306 = ~n13706 ;
  assign y3307 = ~n13710 ;
  assign y3308 = ~n13719 ;
  assign y3309 = ~n13726 ;
  assign y3310 = ~1'b0 ;
  assign y3311 = ~n13733 ;
  assign y3312 = n13745 ;
  assign y3313 = n13748 ;
  assign y3314 = n13755 ;
  assign y3315 = n13760 ;
  assign y3316 = ~n13765 ;
  assign y3317 = ~n13771 ;
  assign y3318 = n13774 ;
  assign y3319 = n13775 ;
  assign y3320 = ~n13776 ;
  assign y3321 = ~1'b0 ;
  assign y3322 = n13779 ;
  assign y3323 = ~n13781 ;
  assign y3324 = n13782 ;
  assign y3325 = ~1'b0 ;
  assign y3326 = ~n13786 ;
  assign y3327 = ~n13787 ;
  assign y3328 = ~n13792 ;
  assign y3329 = ~n1108 ;
  assign y3330 = ~1'b0 ;
  assign y3331 = ~1'b0 ;
  assign y3332 = n13793 ;
  assign y3333 = ~n13798 ;
  assign y3334 = n13806 ;
  assign y3335 = ~n13818 ;
  assign y3336 = ~n13838 ;
  assign y3337 = ~n13846 ;
  assign y3338 = ~n13850 ;
  assign y3339 = n13851 ;
  assign y3340 = ~n13853 ;
  assign y3341 = ~n13855 ;
  assign y3342 = ~n13858 ;
  assign y3343 = n13859 ;
  assign y3344 = n13861 ;
  assign y3345 = n13871 ;
  assign y3346 = ~1'b0 ;
  assign y3347 = n13874 ;
  assign y3348 = ~n13884 ;
  assign y3349 = ~n13885 ;
  assign y3350 = ~n13888 ;
  assign y3351 = ~n13890 ;
  assign y3352 = ~n13896 ;
  assign y3353 = n13898 ;
  assign y3354 = ~n13902 ;
  assign y3355 = ~n13905 ;
  assign y3356 = ~n13907 ;
  assign y3357 = n13910 ;
  assign y3358 = ~n13912 ;
  assign y3359 = n13924 ;
  assign y3360 = n13925 ;
  assign y3361 = ~n13930 ;
  assign y3362 = n13937 ;
  assign y3363 = ~n13940 ;
  assign y3364 = ~1'b0 ;
  assign y3365 = ~n13943 ;
  assign y3366 = n13944 ;
  assign y3367 = n13949 ;
  assign y3368 = ~n13952 ;
  assign y3369 = ~n13954 ;
  assign y3370 = ~1'b0 ;
  assign y3371 = n13958 ;
  assign y3372 = ~n13963 ;
  assign y3373 = n13974 ;
  assign y3374 = n13980 ;
  assign y3375 = ~n13985 ;
  assign y3376 = ~n13986 ;
  assign y3377 = ~n13987 ;
  assign y3378 = ~n13988 ;
  assign y3379 = n13992 ;
  assign y3380 = n13994 ;
  assign y3381 = ~n13998 ;
  assign y3382 = n14002 ;
  assign y3383 = n14009 ;
  assign y3384 = ~n14010 ;
  assign y3385 = n14014 ;
  assign y3386 = ~n14018 ;
  assign y3387 = ~n14023 ;
  assign y3388 = n14029 ;
  assign y3389 = n14032 ;
  assign y3390 = ~n14037 ;
  assign y3391 = ~n14038 ;
  assign y3392 = n14050 ;
  assign y3393 = n14054 ;
  assign y3394 = n14057 ;
  assign y3395 = ~n14062 ;
  assign y3396 = ~n14066 ;
  assign y3397 = n14072 ;
  assign y3398 = ~n14075 ;
  assign y3399 = n14080 ;
  assign y3400 = n14081 ;
  assign y3401 = n14082 ;
  assign y3402 = n14084 ;
  assign y3403 = n14087 ;
  assign y3404 = ~n14091 ;
  assign y3405 = ~n14093 ;
  assign y3406 = ~n14095 ;
  assign y3407 = n14105 ;
  assign y3408 = n14107 ;
  assign y3409 = n14111 ;
  assign y3410 = ~n14114 ;
  assign y3411 = ~n14119 ;
  assign y3412 = ~n14120 ;
  assign y3413 = ~n14122 ;
  assign y3414 = n14126 ;
  assign y3415 = ~n14132 ;
  assign y3416 = n14137 ;
  assign y3417 = n14138 ;
  assign y3418 = n14140 ;
  assign y3419 = ~n14142 ;
  assign y3420 = n14152 ;
  assign y3421 = ~n14160 ;
  assign y3422 = n14162 ;
  assign y3423 = ~n14163 ;
  assign y3424 = ~1'b0 ;
  assign y3425 = ~n14164 ;
  assign y3426 = n14166 ;
  assign y3427 = ~n14169 ;
  assign y3428 = n14171 ;
  assign y3429 = n14172 ;
  assign y3430 = n14175 ;
  assign y3431 = n14176 ;
  assign y3432 = ~n14179 ;
  assign y3433 = n14186 ;
  assign y3434 = n14199 ;
  assign y3435 = ~n14200 ;
  assign y3436 = ~n14202 ;
  assign y3437 = ~n14204 ;
  assign y3438 = ~n14207 ;
  assign y3439 = ~n14213 ;
  assign y3440 = ~n14217 ;
  assign y3441 = ~n14230 ;
  assign y3442 = n14234 ;
  assign y3443 = ~n14236 ;
  assign y3444 = n14238 ;
  assign y3445 = n14242 ;
  assign y3446 = ~1'b0 ;
  assign y3447 = n14247 ;
  assign y3448 = ~n14248 ;
  assign y3449 = ~n14252 ;
  assign y3450 = n14257 ;
  assign y3451 = n14259 ;
  assign y3452 = ~n14262 ;
  assign y3453 = ~n14263 ;
  assign y3454 = n14270 ;
  assign y3455 = ~n14275 ;
  assign y3456 = ~n14280 ;
  assign y3457 = ~n14283 ;
  assign y3458 = n14285 ;
  assign y3459 = n14295 ;
  assign y3460 = n14296 ;
  assign y3461 = n14302 ;
  assign y3462 = ~n14305 ;
  assign y3463 = ~n14307 ;
  assign y3464 = n14309 ;
  assign y3465 = n14310 ;
  assign y3466 = n14315 ;
  assign y3467 = n14321 ;
  assign y3468 = ~1'b0 ;
  assign y3469 = ~n14322 ;
  assign y3470 = n14323 ;
  assign y3471 = n14324 ;
  assign y3472 = n14325 ;
  assign y3473 = ~n14327 ;
  assign y3474 = ~n14330 ;
  assign y3475 = n14335 ;
  assign y3476 = n14338 ;
  assign y3477 = ~n14341 ;
  assign y3478 = ~n14343 ;
  assign y3479 = ~n14345 ;
  assign y3480 = ~n14349 ;
  assign y3481 = ~n14350 ;
  assign y3482 = ~n14351 ;
  assign y3483 = ~1'b0 ;
  assign y3484 = ~n14353 ;
  assign y3485 = n14356 ;
  assign y3486 = ~n14364 ;
  assign y3487 = ~n14365 ;
  assign y3488 = n14366 ;
  assign y3489 = n14367 ;
  assign y3490 = n9504 ;
  assign y3491 = ~n14369 ;
  assign y3492 = n14371 ;
  assign y3493 = ~1'b0 ;
  assign y3494 = ~n14374 ;
  assign y3495 = ~n14375 ;
  assign y3496 = ~n14377 ;
  assign y3497 = ~n14381 ;
  assign y3498 = ~n14383 ;
  assign y3499 = n14391 ;
  assign y3500 = ~n14395 ;
  assign y3501 = ~n14396 ;
  assign y3502 = ~n14399 ;
  assign y3503 = ~1'b0 ;
  assign y3504 = n14404 ;
  assign y3505 = ~n14407 ;
  assign y3506 = ~n14412 ;
  assign y3507 = n14419 ;
  assign y3508 = n14427 ;
  assign y3509 = ~n14430 ;
  assign y3510 = ~n14433 ;
  assign y3511 = ~1'b0 ;
  assign y3512 = n14439 ;
  assign y3513 = ~n14440 ;
  assign y3514 = ~1'b0 ;
  assign y3515 = ~n14446 ;
  assign y3516 = n14454 ;
  assign y3517 = n14455 ;
  assign y3518 = ~n14457 ;
  assign y3519 = n14458 ;
  assign y3520 = ~n14461 ;
  assign y3521 = ~n14466 ;
  assign y3522 = ~n14468 ;
  assign y3523 = ~n14472 ;
  assign y3524 = n14473 ;
  assign y3525 = ~1'b0 ;
  assign y3526 = n14477 ;
  assign y3527 = ~n14481 ;
  assign y3528 = ~n14482 ;
  assign y3529 = ~n14483 ;
  assign y3530 = ~n14488 ;
  assign y3531 = ~n14493 ;
  assign y3532 = ~n14502 ;
  assign y3533 = n14506 ;
  assign y3534 = ~1'b0 ;
  assign y3535 = n14511 ;
  assign y3536 = ~n14513 ;
  assign y3537 = ~n14525 ;
  assign y3538 = ~n14526 ;
  assign y3539 = ~1'b0 ;
  assign y3540 = ~n14528 ;
  assign y3541 = n14532 ;
  assign y3542 = n14533 ;
  assign y3543 = ~1'b0 ;
  assign y3544 = ~n14535 ;
  assign y3545 = n14538 ;
  assign y3546 = ~n14544 ;
  assign y3547 = n14546 ;
  assign y3548 = ~n14548 ;
  assign y3549 = n14556 ;
  assign y3550 = ~1'b0 ;
  assign y3551 = ~n14559 ;
  assign y3552 = ~n14563 ;
  assign y3553 = ~n14569 ;
  assign y3554 = ~n14570 ;
  assign y3555 = n14573 ;
  assign y3556 = ~n14578 ;
  assign y3557 = n14579 ;
  assign y3558 = n14581 ;
  assign y3559 = n14582 ;
  assign y3560 = ~n14585 ;
  assign y3561 = n14586 ;
  assign y3562 = n14587 ;
  assign y3563 = n14592 ;
  assign y3564 = n14597 ;
  assign y3565 = ~n14599 ;
  assign y3566 = n14604 ;
  assign y3567 = ~n14609 ;
  assign y3568 = ~n14617 ;
  assign y3569 = n14621 ;
  assign y3570 = ~n14623 ;
  assign y3571 = ~1'b0 ;
  assign y3572 = n14629 ;
  assign y3573 = n14634 ;
  assign y3574 = ~n14635 ;
  assign y3575 = n14643 ;
  assign y3576 = n14650 ;
  assign y3577 = ~n14655 ;
  assign y3578 = n14658 ;
  assign y3579 = ~n14666 ;
  assign y3580 = n14667 ;
  assign y3581 = ~n14680 ;
  assign y3582 = ~1'b0 ;
  assign y3583 = n14681 ;
  assign y3584 = ~n14683 ;
  assign y3585 = n14684 ;
  assign y3586 = ~n14691 ;
  assign y3587 = ~1'b0 ;
  assign y3588 = n14694 ;
  assign y3589 = ~n14697 ;
  assign y3590 = n14698 ;
  assign y3591 = n14701 ;
  assign y3592 = ~n14703 ;
  assign y3593 = n14707 ;
  assign y3594 = ~n14709 ;
  assign y3595 = ~1'b0 ;
  assign y3596 = ~n14710 ;
  assign y3597 = n14722 ;
  assign y3598 = n14728 ;
  assign y3599 = n14733 ;
  assign y3600 = n14737 ;
  assign y3601 = ~n14738 ;
  assign y3602 = ~n14742 ;
  assign y3603 = n14744 ;
  assign y3604 = ~n14746 ;
  assign y3605 = ~n14747 ;
  assign y3606 = ~n14751 ;
  assign y3607 = n14758 ;
  assign y3608 = ~n14764 ;
  assign y3609 = n14770 ;
  assign y3610 = n14774 ;
  assign y3611 = ~n14784 ;
  assign y3612 = ~n14789 ;
  assign y3613 = ~n14795 ;
  assign y3614 = ~1'b0 ;
  assign y3615 = n14804 ;
  assign y3616 = ~n14807 ;
  assign y3617 = ~n14809 ;
  assign y3618 = n14811 ;
  assign y3619 = n14813 ;
  assign y3620 = ~n14817 ;
  assign y3621 = ~n14825 ;
  assign y3622 = n14830 ;
  assign y3623 = ~1'b0 ;
  assign y3624 = n14833 ;
  assign y3625 = n14836 ;
  assign y3626 = ~n14837 ;
  assign y3627 = ~n14842 ;
  assign y3628 = ~1'b0 ;
  assign y3629 = ~n14851 ;
  assign y3630 = ~n14853 ;
  assign y3631 = ~n14857 ;
  assign y3632 = ~n14861 ;
  assign y3633 = ~n14863 ;
  assign y3634 = ~n14864 ;
  assign y3635 = ~n14865 ;
  assign y3636 = ~n14866 ;
  assign y3637 = n14870 ;
  assign y3638 = n14871 ;
  assign y3639 = n6219 ;
  assign y3640 = ~n14879 ;
  assign y3641 = ~1'b0 ;
  assign y3642 = ~n14881 ;
  assign y3643 = n14884 ;
  assign y3644 = ~n14887 ;
  assign y3645 = n14888 ;
  assign y3646 = n14890 ;
  assign y3647 = ~n14894 ;
  assign y3648 = n14898 ;
  assign y3649 = n14901 ;
  assign y3650 = ~n14905 ;
  assign y3651 = ~1'b0 ;
  assign y3652 = n14916 ;
  assign y3653 = ~n14917 ;
  assign y3654 = ~n14920 ;
  assign y3655 = n14926 ;
  assign y3656 = ~n14929 ;
  assign y3657 = n14934 ;
  assign y3658 = ~1'b0 ;
  assign y3659 = ~n14935 ;
  assign y3660 = ~n14940 ;
  assign y3661 = n14953 ;
  assign y3662 = n14954 ;
  assign y3663 = n14962 ;
  assign y3664 = n14967 ;
  assign y3665 = n14968 ;
  assign y3666 = n14970 ;
  assign y3667 = ~n14971 ;
  assign y3668 = ~n14976 ;
  assign y3669 = n14978 ;
  assign y3670 = ~1'b0 ;
  assign y3671 = n14980 ;
  assign y3672 = ~1'b0 ;
  assign y3673 = ~n14982 ;
  assign y3674 = ~n14984 ;
  assign y3675 = n14989 ;
  assign y3676 = ~n14992 ;
  assign y3677 = n14994 ;
  assign y3678 = ~n14999 ;
  assign y3679 = ~n15000 ;
  assign y3680 = n15005 ;
  assign y3681 = ~n15006 ;
  assign y3682 = ~n15015 ;
  assign y3683 = ~n15019 ;
  assign y3684 = n15022 ;
  assign y3685 = ~n15027 ;
  assign y3686 = ~n15030 ;
  assign y3687 = n15032 ;
  assign y3688 = n15038 ;
  assign y3689 = n15044 ;
  assign y3690 = ~n15045 ;
  assign y3691 = n15047 ;
  assign y3692 = n15052 ;
  assign y3693 = ~n15054 ;
  assign y3694 = n15055 ;
  assign y3695 = n15058 ;
  assign y3696 = n15068 ;
  assign y3697 = n15070 ;
  assign y3698 = n15073 ;
  assign y3699 = ~1'b0 ;
  assign y3700 = n15075 ;
  assign y3701 = n15081 ;
  assign y3702 = n15082 ;
  assign y3703 = ~n15089 ;
  assign y3704 = n15092 ;
  assign y3705 = n15093 ;
  assign y3706 = ~n15098 ;
  assign y3707 = ~n15100 ;
  assign y3708 = ~1'b0 ;
  assign y3709 = n15102 ;
  assign y3710 = ~n15103 ;
  assign y3711 = n15104 ;
  assign y3712 = n15106 ;
  assign y3713 = ~1'b0 ;
  assign y3714 = ~1'b0 ;
  assign y3715 = ~n15107 ;
  assign y3716 = n15109 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = n15117 ;
  assign y3719 = ~n15119 ;
  assign y3720 = ~n15120 ;
  assign y3721 = n15122 ;
  assign y3722 = n15126 ;
  assign y3723 = n15129 ;
  assign y3724 = ~n15130 ;
  assign y3725 = n15131 ;
  assign y3726 = n15135 ;
  assign y3727 = n15137 ;
  assign y3728 = ~n15138 ;
  assign y3729 = ~n15150 ;
  assign y3730 = n15153 ;
  assign y3731 = ~n15158 ;
  assign y3732 = n15160 ;
  assign y3733 = ~n15174 ;
  assign y3734 = ~n15180 ;
  assign y3735 = ~n15182 ;
  assign y3736 = ~n9426 ;
  assign y3737 = ~n15185 ;
  assign y3738 = ~n15189 ;
  assign y3739 = ~n15190 ;
  assign y3740 = ~n15192 ;
  assign y3741 = ~n15197 ;
  assign y3742 = ~n15198 ;
  assign y3743 = n15201 ;
  assign y3744 = ~n15205 ;
  assign y3745 = ~n15207 ;
  assign y3746 = ~1'b0 ;
  assign y3747 = n15215 ;
  assign y3748 = ~n15216 ;
  assign y3749 = n15219 ;
  assign y3750 = n15222 ;
  assign y3751 = ~n15223 ;
  assign y3752 = ~n15225 ;
  assign y3753 = ~n15227 ;
  assign y3754 = n15229 ;
  assign y3755 = n15233 ;
  assign y3756 = n15235 ;
  assign y3757 = ~n15240 ;
  assign y3758 = ~1'b0 ;
  assign y3759 = ~n15243 ;
  assign y3760 = n15245 ;
  assign y3761 = ~n15252 ;
  assign y3762 = n15257 ;
  assign y3763 = ~n15266 ;
  assign y3764 = ~n15275 ;
  assign y3765 = n15279 ;
  assign y3766 = ~n15280 ;
  assign y3767 = ~n15284 ;
  assign y3768 = ~1'b0 ;
  assign y3769 = ~n15286 ;
  assign y3770 = ~n15290 ;
  assign y3771 = ~n15292 ;
  assign y3772 = n15294 ;
  assign y3773 = n15297 ;
  assign y3774 = ~n15299 ;
  assign y3775 = n15302 ;
  assign y3776 = ~n15305 ;
  assign y3777 = n15308 ;
  assign y3778 = ~n15313 ;
  assign y3779 = ~1'b0 ;
  assign y3780 = ~n15315 ;
  assign y3781 = n15317 ;
  assign y3782 = n15329 ;
  assign y3783 = ~1'b0 ;
  assign y3784 = ~1'b0 ;
  assign y3785 = ~n15339 ;
  assign y3786 = ~n1416 ;
  assign y3787 = ~n15340 ;
  assign y3788 = n15342 ;
  assign y3789 = ~n15343 ;
  assign y3790 = n15346 ;
  assign y3791 = n15348 ;
  assign y3792 = ~n15354 ;
  assign y3793 = n15355 ;
  assign y3794 = ~n15366 ;
  assign y3795 = ~1'b0 ;
  assign y3796 = ~n15371 ;
  assign y3797 = n15372 ;
  assign y3798 = ~n15373 ;
  assign y3799 = ~n15383 ;
  assign y3800 = ~1'b0 ;
  assign y3801 = n15385 ;
  assign y3802 = ~n15389 ;
  assign y3803 = ~n15393 ;
  assign y3804 = n15400 ;
  assign y3805 = ~n15402 ;
  assign y3806 = ~n15404 ;
  assign y3807 = n15411 ;
  assign y3808 = ~1'b0 ;
  assign y3809 = ~n15414 ;
  assign y3810 = ~n15417 ;
  assign y3811 = n15422 ;
  assign y3812 = n15427 ;
  assign y3813 = n15431 ;
  assign y3814 = n15436 ;
  assign y3815 = ~n15437 ;
  assign y3816 = ~n15438 ;
  assign y3817 = n15442 ;
  assign y3818 = ~n15445 ;
  assign y3819 = n15447 ;
  assign y3820 = ~n15457 ;
  assign y3821 = ~n15463 ;
  assign y3822 = ~1'b0 ;
  assign y3823 = ~n15466 ;
  assign y3824 = n15471 ;
  assign y3825 = n15478 ;
  assign y3826 = n15481 ;
  assign y3827 = ~n15482 ;
  assign y3828 = ~n15490 ;
  assign y3829 = n15491 ;
  assign y3830 = n15492 ;
  assign y3831 = ~n15506 ;
  assign y3832 = n15514 ;
  assign y3833 = n15516 ;
  assign y3834 = n15517 ;
  assign y3835 = n15527 ;
  assign y3836 = ~n15531 ;
  assign y3837 = ~n15534 ;
  assign y3838 = ~n15536 ;
  assign y3839 = n15546 ;
  assign y3840 = ~n15547 ;
  assign y3841 = n15551 ;
  assign y3842 = n15557 ;
  assign y3843 = n15558 ;
  assign y3844 = n15561 ;
  assign y3845 = ~n15562 ;
  assign y3846 = ~n15569 ;
  assign y3847 = ~n15575 ;
  assign y3848 = ~n15577 ;
  assign y3849 = n15580 ;
  assign y3850 = ~n15586 ;
  assign y3851 = ~n15590 ;
  assign y3852 = n15592 ;
  assign y3853 = ~n15597 ;
  assign y3854 = n15598 ;
  assign y3855 = n15602 ;
  assign y3856 = n15605 ;
  assign y3857 = n15608 ;
  assign y3858 = ~n15609 ;
  assign y3859 = ~1'b0 ;
  assign y3860 = ~1'b0 ;
  assign y3861 = n15611 ;
  assign y3862 = ~n15616 ;
  assign y3863 = ~n15618 ;
  assign y3864 = n15620 ;
  assign y3865 = ~n15621 ;
  assign y3866 = n15627 ;
  assign y3867 = n15629 ;
  assign y3868 = ~n15636 ;
  assign y3869 = ~1'b0 ;
  assign y3870 = ~n15645 ;
  assign y3871 = ~n15648 ;
  assign y3872 = n15650 ;
  assign y3873 = n15652 ;
  assign y3874 = ~n15656 ;
  assign y3875 = n15663 ;
  assign y3876 = n15668 ;
  assign y3877 = ~n15673 ;
  assign y3878 = ~n15679 ;
  assign y3879 = n15682 ;
  assign y3880 = ~n15687 ;
  assign y3881 = ~1'b0 ;
  assign y3882 = n15692 ;
  assign y3883 = n15695 ;
  assign y3884 = ~n15705 ;
  assign y3885 = ~n15709 ;
  assign y3886 = ~n15712 ;
  assign y3887 = ~n15713 ;
  assign y3888 = ~1'b0 ;
  assign y3889 = n15715 ;
  assign y3890 = n15724 ;
  assign y3891 = ~n15732 ;
  assign y3892 = n15737 ;
  assign y3893 = ~n15743 ;
  assign y3894 = n15747 ;
  assign y3895 = n15751 ;
  assign y3896 = ~n15753 ;
  assign y3897 = ~n15756 ;
  assign y3898 = ~n15760 ;
  assign y3899 = n15762 ;
  assign y3900 = ~n15764 ;
  assign y3901 = n15775 ;
  assign y3902 = n15779 ;
  assign y3903 = ~n15780 ;
  assign y3904 = ~n15792 ;
  assign y3905 = ~n15796 ;
  assign y3906 = n15799 ;
  assign y3907 = n15810 ;
  assign y3908 = ~n15821 ;
  assign y3909 = ~1'b0 ;
  assign y3910 = ~n15832 ;
  assign y3911 = n15833 ;
  assign y3912 = ~1'b0 ;
  assign y3913 = ~n15834 ;
  assign y3914 = ~n15835 ;
  assign y3915 = n15837 ;
  assign y3916 = ~n15844 ;
  assign y3917 = n15848 ;
  assign y3918 = ~1'b0 ;
  assign y3919 = ~1'b0 ;
  assign y3920 = ~1'b0 ;
  assign y3921 = n15852 ;
  assign y3922 = ~n15860 ;
  assign y3923 = ~n15862 ;
  assign y3924 = n15867 ;
  assign y3925 = n15868 ;
  assign y3926 = ~1'b0 ;
  assign y3927 = ~n15872 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = ~1'b0 ;
  assign y3930 = n15878 ;
  assign y3931 = n15881 ;
  assign y3932 = ~n15884 ;
  assign y3933 = ~1'b0 ;
  assign y3934 = ~n15892 ;
  assign y3935 = n15895 ;
  assign y3936 = ~n15897 ;
  assign y3937 = n15899 ;
  assign y3938 = ~n15902 ;
  assign y3939 = n15913 ;
  assign y3940 = ~n15915 ;
  assign y3941 = ~1'b0 ;
  assign y3942 = ~n15918 ;
  assign y3943 = ~1'b0 ;
  assign y3944 = ~n15921 ;
  assign y3945 = ~n14035 ;
  assign y3946 = ~n15922 ;
  assign y3947 = ~n15923 ;
  assign y3948 = ~n15924 ;
  assign y3949 = n15931 ;
  assign y3950 = n15936 ;
  assign y3951 = ~n15937 ;
  assign y3952 = ~n15941 ;
  assign y3953 = ~n15942 ;
  assign y3954 = ~n15943 ;
  assign y3955 = ~n15946 ;
  assign y3956 = n15952 ;
  assign y3957 = ~n15954 ;
  assign y3958 = ~n7638 ;
  assign y3959 = n15966 ;
  assign y3960 = ~1'b0 ;
  assign y3961 = ~n15967 ;
  assign y3962 = n15973 ;
  assign y3963 = ~1'b0 ;
  assign y3964 = n15976 ;
  assign y3965 = ~n15985 ;
  assign y3966 = n15992 ;
  assign y3967 = ~n15996 ;
  assign y3968 = n15998 ;
  assign y3969 = ~n16001 ;
  assign y3970 = ~n16004 ;
  assign y3971 = n16006 ;
  assign y3972 = n16010 ;
  assign y3973 = n16013 ;
  assign y3974 = n16018 ;
  assign y3975 = ~n16022 ;
  assign y3976 = ~n16025 ;
  assign y3977 = ~n16028 ;
  assign y3978 = n16032 ;
  assign y3979 = ~n16034 ;
  assign y3980 = ~n16036 ;
  assign y3981 = ~1'b0 ;
  assign y3982 = n16040 ;
  assign y3983 = n16043 ;
  assign y3984 = n16053 ;
  assign y3985 = n16057 ;
  assign y3986 = ~n16058 ;
  assign y3987 = ~1'b0 ;
  assign y3988 = ~n16068 ;
  assign y3989 = n16072 ;
  assign y3990 = n16073 ;
  assign y3991 = ~n16075 ;
  assign y3992 = n16076 ;
  assign y3993 = ~n16077 ;
  assign y3994 = ~n16078 ;
  assign y3995 = n16080 ;
  assign y3996 = n16084 ;
  assign y3997 = ~n16085 ;
  assign y3998 = n16088 ;
  assign y3999 = ~n16089 ;
  assign y4000 = ~n16090 ;
  assign y4001 = n16093 ;
  assign y4002 = n16094 ;
  assign y4003 = n16097 ;
  assign y4004 = ~n16100 ;
  assign y4005 = n16105 ;
  assign y4006 = ~n16108 ;
  assign y4007 = ~n16113 ;
  assign y4008 = n16121 ;
  assign y4009 = ~n16129 ;
  assign y4010 = ~n16130 ;
  assign y4011 = n16132 ;
  assign y4012 = n16133 ;
  assign y4013 = n16138 ;
  assign y4014 = ~1'b0 ;
  assign y4015 = n16141 ;
  assign y4016 = ~n16144 ;
  assign y4017 = ~n16146 ;
  assign y4018 = ~n16153 ;
  assign y4019 = ~n16161 ;
  assign y4020 = ~n16162 ;
  assign y4021 = ~n16169 ;
  assign y4022 = ~n16171 ;
  assign y4023 = ~n16172 ;
  assign y4024 = n16178 ;
  assign y4025 = n16179 ;
  assign y4026 = n16180 ;
  assign y4027 = n16182 ;
  assign y4028 = n16183 ;
  assign y4029 = ~n16185 ;
  assign y4030 = ~n16191 ;
  assign y4031 = n16192 ;
  assign y4032 = ~n16197 ;
  assign y4033 = ~n16199 ;
  assign y4034 = ~n16202 ;
  assign y4035 = n16204 ;
  assign y4036 = ~n16206 ;
  assign y4037 = ~n16212 ;
  assign y4038 = n16222 ;
  assign y4039 = n16223 ;
  assign y4040 = ~1'b0 ;
  assign y4041 = n16233 ;
  assign y4042 = ~n16239 ;
  assign y4043 = ~n16247 ;
  assign y4044 = n16248 ;
  assign y4045 = ~1'b0 ;
  assign y4046 = ~n16251 ;
  assign y4047 = ~n16257 ;
  assign y4048 = n16258 ;
  assign y4049 = ~1'b0 ;
  assign y4050 = ~1'b0 ;
  assign y4051 = ~1'b0 ;
  assign y4052 = ~n16263 ;
  assign y4053 = n16268 ;
  assign y4054 = n16271 ;
  assign y4055 = n16279 ;
  assign y4056 = n16294 ;
  assign y4057 = n16303 ;
  assign y4058 = ~n16316 ;
  assign y4059 = n16324 ;
  assign y4060 = n16325 ;
  assign y4061 = ~n16328 ;
  assign y4062 = n16330 ;
  assign y4063 = n16332 ;
  assign y4064 = n16333 ;
  assign y4065 = ~n16341 ;
  assign y4066 = ~n16343 ;
  assign y4067 = ~n16348 ;
  assign y4068 = ~n16355 ;
  assign y4069 = n16356 ;
  assign y4070 = n16360 ;
  assign y4071 = n16362 ;
  assign y4072 = n16366 ;
  assign y4073 = n16367 ;
  assign y4074 = ~n16370 ;
  assign y4075 = n16372 ;
  assign y4076 = ~n16380 ;
  assign y4077 = ~n16381 ;
  assign y4078 = ~n16383 ;
  assign y4079 = ~n16387 ;
  assign y4080 = ~n16394 ;
  assign y4081 = n16395 ;
  assign y4082 = n16396 ;
  assign y4083 = n16398 ;
  assign y4084 = n16401 ;
  assign y4085 = n16402 ;
  assign y4086 = n16407 ;
  assign y4087 = ~1'b0 ;
  assign y4088 = ~1'b0 ;
  assign y4089 = ~n16409 ;
  assign y4090 = n16411 ;
  assign y4091 = ~n16412 ;
  assign y4092 = n16414 ;
  assign y4093 = ~n16418 ;
  assign y4094 = ~n16422 ;
  assign y4095 = ~n16423 ;
  assign y4096 = ~n16431 ;
  assign y4097 = ~1'b0 ;
  assign y4098 = n16432 ;
  assign y4099 = n16433 ;
  assign y4100 = n16442 ;
  assign y4101 = n16446 ;
  assign y4102 = n16448 ;
  assign y4103 = ~n16454 ;
  assign y4104 = ~n16455 ;
  assign y4105 = n16459 ;
  assign y4106 = ~n16460 ;
  assign y4107 = n16465 ;
  assign y4108 = ~n16469 ;
  assign y4109 = n16470 ;
  assign y4110 = ~n16472 ;
  assign y4111 = n16474 ;
  assign y4112 = ~n16480 ;
  assign y4113 = n16484 ;
  assign y4114 = n16486 ;
  assign y4115 = n16489 ;
  assign y4116 = n16492 ;
  assign y4117 = ~n16498 ;
  assign y4118 = ~1'b0 ;
  assign y4119 = n16504 ;
  assign y4120 = ~n16505 ;
  assign y4121 = n16511 ;
  assign y4122 = ~n16519 ;
  assign y4123 = ~n16522 ;
  assign y4124 = ~n16525 ;
  assign y4125 = ~n16529 ;
  assign y4126 = ~n16536 ;
  assign y4127 = ~n16539 ;
  assign y4128 = ~1'b0 ;
  assign y4129 = ~n16540 ;
  assign y4130 = n16542 ;
  assign y4131 = ~1'b0 ;
  assign y4132 = ~n16551 ;
  assign y4133 = ~n16556 ;
  assign y4134 = ~n16561 ;
  assign y4135 = n16566 ;
  assign y4136 = n16568 ;
  assign y4137 = ~1'b0 ;
  assign y4138 = ~n11334 ;
  assign y4139 = ~n16578 ;
  assign y4140 = n16579 ;
  assign y4141 = n16581 ;
  assign y4142 = n16585 ;
  assign y4143 = ~1'b0 ;
  assign y4144 = ~n16588 ;
  assign y4145 = ~n16589 ;
  assign y4146 = ~1'b0 ;
  assign y4147 = ~n16601 ;
  assign y4148 = n16602 ;
  assign y4149 = ~n16603 ;
  assign y4150 = n16605 ;
  assign y4151 = n16609 ;
  assign y4152 = n16617 ;
  assign y4153 = n16618 ;
  assign y4154 = ~n16623 ;
  assign y4155 = ~n16627 ;
  assign y4156 = ~n16628 ;
  assign y4157 = n16630 ;
  assign y4158 = n16634 ;
  assign y4159 = ~n16638 ;
  assign y4160 = ~n12823 ;
  assign y4161 = n16640 ;
  assign y4162 = ~n16644 ;
  assign y4163 = ~n16645 ;
  assign y4164 = n16647 ;
  assign y4165 = n16651 ;
  assign y4166 = ~n16657 ;
  assign y4167 = ~n16660 ;
  assign y4168 = ~n16663 ;
  assign y4169 = ~n16666 ;
  assign y4170 = ~1'b0 ;
  assign y4171 = ~n16668 ;
  assign y4172 = n16669 ;
  assign y4173 = ~n16671 ;
  assign y4174 = ~n16679 ;
  assign y4175 = ~n16680 ;
  assign y4176 = ~n16682 ;
  assign y4177 = ~n16685 ;
  assign y4178 = ~n16688 ;
  assign y4179 = ~n16690 ;
  assign y4180 = n16695 ;
  assign y4181 = ~n16698 ;
  assign y4182 = ~n16700 ;
  assign y4183 = ~n16706 ;
  assign y4184 = n16707 ;
  assign y4185 = ~n16710 ;
  assign y4186 = ~n16712 ;
  assign y4187 = n16716 ;
  assign y4188 = n16732 ;
  assign y4189 = ~1'b0 ;
  assign y4190 = ~n16734 ;
  assign y4191 = ~n16737 ;
  assign y4192 = ~n16742 ;
  assign y4193 = n16752 ;
  assign y4194 = ~n16763 ;
  assign y4195 = n16765 ;
  assign y4196 = n16769 ;
  assign y4197 = ~n16771 ;
  assign y4198 = n16772 ;
  assign y4199 = n16773 ;
  assign y4200 = n16774 ;
  assign y4201 = n16782 ;
  assign y4202 = ~n16788 ;
  assign y4203 = n16792 ;
  assign y4204 = ~n16793 ;
  assign y4205 = n16795 ;
  assign y4206 = ~1'b0 ;
  assign y4207 = n16798 ;
  assign y4208 = n16801 ;
  assign y4209 = n16802 ;
  assign y4210 = ~n16804 ;
  assign y4211 = n16805 ;
  assign y4212 = ~n16807 ;
  assign y4213 = n16809 ;
  assign y4214 = ~n16810 ;
  assign y4215 = ~n16813 ;
  assign y4216 = ~1'b0 ;
  assign y4217 = ~n16815 ;
  assign y4218 = n16822 ;
  assign y4219 = n16823 ;
  assign y4220 = ~n16825 ;
  assign y4221 = ~n16831 ;
  assign y4222 = n16837 ;
  assign y4223 = ~n16839 ;
  assign y4224 = ~n16841 ;
  assign y4225 = n16843 ;
  assign y4226 = ~1'b0 ;
  assign y4227 = n16845 ;
  assign y4228 = ~n16849 ;
  assign y4229 = ~n16850 ;
  assign y4230 = ~1'b0 ;
  assign y4231 = ~1'b0 ;
  assign y4232 = n16852 ;
  assign y4233 = n16858 ;
  assign y4234 = ~n16860 ;
  assign y4235 = n16864 ;
  assign y4236 = ~n16869 ;
  assign y4237 = n16871 ;
  assign y4238 = n16872 ;
  assign y4239 = ~n16875 ;
  assign y4240 = ~n16878 ;
  assign y4241 = ~n16879 ;
  assign y4242 = ~n16885 ;
  assign y4243 = ~n16903 ;
  assign y4244 = ~n16906 ;
  assign y4245 = ~n16907 ;
  assign y4246 = n16909 ;
  assign y4247 = ~1'b0 ;
  assign y4248 = n16912 ;
  assign y4249 = ~n16922 ;
  assign y4250 = ~n16925 ;
  assign y4251 = ~n16928 ;
  assign y4252 = ~1'b0 ;
  assign y4253 = ~1'b0 ;
  assign y4254 = n16929 ;
  assign y4255 = ~n16934 ;
  assign y4256 = ~n16938 ;
  assign y4257 = ~n16940 ;
  assign y4258 = n16942 ;
  assign y4259 = ~1'b0 ;
  assign y4260 = n16946 ;
  assign y4261 = ~n16947 ;
  assign y4262 = n16949 ;
  assign y4263 = ~n16950 ;
  assign y4264 = ~1'b0 ;
  assign y4265 = n16952 ;
  assign y4266 = ~n16956 ;
  assign y4267 = ~n16959 ;
  assign y4268 = n16960 ;
  assign y4269 = n16961 ;
  assign y4270 = n16963 ;
  assign y4271 = ~n16976 ;
  assign y4272 = n16977 ;
  assign y4273 = ~1'b0 ;
  assign y4274 = ~n16978 ;
  assign y4275 = ~n16981 ;
  assign y4276 = ~n16982 ;
  assign y4277 = ~n16991 ;
  assign y4278 = ~1'b0 ;
  assign y4279 = ~n16999 ;
  assign y4280 = ~n17003 ;
  assign y4281 = ~n17004 ;
  assign y4282 = ~n17006 ;
  assign y4283 = ~n17011 ;
  assign y4284 = n17017 ;
  assign y4285 = n17022 ;
  assign y4286 = ~n17023 ;
  assign y4287 = ~n17024 ;
  assign y4288 = ~n17027 ;
  assign y4289 = ~n17029 ;
  assign y4290 = ~n17030 ;
  assign y4291 = n17034 ;
  assign y4292 = n17035 ;
  assign y4293 = n17043 ;
  assign y4294 = ~n17044 ;
  assign y4295 = n17048 ;
  assign y4296 = ~n17049 ;
  assign y4297 = ~n17051 ;
  assign y4298 = ~n17054 ;
  assign y4299 = ~1'b0 ;
  assign y4300 = n17057 ;
  assign y4301 = ~n17060 ;
  assign y4302 = n17064 ;
  assign y4303 = n17065 ;
  assign y4304 = n17068 ;
  assign y4305 = ~n17071 ;
  assign y4306 = ~n17073 ;
  assign y4307 = ~n17074 ;
  assign y4308 = ~n17077 ;
  assign y4309 = n17080 ;
  assign y4310 = ~n17083 ;
  assign y4311 = n17086 ;
  assign y4312 = ~n17089 ;
  assign y4313 = n17095 ;
  assign y4314 = ~n17097 ;
  assign y4315 = ~n17099 ;
  assign y4316 = n17101 ;
  assign y4317 = n17103 ;
  assign y4318 = n17109 ;
  assign y4319 = ~n17114 ;
  assign y4320 = ~n17115 ;
  assign y4321 = ~n17118 ;
  assign y4322 = ~n17124 ;
  assign y4323 = n17125 ;
  assign y4324 = ~n17126 ;
  assign y4325 = ~n17128 ;
  assign y4326 = ~n17133 ;
  assign y4327 = ~n17136 ;
  assign y4328 = ~1'b0 ;
  assign y4329 = n17140 ;
  assign y4330 = ~n17141 ;
  assign y4331 = ~n17146 ;
  assign y4332 = ~n17147 ;
  assign y4333 = ~n17149 ;
  assign y4334 = n17150 ;
  assign y4335 = ~n17152 ;
  assign y4336 = ~n17155 ;
  assign y4337 = n17159 ;
  assign y4338 = ~1'b0 ;
  assign y4339 = ~n17164 ;
  assign y4340 = ~n17167 ;
  assign y4341 = n17170 ;
  assign y4342 = ~1'b0 ;
  assign y4343 = ~n17172 ;
  assign y4344 = ~n17173 ;
  assign y4345 = n17177 ;
  assign y4346 = ~1'b0 ;
  assign y4347 = ~n17182 ;
  assign y4348 = ~n17183 ;
  assign y4349 = ~n17189 ;
  assign y4350 = n17190 ;
  assign y4351 = ~n17191 ;
  assign y4352 = n17194 ;
  assign y4353 = ~1'b0 ;
  assign y4354 = ~n17204 ;
  assign y4355 = ~n17210 ;
  assign y4356 = ~n17217 ;
  assign y4357 = ~1'b0 ;
  assign y4358 = ~n17218 ;
  assign y4359 = ~n17219 ;
  assign y4360 = n17220 ;
  assign y4361 = n17223 ;
  assign y4362 = ~n17229 ;
  assign y4363 = ~n10831 ;
  assign y4364 = ~n17230 ;
  assign y4365 = n17232 ;
  assign y4366 = n17233 ;
  assign y4367 = ~1'b0 ;
  assign y4368 = n17236 ;
  assign y4369 = ~n17243 ;
  assign y4370 = ~n17246 ;
  assign y4371 = n17255 ;
  assign y4372 = ~n17256 ;
  assign y4373 = ~n17257 ;
  assign y4374 = ~n17259 ;
  assign y4375 = ~n17260 ;
  assign y4376 = n17270 ;
  assign y4377 = ~n17274 ;
  assign y4378 = n17281 ;
  assign y4379 = ~1'b0 ;
  assign y4380 = n17286 ;
  assign y4381 = ~n17290 ;
  assign y4382 = n17292 ;
  assign y4383 = n17297 ;
  assign y4384 = n17298 ;
  assign y4385 = n17303 ;
  assign y4386 = ~n17308 ;
  assign y4387 = n17310 ;
  assign y4388 = ~n17312 ;
  assign y4389 = n17314 ;
  assign y4390 = n17322 ;
  assign y4391 = ~1'b0 ;
  assign y4392 = ~n17325 ;
  assign y4393 = ~n17328 ;
  assign y4394 = ~n17329 ;
  assign y4395 = ~n17333 ;
  assign y4396 = ~n17342 ;
  assign y4397 = ~n17343 ;
  assign y4398 = n17348 ;
  assign y4399 = ~n17353 ;
  assign y4400 = ~1'b0 ;
  assign y4401 = ~n17356 ;
  assign y4402 = ~n17359 ;
  assign y4403 = ~1'b0 ;
  assign y4404 = ~n17361 ;
  assign y4405 = n17362 ;
  assign y4406 = n17365 ;
  assign y4407 = ~n17367 ;
  assign y4408 = ~1'b0 ;
  assign y4409 = n17369 ;
  assign y4410 = n17371 ;
  assign y4411 = ~n17374 ;
  assign y4412 = n17380 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = ~1'b0 ;
  assign y4415 = n17384 ;
  assign y4416 = ~n17385 ;
  assign y4417 = ~n17386 ;
  assign y4418 = n17389 ;
  assign y4419 = ~1'b0 ;
  assign y4420 = ~n17396 ;
  assign y4421 = ~n17398 ;
  assign y4422 = n17409 ;
  assign y4423 = ~n17416 ;
  assign y4424 = ~n17417 ;
  assign y4425 = n17421 ;
  assign y4426 = n17424 ;
  assign y4427 = n17427 ;
  assign y4428 = ~n17428 ;
  assign y4429 = n17437 ;
  assign y4430 = ~n17445 ;
  assign y4431 = ~n17446 ;
  assign y4432 = n17456 ;
  assign y4433 = ~n17457 ;
  assign y4434 = n17461 ;
  assign y4435 = n17462 ;
  assign y4436 = ~n17467 ;
  assign y4437 = n17472 ;
  assign y4438 = ~n17476 ;
  assign y4439 = n17485 ;
  assign y4440 = ~n17490 ;
  assign y4441 = n17497 ;
  assign y4442 = ~1'b0 ;
  assign y4443 = ~1'b0 ;
  assign y4444 = n17498 ;
  assign y4445 = ~n17501 ;
  assign y4446 = n17503 ;
  assign y4447 = n17505 ;
  assign y4448 = ~n6884 ;
  assign y4449 = n17508 ;
  assign y4450 = n17511 ;
  assign y4451 = ~n17513 ;
  assign y4452 = ~n17520 ;
  assign y4453 = n17521 ;
  assign y4454 = ~n17522 ;
  assign y4455 = n17524 ;
  assign y4456 = n17532 ;
  assign y4457 = n17533 ;
  assign y4458 = ~n17537 ;
  assign y4459 = ~1'b0 ;
  assign y4460 = ~n17550 ;
  assign y4461 = n17559 ;
  assign y4462 = ~n17560 ;
  assign y4463 = ~n15557 ;
  assign y4464 = ~n17564 ;
  assign y4465 = n17566 ;
  assign y4466 = ~n17567 ;
  assign y4467 = n17569 ;
  assign y4468 = n17570 ;
  assign y4469 = n17571 ;
  assign y4470 = n17572 ;
  assign y4471 = n17574 ;
  assign y4472 = ~n17576 ;
  assign y4473 = ~n17577 ;
  assign y4474 = ~n17578 ;
  assign y4475 = ~n17580 ;
  assign y4476 = n17585 ;
  assign y4477 = ~n17592 ;
  assign y4478 = ~n17595 ;
  assign y4479 = ~n17602 ;
  assign y4480 = n17611 ;
  assign y4481 = n17614 ;
  assign y4482 = n17617 ;
  assign y4483 = ~n17620 ;
  assign y4484 = ~n17621 ;
  assign y4485 = ~n17622 ;
  assign y4486 = ~1'b0 ;
  assign y4487 = ~n17626 ;
  assign y4488 = n17627 ;
  assign y4489 = ~n17634 ;
  assign y4490 = ~1'b0 ;
  assign y4491 = n17638 ;
  assign y4492 = n17639 ;
  assign y4493 = ~n17641 ;
  assign y4494 = n17649 ;
  assign y4495 = ~1'b0 ;
  assign y4496 = ~n17653 ;
  assign y4497 = n17659 ;
  assign y4498 = n17660 ;
  assign y4499 = n17664 ;
  assign y4500 = ~n17668 ;
  assign y4501 = ~n17673 ;
  assign y4502 = n17679 ;
  assign y4503 = ~n17683 ;
  assign y4504 = n17684 ;
  assign y4505 = ~n17687 ;
  assign y4506 = n17689 ;
  assign y4507 = ~n17691 ;
  assign y4508 = n17692 ;
  assign y4509 = n17693 ;
  assign y4510 = n17696 ;
  assign y4511 = n17705 ;
  assign y4512 = ~n17712 ;
  assign y4513 = ~1'b0 ;
  assign y4514 = ~1'b0 ;
  assign y4515 = n17714 ;
  assign y4516 = n17717 ;
  assign y4517 = ~n17719 ;
  assign y4518 = n17721 ;
  assign y4519 = ~n17722 ;
  assign y4520 = ~1'b0 ;
  assign y4521 = ~1'b0 ;
  assign y4522 = n17730 ;
  assign y4523 = n17732 ;
  assign y4524 = n17734 ;
  assign y4525 = n17740 ;
  assign y4526 = ~n17741 ;
  assign y4527 = ~n17747 ;
  assign y4528 = ~n17748 ;
  assign y4529 = n17750 ;
  assign y4530 = ~n17751 ;
  assign y4531 = ~1'b0 ;
  assign y4532 = ~1'b0 ;
  assign y4533 = n17757 ;
  assign y4534 = n17763 ;
  assign y4535 = n17764 ;
  assign y4536 = n17773 ;
  assign y4537 = n17774 ;
  assign y4538 = ~n17779 ;
  assign y4539 = ~n17780 ;
  assign y4540 = ~n17782 ;
  assign y4541 = 1'b0 ;
  assign y4542 = n17784 ;
  assign y4543 = n17790 ;
  assign y4544 = n17793 ;
  assign y4545 = n17794 ;
  assign y4546 = n17804 ;
  assign y4547 = ~n17805 ;
  assign y4548 = n17806 ;
  assign y4549 = n17812 ;
  assign y4550 = n2057 ;
  assign y4551 = ~n17815 ;
  assign y4552 = n17818 ;
  assign y4553 = n17820 ;
  assign y4554 = n17824 ;
  assign y4555 = ~n17829 ;
  assign y4556 = n17832 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = ~1'b0 ;
  assign y4559 = n17833 ;
  assign y4560 = ~n17838 ;
  assign y4561 = ~n17840 ;
  assign y4562 = ~n17847 ;
  assign y4563 = ~n17848 ;
  assign y4564 = n17849 ;
  assign y4565 = ~n17858 ;
  assign y4566 = ~n17862 ;
  assign y4567 = n17869 ;
  assign y4568 = n17876 ;
  assign y4569 = ~n17878 ;
  assign y4570 = ~1'b0 ;
  assign y4571 = ~1'b0 ;
  assign y4572 = ~1'b0 ;
  assign y4573 = ~n17881 ;
  assign y4574 = n17885 ;
  assign y4575 = n17890 ;
  assign y4576 = n17894 ;
  assign y4577 = ~n17896 ;
  assign y4578 = ~n17899 ;
  assign y4579 = ~1'b0 ;
  assign y4580 = ~n17902 ;
  assign y4581 = ~n17903 ;
  assign y4582 = ~n17906 ;
  assign y4583 = n17907 ;
  assign y4584 = ~n17908 ;
  assign y4585 = ~n17909 ;
  assign y4586 = ~n17913 ;
  assign y4587 = ~n17924 ;
  assign y4588 = n17927 ;
  assign y4589 = ~n17930 ;
  assign y4590 = ~n17938 ;
  assign y4591 = n17940 ;
  assign y4592 = ~n17942 ;
  assign y4593 = n17944 ;
  assign y4594 = ~n17946 ;
  assign y4595 = n17952 ;
  assign y4596 = ~n17956 ;
  assign y4597 = n17960 ;
  assign y4598 = ~n17964 ;
  assign y4599 = ~1'b0 ;
  assign y4600 = n17968 ;
  assign y4601 = n17970 ;
  assign y4602 = n17974 ;
  assign y4603 = ~n17976 ;
  assign y4604 = ~n17980 ;
  assign y4605 = ~1'b0 ;
  assign y4606 = ~n17981 ;
  assign y4607 = ~1'b0 ;
  assign y4608 = n17983 ;
  assign y4609 = ~n17987 ;
  assign y4610 = n17989 ;
  assign y4611 = ~n17995 ;
  assign y4612 = n17998 ;
  assign y4613 = ~n17999 ;
  assign y4614 = n18004 ;
  assign y4615 = ~1'b0 ;
  assign y4616 = ~n18007 ;
  assign y4617 = ~n18009 ;
  assign y4618 = ~1'b0 ;
  assign y4619 = ~n18012 ;
  assign y4620 = ~n18014 ;
  assign y4621 = n18017 ;
  assign y4622 = n18023 ;
  assign y4623 = n18027 ;
  assign y4624 = ~1'b0 ;
  assign y4625 = ~n18031 ;
  assign y4626 = n18033 ;
  assign y4627 = n18035 ;
  assign y4628 = ~n18036 ;
  assign y4629 = ~1'b0 ;
  assign y4630 = n18039 ;
  assign y4631 = ~n18041 ;
  assign y4632 = n18042 ;
  assign y4633 = n18043 ;
  assign y4634 = ~n18044 ;
  assign y4635 = ~n18045 ;
  assign y4636 = ~n18046 ;
  assign y4637 = ~n18047 ;
  assign y4638 = n18050 ;
  assign y4639 = n18051 ;
  assign y4640 = ~n18053 ;
  assign y4641 = ~n18055 ;
  assign y4642 = ~n18056 ;
  assign y4643 = n18057 ;
  assign y4644 = n18058 ;
  assign y4645 = n18061 ;
  assign y4646 = ~n18064 ;
  assign y4647 = ~n18066 ;
  assign y4648 = ~1'b0 ;
  assign y4649 = ~1'b0 ;
  assign y4650 = ~n18067 ;
  assign y4651 = n18074 ;
  assign y4652 = n18078 ;
  assign y4653 = n18079 ;
  assign y4654 = ~n18086 ;
  assign y4655 = ~1'b0 ;
  assign y4656 = n18087 ;
  assign y4657 = ~n18094 ;
  assign y4658 = n18098 ;
  assign y4659 = ~n18099 ;
  assign y4660 = n18100 ;
  assign y4661 = ~n18101 ;
  assign y4662 = ~n18102 ;
  assign y4663 = n18103 ;
  assign y4664 = n18105 ;
  assign y4665 = ~n18109 ;
  assign y4666 = n18112 ;
  assign y4667 = ~n18114 ;
  assign y4668 = ~n18115 ;
  assign y4669 = ~n18116 ;
  assign y4670 = ~n18117 ;
  assign y4671 = ~1'b0 ;
  assign y4672 = ~1'b0 ;
  assign y4673 = n18118 ;
  assign y4674 = n18135 ;
  assign y4675 = ~n18139 ;
  assign y4676 = ~n18141 ;
  assign y4677 = ~n18145 ;
  assign y4678 = n18147 ;
  assign y4679 = n18150 ;
  assign y4680 = n18152 ;
  assign y4681 = n18160 ;
  assign y4682 = ~n7843 ;
  assign y4683 = ~n18163 ;
  assign y4684 = ~n18167 ;
  assign y4685 = ~n18172 ;
  assign y4686 = n18177 ;
  assign y4687 = ~n18186 ;
  assign y4688 = n18188 ;
  assign y4689 = ~n18189 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = ~n18190 ;
  assign y4692 = ~n18196 ;
  assign y4693 = n18199 ;
  assign y4694 = n18205 ;
  assign y4695 = ~n18209 ;
  assign y4696 = ~n18211 ;
  assign y4697 = ~n18212 ;
  assign y4698 = ~1'b0 ;
  assign y4699 = n18219 ;
  assign y4700 = ~n18224 ;
  assign y4701 = ~1'b0 ;
  assign y4702 = ~n18227 ;
  assign y4703 = ~n18228 ;
  assign y4704 = ~n18229 ;
  assign y4705 = ~1'b0 ;
  assign y4706 = n18248 ;
  assign y4707 = n18249 ;
  assign y4708 = ~n18252 ;
  assign y4709 = ~n4888 ;
  assign y4710 = ~n18253 ;
  assign y4711 = ~n18257 ;
  assign y4712 = n18258 ;
  assign y4713 = ~n18262 ;
  assign y4714 = ~1'b0 ;
  assign y4715 = ~1'b0 ;
  assign y4716 = n18265 ;
  assign y4717 = ~n18269 ;
  assign y4718 = ~n18272 ;
  assign y4719 = ~n18276 ;
  assign y4720 = ~n18277 ;
  assign y4721 = ~1'b0 ;
  assign y4722 = ~1'b0 ;
  assign y4723 = n18279 ;
  assign y4724 = n18281 ;
  assign y4725 = n18293 ;
  assign y4726 = ~1'b0 ;
  assign y4727 = n18295 ;
  assign y4728 = n18299 ;
  assign y4729 = ~n18300 ;
  assign y4730 = ~n18301 ;
  assign y4731 = ~n18304 ;
  assign y4732 = n18308 ;
  assign y4733 = ~n18311 ;
  assign y4734 = n18316 ;
  assign y4735 = ~1'b0 ;
  assign y4736 = ~1'b0 ;
  assign y4737 = ~n18321 ;
  assign y4738 = ~n18323 ;
  assign y4739 = ~1'b0 ;
  assign y4740 = ~1'b0 ;
  assign y4741 = ~n18327 ;
  assign y4742 = n18332 ;
  assign y4743 = n18335 ;
  assign y4744 = ~n18340 ;
  assign y4745 = ~n18346 ;
  assign y4746 = n18348 ;
  assign y4747 = ~1'b0 ;
  assign y4748 = n18351 ;
  assign y4749 = n18354 ;
  assign y4750 = n18356 ;
  assign y4751 = ~n18365 ;
  assign y4752 = n18369 ;
  assign y4753 = ~n18371 ;
  assign y4754 = ~n18373 ;
  assign y4755 = ~n18376 ;
  assign y4756 = ~1'b0 ;
  assign y4757 = ~n18377 ;
  assign y4758 = ~n18379 ;
  assign y4759 = ~n18380 ;
  assign y4760 = n18389 ;
  assign y4761 = n18396 ;
  assign y4762 = ~n18399 ;
  assign y4763 = ~n18405 ;
  assign y4764 = n18411 ;
  assign y4765 = ~n18417 ;
  assign y4766 = ~n18419 ;
  assign y4767 = ~n18421 ;
  assign y4768 = ~n18426 ;
  assign y4769 = ~n18430 ;
  assign y4770 = n18435 ;
  assign y4771 = ~n18438 ;
  assign y4772 = ~n18439 ;
  assign y4773 = n18446 ;
  assign y4774 = ~n18448 ;
  assign y4775 = n18450 ;
  assign y4776 = ~n18457 ;
  assign y4777 = n18460 ;
  assign y4778 = ~n18462 ;
  assign y4779 = ~n18463 ;
  assign y4780 = ~n18464 ;
  assign y4781 = n18465 ;
  assign y4782 = ~1'b0 ;
  assign y4783 = n18468 ;
  assign y4784 = ~n18470 ;
  assign y4785 = n18473 ;
  assign y4786 = n18476 ;
  assign y4787 = ~n18480 ;
  assign y4788 = n18481 ;
  assign y4789 = n18482 ;
  assign y4790 = n18487 ;
  assign y4791 = ~n18488 ;
  assign y4792 = ~1'b0 ;
  assign y4793 = ~n18496 ;
  assign y4794 = n18497 ;
  assign y4795 = n18499 ;
  assign y4796 = ~n18504 ;
  assign y4797 = n18508 ;
  assign y4798 = ~n18512 ;
  assign y4799 = ~n18513 ;
  assign y4800 = ~1'b0 ;
  assign y4801 = n18518 ;
  assign y4802 = ~n18524 ;
  assign y4803 = n18525 ;
  assign y4804 = n18527 ;
  assign y4805 = n18532 ;
  assign y4806 = n18533 ;
  assign y4807 = n18537 ;
  assign y4808 = n18545 ;
  assign y4809 = n18548 ;
  assign y4810 = ~n18550 ;
  assign y4811 = n18551 ;
  assign y4812 = ~1'b0 ;
  assign y4813 = ~n18554 ;
  assign y4814 = ~n18555 ;
  assign y4815 = ~n18558 ;
  assign y4816 = n18559 ;
  assign y4817 = ~n18560 ;
  assign y4818 = ~n18564 ;
  assign y4819 = n18570 ;
  assign y4820 = n18573 ;
  assign y4821 = n18575 ;
  assign y4822 = n18577 ;
  assign y4823 = n18579 ;
  assign y4824 = n18582 ;
  assign y4825 = ~n18584 ;
  assign y4826 = n18590 ;
  assign y4827 = ~1'b0 ;
  assign y4828 = n18593 ;
  assign y4829 = ~n18596 ;
  assign y4830 = ~n18605 ;
  assign y4831 = n18606 ;
  assign y4832 = n18607 ;
  assign y4833 = n18609 ;
  assign y4834 = ~1'b0 ;
  assign y4835 = n18610 ;
  assign y4836 = n18616 ;
  assign y4837 = n18617 ;
  assign y4838 = n18619 ;
  assign y4839 = ~n18620 ;
  assign y4840 = ~n18621 ;
  assign y4841 = ~n18624 ;
  assign y4842 = ~n18626 ;
  assign y4843 = ~n18627 ;
  assign y4844 = ~n18631 ;
  assign y4845 = ~1'b0 ;
  assign y4846 = ~n18633 ;
  assign y4847 = n18634 ;
  assign y4848 = n18636 ;
  assign y4849 = n18643 ;
  assign y4850 = n18644 ;
  assign y4851 = ~n18647 ;
  assign y4852 = n18649 ;
  assign y4853 = n18651 ;
  assign y4854 = n18654 ;
  assign y4855 = ~n18656 ;
  assign y4856 = ~n18658 ;
  assign y4857 = ~n18661 ;
  assign y4858 = n18663 ;
  assign y4859 = n18665 ;
  assign y4860 = ~n18668 ;
  assign y4861 = n18669 ;
  assign y4862 = ~n18670 ;
  assign y4863 = ~1'b0 ;
  assign y4864 = ~n18672 ;
  assign y4865 = 1'b0 ;
  assign y4866 = ~n18675 ;
  assign y4867 = n18676 ;
  assign y4868 = ~n18680 ;
  assign y4869 = ~n18682 ;
  assign y4870 = n18613 ;
  assign y4871 = ~n18685 ;
  assign y4872 = n18688 ;
  assign y4873 = n18690 ;
  assign y4874 = ~1'b0 ;
  assign y4875 = n18695 ;
  assign y4876 = n18696 ;
  assign y4877 = ~n18700 ;
  assign y4878 = n18704 ;
  assign y4879 = ~n18708 ;
  assign y4880 = ~n18710 ;
  assign y4881 = n18716 ;
  assign y4882 = n18717 ;
  assign y4883 = n18722 ;
  assign y4884 = ~n18726 ;
  assign y4885 = ~n18732 ;
  assign y4886 = n15872 ;
  assign y4887 = ~n18737 ;
  assign y4888 = n18738 ;
  assign y4889 = ~1'b0 ;
  assign y4890 = ~n18739 ;
  assign y4891 = ~n18742 ;
  assign y4892 = n18743 ;
  assign y4893 = n18746 ;
  assign y4894 = ~n18747 ;
  assign y4895 = ~n18750 ;
  assign y4896 = n18757 ;
  assign y4897 = ~n18760 ;
  assign y4898 = ~n18762 ;
  assign y4899 = ~n18764 ;
  assign y4900 = n18766 ;
  assign y4901 = ~1'b0 ;
  assign y4902 = ~n18769 ;
  assign y4903 = ~n18770 ;
  assign y4904 = ~n18771 ;
  assign y4905 = ~n18772 ;
  assign y4906 = ~n18773 ;
  assign y4907 = ~n18775 ;
  assign y4908 = n18777 ;
  assign y4909 = ~n18781 ;
  assign y4910 = ~n18784 ;
  assign y4911 = ~n18786 ;
  assign y4912 = ~n18788 ;
  assign y4913 = ~n18790 ;
  assign y4914 = n18792 ;
  assign y4915 = n18793 ;
  assign y4916 = n18796 ;
  assign y4917 = ~n18798 ;
  assign y4918 = n18799 ;
  assign y4919 = n18802 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = ~1'b0 ;
  assign y4922 = n18808 ;
  assign y4923 = ~n18809 ;
  assign y4924 = ~n18812 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = ~n18816 ;
  assign y4927 = ~n18817 ;
  assign y4928 = n18818 ;
  assign y4929 = ~n18821 ;
  assign y4930 = n18822 ;
  assign y4931 = ~1'b0 ;
  assign y4932 = ~n18823 ;
  assign y4933 = n18824 ;
  assign y4934 = ~n17921 ;
  assign y4935 = ~n18826 ;
  assign y4936 = ~n18828 ;
  assign y4937 = n18833 ;
  assign y4938 = n18835 ;
  assign y4939 = n18839 ;
  assign y4940 = ~n18841 ;
  assign y4941 = ~n18842 ;
  assign y4942 = ~1'b0 ;
  assign y4943 = n18848 ;
  assign y4944 = ~n18853 ;
  assign y4945 = ~n18856 ;
  assign y4946 = n18858 ;
  assign y4947 = ~1'b0 ;
  assign y4948 = n18860 ;
  assign y4949 = n18866 ;
  assign y4950 = n18869 ;
  assign y4951 = ~1'b0 ;
  assign y4952 = ~n18873 ;
  assign y4953 = ~n18874 ;
  assign y4954 = n18887 ;
  assign y4955 = n18896 ;
  assign y4956 = ~n18897 ;
  assign y4957 = ~n18906 ;
  assign y4958 = ~n18907 ;
  assign y4959 = n18908 ;
  assign y4960 = ~n18909 ;
  assign y4961 = ~n18911 ;
  assign y4962 = ~1'b0 ;
  assign y4963 = n18915 ;
  assign y4964 = ~1'b0 ;
  assign y4965 = n18924 ;
  assign y4966 = n18925 ;
  assign y4967 = n18931 ;
  assign y4968 = ~n18937 ;
  assign y4969 = ~n18939 ;
  assign y4970 = ~n18940 ;
  assign y4971 = n18943 ;
  assign y4972 = ~1'b0 ;
  assign y4973 = ~n18947 ;
  assign y4974 = n18949 ;
  assign y4975 = ~1'b0 ;
  assign y4976 = ~n18954 ;
  assign y4977 = n18955 ;
  assign y4978 = ~n18959 ;
  assign y4979 = n18963 ;
  assign y4980 = ~n18965 ;
  assign y4981 = ~n18968 ;
  assign y4982 = n18970 ;
  assign y4983 = n3747 ;
  assign y4984 = ~n18973 ;
  assign y4985 = n18974 ;
  assign y4986 = ~1'b0 ;
  assign y4987 = n18978 ;
  assign y4988 = n18985 ;
  assign y4989 = n18986 ;
  assign y4990 = n18987 ;
  assign y4991 = ~n18996 ;
  assign y4992 = ~n18997 ;
  assign y4993 = n19003 ;
  assign y4994 = ~1'b0 ;
  assign y4995 = ~n19004 ;
  assign y4996 = ~n19009 ;
  assign y4997 = ~n19011 ;
  assign y4998 = n19012 ;
  assign y4999 = ~n19016 ;
  assign y5000 = ~n19019 ;
  assign y5001 = ~n19020 ;
  assign y5002 = ~n19024 ;
  assign y5003 = n19025 ;
  assign y5004 = n19029 ;
  assign y5005 = n19030 ;
  assign y5006 = ~n19033 ;
  assign y5007 = ~n19035 ;
  assign y5008 = ~n19038 ;
  assign y5009 = n19051 ;
  assign y5010 = ~n19052 ;
  assign y5011 = ~n19057 ;
  assign y5012 = n19060 ;
  assign y5013 = ~n19061 ;
  assign y5014 = n19066 ;
  assign y5015 = ~1'b0 ;
  assign y5016 = ~n19071 ;
  assign y5017 = ~n19073 ;
  assign y5018 = n19075 ;
  assign y5019 = ~n19079 ;
  assign y5020 = ~n19081 ;
  assign y5021 = n19082 ;
  assign y5022 = n19089 ;
  assign y5023 = ~1'b0 ;
  assign y5024 = ~n19096 ;
  assign y5025 = n19102 ;
  assign y5026 = n19108 ;
  assign y5027 = n19109 ;
  assign y5028 = n19110 ;
  assign y5029 = ~1'b0 ;
  assign y5030 = n19113 ;
  assign y5031 = ~n19114 ;
  assign y5032 = n19119 ;
  assign y5033 = ~n19121 ;
  assign y5034 = n19123 ;
  assign y5035 = ~n19124 ;
  assign y5036 = n18811 ;
  assign y5037 = ~n19125 ;
  assign y5038 = n19130 ;
  assign y5039 = ~n19131 ;
  assign y5040 = ~n19134 ;
  assign y5041 = ~n19146 ;
  assign y5042 = ~n19147 ;
  assign y5043 = ~n19148 ;
  assign y5044 = n19149 ;
  assign y5045 = ~n19151 ;
  assign y5046 = ~1'b0 ;
  assign y5047 = ~n19164 ;
  assign y5048 = n19167 ;
  assign y5049 = n19170 ;
  assign y5050 = n19176 ;
  assign y5051 = ~n19177 ;
  assign y5052 = n19180 ;
  assign y5053 = ~n19184 ;
  assign y5054 = ~n19188 ;
  assign y5055 = n19190 ;
  assign y5056 = ~n19194 ;
  assign y5057 = ~n19195 ;
  assign y5058 = ~n19197 ;
  assign y5059 = ~n19200 ;
  assign y5060 = ~n19203 ;
  assign y5061 = ~n19206 ;
  assign y5062 = n19212 ;
  assign y5063 = ~n19213 ;
  assign y5064 = n19216 ;
  assign y5065 = n19217 ;
  assign y5066 = ~n19218 ;
  assign y5067 = n19221 ;
  assign y5068 = n19227 ;
  assign y5069 = ~1'b0 ;
  assign y5070 = n19231 ;
  assign y5071 = n19235 ;
  assign y5072 = ~n19237 ;
  assign y5073 = n19238 ;
  assign y5074 = ~n19239 ;
  assign y5075 = n19244 ;
  assign y5076 = ~n19248 ;
  assign y5077 = ~n19250 ;
  assign y5078 = n19251 ;
  assign y5079 = ~n19255 ;
  assign y5080 = ~n19260 ;
  assign y5081 = ~n19267 ;
  assign y5082 = n19269 ;
  assign y5083 = ~n19274 ;
  assign y5084 = ~n19278 ;
  assign y5085 = n19285 ;
  assign y5086 = n19286 ;
  assign y5087 = n19288 ;
  assign y5088 = n19290 ;
  assign y5089 = n19292 ;
  assign y5090 = ~n19299 ;
  assign y5091 = n19302 ;
  assign y5092 = n19303 ;
  assign y5093 = n19305 ;
  assign y5094 = n19306 ;
  assign y5095 = ~n19308 ;
  assign y5096 = n19312 ;
  assign y5097 = ~n19313 ;
  assign y5098 = ~n19319 ;
  assign y5099 = ~1'b0 ;
  assign y5100 = n19320 ;
  assign y5101 = n19321 ;
  assign y5102 = n19323 ;
  assign y5103 = ~n19324 ;
  assign y5104 = n19326 ;
  assign y5105 = n19333 ;
  assign y5106 = ~n19337 ;
  assign y5107 = n19347 ;
  assign y5108 = n19349 ;
  assign y5109 = ~n19352 ;
  assign y5110 = ~1'b0 ;
  assign y5111 = n19353 ;
  assign y5112 = ~n19354 ;
  assign y5113 = ~n19359 ;
  assign y5114 = n19361 ;
  assign y5115 = ~n19364 ;
  assign y5116 = n19367 ;
  assign y5117 = n19372 ;
  assign y5118 = n19379 ;
  assign y5119 = n19381 ;
  assign y5120 = n19383 ;
  assign y5121 = n19389 ;
  assign y5122 = ~n19390 ;
  assign y5123 = n19393 ;
  assign y5124 = ~n19396 ;
  assign y5125 = ~n19398 ;
  assign y5126 = ~n19403 ;
  assign y5127 = ~n19406 ;
  assign y5128 = ~n19410 ;
  assign y5129 = ~1'b0 ;
  assign y5130 = ~n19413 ;
  assign y5131 = n19417 ;
  assign y5132 = ~n19423 ;
  assign y5133 = ~n19427 ;
  assign y5134 = ~n19428 ;
  assign y5135 = ~n19429 ;
  assign y5136 = ~n19431 ;
  assign y5137 = ~n19438 ;
  assign y5138 = n19443 ;
  assign y5139 = n19445 ;
  assign y5140 = n19446 ;
  assign y5141 = n19450 ;
  assign y5142 = n19451 ;
  assign y5143 = n19455 ;
  assign y5144 = ~n19458 ;
  assign y5145 = ~1'b0 ;
  assign y5146 = n19460 ;
  assign y5147 = n19466 ;
  assign y5148 = ~n19469 ;
  assign y5149 = ~n19470 ;
  assign y5150 = ~n19474 ;
  assign y5151 = n19480 ;
  assign y5152 = ~n19484 ;
  assign y5153 = n19485 ;
  assign y5154 = ~n19486 ;
  assign y5155 = n19488 ;
  assign y5156 = n19493 ;
  assign y5157 = n19497 ;
  assign y5158 = ~n19498 ;
  assign y5159 = ~n19500 ;
  assign y5160 = ~n19505 ;
  assign y5161 = n19506 ;
  assign y5162 = n19508 ;
  assign y5163 = ~n19509 ;
  assign y5164 = ~n19510 ;
  assign y5165 = ~1'b0 ;
  assign y5166 = n19518 ;
  assign y5167 = ~n19520 ;
  assign y5168 = ~n19521 ;
  assign y5169 = ~n19526 ;
  assign y5170 = n19527 ;
  assign y5171 = n19528 ;
  assign y5172 = ~n19531 ;
  assign y5173 = ~n19538 ;
  assign y5174 = n19543 ;
  assign y5175 = ~n19552 ;
  assign y5176 = n19553 ;
  assign y5177 = ~n19556 ;
  assign y5178 = ~n19558 ;
  assign y5179 = ~n19562 ;
  assign y5180 = ~n19563 ;
  assign y5181 = ~1'b0 ;
  assign y5182 = ~n19565 ;
  assign y5183 = n19566 ;
  assign y5184 = ~n19567 ;
  assign y5185 = n19571 ;
  assign y5186 = ~1'b0 ;
  assign y5187 = n19572 ;
  assign y5188 = ~n19581 ;
  assign y5189 = n19582 ;
  assign y5190 = ~1'b0 ;
  assign y5191 = n19586 ;
  assign y5192 = n19587 ;
  assign y5193 = ~n19588 ;
  assign y5194 = ~n19590 ;
  assign y5195 = n19592 ;
  assign y5196 = ~n19594 ;
  assign y5197 = ~n19596 ;
  assign y5198 = ~n19602 ;
  assign y5199 = ~n19603 ;
  assign y5200 = ~n19604 ;
  assign y5201 = ~n19605 ;
  assign y5202 = n19609 ;
  assign y5203 = n19611 ;
  assign y5204 = n19614 ;
  assign y5205 = ~n19623 ;
  assign y5206 = ~1'b0 ;
  assign y5207 = n19625 ;
  assign y5208 = n19629 ;
  assign y5209 = n19630 ;
  assign y5210 = ~n19631 ;
  assign y5211 = ~n19634 ;
  assign y5212 = ~n19636 ;
  assign y5213 = ~1'b0 ;
  assign y5214 = n19639 ;
  assign y5215 = ~n19650 ;
  assign y5216 = n19651 ;
  assign y5217 = ~n19654 ;
  assign y5218 = ~1'b0 ;
  assign y5219 = n19657 ;
  assign y5220 = ~n19660 ;
  assign y5221 = ~n19661 ;
  assign y5222 = ~n19662 ;
  assign y5223 = ~n19663 ;
  assign y5224 = ~n19665 ;
  assign y5225 = ~n19669 ;
  assign y5226 = n19675 ;
  assign y5227 = ~n19676 ;
  assign y5228 = n19677 ;
  assign y5229 = ~n19679 ;
  assign y5230 = n19685 ;
  assign y5231 = ~1'b0 ;
  assign y5232 = n19688 ;
  assign y5233 = ~n19689 ;
  assign y5234 = n19691 ;
  assign y5235 = n19701 ;
  assign y5236 = n19703 ;
  assign y5237 = ~1'b0 ;
  assign y5238 = n19707 ;
  assign y5239 = n19709 ;
  assign y5240 = n19711 ;
  assign y5241 = ~n19716 ;
  assign y5242 = ~n19717 ;
  assign y5243 = ~n19721 ;
  assign y5244 = ~n19723 ;
  assign y5245 = ~n19727 ;
  assign y5246 = n19729 ;
  assign y5247 = ~n19731 ;
  assign y5248 = ~n19734 ;
  assign y5249 = n19738 ;
  assign y5250 = n19740 ;
  assign y5251 = ~n19741 ;
  assign y5252 = n19744 ;
  assign y5253 = n19747 ;
  assign y5254 = ~n19750 ;
  assign y5255 = ~n19754 ;
  assign y5256 = n19756 ;
  assign y5257 = ~n19771 ;
  assign y5258 = n19772 ;
  assign y5259 = ~n19775 ;
  assign y5260 = n19778 ;
  assign y5261 = n19780 ;
  assign y5262 = ~1'b0 ;
  assign y5263 = ~1'b0 ;
  assign y5264 = n19781 ;
  assign y5265 = n19783 ;
  assign y5266 = ~n19784 ;
  assign y5267 = ~n19790 ;
  assign y5268 = n19545 ;
  assign y5269 = ~n19792 ;
  assign y5270 = ~1'b0 ;
  assign y5271 = ~n19799 ;
  assign y5272 = n19800 ;
  assign y5273 = ~n19803 ;
  assign y5274 = ~n19804 ;
  assign y5275 = n19806 ;
  assign y5276 = ~n19807 ;
  assign y5277 = n19811 ;
  assign y5278 = n19813 ;
  assign y5279 = ~n19814 ;
  assign y5280 = n19817 ;
  assign y5281 = ~n19819 ;
  assign y5282 = ~n19820 ;
  assign y5283 = ~1'b0 ;
  assign y5284 = ~n19822 ;
  assign y5285 = n19823 ;
  assign y5286 = ~n19825 ;
  assign y5287 = ~n19826 ;
  assign y5288 = n19827 ;
  assign y5289 = ~1'b0 ;
  assign y5290 = ~1'b0 ;
  assign y5291 = ~n19831 ;
  assign y5292 = ~n19833 ;
  assign y5293 = ~n19836 ;
  assign y5294 = ~n19843 ;
  assign y5295 = n19847 ;
  assign y5296 = ~n19848 ;
  assign y5297 = ~1'b0 ;
  assign y5298 = ~n19850 ;
  assign y5299 = ~n14039 ;
  assign y5300 = n19851 ;
  assign y5301 = ~n19853 ;
  assign y5302 = n19855 ;
  assign y5303 = ~n19856 ;
  assign y5304 = ~n19858 ;
  assign y5305 = n19859 ;
  assign y5306 = ~n19863 ;
  assign y5307 = n19865 ;
  assign y5308 = n19870 ;
  assign y5309 = ~n19877 ;
  assign y5310 = n19886 ;
  assign y5311 = n19887 ;
  assign y5312 = n19891 ;
  assign y5313 = ~n19895 ;
  assign y5314 = n19898 ;
  assign y5315 = ~n19900 ;
  assign y5316 = ~1'b0 ;
  assign y5317 = n19901 ;
  assign y5318 = ~n19907 ;
  assign y5319 = ~n19909 ;
  assign y5320 = n19912 ;
  assign y5321 = ~n19916 ;
  assign y5322 = ~n19917 ;
  assign y5323 = n19918 ;
  assign y5324 = ~1'b0 ;
  assign y5325 = n19921 ;
  assign y5326 = ~n19925 ;
  assign y5327 = n19927 ;
  assign y5328 = ~n19936 ;
  assign y5329 = ~n19940 ;
  assign y5330 = n19943 ;
  assign y5331 = ~n19946 ;
  assign y5332 = n19954 ;
  assign y5333 = n19957 ;
  assign y5334 = n19960 ;
  assign y5335 = n19961 ;
  assign y5336 = ~n19962 ;
  assign y5337 = ~n19965 ;
  assign y5338 = ~n19968 ;
  assign y5339 = n19973 ;
  assign y5340 = ~1'b0 ;
  assign y5341 = n19974 ;
  assign y5342 = n19977 ;
  assign y5343 = ~n19980 ;
  assign y5344 = n19981 ;
  assign y5345 = ~1'b0 ;
  assign y5346 = ~n19982 ;
  assign y5347 = ~n19986 ;
  assign y5348 = n19989 ;
  assign y5349 = ~n19996 ;
  assign y5350 = ~n19998 ;
  assign y5351 = ~1'b0 ;
  assign y5352 = ~1'b0 ;
  assign y5353 = ~n7335 ;
  assign y5354 = n19999 ;
  assign y5355 = n20000 ;
  assign y5356 = n20001 ;
  assign y5357 = n20002 ;
  assign y5358 = n20004 ;
  assign y5359 = ~n20008 ;
  assign y5360 = n20012 ;
  assign y5361 = ~n20017 ;
  assign y5362 = ~n20018 ;
  assign y5363 = n20019 ;
  assign y5364 = ~1'b0 ;
  assign y5365 = ~n20020 ;
  assign y5366 = n20025 ;
  assign y5367 = n20028 ;
  assign y5368 = ~n20029 ;
  assign y5369 = n20033 ;
  assign y5370 = ~n20035 ;
  assign y5371 = ~n20037 ;
  assign y5372 = ~n20039 ;
  assign y5373 = n20041 ;
  assign y5374 = n20045 ;
  assign y5375 = ~n20047 ;
  assign y5376 = n20048 ;
  assign y5377 = n20049 ;
  assign y5378 = n20060 ;
  assign y5379 = ~1'b0 ;
  assign y5380 = n20063 ;
  assign y5381 = ~n20064 ;
  assign y5382 = ~n20065 ;
  assign y5383 = n20067 ;
  assign y5384 = n20070 ;
  assign y5385 = n20071 ;
  assign y5386 = ~n20075 ;
  assign y5387 = ~n20081 ;
  assign y5388 = ~n20083 ;
  assign y5389 = n20084 ;
  assign y5390 = ~n20088 ;
  assign y5391 = n20090 ;
  assign y5392 = ~n20095 ;
  assign y5393 = ~n20097 ;
  assign y5394 = n20106 ;
  assign y5395 = n20116 ;
  assign y5396 = ~n20121 ;
  assign y5397 = ~n20122 ;
  assign y5398 = ~n20127 ;
  assign y5399 = n20128 ;
  assign y5400 = ~n20130 ;
  assign y5401 = ~n20131 ;
  assign y5402 = ~n20132 ;
  assign y5403 = ~n17680 ;
  assign y5404 = ~n20134 ;
  assign y5405 = ~n20137 ;
  assign y5406 = ~n20138 ;
  assign y5407 = ~n20139 ;
  assign y5408 = ~n20140 ;
  assign y5409 = ~n20144 ;
  assign y5410 = ~n20145 ;
  assign y5411 = ~1'b0 ;
  assign y5412 = ~1'b0 ;
  assign y5413 = n20147 ;
  assign y5414 = n20153 ;
  assign y5415 = ~n20156 ;
  assign y5416 = ~n20158 ;
  assign y5417 = ~1'b0 ;
  assign y5418 = n20161 ;
  assign y5419 = n20166 ;
  assign y5420 = n20171 ;
  assign y5421 = ~n15368 ;
  assign y5422 = n20177 ;
  assign y5423 = ~1'b0 ;
  assign y5424 = ~n20179 ;
  assign y5425 = ~1'b0 ;
  assign y5426 = ~n20182 ;
  assign y5427 = ~n20183 ;
  assign y5428 = n20192 ;
  assign y5429 = n20195 ;
  assign y5430 = n20196 ;
  assign y5431 = n20200 ;
  assign y5432 = n20203 ;
  assign y5433 = n20205 ;
  assign y5434 = ~n18736 ;
  assign y5435 = ~1'b0 ;
  assign y5436 = ~n20207 ;
  assign y5437 = ~1'b0 ;
  assign y5438 = ~n20208 ;
  assign y5439 = ~n20210 ;
  assign y5440 = ~n20213 ;
  assign y5441 = n20217 ;
  assign y5442 = n20223 ;
  assign y5443 = ~n20229 ;
  assign y5444 = ~1'b0 ;
  assign y5445 = n20239 ;
  assign y5446 = n20241 ;
  assign y5447 = ~n20246 ;
  assign y5448 = n20254 ;
  assign y5449 = ~n20256 ;
  assign y5450 = ~n20262 ;
  assign y5451 = n20264 ;
  assign y5452 = ~n20265 ;
  assign y5453 = ~n20270 ;
  assign y5454 = n20273 ;
  assign y5455 = n20276 ;
  assign y5456 = n20279 ;
  assign y5457 = ~n20281 ;
  assign y5458 = ~n20284 ;
  assign y5459 = ~n20287 ;
  assign y5460 = n20289 ;
  assign y5461 = ~n20291 ;
  assign y5462 = n20296 ;
  assign y5463 = n20297 ;
  assign y5464 = ~n20300 ;
  assign y5465 = ~1'b0 ;
  assign y5466 = ~1'b0 ;
  assign y5467 = ~n20302 ;
  assign y5468 = ~n20303 ;
  assign y5469 = ~n20304 ;
  assign y5470 = ~n20307 ;
  assign y5471 = n20308 ;
  assign y5472 = n20309 ;
  assign y5473 = n20311 ;
  assign y5474 = n20316 ;
  assign y5475 = n20318 ;
  assign y5476 = n20323 ;
  assign y5477 = ~n20326 ;
  assign y5478 = n20330 ;
  assign y5479 = ~n20336 ;
  assign y5480 = ~n20338 ;
  assign y5481 = n20342 ;
  assign y5482 = ~1'b0 ;
  assign y5483 = n20344 ;
  assign y5484 = n20345 ;
  assign y5485 = n20346 ;
  assign y5486 = n20347 ;
  assign y5487 = ~n20348 ;
  assign y5488 = n20350 ;
  assign y5489 = n20353 ;
  assign y5490 = n20357 ;
  assign y5491 = ~n20365 ;
  assign y5492 = ~n20367 ;
  assign y5493 = n20369 ;
  assign y5494 = n20373 ;
  assign y5495 = n20374 ;
  assign y5496 = ~n20378 ;
  assign y5497 = ~1'b0 ;
  assign y5498 = ~n20379 ;
  assign y5499 = n20388 ;
  assign y5500 = ~1'b0 ;
  assign y5501 = ~n20389 ;
  assign y5502 = ~n20392 ;
  assign y5503 = n20394 ;
  assign y5504 = n20404 ;
  assign y5505 = ~n20406 ;
  assign y5506 = n20408 ;
  assign y5507 = ~n20409 ;
  assign y5508 = ~n20411 ;
  assign y5509 = n20415 ;
  assign y5510 = ~n20422 ;
  assign y5511 = ~n20423 ;
  assign y5512 = ~n20427 ;
  assign y5513 = ~n20428 ;
  assign y5514 = ~n20432 ;
  assign y5515 = ~1'b0 ;
  assign y5516 = n20435 ;
  assign y5517 = ~n20437 ;
  assign y5518 = n20450 ;
  assign y5519 = n20452 ;
  assign y5520 = ~n20455 ;
  assign y5521 = n20458 ;
  assign y5522 = ~n20459 ;
  assign y5523 = ~n20460 ;
  assign y5524 = ~n20463 ;
  assign y5525 = ~n20466 ;
  assign y5526 = ~n20472 ;
  assign y5527 = n20476 ;
  assign y5528 = n20480 ;
  assign y5529 = ~n20487 ;
  assign y5530 = n20489 ;
  assign y5531 = ~n20491 ;
  assign y5532 = n20496 ;
  assign y5533 = n20500 ;
  assign y5534 = n20501 ;
  assign y5535 = n20504 ;
  assign y5536 = ~n20505 ;
  assign y5537 = ~n20507 ;
  assign y5538 = ~n20515 ;
  assign y5539 = ~n20520 ;
  assign y5540 = ~n20521 ;
  assign y5541 = ~n20525 ;
  assign y5542 = ~n20526 ;
  assign y5543 = ~1'b0 ;
  assign y5544 = ~n20528 ;
  assign y5545 = n20534 ;
  assign y5546 = ~n20536 ;
  assign y5547 = ~n20542 ;
  assign y5548 = ~n20547 ;
  assign y5549 = ~n20552 ;
  assign y5550 = n20553 ;
  assign y5551 = n20556 ;
  assign y5552 = ~n20563 ;
  assign y5553 = n20570 ;
  assign y5554 = ~n20574 ;
  assign y5555 = ~n20581 ;
  assign y5556 = ~n20582 ;
  assign y5557 = ~n20585 ;
  assign y5558 = n20588 ;
  assign y5559 = ~n20592 ;
  assign y5560 = ~1'b0 ;
  assign y5561 = ~n20597 ;
  assign y5562 = ~n20604 ;
  assign y5563 = ~n20605 ;
  assign y5564 = ~n20607 ;
  assign y5565 = n20625 ;
  assign y5566 = ~1'b0 ;
  assign y5567 = ~n20630 ;
  assign y5568 = n20631 ;
  assign y5569 = n20636 ;
  assign y5570 = ~n20637 ;
  assign y5571 = n20638 ;
  assign y5572 = ~n20640 ;
  assign y5573 = n20646 ;
  assign y5574 = ~n20648 ;
  assign y5575 = n20652 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = n20657 ;
  assign y5578 = n20663 ;
  assign y5579 = n20667 ;
  assign y5580 = n20671 ;
  assign y5581 = n20672 ;
  assign y5582 = n20676 ;
  assign y5583 = n20680 ;
  assign y5584 = n20683 ;
  assign y5585 = ~n20688 ;
  assign y5586 = n20689 ;
  assign y5587 = ~n20693 ;
  assign y5588 = ~1'b0 ;
  assign y5589 = ~n20695 ;
  assign y5590 = ~n20697 ;
  assign y5591 = ~n20698 ;
  assign y5592 = ~n20705 ;
  assign y5593 = n20708 ;
  assign y5594 = n20709 ;
  assign y5595 = ~n20711 ;
  assign y5596 = n20719 ;
  assign y5597 = n20724 ;
  assign y5598 = ~n20728 ;
  assign y5599 = n20729 ;
  assign y5600 = ~n20732 ;
  assign y5601 = ~n20734 ;
  assign y5602 = ~1'b0 ;
  assign y5603 = ~n20737 ;
  assign y5604 = ~n20738 ;
  assign y5605 = n20740 ;
  assign y5606 = ~1'b0 ;
  assign y5607 = ~n20744 ;
  assign y5608 = ~n20746 ;
  assign y5609 = ~n20747 ;
  assign y5610 = n20751 ;
  assign y5611 = n20755 ;
  assign y5612 = ~n20759 ;
  assign y5613 = n10254 ;
  assign y5614 = ~n20761 ;
  assign y5615 = n20763 ;
  assign y5616 = ~1'b0 ;
  assign y5617 = ~n20768 ;
  assign y5618 = n20769 ;
  assign y5619 = ~n20774 ;
  assign y5620 = n20777 ;
  assign y5621 = n20779 ;
  assign y5622 = ~n20781 ;
  assign y5623 = ~n20783 ;
  assign y5624 = n20785 ;
  assign y5625 = n20787 ;
  assign y5626 = ~n20788 ;
  assign y5627 = ~n20791 ;
  assign y5628 = n20793 ;
  assign y5629 = ~n20795 ;
  assign y5630 = ~1'b0 ;
  assign y5631 = n20800 ;
  assign y5632 = ~n20802 ;
  assign y5633 = ~n20814 ;
  assign y5634 = ~1'b0 ;
  assign y5635 = ~n20816 ;
  assign y5636 = n20822 ;
  assign y5637 = n20823 ;
  assign y5638 = ~n20826 ;
  assign y5639 = ~n20831 ;
  assign y5640 = ~n20833 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = ~1'b0 ;
  assign y5643 = n20834 ;
  assign y5644 = ~n20835 ;
  assign y5645 = ~n20836 ;
  assign y5646 = n20839 ;
  assign y5647 = n20840 ;
  assign y5648 = n20841 ;
  assign y5649 = ~n20846 ;
  assign y5650 = ~n20849 ;
  assign y5651 = n20852 ;
  assign y5652 = ~n20853 ;
  assign y5653 = n20857 ;
  assign y5654 = ~n20861 ;
  assign y5655 = ~n20875 ;
  assign y5656 = n20876 ;
  assign y5657 = ~n20880 ;
  assign y5658 = 1'b0 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = ~n20886 ;
  assign y5661 = n20894 ;
  assign y5662 = n20896 ;
  assign y5663 = n20899 ;
  assign y5664 = n20900 ;
  assign y5665 = ~1'b0 ;
  assign y5666 = ~1'b0 ;
  assign y5667 = ~1'b0 ;
  assign y5668 = ~n20901 ;
  assign y5669 = ~n20902 ;
  assign y5670 = ~n20904 ;
  assign y5671 = n20905 ;
  assign y5672 = ~n20906 ;
  assign y5673 = n20915 ;
  assign y5674 = ~n20916 ;
  assign y5675 = n20920 ;
  assign y5676 = ~n20921 ;
  assign y5677 = ~n20924 ;
  assign y5678 = n20932 ;
  assign y5679 = ~n20934 ;
  assign y5680 = ~n20936 ;
  assign y5681 = ~n20938 ;
  assign y5682 = n20945 ;
  assign y5683 = n20948 ;
  assign y5684 = ~n20953 ;
  assign y5685 = ~n20954 ;
  assign y5686 = n20961 ;
  assign y5687 = n20962 ;
  assign y5688 = ~n20965 ;
  assign y5689 = n20969 ;
  assign y5690 = ~n20970 ;
  assign y5691 = ~n20980 ;
  assign y5692 = n20983 ;
  assign y5693 = n20988 ;
  assign y5694 = ~n20996 ;
  assign y5695 = ~n20998 ;
  assign y5696 = ~n21004 ;
  assign y5697 = n21006 ;
  assign y5698 = n21010 ;
  assign y5699 = n21011 ;
  assign y5700 = n21014 ;
  assign y5701 = ~1'b0 ;
  assign y5702 = ~n21019 ;
  assign y5703 = n21025 ;
  assign y5704 = n21027 ;
  assign y5705 = n21031 ;
  assign y5706 = n21033 ;
  assign y5707 = n21034 ;
  assign y5708 = ~n21040 ;
  assign y5709 = ~n21042 ;
  assign y5710 = n21049 ;
  assign y5711 = ~n21055 ;
  assign y5712 = ~n21059 ;
  assign y5713 = ~1'b0 ;
  assign y5714 = ~1'b0 ;
  assign y5715 = n21060 ;
  assign y5716 = ~n21064 ;
  assign y5717 = ~n21068 ;
  assign y5718 = ~n21069 ;
  assign y5719 = ~n21071 ;
  assign y5720 = ~1'b0 ;
  assign y5721 = ~1'b0 ;
  assign y5722 = n21074 ;
  assign y5723 = ~n21077 ;
  assign y5724 = n21078 ;
  assign y5725 = ~n21086 ;
  assign y5726 = ~n21088 ;
  assign y5727 = n21090 ;
  assign y5728 = n21093 ;
  assign y5729 = n21096 ;
  assign y5730 = ~1'b0 ;
  assign y5731 = ~1'b0 ;
  assign y5732 = n21098 ;
  assign y5733 = n21099 ;
  assign y5734 = ~n21100 ;
  assign y5735 = ~n21104 ;
  assign y5736 = ~n21107 ;
  assign y5737 = n21108 ;
  assign y5738 = ~n21110 ;
  assign y5739 = ~n21111 ;
  assign y5740 = ~n21113 ;
  assign y5741 = ~1'b0 ;
  assign y5742 = ~1'b0 ;
  assign y5743 = n21120 ;
  assign y5744 = n21125 ;
  assign y5745 = n21128 ;
  assign y5746 = ~n21129 ;
  assign y5747 = ~n21136 ;
  assign y5748 = ~1'b0 ;
  assign y5749 = n21137 ;
  assign y5750 = n21139 ;
  assign y5751 = ~n21143 ;
  assign y5752 = ~n21154 ;
  assign y5753 = n21157 ;
  assign y5754 = ~n21162 ;
  assign y5755 = ~1'b0 ;
  assign y5756 = n21163 ;
  assign y5757 = n21164 ;
  assign y5758 = n21166 ;
  assign y5759 = ~n21167 ;
  assign y5760 = ~n21169 ;
  assign y5761 = n21171 ;
  assign y5762 = n21177 ;
  assign y5763 = ~1'b0 ;
  assign y5764 = ~n21183 ;
  assign y5765 = ~n21185 ;
  assign y5766 = n21186 ;
  assign y5767 = ~1'b0 ;
  assign y5768 = ~n21188 ;
  assign y5769 = ~1'b0 ;
  assign y5770 = ~n21194 ;
  assign y5771 = ~n21196 ;
  assign y5772 = ~n21197 ;
  assign y5773 = n21198 ;
  assign y5774 = n21199 ;
  assign y5775 = ~n21203 ;
  assign y5776 = ~n21209 ;
  assign y5777 = ~n21210 ;
  assign y5778 = n20621 ;
  assign y5779 = ~n21213 ;
  assign y5780 = n21214 ;
  assign y5781 = ~n21217 ;
  assign y5782 = n21221 ;
  assign y5783 = ~n21222 ;
  assign y5784 = n21225 ;
  assign y5785 = ~n21228 ;
  assign y5786 = n21234 ;
  assign y5787 = ~n21236 ;
  assign y5788 = n21237 ;
  assign y5789 = n21238 ;
  assign y5790 = ~1'b0 ;
  assign y5791 = n21240 ;
  assign y5792 = ~n21242 ;
  assign y5793 = ~n21250 ;
  assign y5794 = ~n21251 ;
  assign y5795 = ~n21252 ;
  assign y5796 = ~n21253 ;
  assign y5797 = ~n21254 ;
  assign y5798 = n21260 ;
  assign y5799 = ~1'b0 ;
  assign y5800 = n21262 ;
  assign y5801 = ~n21266 ;
  assign y5802 = ~n21269 ;
  assign y5803 = ~n21273 ;
  assign y5804 = n21277 ;
  assign y5805 = n21278 ;
  assign y5806 = ~n21279 ;
  assign y5807 = n21281 ;
  assign y5808 = ~n21284 ;
  assign y5809 = ~n21287 ;
  assign y5810 = ~1'b0 ;
  assign y5811 = ~n21289 ;
  assign y5812 = ~n21294 ;
  assign y5813 = ~n458 ;
  assign y5814 = n21295 ;
  assign y5815 = ~n21296 ;
  assign y5816 = n21304 ;
  assign y5817 = ~n21309 ;
  assign y5818 = n21311 ;
  assign y5819 = n21314 ;
  assign y5820 = n21319 ;
  assign y5821 = n21321 ;
  assign y5822 = n21322 ;
  assign y5823 = ~n21325 ;
  assign y5824 = ~1'b0 ;
  assign y5825 = ~n21327 ;
  assign y5826 = n21332 ;
  assign y5827 = n21333 ;
  assign y5828 = ~n21337 ;
  assign y5829 = ~n21340 ;
  assign y5830 = ~n21343 ;
  assign y5831 = ~n21345 ;
  assign y5832 = ~n21347 ;
  assign y5833 = n21351 ;
  assign y5834 = n21358 ;
  assign y5835 = n21364 ;
  assign y5836 = n21365 ;
  assign y5837 = n21369 ;
  assign y5838 = ~n21372 ;
  assign y5839 = ~1'b0 ;
  assign y5840 = n21373 ;
  assign y5841 = n21375 ;
  assign y5842 = n21377 ;
  assign y5843 = n21379 ;
  assign y5844 = ~n21381 ;
  assign y5845 = n21385 ;
  assign y5846 = ~n21387 ;
  assign y5847 = n21389 ;
  assign y5848 = n21392 ;
  assign y5849 = n21395 ;
  assign y5850 = n21397 ;
  assign y5851 = n21400 ;
  assign y5852 = ~1'b0 ;
  assign y5853 = n21401 ;
  assign y5854 = n21403 ;
  assign y5855 = ~n21406 ;
  assign y5856 = ~n21410 ;
  assign y5857 = n21411 ;
  assign y5858 = ~n21413 ;
  assign y5859 = n21414 ;
  assign y5860 = n21416 ;
  assign y5861 = n21419 ;
  assign y5862 = ~n21423 ;
  assign y5863 = n21424 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = ~n21433 ;
  assign y5866 = n21434 ;
  assign y5867 = n21439 ;
  assign y5868 = ~n21440 ;
  assign y5869 = n21446 ;
  assign y5870 = ~n21449 ;
  assign y5871 = ~n21450 ;
  assign y5872 = n21451 ;
  assign y5873 = ~n21457 ;
  assign y5874 = n21459 ;
  assign y5875 = ~1'b0 ;
  assign y5876 = n21462 ;
  assign y5877 = ~n21468 ;
  assign y5878 = n21469 ;
  assign y5879 = n21480 ;
  assign y5880 = n21482 ;
  assign y5881 = n21483 ;
  assign y5882 = ~n21485 ;
  assign y5883 = ~n21491 ;
  assign y5884 = ~n21492 ;
  assign y5885 = n21493 ;
  assign y5886 = n21495 ;
  assign y5887 = ~n21496 ;
  assign y5888 = n21498 ;
  assign y5889 = ~1'b0 ;
  assign y5890 = ~n21506 ;
  assign y5891 = ~n21509 ;
  assign y5892 = ~n21510 ;
  assign y5893 = ~n21515 ;
  assign y5894 = n21516 ;
  assign y5895 = ~n21520 ;
  assign y5896 = ~n21522 ;
  assign y5897 = n21524 ;
  assign y5898 = ~n21526 ;
  assign y5899 = ~1'b0 ;
  assign y5900 = n15218 ;
  assign y5901 = ~n21528 ;
  assign y5902 = ~n21531 ;
  assign y5903 = ~n21536 ;
  assign y5904 = ~n21538 ;
  assign y5905 = ~1'b0 ;
  assign y5906 = ~n21542 ;
  assign y5907 = n21545 ;
  assign y5908 = ~n21549 ;
  assign y5909 = n21552 ;
  assign y5910 = ~n21555 ;
  assign y5911 = ~n21559 ;
  assign y5912 = ~1'b0 ;
  assign y5913 = ~1'b0 ;
  assign y5914 = ~n21561 ;
  assign y5915 = ~n21563 ;
  assign y5916 = n21564 ;
  assign y5917 = ~1'b0 ;
  assign y5918 = ~1'b0 ;
  assign y5919 = n21566 ;
  assign y5920 = ~n21569 ;
  assign y5921 = n21574 ;
  assign y5922 = n21579 ;
  assign y5923 = ~n21580 ;
  assign y5924 = n21581 ;
  assign y5925 = ~n21585 ;
  assign y5926 = ~n21587 ;
  assign y5927 = n21589 ;
  assign y5928 = ~n21596 ;
  assign y5929 = ~n21601 ;
  assign y5930 = ~n21604 ;
  assign y5931 = ~n21605 ;
  assign y5932 = n21609 ;
  assign y5933 = ~n21614 ;
  assign y5934 = ~n21625 ;
  assign y5935 = ~n21628 ;
  assign y5936 = ~n21630 ;
  assign y5937 = ~n21634 ;
  assign y5938 = n21636 ;
  assign y5939 = n21637 ;
  assign y5940 = ~n21644 ;
  assign y5941 = n21645 ;
  assign y5942 = n21647 ;
  assign y5943 = n21650 ;
  assign y5944 = ~n21655 ;
  assign y5945 = n21659 ;
  assign y5946 = ~n21660 ;
  assign y5947 = n21666 ;
  assign y5948 = n21668 ;
  assign y5949 = n21671 ;
  assign y5950 = n2578 ;
  assign y5951 = n21675 ;
  assign y5952 = n21681 ;
  assign y5953 = ~n7627 ;
  assign y5954 = n21682 ;
  assign y5955 = ~1'b0 ;
  assign y5956 = n21684 ;
  assign y5957 = n21691 ;
  assign y5958 = ~n21693 ;
  assign y5959 = ~n21696 ;
  assign y5960 = ~n21697 ;
  assign y5961 = n21699 ;
  assign y5962 = n21705 ;
  assign y5963 = n21707 ;
  assign y5964 = ~n21709 ;
  assign y5965 = n21723 ;
  assign y5966 = n21725 ;
  assign y5967 = ~n21727 ;
  assign y5968 = ~n21729 ;
  assign y5969 = n21730 ;
  assign y5970 = n21735 ;
  assign y5971 = n21739 ;
  assign y5972 = ~n21740 ;
  assign y5973 = ~1'b0 ;
  assign y5974 = ~n21747 ;
  assign y5975 = ~n21749 ;
  assign y5976 = n21752 ;
  assign y5977 = ~n21758 ;
  assign y5978 = ~1'b0 ;
  assign y5979 = ~n21759 ;
  assign y5980 = ~n21760 ;
  assign y5981 = n21764 ;
  assign y5982 = n21769 ;
  assign y5983 = n21779 ;
  assign y5984 = n21782 ;
  assign y5985 = ~1'b0 ;
  assign y5986 = ~n21794 ;
  assign y5987 = ~n21796 ;
  assign y5988 = ~n21799 ;
  assign y5989 = ~n21804 ;
  assign y5990 = ~n21809 ;
  assign y5991 = n21813 ;
  assign y5992 = ~n21814 ;
  assign y5993 = ~n21817 ;
  assign y5994 = ~n21818 ;
  assign y5995 = ~1'b0 ;
  assign y5996 = n21820 ;
  assign y5997 = ~n21822 ;
  assign y5998 = ~n21824 ;
  assign y5999 = n21825 ;
  assign y6000 = ~n2909 ;
  assign y6001 = ~n21826 ;
  assign y6002 = ~n21827 ;
  assign y6003 = n21830 ;
  assign y6004 = ~n21832 ;
  assign y6005 = ~n21836 ;
  assign y6006 = ~n21841 ;
  assign y6007 = ~n21843 ;
  assign y6008 = ~1'b0 ;
  assign y6009 = n21846 ;
  assign y6010 = n21851 ;
  assign y6011 = n21852 ;
  assign y6012 = n21855 ;
  assign y6013 = ~n21857 ;
  assign y6014 = ~n21860 ;
  assign y6015 = n21862 ;
  assign y6016 = ~n21864 ;
  assign y6017 = n21865 ;
  assign y6018 = ~n21871 ;
  assign y6019 = n21877 ;
  assign y6020 = n21882 ;
  assign y6021 = ~n21884 ;
  assign y6022 = n21887 ;
  assign y6023 = ~n21888 ;
  assign y6024 = ~n21889 ;
  assign y6025 = ~n21891 ;
  assign y6026 = n21895 ;
  assign y6027 = ~n21897 ;
  assign y6028 = n21899 ;
  assign y6029 = n21904 ;
  assign y6030 = n21906 ;
  assign y6031 = ~1'b0 ;
  assign y6032 = n21908 ;
  assign y6033 = n21910 ;
  assign y6034 = ~n21912 ;
  assign y6035 = n21914 ;
  assign y6036 = n21917 ;
  assign y6037 = n21921 ;
  assign y6038 = ~1'b0 ;
  assign y6039 = ~1'b0 ;
  assign y6040 = ~n21923 ;
  assign y6041 = ~n21927 ;
  assign y6042 = ~n21928 ;
  assign y6043 = n21929 ;
  assign y6044 = ~n21933 ;
  assign y6045 = ~n21934 ;
  assign y6046 = ~n21940 ;
  assign y6047 = ~n21941 ;
  assign y6048 = ~n21944 ;
  assign y6049 = n21949 ;
  assign y6050 = ~n21950 ;
  assign y6051 = n21953 ;
  assign y6052 = n12694 ;
  assign y6053 = ~n21954 ;
  assign y6054 = ~1'b0 ;
  assign y6055 = ~1'b0 ;
  assign y6056 = ~n21956 ;
  assign y6057 = ~n21958 ;
  assign y6058 = ~n21959 ;
  assign y6059 = n21960 ;
  assign y6060 = ~n21961 ;
  assign y6061 = n21962 ;
  assign y6062 = ~n21964 ;
  assign y6063 = ~n21966 ;
  assign y6064 = ~n21969 ;
  assign y6065 = ~n21971 ;
  assign y6066 = ~n21974 ;
  assign y6067 = n21975 ;
  assign y6068 = ~n21977 ;
  assign y6069 = ~n21978 ;
  assign y6070 = ~n21980 ;
  assign y6071 = ~n21990 ;
  assign y6072 = n21994 ;
  assign y6073 = ~1'b0 ;
  assign y6074 = n21996 ;
  assign y6075 = ~n21997 ;
  assign y6076 = n21998 ;
  assign y6077 = ~n22000 ;
  assign y6078 = ~n22001 ;
  assign y6079 = ~n22004 ;
  assign y6080 = ~n22008 ;
  assign y6081 = n22010 ;
  assign y6082 = ~n22012 ;
  assign y6083 = ~n22013 ;
  assign y6084 = ~n22014 ;
  assign y6085 = n22017 ;
  assign y6086 = ~n22018 ;
  assign y6087 = n22019 ;
  assign y6088 = n22020 ;
  assign y6089 = ~n22024 ;
  assign y6090 = n22028 ;
  assign y6091 = n22032 ;
  assign y6092 = n22033 ;
  assign y6093 = ~n22036 ;
  assign y6094 = ~n22038 ;
  assign y6095 = ~1'b0 ;
  assign y6096 = ~n22042 ;
  assign y6097 = n22044 ;
  assign y6098 = n22046 ;
  assign y6099 = ~n22048 ;
  assign y6100 = ~n22049 ;
  assign y6101 = n22051 ;
  assign y6102 = n22053 ;
  assign y6103 = ~n22058 ;
  assign y6104 = ~1'b0 ;
  assign y6105 = n22059 ;
  assign y6106 = n22062 ;
  assign y6107 = ~n22064 ;
  assign y6108 = n22067 ;
  assign y6109 = n22069 ;
  assign y6110 = ~n15881 ;
  assign y6111 = ~n22073 ;
  assign y6112 = n22074 ;
  assign y6113 = ~n22075 ;
  assign y6114 = n22077 ;
  assign y6115 = n22081 ;
  assign y6116 = n22083 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = ~n22086 ;
  assign y6119 = n22088 ;
  assign y6120 = n22090 ;
  assign y6121 = n22096 ;
  assign y6122 = ~n22097 ;
  assign y6123 = ~n22099 ;
  assign y6124 = ~n22100 ;
  assign y6125 = n22102 ;
  assign y6126 = ~1'b0 ;
  assign y6127 = ~n22107 ;
  assign y6128 = ~n22109 ;
  assign y6129 = n22111 ;
  assign y6130 = ~n22115 ;
  assign y6131 = ~n22116 ;
  assign y6132 = ~1'b0 ;
  assign y6133 = ~1'b0 ;
  assign y6134 = n22122 ;
  assign y6135 = n22123 ;
  assign y6136 = n22127 ;
  assign y6137 = n22133 ;
  assign y6138 = ~n22138 ;
  assign y6139 = n22139 ;
  assign y6140 = ~n22142 ;
  assign y6141 = n22143 ;
  assign y6142 = ~n22144 ;
  assign y6143 = n22145 ;
  assign y6144 = ~n22148 ;
  assign y6145 = n22152 ;
  assign y6146 = ~1'b0 ;
  assign y6147 = ~n22154 ;
  assign y6148 = ~n22158 ;
  assign y6149 = ~n22167 ;
  assign y6150 = n22173 ;
  assign y6151 = n22176 ;
  assign y6152 = ~n22177 ;
  assign y6153 = n22182 ;
  assign y6154 = ~n22186 ;
  assign y6155 = n22189 ;
  assign y6156 = ~n22192 ;
  assign y6157 = ~n22195 ;
  assign y6158 = ~n22196 ;
  assign y6159 = n22197 ;
  assign y6160 = n22202 ;
  assign y6161 = ~n22208 ;
  assign y6162 = n22210 ;
  assign y6163 = ~n22213 ;
  assign y6164 = ~n2169 ;
  assign y6165 = n22214 ;
  assign y6166 = ~n22215 ;
  assign y6167 = ~n22217 ;
  assign y6168 = n22218 ;
  assign y6169 = ~n22219 ;
  assign y6170 = n22229 ;
  assign y6171 = ~n22232 ;
  assign y6172 = ~n22240 ;
  assign y6173 = ~n22243 ;
  assign y6174 = ~n22244 ;
  assign y6175 = n22245 ;
  assign y6176 = ~n22248 ;
  assign y6177 = n22249 ;
  assign y6178 = ~n22252 ;
  assign y6179 = n22253 ;
  assign y6180 = n22254 ;
  assign y6181 = n22261 ;
  assign y6182 = ~n22263 ;
  assign y6183 = ~n22265 ;
  assign y6184 = ~n22266 ;
  assign y6185 = n22271 ;
  assign y6186 = ~1'b0 ;
  assign y6187 = ~n22275 ;
  assign y6188 = n22277 ;
  assign y6189 = ~n22279 ;
  assign y6190 = n17588 ;
  assign y6191 = ~n22280 ;
  assign y6192 = ~n22289 ;
  assign y6193 = n22298 ;
  assign y6194 = ~1'b0 ;
  assign y6195 = n22307 ;
  assign y6196 = ~n22310 ;
  assign y6197 = n22311 ;
  assign y6198 = ~n22314 ;
  assign y6199 = ~n22318 ;
  assign y6200 = ~n22322 ;
  assign y6201 = ~n22325 ;
  assign y6202 = n22329 ;
  assign y6203 = ~n22330 ;
  assign y6204 = n22331 ;
  assign y6205 = n22337 ;
  assign y6206 = ~n22338 ;
  assign y6207 = ~n22340 ;
  assign y6208 = ~n22348 ;
  assign y6209 = n22350 ;
  assign y6210 = ~1'b0 ;
  assign y6211 = n22352 ;
  assign y6212 = n22353 ;
  assign y6213 = n22354 ;
  assign y6214 = n22355 ;
  assign y6215 = ~n22358 ;
  assign y6216 = n22360 ;
  assign y6217 = ~n22361 ;
  assign y6218 = ~1'b0 ;
  assign y6219 = ~n22362 ;
  assign y6220 = ~n22363 ;
  assign y6221 = ~n22364 ;
  assign y6222 = n22367 ;
  assign y6223 = n22375 ;
  assign y6224 = ~n22377 ;
  assign y6225 = ~1'b0 ;
  assign y6226 = ~n22379 ;
  assign y6227 = ~n22382 ;
  assign y6228 = n22384 ;
  assign y6229 = ~n22387 ;
  assign y6230 = ~n22393 ;
  assign y6231 = n22394 ;
  assign y6232 = ~n22408 ;
  assign y6233 = ~1'b0 ;
  assign y6234 = ~1'b0 ;
  assign y6235 = n22411 ;
  assign y6236 = n22416 ;
  assign y6237 = ~n22417 ;
  assign y6238 = ~n22418 ;
  assign y6239 = n22419 ;
  assign y6240 = ~n22422 ;
  assign y6241 = n22428 ;
  assign y6242 = ~n22430 ;
  assign y6243 = ~n22431 ;
  assign y6244 = n22432 ;
  assign y6245 = n22433 ;
  assign y6246 = ~n22435 ;
  assign y6247 = n22436 ;
  assign y6248 = ~n22438 ;
  assign y6249 = ~n22439 ;
  assign y6250 = ~1'b0 ;
  assign y6251 = ~1'b0 ;
  assign y6252 = ~1'b0 ;
  assign y6253 = ~n22441 ;
  assign y6254 = n22446 ;
  assign y6255 = n22450 ;
  assign y6256 = ~n22453 ;
  assign y6257 = n22457 ;
  assign y6258 = n22458 ;
  assign y6259 = n22459 ;
  assign y6260 = ~n22460 ;
  assign y6261 = ~n22468 ;
  assign y6262 = n22471 ;
  assign y6263 = n22477 ;
  assign y6264 = ~1'b0 ;
  assign y6265 = ~n22481 ;
  assign y6266 = n22483 ;
  assign y6267 = ~n22492 ;
  assign y6268 = ~n22496 ;
  assign y6269 = n22497 ;
  assign y6270 = ~n22499 ;
  assign y6271 = ~1'b0 ;
  assign y6272 = ~1'b0 ;
  assign y6273 = ~n22500 ;
  assign y6274 = n22504 ;
  assign y6275 = n22505 ;
  assign y6276 = ~n22508 ;
  assign y6277 = ~n22511 ;
  assign y6278 = ~n22520 ;
  assign y6279 = n22522 ;
  assign y6280 = ~1'b0 ;
  assign y6281 = ~n22525 ;
  assign y6282 = ~n22526 ;
  assign y6283 = n22528 ;
  assign y6284 = n22529 ;
  assign y6285 = ~n22531 ;
  assign y6286 = ~n22532 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = n22534 ;
  assign y6289 = ~n22537 ;
  assign y6290 = ~n22539 ;
  assign y6291 = ~n22542 ;
  assign y6292 = ~1'b0 ;
  assign y6293 = ~1'b0 ;
  assign y6294 = ~n22544 ;
  assign y6295 = ~n22545 ;
  assign y6296 = n22548 ;
  assign y6297 = n22550 ;
  assign y6298 = n22554 ;
  assign y6299 = ~1'b0 ;
  assign y6300 = n22557 ;
  assign y6301 = ~n22558 ;
  assign y6302 = n22566 ;
  assign y6303 = n22570 ;
  assign y6304 = ~n22571 ;
  assign y6305 = ~n22575 ;
  assign y6306 = ~n22579 ;
  assign y6307 = ~n22580 ;
  assign y6308 = n22582 ;
  assign y6309 = ~n22588 ;
  assign y6310 = n22590 ;
  assign y6311 = ~n22591 ;
  assign y6312 = n22594 ;
  assign y6313 = n22604 ;
  assign y6314 = ~n22607 ;
  assign y6315 = ~n22608 ;
  assign y6316 = ~n22610 ;
  assign y6317 = n22616 ;
  assign y6318 = ~n22619 ;
  assign y6319 = n22629 ;
  assign y6320 = n22630 ;
  assign y6321 = n22633 ;
  assign y6322 = ~n22638 ;
  assign y6323 = ~1'b0 ;
  assign y6324 = n22639 ;
  assign y6325 = n22647 ;
  assign y6326 = ~n22648 ;
  assign y6327 = ~n22650 ;
  assign y6328 = n22653 ;
  assign y6329 = n22654 ;
  assign y6330 = ~n22655 ;
  assign y6331 = ~n22657 ;
  assign y6332 = ~n22660 ;
  assign y6333 = ~n22664 ;
  assign y6334 = ~n22668 ;
  assign y6335 = ~n22671 ;
  assign y6336 = n22676 ;
  assign y6337 = n22684 ;
  assign y6338 = n22689 ;
  assign y6339 = ~n22697 ;
  assign y6340 = ~n22699 ;
  assign y6341 = ~1'b0 ;
  assign y6342 = n22702 ;
  assign y6343 = n22705 ;
  assign y6344 = ~n22713 ;
  assign y6345 = n22717 ;
  assign y6346 = n22718 ;
  assign y6347 = n22719 ;
  assign y6348 = ~n22722 ;
  assign y6349 = n22727 ;
  assign y6350 = n22731 ;
  assign y6351 = n22734 ;
  assign y6352 = n22737 ;
  assign y6353 = n22740 ;
  assign y6354 = ~1'b0 ;
  assign y6355 = n22744 ;
  assign y6356 = n22746 ;
  assign y6357 = ~n22749 ;
  assign y6358 = n22751 ;
  assign y6359 = ~n22753 ;
  assign y6360 = n22755 ;
  assign y6361 = ~n22758 ;
  assign y6362 = ~n22764 ;
  assign y6363 = ~n22765 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = ~n22770 ;
  assign y6366 = n22776 ;
  assign y6367 = ~n22783 ;
  assign y6368 = n22784 ;
  assign y6369 = n22785 ;
  assign y6370 = ~1'b0 ;
  assign y6371 = ~n22790 ;
  assign y6372 = n22793 ;
  assign y6373 = ~n22798 ;
  assign y6374 = ~n22803 ;
  assign y6375 = ~n22806 ;
  assign y6376 = n22807 ;
  assign y6377 = n22808 ;
  assign y6378 = n22811 ;
  assign y6379 = ~n22813 ;
  assign y6380 = ~n22823 ;
  assign y6381 = n22826 ;
  assign y6382 = ~n22829 ;
  assign y6383 = ~n22835 ;
  assign y6384 = ~n22836 ;
  assign y6385 = n22838 ;
  assign y6386 = ~n22841 ;
  assign y6387 = ~n22842 ;
  assign y6388 = ~1'b0 ;
  assign y6389 = n22843 ;
  assign y6390 = ~n22848 ;
  assign y6391 = n22849 ;
  assign y6392 = n22851 ;
  assign y6393 = n22852 ;
  assign y6394 = ~1'b0 ;
  assign y6395 = ~1'b0 ;
  assign y6396 = ~n22856 ;
  assign y6397 = ~n22857 ;
  assign y6398 = ~n22872 ;
  assign y6399 = ~n22874 ;
  assign y6400 = ~n22875 ;
  assign y6401 = ~1'b0 ;
  assign y6402 = ~n22878 ;
  assign y6403 = n22879 ;
  assign y6404 = n22882 ;
  assign y6405 = n22883 ;
  assign y6406 = n22892 ;
  assign y6407 = ~1'b0 ;
  assign y6408 = ~n22894 ;
  assign y6409 = n22895 ;
  assign y6410 = n22897 ;
  assign y6411 = ~n22901 ;
  assign y6412 = ~n22904 ;
  assign y6413 = ~n22905 ;
  assign y6414 = n22906 ;
  assign y6415 = ~n22913 ;
  assign y6416 = n22916 ;
  assign y6417 = ~n22918 ;
  assign y6418 = ~n22921 ;
  assign y6419 = ~1'b0 ;
  assign y6420 = ~n22922 ;
  assign y6421 = ~n22924 ;
  assign y6422 = ~n22925 ;
  assign y6423 = n22927 ;
  assign y6424 = ~n22933 ;
  assign y6425 = ~n22939 ;
  assign y6426 = ~1'b0 ;
  assign y6427 = n22942 ;
  assign y6428 = n22946 ;
  assign y6429 = n22948 ;
  assign y6430 = ~n22953 ;
  assign y6431 = n22956 ;
  assign y6432 = ~n22957 ;
  assign y6433 = ~1'b0 ;
  assign y6434 = n22958 ;
  assign y6435 = n22959 ;
  assign y6436 = ~n22961 ;
  assign y6437 = n22966 ;
  assign y6438 = n22967 ;
  assign y6439 = ~n22973 ;
  assign y6440 = n22974 ;
  assign y6441 = ~1'b0 ;
  assign y6442 = n22975 ;
  assign y6443 = ~n22976 ;
  assign y6444 = n22979 ;
  assign y6445 = ~n22981 ;
  assign y6446 = ~1'b0 ;
  assign y6447 = ~n22983 ;
  assign y6448 = n22984 ;
  assign y6449 = n22986 ;
  assign y6450 = n22989 ;
  assign y6451 = n22990 ;
  assign y6452 = ~n22993 ;
  assign y6453 = ~1'b0 ;
  assign y6454 = ~n22996 ;
  assign y6455 = ~n23000 ;
  assign y6456 = ~n23010 ;
  assign y6457 = ~n23012 ;
  assign y6458 = ~n23016 ;
  assign y6459 = ~n23019 ;
  assign y6460 = ~n23020 ;
  assign y6461 = ~n23022 ;
  assign y6462 = ~n23027 ;
  assign y6463 = ~n23028 ;
  assign y6464 = n23032 ;
  assign y6465 = ~n23035 ;
  assign y6466 = n23037 ;
  assign y6467 = n23041 ;
  assign y6468 = ~n23042 ;
  assign y6469 = ~n23043 ;
  assign y6470 = ~n23056 ;
  assign y6471 = ~n23059 ;
  assign y6472 = ~n23063 ;
  assign y6473 = n23065 ;
  assign y6474 = n23066 ;
  assign y6475 = n23067 ;
  assign y6476 = n23070 ;
  assign y6477 = n23071 ;
  assign y6478 = ~1'b0 ;
  assign y6479 = ~n23076 ;
  assign y6480 = n23080 ;
  assign y6481 = n23082 ;
  assign y6482 = ~n23084 ;
  assign y6483 = ~n23090 ;
  assign y6484 = ~n23091 ;
  assign y6485 = ~n23097 ;
  assign y6486 = ~1'b0 ;
  assign y6487 = ~n23099 ;
  assign y6488 = n23100 ;
  assign y6489 = ~n23105 ;
  assign y6490 = ~n23106 ;
  assign y6491 = ~n10399 ;
  assign y6492 = ~n23109 ;
  assign y6493 = n23110 ;
  assign y6494 = ~n23112 ;
  assign y6495 = n23113 ;
  assign y6496 = ~n23114 ;
  assign y6497 = ~n23115 ;
  assign y6498 = ~n23116 ;
  assign y6499 = ~n23117 ;
  assign y6500 = n23122 ;
  assign y6501 = ~n23124 ;
  assign y6502 = n23126 ;
  assign y6503 = n23128 ;
  assign y6504 = ~n23129 ;
  assign y6505 = n23132 ;
  assign y6506 = ~n23136 ;
  assign y6507 = n23137 ;
  assign y6508 = n23140 ;
  assign y6509 = n23147 ;
  assign y6510 = ~n23151 ;
  assign y6511 = n23155 ;
  assign y6512 = ~n23157 ;
  assign y6513 = n23158 ;
  assign y6514 = ~n23159 ;
  assign y6515 = n23161 ;
  assign y6516 = ~n23162 ;
  assign y6517 = ~1'b0 ;
  assign y6518 = ~n23164 ;
  assign y6519 = ~1'b0 ;
  assign y6520 = ~n23170 ;
  assign y6521 = n23171 ;
  assign y6522 = n23174 ;
  assign y6523 = ~n23176 ;
  assign y6524 = ~n23178 ;
  assign y6525 = ~1'b0 ;
  assign y6526 = ~n23179 ;
  assign y6527 = ~n23180 ;
  assign y6528 = n23182 ;
  assign y6529 = ~1'b0 ;
  assign y6530 = n23183 ;
  assign y6531 = n23186 ;
  assign y6532 = n23187 ;
  assign y6533 = ~n23188 ;
  assign y6534 = ~n23192 ;
  assign y6535 = ~n23193 ;
  assign y6536 = n23206 ;
  assign y6537 = ~n23209 ;
  assign y6538 = n23210 ;
  assign y6539 = n23219 ;
  assign y6540 = ~n23220 ;
  assign y6541 = n23224 ;
  assign y6542 = ~1'b0 ;
  assign y6543 = ~n23226 ;
  assign y6544 = n23229 ;
  assign y6545 = n23232 ;
  assign y6546 = ~n23234 ;
  assign y6547 = ~n23238 ;
  assign y6548 = ~n23242 ;
  assign y6549 = n23249 ;
  assign y6550 = n23253 ;
  assign y6551 = n23257 ;
  assign y6552 = ~n23258 ;
  assign y6553 = n23262 ;
  assign y6554 = n23264 ;
  assign y6555 = n23266 ;
  assign y6556 = n23267 ;
  assign y6557 = ~n23271 ;
  assign y6558 = ~1'b0 ;
  assign y6559 = ~n23273 ;
  assign y6560 = ~n23278 ;
  assign y6561 = n23281 ;
  assign y6562 = n23287 ;
  assign y6563 = ~n23288 ;
  assign y6564 = n23289 ;
  assign y6565 = ~n23291 ;
  assign y6566 = n23293 ;
  assign y6567 = n23295 ;
  assign y6568 = ~n23297 ;
  assign y6569 = n23303 ;
  assign y6570 = n23304 ;
  assign y6571 = n23309 ;
  assign y6572 = ~n23311 ;
  assign y6573 = n23313 ;
  assign y6574 = ~n23317 ;
  assign y6575 = n23320 ;
  assign y6576 = ~n23321 ;
  assign y6577 = n23323 ;
  assign y6578 = n3966 ;
  assign y6579 = ~n23326 ;
  assign y6580 = ~n23328 ;
  assign y6581 = ~n23329 ;
  assign y6582 = ~n23331 ;
  assign y6583 = n23334 ;
  assign y6584 = ~n23335 ;
  assign y6585 = ~n23339 ;
  assign y6586 = ~n23343 ;
  assign y6587 = n23344 ;
  assign y6588 = ~1'b0 ;
  assign y6589 = ~n23349 ;
  assign y6590 = ~n23352 ;
  assign y6591 = n23355 ;
  assign y6592 = ~n23356 ;
  assign y6593 = ~n23360 ;
  assign y6594 = n23361 ;
  assign y6595 = ~n23362 ;
  assign y6596 = ~1'b0 ;
  assign y6597 = ~n23364 ;
  assign y6598 = ~n23367 ;
  assign y6599 = ~n23371 ;
  assign y6600 = ~n23372 ;
  assign y6601 = n23373 ;
  assign y6602 = ~n23374 ;
  assign y6603 = n23375 ;
  assign y6604 = ~1'b0 ;
  assign y6605 = ~n23376 ;
  assign y6606 = ~1'b0 ;
  assign y6607 = ~1'b0 ;
  assign y6608 = ~n23379 ;
  assign y6609 = ~n23380 ;
  assign y6610 = n23382 ;
  assign y6611 = ~n23389 ;
  assign y6612 = ~n23390 ;
  assign y6613 = ~1'b0 ;
  assign y6614 = ~n23392 ;
  assign y6615 = n23394 ;
  assign y6616 = ~n23396 ;
  assign y6617 = n23397 ;
  assign y6618 = ~n23399 ;
  assign y6619 = ~n23400 ;
  assign y6620 = ~n23401 ;
  assign y6621 = n23405 ;
  assign y6622 = ~n23413 ;
  assign y6623 = n23416 ;
  assign y6624 = n23421 ;
  assign y6625 = n23424 ;
  assign y6626 = n23426 ;
  assign y6627 = ~n23427 ;
  assign y6628 = ~n23431 ;
  assign y6629 = ~n23435 ;
  assign y6630 = ~1'b0 ;
  assign y6631 = ~n23439 ;
  assign y6632 = n23441 ;
  assign y6633 = n23445 ;
  assign y6634 = n23447 ;
  assign y6635 = ~n23452 ;
  assign y6636 = ~n23455 ;
  assign y6637 = ~n23460 ;
  assign y6638 = ~1'b0 ;
  assign y6639 = ~n23461 ;
  assign y6640 = ~n23466 ;
  assign y6641 = ~1'b0 ;
  assign y6642 = ~n23470 ;
  assign y6643 = ~n23473 ;
  assign y6644 = ~n2221 ;
  assign y6645 = ~n23476 ;
  assign y6646 = ~n761 ;
  assign y6647 = ~n23479 ;
  assign y6648 = ~n23484 ;
  assign y6649 = ~1'b0 ;
  assign y6650 = ~n23492 ;
  assign y6651 = n23493 ;
  assign y6652 = n23498 ;
  assign y6653 = n23502 ;
  assign y6654 = ~n23503 ;
  assign y6655 = n23512 ;
  assign y6656 = n23513 ;
  assign y6657 = n23515 ;
  assign y6658 = n23520 ;
  assign y6659 = ~1'b0 ;
  assign y6660 = ~n23526 ;
  assign y6661 = n23530 ;
  assign y6662 = n23533 ;
  assign y6663 = n23534 ;
  assign y6664 = ~n23536 ;
  assign y6665 = ~n23537 ;
  assign y6666 = n23538 ;
  assign y6667 = ~n23539 ;
  assign y6668 = ~n23544 ;
  assign y6669 = n23545 ;
  assign y6670 = n23547 ;
  assign y6671 = ~n23548 ;
  assign y6672 = ~n23550 ;
  assign y6673 = ~n23553 ;
  assign y6674 = ~1'b0 ;
  assign y6675 = ~n23557 ;
  assign y6676 = ~n23558 ;
  assign y6677 = n23559 ;
  assign y6678 = n23561 ;
  assign y6679 = n23577 ;
  assign y6680 = ~n23578 ;
  assign y6681 = ~1'b0 ;
  assign y6682 = ~n23580 ;
  assign y6683 = ~n23583 ;
  assign y6684 = ~n23584 ;
  assign y6685 = n23586 ;
  assign y6686 = ~n23591 ;
  assign y6687 = ~n23595 ;
  assign y6688 = n23598 ;
  assign y6689 = ~n23602 ;
  assign y6690 = ~n23604 ;
  assign y6691 = ~n23608 ;
  assign y6692 = n23612 ;
  assign y6693 = n23615 ;
  assign y6694 = ~1'b0 ;
  assign y6695 = ~n23620 ;
  assign y6696 = n23624 ;
  assign y6697 = ~n23627 ;
  assign y6698 = ~n23630 ;
  assign y6699 = n23631 ;
  assign y6700 = ~n23637 ;
  assign y6701 = n23642 ;
  assign y6702 = ~1'b0 ;
  assign y6703 = ~n23648 ;
  assign y6704 = n23650 ;
  assign y6705 = n23654 ;
  assign y6706 = ~n23661 ;
  assign y6707 = n23662 ;
  assign y6708 = ~1'b0 ;
  assign y6709 = n23664 ;
  assign y6710 = n23666 ;
  assign y6711 = ~n23668 ;
  assign y6712 = n23672 ;
  assign y6713 = ~1'b0 ;
  assign y6714 = n23676 ;
  assign y6715 = n23685 ;
  assign y6716 = n23688 ;
  assign y6717 = ~n23691 ;
  assign y6718 = ~1'b0 ;
  assign y6719 = ~n23695 ;
  assign y6720 = ~n23700 ;
  assign y6721 = ~n23703 ;
  assign y6722 = ~n23706 ;
  assign y6723 = ~n23709 ;
  assign y6724 = ~n23711 ;
  assign y6725 = ~1'b0 ;
  assign y6726 = ~n23714 ;
  assign y6727 = ~n23715 ;
  assign y6728 = ~n23717 ;
  assign y6729 = ~n23718 ;
  assign y6730 = n23719 ;
  assign y6731 = n23721 ;
  assign y6732 = ~1'b0 ;
  assign y6733 = ~n23722 ;
  assign y6734 = ~n23726 ;
  assign y6735 = ~n23732 ;
  assign y6736 = ~n23737 ;
  assign y6737 = n23742 ;
  assign y6738 = ~n23744 ;
  assign y6739 = n23747 ;
  assign y6740 = ~n23749 ;
  assign y6741 = n23752 ;
  assign y6742 = ~n23753 ;
  assign y6743 = ~n23756 ;
  assign y6744 = n23757 ;
  assign y6745 = ~n23762 ;
  assign y6746 = n23766 ;
  assign y6747 = ~1'b0 ;
  assign y6748 = ~n23774 ;
  assign y6749 = ~n23777 ;
  assign y6750 = n23781 ;
  assign y6751 = ~n23784 ;
  assign y6752 = ~n23791 ;
  assign y6753 = n23794 ;
  assign y6754 = ~n23796 ;
  assign y6755 = ~n23798 ;
  assign y6756 = ~n23799 ;
  assign y6757 = n23801 ;
  assign y6758 = ~n23803 ;
  assign y6759 = ~n23807 ;
  assign y6760 = ~n23814 ;
  assign y6761 = ~n23815 ;
  assign y6762 = n23816 ;
  assign y6763 = ~n23818 ;
  assign y6764 = n23819 ;
  assign y6765 = ~n23825 ;
  assign y6766 = ~n23828 ;
  assign y6767 = n23830 ;
  assign y6768 = ~n23832 ;
  assign y6769 = ~n23837 ;
  assign y6770 = n23840 ;
  assign y6771 = ~n23841 ;
  assign y6772 = n23842 ;
  assign y6773 = n23843 ;
  assign y6774 = n11316 ;
  assign y6775 = n23846 ;
  assign y6776 = ~1'b0 ;
  assign y6777 = ~n23851 ;
  assign y6778 = ~n23855 ;
  assign y6779 = n23857 ;
  assign y6780 = n23866 ;
  assign y6781 = n23868 ;
  assign y6782 = ~n23870 ;
  assign y6783 = ~n23871 ;
  assign y6784 = n23873 ;
  assign y6785 = ~n23875 ;
  assign y6786 = ~n23876 ;
  assign y6787 = ~n23882 ;
  assign y6788 = ~n23890 ;
  assign y6789 = n23893 ;
  assign y6790 = ~n23895 ;
  assign y6791 = n23902 ;
  assign y6792 = ~1'b0 ;
  assign y6793 = n23904 ;
  assign y6794 = ~n23906 ;
  assign y6795 = n23908 ;
  assign y6796 = n23909 ;
  assign y6797 = ~n23910 ;
  assign y6798 = n23911 ;
  assign y6799 = n23913 ;
  assign y6800 = ~n23914 ;
  assign y6801 = n23916 ;
  assign y6802 = n23917 ;
  assign y6803 = ~1'b0 ;
  assign y6804 = ~n23918 ;
  assign y6805 = n23921 ;
  assign y6806 = n23923 ;
  assign y6807 = ~n23929 ;
  assign y6808 = n23930 ;
  assign y6809 = ~n23932 ;
  assign y6810 = n23934 ;
  assign y6811 = ~n23936 ;
  assign y6812 = ~1'b0 ;
  assign y6813 = n23937 ;
  assign y6814 = ~n23938 ;
  assign y6815 = ~n23939 ;
  assign y6816 = ~n23945 ;
  assign y6817 = n23946 ;
  assign y6818 = ~n23950 ;
  assign y6819 = ~1'b0 ;
  assign y6820 = ~1'b0 ;
  assign y6821 = ~n8695 ;
  assign y6822 = n23953 ;
  assign y6823 = ~n23954 ;
  assign y6824 = n23959 ;
  assign y6825 = ~n23966 ;
  assign y6826 = n23968 ;
  assign y6827 = n23974 ;
  assign y6828 = ~1'b0 ;
  assign y6829 = ~n23976 ;
  assign y6830 = n23977 ;
  assign y6831 = ~n23978 ;
  assign y6832 = ~n23981 ;
  assign y6833 = ~n23982 ;
  assign y6834 = n23983 ;
  assign y6835 = ~n23990 ;
  assign y6836 = ~n23997 ;
  assign y6837 = ~n24005 ;
  assign y6838 = n24011 ;
  assign y6839 = ~1'b0 ;
  assign y6840 = n24018 ;
  assign y6841 = n24019 ;
  assign y6842 = ~n24021 ;
  assign y6843 = n24022 ;
  assign y6844 = ~n24024 ;
  assign y6845 = n24026 ;
  assign y6846 = ~n10297 ;
  assign y6847 = n24033 ;
  assign y6848 = ~n24034 ;
  assign y6849 = ~n24038 ;
  assign y6850 = ~n24044 ;
  assign y6851 = ~n24047 ;
  assign y6852 = n24048 ;
  assign y6853 = n24051 ;
  assign y6854 = n24053 ;
  assign y6855 = ~1'b0 ;
  assign y6856 = n24056 ;
  assign y6857 = ~n24057 ;
  assign y6858 = n24062 ;
  assign y6859 = ~n24066 ;
  assign y6860 = ~n24069 ;
  assign y6861 = ~n24071 ;
  assign y6862 = n24072 ;
  assign y6863 = ~n24074 ;
  assign y6864 = 1'b0 ;
  assign y6865 = ~1'b0 ;
  assign y6866 = n24075 ;
  assign y6867 = n24078 ;
  assign y6868 = n24081 ;
  assign y6869 = n24082 ;
  assign y6870 = ~1'b0 ;
  assign y6871 = ~n24084 ;
  assign y6872 = n24086 ;
  assign y6873 = n24087 ;
  assign y6874 = ~n24089 ;
  assign y6875 = n24092 ;
  assign y6876 = ~n24103 ;
  assign y6877 = n24104 ;
  assign y6878 = n24108 ;
  assign y6879 = ~n24110 ;
  assign y6880 = n24114 ;
  assign y6881 = ~n24118 ;
  assign y6882 = n24121 ;
  assign y6883 = ~n24128 ;
  assign y6884 = ~n24129 ;
  assign y6885 = ~n24134 ;
  assign y6886 = ~n24137 ;
  assign y6887 = ~n24138 ;
  assign y6888 = ~n24139 ;
  assign y6889 = ~n24140 ;
  assign y6890 = ~n24141 ;
  assign y6891 = ~n24145 ;
  assign y6892 = ~n24152 ;
  assign y6893 = ~1'b0 ;
  assign y6894 = ~1'b0 ;
  assign y6895 = ~1'b0 ;
  assign y6896 = ~n24154 ;
  assign y6897 = n24155 ;
  assign y6898 = n24158 ;
  assign y6899 = ~n24161 ;
  assign y6900 = n24163 ;
  assign y6901 = ~n24166 ;
  assign y6902 = ~n24169 ;
  assign y6903 = ~n24172 ;
  assign y6904 = ~n24187 ;
  assign y6905 = n24189 ;
  assign y6906 = ~n24193 ;
  assign y6907 = n24194 ;
  assign y6908 = n24197 ;
  assign y6909 = ~n24199 ;
  assign y6910 = ~n24200 ;
  assign y6911 = ~n24202 ;
  assign y6912 = ~n24205 ;
  assign y6913 = n24206 ;
  assign y6914 = ~n24210 ;
  assign y6915 = ~n24211 ;
  assign y6916 = ~n24219 ;
  assign y6917 = ~n24221 ;
  assign y6918 = ~n24222 ;
  assign y6919 = n24227 ;
  assign y6920 = ~n24231 ;
  assign y6921 = n24240 ;
  assign y6922 = ~n24242 ;
  assign y6923 = ~n24245 ;
  assign y6924 = ~1'b0 ;
  assign y6925 = ~n24249 ;
  assign y6926 = n24253 ;
  assign y6927 = ~n24256 ;
  assign y6928 = ~n24257 ;
  assign y6929 = n24258 ;
  assign y6930 = n24259 ;
  assign y6931 = ~n24264 ;
  assign y6932 = ~n24266 ;
  assign y6933 = n24270 ;
  assign y6934 = ~n24273 ;
  assign y6935 = ~n6488 ;
  assign y6936 = n24274 ;
  assign y6937 = n24275 ;
  assign y6938 = ~n24277 ;
  assign y6939 = n24279 ;
  assign y6940 = ~n24281 ;
  assign y6941 = n24285 ;
  assign y6942 = ~1'b0 ;
  assign y6943 = ~n24291 ;
  assign y6944 = ~n24296 ;
  assign y6945 = n24297 ;
  assign y6946 = ~n24300 ;
  assign y6947 = ~n24303 ;
  assign y6948 = ~n24307 ;
  assign y6949 = n24311 ;
  assign y6950 = ~1'b0 ;
  assign y6951 = ~1'b0 ;
  assign y6952 = n24314 ;
  assign y6953 = n24321 ;
  assign y6954 = n24326 ;
  assign y6955 = n24329 ;
  assign y6956 = n24337 ;
  assign y6957 = ~n24338 ;
  assign y6958 = ~n24341 ;
  assign y6959 = ~n24345 ;
  assign y6960 = ~1'b0 ;
  assign y6961 = ~n24347 ;
  assign y6962 = n24350 ;
  assign y6963 = n24352 ;
  assign y6964 = n24359 ;
  assign y6965 = ~n24361 ;
  assign y6966 = ~n24365 ;
  assign y6967 = n24366 ;
  assign y6968 = ~n24369 ;
  assign y6969 = ~1'b0 ;
  assign y6970 = ~1'b0 ;
  assign y6971 = n24370 ;
  assign y6972 = n24378 ;
  assign y6973 = ~n24381 ;
  assign y6974 = ~n24383 ;
  assign y6975 = ~1'b0 ;
  assign y6976 = ~n24386 ;
  assign y6977 = ~1'b0 ;
  assign y6978 = ~n24393 ;
  assign y6979 = n24394 ;
  assign y6980 = ~n24395 ;
  assign y6981 = n24396 ;
  assign y6982 = n24399 ;
  assign y6983 = n24406 ;
  assign y6984 = n24410 ;
  assign y6985 = n24414 ;
  assign y6986 = ~1'b0 ;
  assign y6987 = n24418 ;
  assign y6988 = n24421 ;
  assign y6989 = n24429 ;
  assign y6990 = ~n24433 ;
  assign y6991 = n24436 ;
  assign y6992 = ~n24440 ;
  assign y6993 = ~n24441 ;
  assign y6994 = n24444 ;
  assign y6995 = ~n24447 ;
  assign y6996 = ~1'b0 ;
  assign y6997 = n24451 ;
  assign y6998 = ~n24460 ;
  assign y6999 = n24467 ;
  assign y7000 = ~n24468 ;
  assign y7001 = ~n24469 ;
  assign y7002 = ~1'b0 ;
  assign y7003 = ~n11583 ;
  assign y7004 = ~n24470 ;
  assign y7005 = ~n24473 ;
  assign y7006 = ~n24480 ;
  assign y7007 = n24482 ;
  assign y7008 = n24487 ;
  assign y7009 = ~n24488 ;
  assign y7010 = ~1'b0 ;
  assign y7011 = n24490 ;
  assign y7012 = ~n24491 ;
  assign y7013 = ~n24494 ;
  assign y7014 = ~n24499 ;
  assign y7015 = ~n24500 ;
  assign y7016 = ~n24501 ;
  assign y7017 = ~n24504 ;
  assign y7018 = ~n24505 ;
  assign y7019 = ~n24507 ;
  assign y7020 = n24509 ;
  assign y7021 = n24517 ;
  assign y7022 = ~n24522 ;
  assign y7023 = n24526 ;
  assign y7024 = ~n24527 ;
  assign y7025 = n24529 ;
  assign y7026 = n24530 ;
  assign y7027 = ~1'b0 ;
  assign y7028 = ~n24534 ;
  assign y7029 = n24537 ;
  assign y7030 = n24541 ;
  assign y7031 = ~n24545 ;
  assign y7032 = ~n24551 ;
  assign y7033 = n24556 ;
  assign y7034 = ~n24565 ;
  assign y7035 = ~n24566 ;
  assign y7036 = n24570 ;
  assign y7037 = n24574 ;
  assign y7038 = ~n24575 ;
  assign y7039 = ~n14762 ;
  assign y7040 = n24580 ;
  assign y7041 = n24581 ;
  assign y7042 = ~n24588 ;
  assign y7043 = n24590 ;
  assign y7044 = n24597 ;
  assign y7045 = n24598 ;
  assign y7046 = ~n24600 ;
  assign y7047 = ~n24602 ;
  assign y7048 = ~n24605 ;
  assign y7049 = ~n24615 ;
  assign y7050 = n24618 ;
  assign y7051 = n24622 ;
  assign y7052 = n24624 ;
  assign y7053 = n24627 ;
  assign y7054 = ~n24628 ;
  assign y7055 = ~1'b0 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = n24630 ;
  assign y7058 = ~n24635 ;
  assign y7059 = n24638 ;
  assign y7060 = ~1'b0 ;
  assign y7061 = ~1'b0 ;
  assign y7062 = n24640 ;
  assign y7063 = ~n24642 ;
  assign y7064 = n24643 ;
  assign y7065 = n24644 ;
  assign y7066 = ~n24645 ;
  assign y7067 = ~n24647 ;
  assign y7068 = ~n24649 ;
  assign y7069 = ~n24651 ;
  assign y7070 = ~n24655 ;
  assign y7071 = n24660 ;
  assign y7072 = n24662 ;
  assign y7073 = ~n24664 ;
  assign y7074 = n24666 ;
  assign y7075 = ~n24669 ;
  assign y7076 = ~n24671 ;
  assign y7077 = ~n24673 ;
  assign y7078 = ~n24679 ;
  assign y7079 = ~n24681 ;
  assign y7080 = ~n24685 ;
  assign y7081 = ~n24688 ;
  assign y7082 = ~n24691 ;
  assign y7083 = 1'b0 ;
  assign y7084 = n24693 ;
  assign y7085 = ~n24694 ;
  assign y7086 = n24695 ;
  assign y7087 = ~n24698 ;
  assign y7088 = n9052 ;
  assign y7089 = n24701 ;
  assign y7090 = ~n24703 ;
  assign y7091 = ~n24705 ;
  assign y7092 = n24706 ;
  assign y7093 = n24707 ;
  assign y7094 = ~n24708 ;
  assign y7095 = ~n24710 ;
  assign y7096 = n24714 ;
  assign y7097 = n24716 ;
  assign y7098 = n24720 ;
  assign y7099 = ~1'b0 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = n24722 ;
  assign y7102 = n24726 ;
  assign y7103 = ~n24729 ;
  assign y7104 = ~n24732 ;
  assign y7105 = ~n24736 ;
  assign y7106 = n24742 ;
  assign y7107 = ~1'b0 ;
  assign y7108 = ~n24746 ;
  assign y7109 = n24748 ;
  assign y7110 = ~n24752 ;
  assign y7111 = ~n24753 ;
  assign y7112 = ~n24761 ;
  assign y7113 = n24765 ;
  assign y7114 = ~n24769 ;
  assign y7115 = ~n24770 ;
  assign y7116 = n24776 ;
  assign y7117 = n24780 ;
  assign y7118 = n24781 ;
  assign y7119 = n24783 ;
  assign y7120 = ~n24785 ;
  assign y7121 = n24786 ;
  assign y7122 = n24792 ;
  assign y7123 = n24793 ;
  assign y7124 = ~n24802 ;
  assign y7125 = ~n24805 ;
  assign y7126 = n24811 ;
  assign y7127 = n24813 ;
  assign y7128 = n24816 ;
  assign y7129 = n24817 ;
  assign y7130 = ~1'b0 ;
  assign y7131 = ~n24820 ;
  assign y7132 = ~n24826 ;
  assign y7133 = n24827 ;
  assign y7134 = n24828 ;
  assign y7135 = n24829 ;
  assign y7136 = n24837 ;
  assign y7137 = ~n24838 ;
  assign y7138 = n24841 ;
  assign y7139 = ~n24842 ;
  assign y7140 = n24843 ;
  assign y7141 = ~n24845 ;
  assign y7142 = n24846 ;
  assign y7143 = n24848 ;
  assign y7144 = n24849 ;
  assign y7145 = ~n24855 ;
  assign y7146 = ~n24861 ;
  assign y7147 = n24863 ;
  assign y7148 = ~1'b0 ;
  assign y7149 = n24866 ;
  assign y7150 = ~n24867 ;
  assign y7151 = ~n24871 ;
  assign y7152 = n24872 ;
  assign y7153 = n24880 ;
  assign y7154 = n24881 ;
  assign y7155 = n24883 ;
  assign y7156 = ~n24885 ;
  assign y7157 = n24887 ;
  assign y7158 = ~n24893 ;
  assign y7159 = ~n24901 ;
  assign y7160 = n24903 ;
  assign y7161 = ~n24904 ;
  assign y7162 = ~n24905 ;
  assign y7163 = n24906 ;
  assign y7164 = n24908 ;
  assign y7165 = ~n24910 ;
  assign y7166 = ~n24915 ;
  assign y7167 = n24916 ;
  assign y7168 = ~n24919 ;
  assign y7169 = ~n24921 ;
  assign y7170 = ~n24923 ;
  assign y7171 = ~n24925 ;
  assign y7172 = ~1'b0 ;
  assign y7173 = n24926 ;
  assign y7174 = ~n24927 ;
  assign y7175 = ~n24928 ;
  assign y7176 = n24929 ;
  assign y7177 = n24930 ;
  assign y7178 = ~n24933 ;
  assign y7179 = n24935 ;
  assign y7180 = n24936 ;
  assign y7181 = ~n24940 ;
  assign y7182 = n24943 ;
  assign y7183 = ~n24945 ;
  assign y7184 = n24946 ;
  assign y7185 = ~n24947 ;
  assign y7186 = n24953 ;
  assign y7187 = n24954 ;
  assign y7188 = ~n24958 ;
  assign y7189 = ~n24961 ;
  assign y7190 = n24964 ;
  assign y7191 = n24965 ;
  assign y7192 = n24967 ;
  assign y7193 = ~1'b0 ;
  assign y7194 = ~1'b0 ;
  assign y7195 = ~n24969 ;
  assign y7196 = n24972 ;
  assign y7197 = n24973 ;
  assign y7198 = n24974 ;
  assign y7199 = ~1'b0 ;
  assign y7200 = ~n24976 ;
  assign y7201 = n24981 ;
  assign y7202 = ~n24982 ;
  assign y7203 = n24983 ;
  assign y7204 = ~n24985 ;
  assign y7205 = ~n24990 ;
  assign y7206 = n24994 ;
  assign y7207 = n24998 ;
  assign y7208 = ~1'b0 ;
  assign y7209 = ~n25003 ;
  assign y7210 = ~n25007 ;
  assign y7211 = ~n25011 ;
  assign y7212 = n25014 ;
  assign y7213 = ~n12723 ;
  assign y7214 = n25016 ;
  assign y7215 = ~n25017 ;
  assign y7216 = ~1'b0 ;
  assign y7217 = n25018 ;
  assign y7218 = n25022 ;
  assign y7219 = ~n25026 ;
  assign y7220 = n25028 ;
  assign y7221 = ~n25034 ;
  assign y7222 = ~n25035 ;
  assign y7223 = n25036 ;
  assign y7224 = ~1'b0 ;
  assign y7225 = n25037 ;
  assign y7226 = n25042 ;
  assign y7227 = ~n25054 ;
  assign y7228 = ~n25056 ;
  assign y7229 = ~n25059 ;
  assign y7230 = ~n25060 ;
  assign y7231 = n25061 ;
  assign y7232 = ~n25069 ;
  assign y7233 = ~1'b0 ;
  assign y7234 = ~1'b0 ;
  assign y7235 = n25070 ;
  assign y7236 = n25073 ;
  assign y7237 = n25080 ;
  assign y7238 = n25081 ;
  assign y7239 = ~n25085 ;
  assign y7240 = ~n25086 ;
  assign y7241 = n25092 ;
  assign y7242 = ~n25095 ;
  assign y7243 = ~n25099 ;
  assign y7244 = n25102 ;
  assign y7245 = n25103 ;
  assign y7246 = ~n25104 ;
  assign y7247 = ~n25106 ;
  assign y7248 = n25107 ;
  assign y7249 = n25108 ;
  assign y7250 = ~n25110 ;
  assign y7251 = n25113 ;
  assign y7252 = n25115 ;
  assign y7253 = ~n25117 ;
  assign y7254 = n25120 ;
  assign y7255 = n25128 ;
  assign y7256 = ~n25130 ;
  assign y7257 = n25133 ;
  assign y7258 = ~1'b0 ;
  assign y7259 = ~n25135 ;
  assign y7260 = n25138 ;
  assign y7261 = ~n25139 ;
  assign y7262 = n25143 ;
  assign y7263 = ~n25147 ;
  assign y7264 = ~n25149 ;
  assign y7265 = n25151 ;
  assign y7266 = n25164 ;
  assign y7267 = ~n25166 ;
  assign y7268 = ~n25169 ;
  assign y7269 = ~n25172 ;
  assign y7270 = n25174 ;
  assign y7271 = ~n25175 ;
  assign y7272 = ~n25176 ;
  assign y7273 = n25180 ;
  assign y7274 = ~n25183 ;
  assign y7275 = ~1'b0 ;
  assign y7276 = n25185 ;
  assign y7277 = ~n25186 ;
  assign y7278 = ~n25187 ;
  assign y7279 = n25190 ;
  assign y7280 = n25191 ;
  assign y7281 = n25193 ;
  assign y7282 = ~1'b0 ;
  assign y7283 = ~n13669 ;
  assign y7284 = n25195 ;
  assign y7285 = ~n25196 ;
  assign y7286 = n25199 ;
  assign y7287 = n25200 ;
  assign y7288 = n25201 ;
  assign y7289 = ~n25203 ;
  assign y7290 = n25206 ;
  assign y7291 = n25211 ;
  assign y7292 = n25214 ;
  assign y7293 = ~n25216 ;
  assign y7294 = n25218 ;
  assign y7295 = ~n25223 ;
  assign y7296 = ~n25224 ;
  assign y7297 = n25225 ;
  assign y7298 = ~n25230 ;
  assign y7299 = ~n25233 ;
  assign y7300 = n25237 ;
  assign y7301 = n25243 ;
  assign y7302 = ~1'b0 ;
  assign y7303 = ~1'b0 ;
  assign y7304 = n25245 ;
  assign y7305 = ~n25250 ;
  assign y7306 = ~n25251 ;
  assign y7307 = ~n25252 ;
  assign y7308 = ~1'b0 ;
  assign y7309 = n25254 ;
  assign y7310 = ~n25256 ;
  assign y7311 = n25257 ;
  assign y7312 = n25260 ;
  assign y7313 = ~n25263 ;
  assign y7314 = ~n25264 ;
  assign y7315 = n25265 ;
  assign y7316 = ~n25267 ;
  assign y7317 = ~n25271 ;
  assign y7318 = ~n25273 ;
  assign y7319 = n25278 ;
  assign y7320 = n25284 ;
  assign y7321 = n25289 ;
  assign y7322 = ~n25290 ;
  assign y7323 = ~n25292 ;
  assign y7324 = ~n25295 ;
  assign y7325 = n25300 ;
  assign y7326 = n25302 ;
  assign y7327 = ~1'b0 ;
  assign y7328 = n25305 ;
  assign y7329 = ~n25306 ;
  assign y7330 = ~n25307 ;
  assign y7331 = ~n25309 ;
  assign y7332 = n25311 ;
  assign y7333 = n25314 ;
  assign y7334 = ~n25322 ;
  assign y7335 = ~n25326 ;
  assign y7336 = ~n25328 ;
  assign y7337 = n25329 ;
  assign y7338 = ~n25333 ;
  assign y7339 = ~n25335 ;
  assign y7340 = ~n25344 ;
  assign y7341 = ~n25345 ;
  assign y7342 = ~n25347 ;
  assign y7343 = n25350 ;
  assign y7344 = n25356 ;
  assign y7345 = ~n25358 ;
  assign y7346 = ~n25362 ;
  assign y7347 = ~1'b0 ;
  assign y7348 = ~n25366 ;
  assign y7349 = ~n25380 ;
  assign y7350 = ~n25381 ;
  assign y7351 = ~n25382 ;
  assign y7352 = ~n24650 ;
  assign y7353 = ~1'b0 ;
  assign y7354 = n25383 ;
  assign y7355 = n25385 ;
  assign y7356 = n25387 ;
  assign y7357 = ~n25396 ;
  assign y7358 = n25397 ;
  assign y7359 = ~n25401 ;
  assign y7360 = ~n25402 ;
  assign y7361 = n25404 ;
  assign y7362 = n25407 ;
  assign y7363 = ~n25408 ;
  assign y7364 = ~n25409 ;
  assign y7365 = ~n25411 ;
  assign y7366 = ~n25412 ;
  assign y7367 = n25414 ;
  assign y7368 = n25417 ;
  assign y7369 = ~n25421 ;
  assign y7370 = ~n25425 ;
  assign y7371 = ~1'b0 ;
  assign y7372 = n25429 ;
  assign y7373 = ~n25434 ;
  assign y7374 = ~n25440 ;
  assign y7375 = ~n25442 ;
  assign y7376 = ~n25444 ;
  assign y7377 = n25446 ;
  assign y7378 = ~n25447 ;
  assign y7379 = ~n25451 ;
  assign y7380 = ~n25453 ;
  assign y7381 = n25455 ;
  assign y7382 = ~1'b0 ;
  assign y7383 = n25456 ;
  assign y7384 = ~n25457 ;
  assign y7385 = ~n25464 ;
  assign y7386 = ~n25465 ;
  assign y7387 = n25467 ;
  assign y7388 = ~n25469 ;
  assign y7389 = ~n25470 ;
  assign y7390 = n25476 ;
  assign y7391 = n25478 ;
  assign y7392 = n25479 ;
  assign y7393 = n25483 ;
  assign y7394 = n25488 ;
  assign y7395 = n25493 ;
  assign y7396 = n25497 ;
  assign y7397 = n25499 ;
  assign y7398 = n25500 ;
  assign y7399 = ~n25503 ;
  assign y7400 = ~n25506 ;
  assign y7401 = n25507 ;
  assign y7402 = ~n25509 ;
  assign y7403 = ~n25511 ;
  assign y7404 = n25514 ;
  assign y7405 = ~n23544 ;
  assign y7406 = ~n25515 ;
  assign y7407 = ~n25516 ;
  assign y7408 = n25518 ;
  assign y7409 = ~1'b0 ;
  assign y7410 = n25520 ;
  assign y7411 = ~n25526 ;
  assign y7412 = n25530 ;
  assign y7413 = n25535 ;
  assign y7414 = n25538 ;
  assign y7415 = ~n25541 ;
  assign y7416 = ~n25542 ;
  assign y7417 = ~1'b0 ;
  assign y7418 = ~n25544 ;
  assign y7419 = n25546 ;
  assign y7420 = n25548 ;
  assign y7421 = n25551 ;
  assign y7422 = ~n25556 ;
  assign y7423 = ~n25557 ;
  assign y7424 = n25562 ;
  assign y7425 = n25564 ;
  assign y7426 = n25565 ;
  assign y7427 = n25568 ;
  assign y7428 = ~n25571 ;
  assign y7429 = n25574 ;
  assign y7430 = n25575 ;
  assign y7431 = n25576 ;
  assign y7432 = ~n25577 ;
  assign y7433 = ~n25578 ;
  assign y7434 = n25585 ;
  assign y7435 = n25586 ;
  assign y7436 = ~n25592 ;
  assign y7437 = ~n25601 ;
  assign y7438 = n25602 ;
  assign y7439 = n25605 ;
  assign y7440 = ~n25608 ;
  assign y7441 = n25611 ;
  assign y7442 = ~n25612 ;
  assign y7443 = ~n25614 ;
  assign y7444 = ~n25616 ;
  assign y7445 = ~n25620 ;
  assign y7446 = n25622 ;
  assign y7447 = ~n25623 ;
  assign y7448 = ~n25624 ;
  assign y7449 = n25626 ;
  assign y7450 = ~n25627 ;
  assign y7451 = n25631 ;
  assign y7452 = n25633 ;
  assign y7453 = ~1'b0 ;
  assign y7454 = n25635 ;
  assign y7455 = n25637 ;
  assign y7456 = n25641 ;
  assign y7457 = ~n25642 ;
  assign y7458 = ~n25643 ;
  assign y7459 = n25644 ;
  assign y7460 = ~n25646 ;
  assign y7461 = n25647 ;
  assign y7462 = ~1'b0 ;
  assign y7463 = n25648 ;
  assign y7464 = ~n25649 ;
  assign y7465 = ~n25650 ;
  assign y7466 = ~n25658 ;
  assign y7467 = ~n25659 ;
  assign y7468 = ~n25662 ;
  assign y7469 = ~1'b0 ;
  assign y7470 = ~1'b0 ;
  assign y7471 = ~n25667 ;
  assign y7472 = ~n25671 ;
  assign y7473 = n25673 ;
  assign y7474 = n25675 ;
  assign y7475 = n25678 ;
  assign y7476 = n25680 ;
  assign y7477 = ~1'b0 ;
  assign y7478 = ~n25682 ;
  assign y7479 = n25683 ;
  assign y7480 = n25684 ;
  assign y7481 = ~n7306 ;
  assign y7482 = n25687 ;
  assign y7483 = n25688 ;
  assign y7484 = ~n25690 ;
  assign y7485 = ~1'b0 ;
  assign y7486 = ~n25693 ;
  assign y7487 = ~1'b0 ;
  assign y7488 = n25696 ;
  assign y7489 = ~n25697 ;
  assign y7490 = n25698 ;
  assign y7491 = n25699 ;
  assign y7492 = ~n25700 ;
  assign y7493 = ~1'b0 ;
  assign y7494 = n25702 ;
  assign y7495 = ~1'b0 ;
  assign y7496 = ~n25703 ;
  assign y7497 = n25704 ;
  assign y7498 = n25707 ;
  assign y7499 = n25709 ;
  assign y7500 = n25710 ;
  assign y7501 = ~n25715 ;
  assign y7502 = n25716 ;
  assign y7503 = ~n25717 ;
  assign y7504 = n25719 ;
  assign y7505 = ~n25722 ;
  assign y7506 = n25723 ;
  assign y7507 = ~n25738 ;
  assign y7508 = ~n25739 ;
  assign y7509 = ~n25740 ;
  assign y7510 = ~1'b0 ;
  assign y7511 = ~n25745 ;
  assign y7512 = ~n25746 ;
  assign y7513 = n25748 ;
  assign y7514 = ~n25749 ;
  assign y7515 = n25751 ;
  assign y7516 = ~n25752 ;
  assign y7517 = ~1'b0 ;
  assign y7518 = n25755 ;
  assign y7519 = n25757 ;
  assign y7520 = n25763 ;
  assign y7521 = ~n25764 ;
  assign y7522 = n25770 ;
  assign y7523 = ~n25772 ;
  assign y7524 = n25773 ;
  assign y7525 = ~n25776 ;
  assign y7526 = n25777 ;
  assign y7527 = ~n25779 ;
  assign y7528 = ~n25781 ;
  assign y7529 = n25783 ;
  assign y7530 = ~n25784 ;
  assign y7531 = n25785 ;
  assign y7532 = ~n25787 ;
  assign y7533 = n25788 ;
  assign y7534 = ~n25790 ;
  assign y7535 = ~n25792 ;
  assign y7536 = ~n25800 ;
  assign y7537 = n25803 ;
  assign y7538 = n168 ;
  assign y7539 = ~n25805 ;
  assign y7540 = n25806 ;
  assign y7541 = ~n25811 ;
  assign y7542 = ~n25813 ;
  assign y7543 = ~n25814 ;
  assign y7544 = n25818 ;
  assign y7545 = n25821 ;
  assign y7546 = n25823 ;
  assign y7547 = ~n25824 ;
  assign y7548 = ~n25825 ;
  assign y7549 = ~n25827 ;
  assign y7550 = ~n25829 ;
  assign y7551 = n25830 ;
  assign y7552 = ~n25832 ;
  assign y7553 = ~n25835 ;
  assign y7554 = n11737 ;
  assign y7555 = n25841 ;
  assign y7556 = ~n25842 ;
  assign y7557 = n25844 ;
  assign y7558 = n25847 ;
  assign y7559 = n25848 ;
  assign y7560 = n25853 ;
  assign y7561 = ~1'b0 ;
  assign y7562 = ~n25854 ;
  assign y7563 = ~n25855 ;
  assign y7564 = ~n25861 ;
  assign y7565 = ~n25862 ;
  assign y7566 = ~n25864 ;
  assign y7567 = ~n25866 ;
  assign y7568 = ~n25870 ;
  assign y7569 = ~1'b0 ;
  assign y7570 = ~n25873 ;
  assign y7571 = ~n25875 ;
  assign y7572 = n25876 ;
  assign y7573 = ~n25877 ;
  assign y7574 = ~n25878 ;
  assign y7575 = ~n25880 ;
  assign y7576 = ~n25882 ;
  assign y7577 = ~1'b0 ;
  assign y7578 = ~n25887 ;
  assign y7579 = ~n25888 ;
  assign y7580 = ~n25892 ;
  assign y7581 = ~n25893 ;
  assign y7582 = ~n25894 ;
  assign y7583 = ~n16458 ;
  assign y7584 = ~n25896 ;
  assign y7585 = n25903 ;
  assign y7586 = n25905 ;
  assign y7587 = n25906 ;
  assign y7588 = n25908 ;
  assign y7589 = ~n25915 ;
  assign y7590 = n25917 ;
  assign y7591 = ~1'b0 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = n25919 ;
  assign y7594 = n25923 ;
  assign y7595 = ~n25926 ;
  assign y7596 = ~n25930 ;
  assign y7597 = ~n25935 ;
  assign y7598 = n25936 ;
  assign y7599 = ~n25939 ;
  assign y7600 = ~n25942 ;
  assign y7601 = ~1'b0 ;
  assign y7602 = ~n3243 ;
  assign y7603 = n25943 ;
  assign y7604 = ~n25946 ;
  assign y7605 = ~n25947 ;
  assign y7606 = ~n25949 ;
  assign y7607 = ~1'b0 ;
  assign y7608 = ~n25951 ;
  assign y7609 = ~n25960 ;
  assign y7610 = n25963 ;
  assign y7611 = ~n25975 ;
  assign y7612 = ~n25979 ;
  assign y7613 = n25981 ;
  assign y7614 = ~1'b0 ;
  assign y7615 = ~n25986 ;
  assign y7616 = ~1'b0 ;
  assign y7617 = n25987 ;
  assign y7618 = n25989 ;
  assign y7619 = ~n25992 ;
  assign y7620 = ~n25995 ;
  assign y7621 = n25998 ;
  assign y7622 = ~n26002 ;
  assign y7623 = ~1'b0 ;
  assign y7624 = ~1'b0 ;
  assign y7625 = n26007 ;
  assign y7626 = n26012 ;
  assign y7627 = n26013 ;
  assign y7628 = ~n26014 ;
  assign y7629 = n26015 ;
  assign y7630 = n26016 ;
  assign y7631 = ~1'b0 ;
  assign y7632 = ~1'b0 ;
  assign y7633 = n26017 ;
  assign y7634 = n26019 ;
  assign y7635 = ~n26020 ;
  assign y7636 = n26021 ;
  assign y7637 = n26023 ;
  assign y7638 = n26025 ;
  assign y7639 = n26026 ;
  assign y7640 = n26034 ;
  assign y7641 = ~n26036 ;
  assign y7642 = n26037 ;
  assign y7643 = n26039 ;
  assign y7644 = n26042 ;
  assign y7645 = n26053 ;
  assign y7646 = ~n26055 ;
  assign y7647 = n26057 ;
  assign y7648 = n26059 ;
  assign y7649 = n26061 ;
  assign y7650 = ~n26062 ;
  assign y7651 = n26064 ;
  assign y7652 = n26065 ;
  assign y7653 = n26066 ;
  assign y7654 = ~n26068 ;
  assign y7655 = n26071 ;
  assign y7656 = ~n26077 ;
  assign y7657 = n26080 ;
  assign y7658 = n26082 ;
  assign y7659 = ~n26088 ;
  assign y7660 = ~n26090 ;
  assign y7661 = ~n26091 ;
  assign y7662 = n26093 ;
  assign y7663 = ~n26097 ;
  assign y7664 = n26100 ;
  assign y7665 = ~n26103 ;
  assign y7666 = n26107 ;
  assign y7667 = n26112 ;
  assign y7668 = ~n26113 ;
  assign y7669 = ~n26115 ;
  assign y7670 = n26118 ;
  assign y7671 = ~n26119 ;
  assign y7672 = ~n26121 ;
  assign y7673 = n26123 ;
  assign y7674 = ~1'b0 ;
  assign y7675 = ~n26125 ;
  assign y7676 = ~1'b0 ;
  assign y7677 = ~n26126 ;
  assign y7678 = ~n26133 ;
  assign y7679 = ~n26135 ;
  assign y7680 = ~n26139 ;
  assign y7681 = ~n26143 ;
  assign y7682 = n26144 ;
  assign y7683 = n26151 ;
  assign y7684 = ~1'b0 ;
  assign y7685 = n26153 ;
  assign y7686 = n26155 ;
  assign y7687 = ~n26157 ;
  assign y7688 = n26167 ;
  assign y7689 = ~n26169 ;
  assign y7690 = ~n26172 ;
  assign y7691 = n26174 ;
  assign y7692 = n21616 ;
  assign y7693 = n26177 ;
  assign y7694 = ~n26182 ;
  assign y7695 = ~n26185 ;
  assign y7696 = ~n26194 ;
  assign y7697 = n3018 ;
  assign y7698 = n26195 ;
  assign y7699 = ~n26197 ;
  assign y7700 = n26204 ;
  assign y7701 = ~1'b0 ;
  assign y7702 = ~n26206 ;
  assign y7703 = ~n26210 ;
  assign y7704 = ~n26213 ;
  assign y7705 = n26214 ;
  assign y7706 = ~n26219 ;
  assign y7707 = n26221 ;
  assign y7708 = n26222 ;
  assign y7709 = n26223 ;
  assign y7710 = ~n26227 ;
  assign y7711 = ~n26230 ;
  assign y7712 = ~n26234 ;
  assign y7713 = ~n26235 ;
  assign y7714 = ~n26237 ;
  assign y7715 = ~n26239 ;
  assign y7716 = n26241 ;
  assign y7717 = ~n26243 ;
  assign y7718 = ~n26245 ;
  assign y7719 = ~n26249 ;
  assign y7720 = ~n26253 ;
  assign y7721 = ~1'b0 ;
  assign y7722 = ~1'b0 ;
  assign y7723 = n26258 ;
  assign y7724 = n26259 ;
  assign y7725 = n26262 ;
  assign y7726 = ~n26263 ;
  assign y7727 = ~n26267 ;
  assign y7728 = ~n26268 ;
  assign y7729 = n26270 ;
  assign y7730 = ~1'b0 ;
  assign y7731 = ~n26275 ;
  assign y7732 = ~n26277 ;
  assign y7733 = ~n26281 ;
  assign y7734 = n26285 ;
  assign y7735 = n26286 ;
  assign y7736 = ~n26287 ;
  assign y7737 = ~1'b0 ;
  assign y7738 = n26291 ;
  assign y7739 = ~1'b0 ;
  assign y7740 = ~n26300 ;
  assign y7741 = ~n26302 ;
  assign y7742 = ~n26309 ;
  assign y7743 = n26310 ;
  assign y7744 = ~n26314 ;
  assign y7745 = n26317 ;
  assign y7746 = n26318 ;
  assign y7747 = ~n26320 ;
  assign y7748 = n26324 ;
  assign y7749 = ~n26325 ;
  assign y7750 = ~n26329 ;
  assign y7751 = ~n26330 ;
  assign y7752 = ~n26332 ;
  assign y7753 = ~1'b0 ;
  assign y7754 = n26333 ;
  assign y7755 = ~n26338 ;
  assign y7756 = ~n26342 ;
  assign y7757 = n26346 ;
  assign y7758 = ~n26347 ;
  assign y7759 = ~n26350 ;
  assign y7760 = ~n26352 ;
  assign y7761 = n26354 ;
  assign y7762 = ~n26355 ;
  assign y7763 = ~n26356 ;
  assign y7764 = ~n26357 ;
  assign y7765 = n26360 ;
  assign y7766 = n26374 ;
  assign y7767 = ~n26375 ;
  assign y7768 = n26379 ;
  assign y7769 = n26385 ;
  assign y7770 = ~1'b0 ;
  assign y7771 = ~n26388 ;
  assign y7772 = ~n26390 ;
  assign y7773 = n26391 ;
  assign y7774 = ~n26393 ;
  assign y7775 = n26396 ;
  assign y7776 = ~n26399 ;
  assign y7777 = ~n26400 ;
  assign y7778 = ~n26401 ;
  assign y7779 = n26405 ;
  assign y7780 = ~n26407 ;
  assign y7781 = ~n26409 ;
  assign y7782 = n26414 ;
  assign y7783 = ~n26415 ;
  assign y7784 = ~n26416 ;
  assign y7785 = n26420 ;
  assign y7786 = ~n26425 ;
  assign y7787 = ~n26429 ;
  assign y7788 = ~n26431 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = n26432 ;
  assign y7791 = n26435 ;
  assign y7792 = ~n26437 ;
  assign y7793 = ~n26439 ;
  assign y7794 = n26440 ;
  assign y7795 = ~1'b0 ;
  assign y7796 = ~n26442 ;
  assign y7797 = n26448 ;
  assign y7798 = n26449 ;
  assign y7799 = n26451 ;
  assign y7800 = ~n26455 ;
  assign y7801 = ~n26457 ;
  assign y7802 = n26459 ;
  assign y7803 = ~n26461 ;
  assign y7804 = n26465 ;
  assign y7805 = ~1'b0 ;
  assign y7806 = ~n26468 ;
  assign y7807 = ~n26478 ;
  assign y7808 = ~n26479 ;
  assign y7809 = n26480 ;
  assign y7810 = n26481 ;
  assign y7811 = ~n26485 ;
  assign y7812 = n26486 ;
  assign y7813 = n26487 ;
  assign y7814 = ~n26489 ;
  assign y7815 = n26493 ;
  assign y7816 = n26495 ;
  assign y7817 = n26496 ;
  assign y7818 = n26500 ;
  assign y7819 = n26501 ;
  assign y7820 = ~n26503 ;
  assign y7821 = n26505 ;
  assign y7822 = n26508 ;
  assign y7823 = ~n26512 ;
  assign y7824 = ~n26514 ;
  assign y7825 = ~1'b0 ;
  assign y7826 = ~n26517 ;
  assign y7827 = ~n26519 ;
  assign y7828 = ~n26101 ;
  assign y7829 = ~n26521 ;
  assign y7830 = n26523 ;
  assign y7831 = n26525 ;
  assign y7832 = n26527 ;
  assign y7833 = n26528 ;
  assign y7834 = ~1'b0 ;
  assign y7835 = n26531 ;
  assign y7836 = n26535 ;
  assign y7837 = ~n26536 ;
  assign y7838 = ~n26538 ;
  assign y7839 = ~n26539 ;
  assign y7840 = ~1'b0 ;
  assign y7841 = n26541 ;
  assign y7842 = ~n26545 ;
  assign y7843 = ~1'b0 ;
  assign y7844 = n26546 ;
  assign y7845 = n26551 ;
  assign y7846 = n26552 ;
  assign y7847 = ~n26556 ;
  assign y7848 = n26558 ;
  assign y7849 = ~n26564 ;
  assign y7850 = ~n26565 ;
  assign y7851 = n26569 ;
  assign y7852 = n26570 ;
  assign y7853 = n26571 ;
  assign y7854 = ~n26572 ;
  assign y7855 = ~n26573 ;
  assign y7856 = ~n26578 ;
  assign y7857 = ~1'b0 ;
  assign y7858 = ~1'b0 ;
  assign y7859 = ~n26579 ;
  assign y7860 = ~n26582 ;
  assign y7861 = n26585 ;
  assign y7862 = n26586 ;
  assign y7863 = n26588 ;
  assign y7864 = ~1'b0 ;
  assign y7865 = ~1'b0 ;
  assign y7866 = n26591 ;
  assign y7867 = n26594 ;
  assign y7868 = ~n26600 ;
  assign y7869 = n26604 ;
  assign y7870 = ~n26609 ;
  assign y7871 = n26612 ;
  assign y7872 = ~n26614 ;
  assign y7873 = n26616 ;
  assign y7874 = ~n26619 ;
  assign y7875 = n26623 ;
  assign y7876 = ~n26624 ;
  assign y7877 = n26629 ;
  assign y7878 = ~n26631 ;
  assign y7879 = n26633 ;
  assign y7880 = ~n26636 ;
  assign y7881 = ~1'b0 ;
  assign y7882 = n26637 ;
  assign y7883 = n26642 ;
  assign y7884 = n26643 ;
  assign y7885 = n26644 ;
  assign y7886 = ~1'b0 ;
  assign y7887 = ~n26645 ;
  assign y7888 = n26652 ;
  assign y7889 = ~n26655 ;
  assign y7890 = ~1'b0 ;
  assign y7891 = n26656 ;
  assign y7892 = ~n26657 ;
  assign y7893 = n26660 ;
  assign y7894 = n26665 ;
  assign y7895 = ~n26670 ;
  assign y7896 = ~1'b0 ;
  assign y7897 = ~1'b0 ;
  assign y7898 = n26671 ;
  assign y7899 = ~n26674 ;
  assign y7900 = ~n26677 ;
  assign y7901 = ~n26684 ;
  assign y7902 = ~n26685 ;
  assign y7903 = ~n26686 ;
  assign y7904 = n26689 ;
  assign y7905 = n26693 ;
  assign y7906 = ~n26698 ;
  assign y7907 = n26701 ;
  assign y7908 = ~n26705 ;
  assign y7909 = ~n26706 ;
  assign y7910 = ~n26707 ;
  assign y7911 = n26713 ;
  assign y7912 = ~n26717 ;
  assign y7913 = ~n26719 ;
  assign y7914 = ~n26721 ;
  assign y7915 = ~n26722 ;
  assign y7916 = ~n26724 ;
  assign y7917 = ~n26728 ;
  assign y7918 = n26732 ;
  assign y7919 = n26736 ;
  assign y7920 = ~n26737 ;
  assign y7921 = n26743 ;
  assign y7922 = ~1'b0 ;
  assign y7923 = ~n26746 ;
  assign y7924 = n26747 ;
  assign y7925 = ~n26748 ;
  assign y7926 = n26751 ;
  assign y7927 = ~n26752 ;
  assign y7928 = ~n26753 ;
  assign y7929 = ~n26755 ;
  assign y7930 = n26758 ;
  assign y7931 = n26759 ;
  assign y7932 = n26763 ;
  assign y7933 = n26765 ;
  assign y7934 = n26766 ;
  assign y7935 = n6461 ;
  assign y7936 = ~n26767 ;
  assign y7937 = ~n26770 ;
  assign y7938 = n26772 ;
  assign y7939 = ~n26773 ;
  assign y7940 = n26776 ;
  assign y7941 = n26781 ;
  assign y7942 = n26784 ;
  assign y7943 = ~n26790 ;
  assign y7944 = ~1'b0 ;
  assign y7945 = ~1'b0 ;
  assign y7946 = ~n26791 ;
  assign y7947 = ~n26792 ;
  assign y7948 = n26795 ;
  assign y7949 = n26796 ;
  assign y7950 = ~n26798 ;
  assign y7951 = n26799 ;
  assign y7952 = n26801 ;
  assign y7953 = n26802 ;
  assign y7954 = ~n26805 ;
  assign y7955 = ~n26806 ;
  assign y7956 = n26807 ;
  assign y7957 = ~n8042 ;
  assign y7958 = n26812 ;
  assign y7959 = n26816 ;
  assign y7960 = ~n26817 ;
  assign y7961 = n26818 ;
  assign y7962 = ~n26819 ;
  assign y7963 = ~n26821 ;
  assign y7964 = n26822 ;
  assign y7965 = ~n26823 ;
  assign y7966 = n26829 ;
  assign y7967 = ~n26833 ;
  assign y7968 = ~n26835 ;
  assign y7969 = n26837 ;
  assign y7970 = ~n26841 ;
  assign y7971 = n26843 ;
  assign y7972 = ~n26845 ;
  assign y7973 = ~n26846 ;
  assign y7974 = ~n26848 ;
  assign y7975 = n26852 ;
  assign y7976 = n26856 ;
  assign y7977 = ~1'b0 ;
  assign y7978 = n26860 ;
  assign y7979 = ~n26864 ;
  assign y7980 = ~n26867 ;
  assign y7981 = n26868 ;
  assign y7982 = ~n26869 ;
  assign y7983 = ~n26872 ;
  assign y7984 = n26876 ;
  assign y7985 = n26878 ;
  assign y7986 = ~n26885 ;
  assign y7987 = n26887 ;
  assign y7988 = ~n26889 ;
  assign y7989 = n26890 ;
  assign y7990 = n26893 ;
  assign y7991 = n26894 ;
  assign y7992 = n26898 ;
  assign y7993 = n26899 ;
  assign y7994 = n26900 ;
  assign y7995 = ~1'b0 ;
  assign y7996 = n26903 ;
  assign y7997 = ~n26906 ;
  assign y7998 = n26908 ;
  assign y7999 = ~n26914 ;
  assign y8000 = n26917 ;
  assign y8001 = ~n26918 ;
  assign y8002 = n26920 ;
  assign y8003 = ~n26922 ;
  assign y8004 = ~n26926 ;
  assign y8005 = ~1'b0 ;
  assign y8006 = ~n26928 ;
  assign y8007 = n26929 ;
  assign y8008 = n26930 ;
  assign y8009 = ~n26934 ;
  assign y8010 = ~1'b0 ;
  assign y8011 = ~n26936 ;
  assign y8012 = n26939 ;
  assign y8013 = ~n26941 ;
  assign y8014 = ~n26943 ;
  assign y8015 = ~n26944 ;
  assign y8016 = ~n26945 ;
  assign y8017 = ~n26947 ;
  assign y8018 = ~n26948 ;
  assign y8019 = ~n26949 ;
  assign y8020 = ~n26950 ;
  assign y8021 = ~1'b0 ;
  assign y8022 = ~1'b0 ;
  assign y8023 = ~n26955 ;
  assign y8024 = n26956 ;
  assign y8025 = ~n26960 ;
  assign y8026 = n26961 ;
  assign y8027 = n26963 ;
  assign y8028 = ~n26965 ;
  assign y8029 = n26968 ;
  assign y8030 = n26971 ;
  assign y8031 = n26972 ;
  assign y8032 = ~n26973 ;
  assign y8033 = ~n26977 ;
  assign y8034 = n26978 ;
  assign y8035 = n26979 ;
  assign y8036 = ~n26980 ;
  assign y8037 = n26981 ;
  assign y8038 = ~n26982 ;
  assign y8039 = n26984 ;
  assign y8040 = n26986 ;
  assign y8041 = ~n26991 ;
  assign y8042 = n26992 ;
  assign y8043 = ~n26998 ;
  assign y8044 = ~n26999 ;
  assign y8045 = n27002 ;
  assign y8046 = ~n27006 ;
  assign y8047 = n27007 ;
  assign y8048 = ~n27008 ;
  assign y8049 = n27009 ;
  assign y8050 = ~n27013 ;
  assign y8051 = ~n27015 ;
  assign y8052 = ~1'b0 ;
  assign y8053 = ~n27018 ;
  assign y8054 = ~1'b0 ;
  assign y8055 = ~n27019 ;
  assign y8056 = n27021 ;
  assign y8057 = ~n27025 ;
  assign y8058 = n27026 ;
  assign y8059 = n27027 ;
  assign y8060 = n27029 ;
  assign y8061 = ~n27032 ;
  assign y8062 = n27035 ;
  assign y8063 = n27036 ;
  assign y8064 = n27037 ;
  assign y8065 = ~n27039 ;
  assign y8066 = n27040 ;
  assign y8067 = ~n27043 ;
  assign y8068 = ~n27045 ;
  assign y8069 = ~1'b0 ;
  assign y8070 = ~n27046 ;
  assign y8071 = n27048 ;
  assign y8072 = ~n27053 ;
  assign y8073 = n27054 ;
  assign y8074 = ~n27062 ;
  assign y8075 = ~n27063 ;
  assign y8076 = ~n27064 ;
  assign y8077 = ~n27066 ;
  assign y8078 = ~n27068 ;
  assign y8079 = n27072 ;
  assign y8080 = ~n27073 ;
  assign y8081 = n27074 ;
  assign y8082 = n27075 ;
  assign y8083 = ~n27077 ;
  assign y8084 = ~n27080 ;
  assign y8085 = n27082 ;
  assign y8086 = ~1'b0 ;
  assign y8087 = n27084 ;
  assign y8088 = n27085 ;
  assign y8089 = n27086 ;
  assign y8090 = n27087 ;
  assign y8091 = n27091 ;
  assign y8092 = n27094 ;
  assign y8093 = ~1'b0 ;
  assign y8094 = ~n27096 ;
  assign y8095 = n27098 ;
  assign y8096 = n27100 ;
  assign y8097 = n27101 ;
  assign y8098 = n27102 ;
  assign y8099 = ~n27104 ;
  assign y8100 = ~n27109 ;
  assign y8101 = n27111 ;
  assign y8102 = ~n27112 ;
  assign y8103 = ~n27117 ;
  assign y8104 = n27119 ;
  assign y8105 = n27121 ;
  assign y8106 = n27127 ;
  assign y8107 = n27128 ;
  assign y8108 = ~n27130 ;
  assign y8109 = n27133 ;
  assign y8110 = ~n27134 ;
  assign y8111 = n27139 ;
  assign y8112 = n27142 ;
  assign y8113 = n27143 ;
  assign y8114 = n27147 ;
  assign y8115 = ~n27149 ;
  assign y8116 = n27152 ;
  assign y8117 = ~n27154 ;
  assign y8118 = n27159 ;
  assign y8119 = n27161 ;
  assign y8120 = n27162 ;
  assign y8121 = n27163 ;
  assign y8122 = n27165 ;
  assign y8123 = n27166 ;
  assign y8124 = n27167 ;
  assign y8125 = n27171 ;
  assign y8126 = ~n27173 ;
  assign y8127 = n27175 ;
  assign y8128 = ~1'b0 ;
  assign y8129 = ~n27177 ;
  assign y8130 = n27178 ;
  assign y8131 = n25733 ;
  assign y8132 = n27183 ;
  assign y8133 = n27187 ;
  assign y8134 = ~n27194 ;
  assign y8135 = ~1'b0 ;
  assign y8136 = ~n27196 ;
  assign y8137 = ~n27199 ;
  assign y8138 = ~n27200 ;
  assign y8139 = ~n27202 ;
  assign y8140 = n27205 ;
  assign y8141 = n27206 ;
  assign y8142 = ~n27207 ;
  assign y8143 = n27214 ;
  assign y8144 = ~n27216 ;
  assign y8145 = n27218 ;
  assign y8146 = ~1'b0 ;
  assign y8147 = ~n27220 ;
  assign y8148 = ~n27227 ;
  assign y8149 = ~n27228 ;
  assign y8150 = ~n27235 ;
  assign y8151 = ~n27243 ;
  assign y8152 = ~n27245 ;
  assign y8153 = ~1'b0 ;
  assign y8154 = n27248 ;
  assign y8155 = n27252 ;
  assign y8156 = ~n27253 ;
  assign y8157 = ~n27254 ;
  assign y8158 = n27257 ;
  assign y8159 = n27258 ;
  assign y8160 = ~n27261 ;
  assign y8161 = ~1'b0 ;
  assign y8162 = n27264 ;
  assign y8163 = ~n27265 ;
  assign y8164 = n27266 ;
  assign y8165 = n27267 ;
  assign y8166 = n27270 ;
  assign y8167 = n27271 ;
  assign y8168 = ~n27274 ;
  assign y8169 = n27276 ;
  assign y8170 = ~n27278 ;
  assign y8171 = n27280 ;
  assign y8172 = ~1'b0 ;
  assign y8173 = ~n27281 ;
  assign y8174 = n27283 ;
  assign y8175 = ~n27287 ;
  assign y8176 = ~n27288 ;
  assign y8177 = n27292 ;
  assign y8178 = n27294 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = n27297 ;
  assign y8181 = ~n27300 ;
  assign y8182 = ~n27302 ;
  assign y8183 = n27303 ;
  assign y8184 = ~n27305 ;
  assign y8185 = ~n27307 ;
  assign y8186 = ~n27309 ;
  assign y8187 = ~n27310 ;
  assign y8188 = n27315 ;
  assign y8189 = n27321 ;
  assign y8190 = ~n27326 ;
  assign y8191 = ~n27327 ;
  assign y8192 = n27328 ;
  assign y8193 = ~n27331 ;
  assign y8194 = n27333 ;
  assign y8195 = ~n27335 ;
  assign y8196 = ~n27337 ;
  assign y8197 = n27338 ;
  assign y8198 = ~n27340 ;
  assign y8199 = n27341 ;
  assign y8200 = ~n27342 ;
  assign y8201 = ~n27344 ;
  assign y8202 = n27346 ;
  assign y8203 = ~n27348 ;
  assign y8204 = n27356 ;
  assign y8205 = n27357 ;
  assign y8206 = n27359 ;
  assign y8207 = n27362 ;
  assign y8208 = ~n27365 ;
  assign y8209 = n27367 ;
  assign y8210 = ~1'b0 ;
  assign y8211 = ~1'b0 ;
  assign y8212 = ~n27369 ;
  assign y8213 = n27373 ;
  assign y8214 = n27374 ;
  assign y8215 = n27375 ;
  assign y8216 = ~n27378 ;
  assign y8217 = ~n27387 ;
  assign y8218 = n27392 ;
  assign y8219 = ~n27395 ;
  assign y8220 = n27399 ;
  assign y8221 = ~n27401 ;
  assign y8222 = ~n27406 ;
  assign y8223 = n27411 ;
  assign y8224 = n27412 ;
  assign y8225 = ~n27416 ;
  assign y8226 = ~n27417 ;
  assign y8227 = n27418 ;
  assign y8228 = ~n27420 ;
  assign y8229 = ~1'b0 ;
  assign y8230 = ~1'b0 ;
  assign y8231 = ~1'b0 ;
  assign y8232 = n27422 ;
  assign y8233 = ~n27423 ;
  assign y8234 = ~n27425 ;
  assign y8235 = n27426 ;
  assign y8236 = n27427 ;
  assign y8237 = ~1'b0 ;
  assign y8238 = n27430 ;
  assign y8239 = ~n27432 ;
  assign y8240 = ~n27435 ;
  assign y8241 = ~n27437 ;
  assign y8242 = n27439 ;
  assign y8243 = n27440 ;
  assign y8244 = n27443 ;
  assign y8245 = ~n27447 ;
  assign y8246 = ~n27449 ;
  assign y8247 = ~1'b0 ;
  assign y8248 = ~n27451 ;
  assign y8249 = n27455 ;
  assign y8250 = ~1'b0 ;
  assign y8251 = n27458 ;
  assign y8252 = n27460 ;
  assign y8253 = n27463 ;
  assign y8254 = ~1'b0 ;
  assign y8255 = ~n27465 ;
  assign y8256 = ~n27466 ;
  assign y8257 = n27469 ;
  assign y8258 = ~n27474 ;
  assign y8259 = ~n27477 ;
  assign y8260 = ~n27480 ;
  assign y8261 = ~n27482 ;
  assign y8262 = n27486 ;
  assign y8263 = ~n27488 ;
  assign y8264 = ~n27493 ;
  assign y8265 = ~n15486 ;
  assign y8266 = n27494 ;
  assign y8267 = n27495 ;
  assign y8268 = n1851 ;
  assign y8269 = n27496 ;
  assign y8270 = n27501 ;
  assign y8271 = n27504 ;
  assign y8272 = ~1'b0 ;
  assign y8273 = ~1'b0 ;
  assign y8274 = ~1'b0 ;
  assign y8275 = n26216 ;
  assign y8276 = ~n27505 ;
  assign y8277 = ~n27508 ;
  assign y8278 = ~n27514 ;
  assign y8279 = n27520 ;
  assign y8280 = n27526 ;
  assign y8281 = ~n27528 ;
  assign y8282 = ~n27530 ;
  assign y8283 = n27533 ;
  assign y8284 = ~n27535 ;
  assign y8285 = ~n27536 ;
  assign y8286 = n27541 ;
  assign y8287 = n27543 ;
  assign y8288 = n27544 ;
  assign y8289 = n27546 ;
  assign y8290 = ~n27550 ;
  assign y8291 = n27551 ;
  assign y8292 = ~n27554 ;
  assign y8293 = ~1'b0 ;
  assign y8294 = ~n27555 ;
  assign y8295 = n27561 ;
  assign y8296 = ~n27562 ;
  assign y8297 = n27563 ;
  assign y8298 = n27567 ;
  assign y8299 = ~n27571 ;
  assign y8300 = ~1'b0 ;
  assign y8301 = n27572 ;
  assign y8302 = n27576 ;
  assign y8303 = n27577 ;
  assign y8304 = ~n27581 ;
  assign y8305 = n27583 ;
  assign y8306 = ~n27584 ;
  assign y8307 = n27586 ;
  assign y8308 = n27588 ;
  assign y8309 = n27590 ;
  assign y8310 = ~1'b0 ;
  assign y8311 = ~n27595 ;
  assign y8312 = ~n27598 ;
  assign y8313 = n27601 ;
  assign y8314 = ~n27604 ;
  assign y8315 = ~n27607 ;
  assign y8316 = ~n27613 ;
  assign y8317 = n27618 ;
  assign y8318 = ~n27622 ;
  assign y8319 = ~n27623 ;
  assign y8320 = ~n27625 ;
  assign y8321 = ~n27626 ;
  assign y8322 = n27627 ;
  assign y8323 = ~n27628 ;
  assign y8324 = ~n27631 ;
  assign y8325 = n27635 ;
  assign y8326 = n27640 ;
  assign y8327 = ~n27642 ;
  assign y8328 = ~n27644 ;
  assign y8329 = n27648 ;
  assign y8330 = ~n27649 ;
  assign y8331 = ~1'b0 ;
  assign y8332 = ~n27651 ;
  assign y8333 = ~n27652 ;
  assign y8334 = ~n27653 ;
  assign y8335 = n27654 ;
  assign y8336 = ~n27655 ;
  assign y8337 = n27661 ;
  assign y8338 = n4641 ;
  assign y8339 = n27662 ;
  assign y8340 = ~n27663 ;
  assign y8341 = n27667 ;
  assign y8342 = n27669 ;
  assign y8343 = n27670 ;
  assign y8344 = ~n27671 ;
  assign y8345 = ~n27673 ;
  assign y8346 = ~n27674 ;
  assign y8347 = ~n27677 ;
  assign y8348 = ~n27683 ;
  assign y8349 = ~n3477 ;
  assign y8350 = n27686 ;
  assign y8351 = ~1'b0 ;
  assign y8352 = n27688 ;
  assign y8353 = ~n27690 ;
  assign y8354 = ~n27695 ;
  assign y8355 = n27698 ;
  assign y8356 = n27700 ;
  assign y8357 = ~n27702 ;
  assign y8358 = n27704 ;
  assign y8359 = ~1'b0 ;
  assign y8360 = n27707 ;
  assign y8361 = n27708 ;
  assign y8362 = ~n27714 ;
  assign y8363 = n27715 ;
  assign y8364 = n27719 ;
  assign y8365 = n27720 ;
  assign y8366 = ~n27724 ;
  assign y8367 = n27727 ;
  assign y8368 = n27731 ;
  assign y8369 = ~n27732 ;
  assign y8370 = ~n27735 ;
  assign y8371 = ~n27736 ;
  assign y8372 = ~n27737 ;
  assign y8373 = ~n27743 ;
  assign y8374 = n27746 ;
  assign y8375 = n27748 ;
  assign y8376 = ~n27750 ;
  assign y8377 = n27753 ;
  assign y8378 = ~n27754 ;
  assign y8379 = n27755 ;
  assign y8380 = ~n27756 ;
  assign y8381 = ~n27758 ;
  assign y8382 = n27765 ;
  assign y8383 = n27766 ;
  assign y8384 = ~n27769 ;
  assign y8385 = n27771 ;
  assign y8386 = ~n27772 ;
  assign y8387 = n27776 ;
  assign y8388 = n27778 ;
  assign y8389 = ~n27781 ;
  assign y8390 = ~n27785 ;
  assign y8391 = n27790 ;
  assign y8392 = ~n27792 ;
  assign y8393 = n27794 ;
  assign y8394 = n27796 ;
  assign y8395 = ~n27799 ;
  assign y8396 = n27803 ;
  assign y8397 = ~n27804 ;
  assign y8398 = n27805 ;
  assign y8399 = n27808 ;
  assign y8400 = ~n27812 ;
  assign y8401 = n27813 ;
  assign y8402 = ~n27816 ;
  assign y8403 = ~n27817 ;
  assign y8404 = ~n27818 ;
  assign y8405 = n27821 ;
  assign y8406 = ~n27824 ;
  assign y8407 = n27826 ;
  assign y8408 = ~n27828 ;
  assign y8409 = ~1'b0 ;
  assign y8410 = n27833 ;
  assign y8411 = n27836 ;
  assign y8412 = ~n27839 ;
  assign y8413 = ~n27840 ;
  assign y8414 = ~n27844 ;
  assign y8415 = n27845 ;
  assign y8416 = ~n27848 ;
  assign y8417 = ~1'b0 ;
  assign y8418 = n27849 ;
  assign y8419 = n27852 ;
  assign y8420 = ~n27855 ;
  assign y8421 = ~n27856 ;
  assign y8422 = ~n27857 ;
  assign y8423 = ~n27860 ;
  assign y8424 = ~1'b0 ;
  assign y8425 = n27863 ;
  assign y8426 = ~n27864 ;
  assign y8427 = ~n27867 ;
  assign y8428 = n27869 ;
  assign y8429 = ~n27872 ;
  assign y8430 = ~n27873 ;
  assign y8431 = n27874 ;
  assign y8432 = n27877 ;
  assign y8433 = n27880 ;
  assign y8434 = ~n27883 ;
  assign y8435 = n27885 ;
  assign y8436 = n27887 ;
  assign y8437 = n27888 ;
  assign y8438 = n27889 ;
  assign y8439 = ~n27893 ;
  assign y8440 = n27895 ;
  assign y8441 = ~n27897 ;
  assign y8442 = n27901 ;
  assign y8443 = ~1'b0 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = n27902 ;
  assign y8446 = ~n27904 ;
  assign y8447 = ~n27905 ;
  assign y8448 = n27907 ;
  assign y8449 = n27910 ;
  assign y8450 = n27911 ;
  assign y8451 = ~n27913 ;
  assign y8452 = ~n27914 ;
  assign y8453 = ~1'b0 ;
  assign y8454 = ~n27915 ;
  assign y8455 = ~n27917 ;
  assign y8456 = ~n27919 ;
  assign y8457 = n27920 ;
  assign y8458 = ~n27922 ;
  assign y8459 = n27923 ;
  assign y8460 = n27924 ;
  assign y8461 = n27927 ;
  assign y8462 = ~1'b0 ;
  assign y8463 = ~n27931 ;
  assign y8464 = ~n27933 ;
  assign y8465 = n27936 ;
  assign y8466 = ~n27938 ;
  assign y8467 = n27942 ;
  assign y8468 = n12533 ;
  assign y8469 = ~n27943 ;
  assign y8470 = ~n27944 ;
  assign y8471 = ~1'b0 ;
  assign y8472 = ~1'b0 ;
  assign y8473 = ~n27948 ;
  assign y8474 = ~n27950 ;
  assign y8475 = n27954 ;
  assign y8476 = ~n27959 ;
  assign y8477 = ~n27964 ;
  assign y8478 = ~n27966 ;
  assign y8479 = n27970 ;
  assign y8480 = ~n27975 ;
  assign y8481 = ~n27983 ;
  assign y8482 = ~n27987 ;
  assign y8483 = ~n27990 ;
  assign y8484 = ~n27993 ;
  assign y8485 = ~n27994 ;
  assign y8486 = ~n27996 ;
  assign y8487 = n28000 ;
  assign y8488 = ~n28004 ;
  assign y8489 = n28010 ;
  assign y8490 = ~1'b0 ;
  assign y8491 = n28011 ;
  assign y8492 = ~n28014 ;
  assign y8493 = ~n28015 ;
  assign y8494 = ~n28016 ;
  assign y8495 = n28017 ;
  assign y8496 = n28018 ;
  assign y8497 = n28019 ;
  assign y8498 = n28024 ;
  assign y8499 = ~n28025 ;
  assign y8500 = ~n28026 ;
  assign y8501 = n28033 ;
  assign y8502 = n28034 ;
  assign y8503 = ~n28038 ;
  assign y8504 = ~n28042 ;
  assign y8505 = ~n28043 ;
  assign y8506 = n28044 ;
  assign y8507 = n28048 ;
  assign y8508 = ~n28058 ;
  assign y8509 = n28062 ;
  assign y8510 = ~1'b0 ;
  assign y8511 = n28066 ;
  assign y8512 = n28068 ;
  assign y8513 = n22255 ;
  assign y8514 = n28071 ;
  assign y8515 = ~n28072 ;
  assign y8516 = n28073 ;
  assign y8517 = ~n28074 ;
  assign y8518 = ~1'b0 ;
  assign y8519 = ~n28077 ;
  assign y8520 = n28079 ;
  assign y8521 = n28085 ;
  assign y8522 = n28087 ;
  assign y8523 = n28096 ;
  assign y8524 = n28097 ;
  assign y8525 = n28099 ;
  assign y8526 = n28100 ;
  assign y8527 = ~n28101 ;
  assign y8528 = ~n28109 ;
  assign y8529 = ~n28113 ;
  assign y8530 = ~1'b0 ;
  assign y8531 = ~1'b0 ;
  assign y8532 = ~n28114 ;
  assign y8533 = n28115 ;
  assign y8534 = n21590 ;
  assign y8535 = ~n28119 ;
  assign y8536 = ~n28121 ;
  assign y8537 = ~n28122 ;
  assign y8538 = n28128 ;
  assign y8539 = ~n28130 ;
  assign y8540 = n28132 ;
  assign y8541 = ~n28137 ;
  assign y8542 = ~n28138 ;
  assign y8543 = n28140 ;
  assign y8544 = n28143 ;
  assign y8545 = ~n28149 ;
  assign y8546 = n28150 ;
  assign y8547 = n28152 ;
  assign y8548 = n28153 ;
  assign y8549 = ~n28155 ;
  assign y8550 = ~1'b0 ;
  assign y8551 = ~n28158 ;
  assign y8552 = n28159 ;
  assign y8553 = n28163 ;
  assign y8554 = n28165 ;
  assign y8555 = n28166 ;
  assign y8556 = n28170 ;
  assign y8557 = ~n28171 ;
  assign y8558 = ~n28173 ;
  assign y8559 = n28178 ;
  assign y8560 = n28179 ;
  assign y8561 = ~1'b0 ;
  assign y8562 = ~n28186 ;
  assign y8563 = ~n28188 ;
  assign y8564 = n28189 ;
  assign y8565 = n28194 ;
  assign y8566 = ~n28195 ;
  assign y8567 = n28198 ;
  assign y8568 = ~1'b0 ;
  assign y8569 = ~1'b0 ;
  assign y8570 = ~1'b0 ;
  assign y8571 = n28199 ;
  assign y8572 = n28201 ;
  assign y8573 = ~n28203 ;
  assign y8574 = n28204 ;
  assign y8575 = n28205 ;
  assign y8576 = ~n28206 ;
  assign y8577 = ~n28208 ;
  assign y8578 = n28211 ;
  assign y8579 = n28213 ;
  assign y8580 = n28214 ;
  assign y8581 = n28215 ;
  assign y8582 = n28220 ;
  assign y8583 = n28221 ;
  assign y8584 = ~n28222 ;
  assign y8585 = n28223 ;
  assign y8586 = n28228 ;
  assign y8587 = ~1'b0 ;
  assign y8588 = ~n28230 ;
  assign y8589 = n28241 ;
  assign y8590 = ~n28242 ;
  assign y8591 = n28244 ;
  assign y8592 = n28245 ;
  assign y8593 = n28248 ;
  assign y8594 = n28252 ;
  assign y8595 = ~n182 ;
  assign y8596 = n28253 ;
  assign y8597 = ~n28256 ;
  assign y8598 = n28258 ;
  assign y8599 = ~n28263 ;
  assign y8600 = n28264 ;
  assign y8601 = n28267 ;
  assign y8602 = n28268 ;
  assign y8603 = ~1'b0 ;
  assign y8604 = ~n28271 ;
  assign y8605 = ~n28276 ;
  assign y8606 = n28284 ;
  assign y8607 = ~n28286 ;
  assign y8608 = ~n28287 ;
  assign y8609 = ~n28288 ;
  assign y8610 = n28289 ;
  assign y8611 = n28296 ;
  assign y8612 = n28297 ;
  assign y8613 = ~1'b0 ;
  assign y8614 = ~n28302 ;
  assign y8615 = ~n28303 ;
  assign y8616 = n28304 ;
  assign y8617 = ~n28307 ;
  assign y8618 = ~n28312 ;
  assign y8619 = n28316 ;
  assign y8620 = ~n28320 ;
  assign y8621 = n28324 ;
  assign y8622 = n28328 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = n28332 ;
  assign y8625 = n28337 ;
  assign y8626 = n28339 ;
  assign y8627 = n28340 ;
  assign y8628 = n28346 ;
  assign y8629 = ~n28349 ;
  assign y8630 = ~n28350 ;
  assign y8631 = n28352 ;
  assign y8632 = ~n28353 ;
  assign y8633 = n28356 ;
  assign y8634 = n28357 ;
  assign y8635 = ~n28361 ;
  assign y8636 = n28362 ;
  assign y8637 = n28364 ;
  assign y8638 = ~n28365 ;
  assign y8639 = ~n28371 ;
  assign y8640 = ~1'b0 ;
  assign y8641 = ~n28375 ;
  assign y8642 = n28380 ;
  assign y8643 = ~n28381 ;
  assign y8644 = n28384 ;
  assign y8645 = n28385 ;
  assign y8646 = ~n28386 ;
  assign y8647 = ~n28389 ;
  assign y8648 = ~n28391 ;
  assign y8649 = ~1'b0 ;
  assign y8650 = ~1'b0 ;
  assign y8651 = ~1'b0 ;
  assign y8652 = ~n28393 ;
  assign y8653 = ~n28394 ;
  assign y8654 = ~n28398 ;
  assign y8655 = ~n28399 ;
  assign y8656 = n28401 ;
  assign y8657 = ~n28402 ;
  assign y8658 = n28403 ;
  assign y8659 = ~n28405 ;
  assign y8660 = n28408 ;
  assign y8661 = ~1'b0 ;
  assign y8662 = ~n28411 ;
  assign y8663 = ~n28418 ;
  assign y8664 = n28420 ;
  assign y8665 = n28421 ;
  assign y8666 = ~n28424 ;
  assign y8667 = n28425 ;
  assign y8668 = ~n28427 ;
  assign y8669 = ~1'b0 ;
  assign y8670 = n28428 ;
  assign y8671 = n28431 ;
  assign y8672 = n28437 ;
  assign y8673 = ~n28438 ;
  assign y8674 = n28439 ;
  assign y8675 = ~n28440 ;
  assign y8676 = ~n28444 ;
  assign y8677 = n28445 ;
  assign y8678 = ~n28447 ;
  assign y8679 = n28451 ;
  assign y8680 = n28452 ;
  assign y8681 = ~1'b0 ;
  assign y8682 = n28455 ;
  assign y8683 = n28458 ;
  assign y8684 = n28459 ;
  assign y8685 = n28460 ;
  assign y8686 = ~n28463 ;
  assign y8687 = n28469 ;
  assign y8688 = n28470 ;
  assign y8689 = ~n28474 ;
  assign y8690 = n28475 ;
  assign y8691 = n28480 ;
  assign y8692 = ~n28481 ;
  assign y8693 = ~n28487 ;
  assign y8694 = ~n28489 ;
  assign y8695 = ~n28490 ;
  assign y8696 = ~n28491 ;
  assign y8697 = ~n28493 ;
  assign y8698 = n28496 ;
  assign y8699 = ~n28501 ;
  assign y8700 = ~n28504 ;
  assign y8701 = ~1'b0 ;
  assign y8702 = ~1'b0 ;
  assign y8703 = n28505 ;
  assign y8704 = n28510 ;
  assign y8705 = ~n28514 ;
  assign y8706 = n28515 ;
  assign y8707 = ~n28517 ;
  assign y8708 = ~n28520 ;
  assign y8709 = ~1'b0 ;
  assign y8710 = ~n28522 ;
  assign y8711 = n28526 ;
  assign y8712 = ~n28534 ;
  assign y8713 = n28538 ;
  assign y8714 = ~n28541 ;
  assign y8715 = ~n28545 ;
  assign y8716 = ~1'b0 ;
  assign y8717 = ~n28548 ;
  assign y8718 = ~n28550 ;
  assign y8719 = n28553 ;
  assign y8720 = n28554 ;
  assign y8721 = ~n28557 ;
  assign y8722 = n28559 ;
  assign y8723 = ~n28562 ;
  assign y8724 = n28565 ;
  assign y8725 = ~n28566 ;
  assign y8726 = ~1'b0 ;
  assign y8727 = ~n28568 ;
  assign y8728 = ~n28569 ;
  assign y8729 = n28573 ;
  assign y8730 = n1037 ;
  assign y8731 = ~n28578 ;
  assign y8732 = ~1'b0 ;
  assign y8733 = ~n28579 ;
  assign y8734 = ~n28581 ;
  assign y8735 = n28586 ;
  assign y8736 = n28589 ;
  assign y8737 = ~n28590 ;
  assign y8738 = ~n28594 ;
  assign y8739 = n28596 ;
  assign y8740 = n28599 ;
  assign y8741 = n28605 ;
  assign y8742 = ~n28606 ;
  assign y8743 = n28608 ;
  assign y8744 = n28611 ;
  assign y8745 = ~n28613 ;
  assign y8746 = ~n28614 ;
  assign y8747 = ~n28615 ;
  assign y8748 = n28618 ;
  assign y8749 = ~1'b0 ;
  assign y8750 = ~n28622 ;
  assign y8751 = ~1'b0 ;
  assign y8752 = n28623 ;
  assign y8753 = ~1'b0 ;
  assign y8754 = n28631 ;
  assign y8755 = n28633 ;
  assign y8756 = ~n28634 ;
  assign y8757 = n28639 ;
  assign y8758 = ~n28641 ;
  assign y8759 = ~n28645 ;
  assign y8760 = ~n28647 ;
  assign y8761 = ~1'b0 ;
  assign y8762 = ~n28650 ;
  assign y8763 = n28653 ;
  assign y8764 = n28656 ;
  assign y8765 = ~n28657 ;
  assign y8766 = n28659 ;
  assign y8767 = n28661 ;
  assign y8768 = ~n28666 ;
  assign y8769 = ~n28668 ;
  assign y8770 = ~1'b0 ;
  assign y8771 = ~1'b0 ;
  assign y8772 = ~n28670 ;
  assign y8773 = n28671 ;
  assign y8774 = ~n28679 ;
  assign y8775 = n28682 ;
  assign y8776 = ~n28684 ;
  assign y8777 = ~1'b0 ;
  assign y8778 = ~1'b0 ;
  assign y8779 = ~n28685 ;
  assign y8780 = ~n28688 ;
  assign y8781 = n28690 ;
  assign y8782 = n28693 ;
  assign y8783 = n28696 ;
  assign y8784 = n28698 ;
  assign y8785 = ~n28702 ;
  assign y8786 = ~1'b0 ;
  assign y8787 = ~n28704 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~n28706 ;
  assign y8790 = n28709 ;
  assign y8791 = n28710 ;
  assign y8792 = n28711 ;
  assign y8793 = ~n28712 ;
  assign y8794 = n28716 ;
  assign y8795 = ~n28717 ;
  assign y8796 = n28724 ;
  assign y8797 = n28727 ;
  assign y8798 = ~n28729 ;
  assign y8799 = ~n28730 ;
  assign y8800 = n28731 ;
  assign y8801 = n28732 ;
  assign y8802 = ~n28734 ;
  assign y8803 = n28735 ;
  assign y8804 = ~n28738 ;
  assign y8805 = ~1'b0 ;
  assign y8806 = ~1'b0 ;
  assign y8807 = n28740 ;
  assign y8808 = ~n28742 ;
  assign y8809 = ~n28745 ;
  assign y8810 = n27609 ;
  assign y8811 = n28746 ;
  assign y8812 = ~n28747 ;
  assign y8813 = ~n28749 ;
  assign y8814 = ~1'b0 ;
  assign y8815 = n28750 ;
  assign y8816 = n28751 ;
  assign y8817 = ~n28753 ;
  assign y8818 = ~n28758 ;
  assign y8819 = ~n28759 ;
  assign y8820 = n28760 ;
  assign y8821 = n28761 ;
  assign y8822 = n28763 ;
  assign y8823 = n28765 ;
  assign y8824 = ~n28767 ;
  assign y8825 = ~1'b0 ;
  assign y8826 = ~n28771 ;
  assign y8827 = ~n28773 ;
  assign y8828 = n28774 ;
  assign y8829 = ~n28779 ;
  assign y8830 = ~n28783 ;
  assign y8831 = ~n28787 ;
  assign y8832 = ~n28789 ;
  assign y8833 = ~n28790 ;
  assign y8834 = ~n1833 ;
  assign y8835 = ~n28791 ;
  assign y8836 = ~n28794 ;
  assign y8837 = ~n28796 ;
  assign y8838 = n28797 ;
  assign y8839 = ~n28798 ;
  assign y8840 = ~n10929 ;
  assign y8841 = ~1'b0 ;
  assign y8842 = ~n28800 ;
  assign y8843 = ~1'b0 ;
  assign y8844 = ~1'b0 ;
  assign y8845 = ~n28801 ;
  assign y8846 = n28803 ;
  assign y8847 = ~n28804 ;
  assign y8848 = ~n28808 ;
  assign y8849 = n28809 ;
  assign y8850 = n28813 ;
  assign y8851 = n28817 ;
  assign y8852 = n28819 ;
  assign y8853 = ~n28821 ;
  assign y8854 = ~n28823 ;
  assign y8855 = ~n26142 ;
  assign y8856 = ~n23347 ;
  assign y8857 = n28824 ;
  assign y8858 = n28826 ;
  assign y8859 = ~1'b0 ;
  assign y8860 = ~1'b0 ;
  assign y8861 = ~n28827 ;
  assign y8862 = ~n28830 ;
  assign y8863 = ~n28832 ;
  assign y8864 = n28834 ;
  assign y8865 = n28837 ;
  assign y8866 = n28839 ;
  assign y8867 = n24437 ;
  assign y8868 = n28841 ;
  assign y8869 = n28843 ;
  assign y8870 = n28850 ;
  assign y8871 = ~n28853 ;
  assign y8872 = n28854 ;
  assign y8873 = n28856 ;
  assign y8874 = ~n28857 ;
  assign y8875 = ~n28858 ;
  assign y8876 = n28859 ;
  assign y8877 = ~n28861 ;
  assign y8878 = n28863 ;
  assign y8879 = ~1'b0 ;
  assign y8880 = n28868 ;
  assign y8881 = ~1'b0 ;
  assign y8882 = ~n28876 ;
  assign y8883 = ~n28877 ;
  assign y8884 = ~n28883 ;
  assign y8885 = ~n28887 ;
  assign y8886 = n28888 ;
  assign y8887 = ~n28891 ;
  assign y8888 = n28893 ;
  assign y8889 = ~n28898 ;
  assign y8890 = ~1'b0 ;
  assign y8891 = ~1'b0 ;
  assign y8892 = ~n28902 ;
  assign y8893 = ~n28904 ;
  assign y8894 = n28906 ;
  assign y8895 = ~n28907 ;
  assign y8896 = ~n28908 ;
  assign y8897 = n28911 ;
  assign y8898 = ~n28913 ;
  assign y8899 = ~n28915 ;
  assign y8900 = ~n28919 ;
  assign y8901 = ~n28923 ;
  assign y8902 = ~n28928 ;
  assign y8903 = ~n28929 ;
  assign y8904 = n28932 ;
  assign y8905 = n28933 ;
  assign y8906 = n28936 ;
  assign y8907 = n28937 ;
  assign y8908 = n28939 ;
  assign y8909 = ~1'b0 ;
  assign y8910 = ~n28941 ;
  assign y8911 = n28943 ;
  assign y8912 = ~n28946 ;
  assign y8913 = n28947 ;
  assign y8914 = ~n28951 ;
  assign y8915 = ~n28954 ;
  assign y8916 = n28955 ;
  assign y8917 = ~n28956 ;
  assign y8918 = ~n28957 ;
  assign y8919 = n28961 ;
  assign y8920 = n28968 ;
  assign y8921 = ~n28970 ;
  assign y8922 = ~1'b0 ;
  assign y8923 = ~n28971 ;
  assign y8924 = n28977 ;
  assign y8925 = ~n28981 ;
  assign y8926 = n28982 ;
  assign y8927 = n28983 ;
  assign y8928 = n28984 ;
  assign y8929 = ~n28992 ;
  assign y8930 = ~n28994 ;
  assign y8931 = ~n28996 ;
  assign y8932 = n28997 ;
  assign y8933 = n29002 ;
  assign y8934 = n29003 ;
  assign y8935 = n29004 ;
  assign y8936 = n29005 ;
  assign y8937 = ~n29008 ;
  assign y8938 = ~n29012 ;
  assign y8939 = ~1'b0 ;
  assign y8940 = ~1'b0 ;
  assign y8941 = ~n29013 ;
  assign y8942 = n29022 ;
  assign y8943 = n29025 ;
  assign y8944 = n29026 ;
  assign y8945 = ~n29027 ;
  assign y8946 = ~n29031 ;
  assign y8947 = ~n29032 ;
  assign y8948 = ~n29035 ;
  assign y8949 = ~n29037 ;
  assign y8950 = n29038 ;
  assign y8951 = ~x111 ;
  assign y8952 = n29039 ;
  assign y8953 = ~n29041 ;
  assign y8954 = ~n29043 ;
  assign y8955 = n29050 ;
  assign y8956 = ~n29054 ;
  assign y8957 = ~1'b0 ;
  assign y8958 = n29056 ;
  assign y8959 = ~n29059 ;
  assign y8960 = n29060 ;
  assign y8961 = ~n29064 ;
  assign y8962 = n29065 ;
  assign y8963 = n29066 ;
  assign y8964 = ~n29069 ;
  assign y8965 = n29071 ;
  assign y8966 = ~1'b0 ;
  assign y8967 = ~1'b0 ;
  assign y8968 = ~n29074 ;
  assign y8969 = ~1'b0 ;
  assign y8970 = ~n29075 ;
  assign y8971 = ~n29077 ;
  assign y8972 = ~n29078 ;
  assign y8973 = n29079 ;
  assign y8974 = n29080 ;
  assign y8975 = ~n29081 ;
  assign y8976 = ~n29086 ;
  assign y8977 = n29087 ;
  assign y8978 = ~n29089 ;
  assign y8979 = n29092 ;
  assign y8980 = ~n29093 ;
  assign y8981 = ~n29096 ;
  assign y8982 = ~n29105 ;
  assign y8983 = n29107 ;
  assign y8984 = n29110 ;
  assign y8985 = n29111 ;
  assign y8986 = n29112 ;
  assign y8987 = ~n29114 ;
  assign y8988 = n29115 ;
  assign y8989 = n29118 ;
  assign y8990 = ~n29119 ;
  assign y8991 = ~n29121 ;
  assign y8992 = ~n29122 ;
  assign y8993 = n29124 ;
  assign y8994 = n29125 ;
  assign y8995 = ~n29126 ;
  assign y8996 = ~n29129 ;
  assign y8997 = ~n29136 ;
  assign y8998 = ~n29139 ;
  assign y8999 = n29142 ;
  assign y9000 = n29144 ;
  assign y9001 = ~n29148 ;
  assign y9002 = ~n29149 ;
  assign y9003 = ~n29150 ;
  assign y9004 = ~n29151 ;
  assign y9005 = ~n29153 ;
  assign y9006 = ~1'b0 ;
  assign y9007 = ~1'b0 ;
  assign y9008 = n29154 ;
  assign y9009 = ~n29156 ;
  assign y9010 = n29159 ;
  assign y9011 = n29160 ;
  assign y9012 = n29162 ;
  assign y9013 = ~n29165 ;
  assign y9014 = ~n29169 ;
  assign y9015 = n29172 ;
  assign y9016 = n29174 ;
  assign y9017 = ~1'b0 ;
  assign y9018 = n29177 ;
  assign y9019 = ~n29179 ;
  assign y9020 = ~n29180 ;
  assign y9021 = ~n29185 ;
  assign y9022 = ~n29187 ;
  assign y9023 = n29189 ;
  assign y9024 = n29192 ;
  assign y9025 = n29195 ;
  assign y9026 = ~1'b0 ;
  assign y9027 = ~1'b0 ;
  assign y9028 = n29196 ;
  assign y9029 = n29197 ;
  assign y9030 = ~n29202 ;
  assign y9031 = ~n29208 ;
  assign y9032 = n29209 ;
  assign y9033 = n29210 ;
  assign y9034 = ~n29211 ;
  assign y9035 = n29216 ;
  assign y9036 = ~n29218 ;
  assign y9037 = ~1'b0 ;
  assign y9038 = ~n29223 ;
  assign y9039 = ~1'b0 ;
  assign y9040 = n29224 ;
  assign y9041 = n29225 ;
  assign y9042 = ~n29226 ;
  assign y9043 = ~n29230 ;
  assign y9044 = n29233 ;
  assign y9045 = n29237 ;
  assign y9046 = ~n29239 ;
  assign y9047 = n29241 ;
  assign y9048 = n29243 ;
  assign y9049 = ~1'b0 ;
  assign y9050 = n29244 ;
  assign y9051 = ~n29245 ;
  assign y9052 = n29247 ;
  assign y9053 = n29252 ;
  assign y9054 = ~n29255 ;
  assign y9055 = ~n29258 ;
  assign y9056 = ~1'b0 ;
  assign y9057 = ~1'b0 ;
  assign y9058 = ~n29259 ;
  assign y9059 = ~1'b0 ;
  assign y9060 = n29266 ;
  assign y9061 = ~n29269 ;
  assign y9062 = ~n29272 ;
  assign y9063 = ~n29273 ;
  assign y9064 = ~n29278 ;
  assign y9065 = ~n29281 ;
  assign y9066 = ~1'b0 ;
  assign y9067 = n29283 ;
  assign y9068 = ~1'b0 ;
  assign y9069 = n29285 ;
  assign y9070 = ~n29286 ;
  assign y9071 = ~n29291 ;
  assign y9072 = n29292 ;
  assign y9073 = n29296 ;
  assign y9074 = n29298 ;
  assign y9075 = n29299 ;
  assign y9076 = n29301 ;
  assign y9077 = ~n29302 ;
  assign y9078 = ~n29305 ;
  assign y9079 = ~1'b0 ;
  assign y9080 = ~n29308 ;
  assign y9081 = ~n29309 ;
  assign y9082 = ~n29310 ;
  assign y9083 = ~n29311 ;
  assign y9084 = ~n29312 ;
  assign y9085 = ~n29315 ;
  assign y9086 = n29318 ;
  assign y9087 = n29320 ;
  assign y9088 = ~1'b0 ;
  assign y9089 = ~1'b0 ;
  assign y9090 = n29323 ;
  assign y9091 = ~n29324 ;
  assign y9092 = n29327 ;
  assign y9093 = ~n29328 ;
  assign y9094 = n29330 ;
  assign y9095 = n29333 ;
  assign y9096 = ~n29334 ;
  assign y9097 = ~1'b0 ;
  assign y9098 = n29335 ;
  assign y9099 = n29337 ;
  assign y9100 = n29340 ;
  assign y9101 = ~n26160 ;
  assign y9102 = ~n29342 ;
  assign y9103 = ~n29348 ;
  assign y9104 = n29350 ;
  assign y9105 = ~n29355 ;
  assign y9106 = n29357 ;
  assign y9107 = ~1'b0 ;
  assign y9108 = ~1'b0 ;
  assign y9109 = ~1'b0 ;
  assign y9110 = ~n29361 ;
  assign y9111 = ~n29364 ;
  assign y9112 = ~n29365 ;
  assign y9113 = ~n29367 ;
  assign y9114 = n29368 ;
  assign y9115 = ~n1202 ;
  assign y9116 = ~n29371 ;
  assign y9117 = ~n29373 ;
  assign y9118 = ~1'b0 ;
  assign y9119 = ~1'b0 ;
  assign y9120 = n29376 ;
  assign y9121 = ~n29380 ;
  assign y9122 = ~n29381 ;
  assign y9123 = ~n29382 ;
  assign y9124 = n29387 ;
  assign y9125 = n29389 ;
  assign y9126 = n29392 ;
  assign y9127 = n29394 ;
  assign y9128 = ~n29396 ;
  assign y9129 = ~n29398 ;
  assign y9130 = n29399 ;
  assign y9131 = n29406 ;
  assign y9132 = n1005 ;
  assign y9133 = ~n29410 ;
  assign y9134 = n29413 ;
  assign y9135 = ~n29414 ;
  assign y9136 = ~n29422 ;
  assign y9137 = ~n29424 ;
  assign y9138 = ~n29426 ;
  assign y9139 = ~n29428 ;
  assign y9140 = ~n29431 ;
  assign y9141 = ~n29432 ;
  assign y9142 = n29433 ;
  assign y9143 = n29435 ;
  assign y9144 = n29437 ;
  assign y9145 = ~n29439 ;
  assign y9146 = ~n29441 ;
  assign y9147 = ~n29444 ;
  assign y9148 = n29451 ;
  assign y9149 = n29453 ;
  assign y9150 = ~n29455 ;
  assign y9151 = n29462 ;
  assign y9152 = ~n29465 ;
  assign y9153 = n18456 ;
  assign y9154 = ~n29466 ;
  assign y9155 = n29468 ;
  assign y9156 = ~n29474 ;
  assign y9157 = ~1'b0 ;
  assign y9158 = ~1'b0 ;
  assign y9159 = ~n29478 ;
  assign y9160 = ~n29479 ;
  assign y9161 = ~n29481 ;
  assign y9162 = ~n29484 ;
  assign y9163 = ~n29485 ;
  assign y9164 = n29488 ;
  assign y9165 = ~n29490 ;
  assign y9166 = ~n29493 ;
  assign y9167 = n29495 ;
  assign y9168 = n29496 ;
  assign y9169 = n29498 ;
  assign y9170 = ~n29499 ;
  assign y9171 = n29500 ;
  assign y9172 = n29503 ;
  assign y9173 = ~n29506 ;
  assign y9174 = ~n29510 ;
  assign y9175 = ~n29513 ;
  assign y9176 = ~n29518 ;
  assign y9177 = n29519 ;
  assign y9178 = ~n29521 ;
  assign y9179 = n29523 ;
  assign y9180 = ~1'b0 ;
  assign y9181 = ~n29525 ;
  assign y9182 = ~n29526 ;
  assign y9183 = n29536 ;
  assign y9184 = n29537 ;
  assign y9185 = ~n29539 ;
  assign y9186 = n29541 ;
  assign y9187 = n29542 ;
  assign y9188 = ~n29551 ;
  assign y9189 = ~n29552 ;
  assign y9190 = n29554 ;
  assign y9191 = ~1'b0 ;
  assign y9192 = n29556 ;
  assign y9193 = ~n29557 ;
  assign y9194 = n29558 ;
  assign y9195 = ~n29559 ;
  assign y9196 = n29560 ;
  assign y9197 = ~n29561 ;
  assign y9198 = ~n29563 ;
  assign y9199 = n29566 ;
  assign y9200 = ~n29570 ;
  assign y9201 = n29572 ;
  assign y9202 = ~n29575 ;
  assign y9203 = n29576 ;
  assign y9204 = ~n29577 ;
  assign y9205 = n29579 ;
  assign y9206 = n29582 ;
  assign y9207 = ~n29588 ;
  assign y9208 = ~n29593 ;
  assign y9209 = ~n29598 ;
  assign y9210 = ~n29600 ;
  assign y9211 = ~n29601 ;
  assign y9212 = ~n29603 ;
  assign y9213 = ~n29604 ;
  assign y9214 = n29605 ;
  assign y9215 = n29607 ;
  assign y9216 = ~n29610 ;
  assign y9217 = ~n29611 ;
  assign y9218 = ~n29613 ;
  assign y9219 = n29614 ;
  assign y9220 = ~1'b0 ;
  assign y9221 = ~n29618 ;
  assign y9222 = n29621 ;
  assign y9223 = ~n29624 ;
  assign y9224 = ~n29626 ;
  assign y9225 = n29629 ;
  assign y9226 = n29637 ;
  assign y9227 = ~n29639 ;
  assign y9228 = n29649 ;
  assign y9229 = ~n29654 ;
  assign y9230 = n29658 ;
  assign y9231 = ~n29660 ;
  assign y9232 = ~n29661 ;
  assign y9233 = ~1'b0 ;
  assign y9234 = ~n29664 ;
  assign y9235 = ~n29666 ;
  assign y9236 = ~n29670 ;
  assign y9237 = n29671 ;
  assign y9238 = ~n29673 ;
  assign y9239 = ~n29678 ;
  assign y9240 = ~n29679 ;
  assign y9241 = ~n29680 ;
  assign y9242 = ~1'b0 ;
  assign y9243 = n29681 ;
  assign y9244 = ~n29687 ;
  assign y9245 = ~n29688 ;
  assign y9246 = ~n29689 ;
  assign y9247 = ~n12617 ;
  assign y9248 = ~n29692 ;
  assign y9249 = n29694 ;
  assign y9250 = ~1'b0 ;
  assign y9251 = n29699 ;
  assign y9252 = ~1'b0 ;
  assign y9253 = ~1'b0 ;
  assign y9254 = n29703 ;
  assign y9255 = ~n29705 ;
  assign y9256 = ~n29706 ;
  assign y9257 = ~n29712 ;
  assign y9258 = ~n29713 ;
  assign y9259 = n29715 ;
  assign y9260 = ~n29717 ;
  assign y9261 = n29721 ;
  assign y9262 = ~n3454 ;
  assign y9263 = n29723 ;
  assign y9264 = ~n29727 ;
  assign y9265 = ~n29730 ;
  assign y9266 = n29739 ;
  assign y9267 = ~n29740 ;
  assign y9268 = n29747 ;
  assign y9269 = n29750 ;
  assign y9270 = n29752 ;
  assign y9271 = ~n29756 ;
  assign y9272 = n29758 ;
  assign y9273 = ~n29760 ;
  assign y9274 = n29763 ;
  assign y9275 = n29767 ;
  assign y9276 = ~n29769 ;
  assign y9277 = n29772 ;
  assign y9278 = ~n29773 ;
  assign y9279 = ~n29779 ;
  assign y9280 = n29781 ;
  assign y9281 = ~n29784 ;
  assign y9282 = n29787 ;
  assign y9283 = n29789 ;
  assign y9284 = ~n29790 ;
  assign y9285 = ~n29791 ;
  assign y9286 = n29793 ;
  assign y9287 = ~n29794 ;
  assign y9288 = n29800 ;
  assign y9289 = n29803 ;
  assign y9290 = n29804 ;
  assign y9291 = n29805 ;
  assign y9292 = ~n29807 ;
  assign y9293 = ~n29809 ;
  assign y9294 = ~n29813 ;
  assign y9295 = n29814 ;
  assign y9296 = n29815 ;
  assign y9297 = n29816 ;
  assign y9298 = ~n29817 ;
  assign y9299 = ~n29818 ;
  assign y9300 = n29822 ;
  assign y9301 = n29824 ;
  assign y9302 = ~n29832 ;
  assign y9303 = ~n29834 ;
  assign y9304 = ~n29836 ;
  assign y9305 = n29840 ;
  assign y9306 = n29841 ;
  assign y9307 = n29844 ;
  assign y9308 = n29845 ;
  assign y9309 = ~n29849 ;
  assign y9310 = n29851 ;
  assign y9311 = ~n29853 ;
  assign y9312 = ~n29855 ;
  assign y9313 = n29858 ;
  assign y9314 = ~n29861 ;
  assign y9315 = n29863 ;
  assign y9316 = ~n29865 ;
  assign y9317 = n29867 ;
  assign y9318 = ~n29871 ;
  assign y9319 = ~1'b0 ;
  assign y9320 = ~n29873 ;
  assign y9321 = n29874 ;
  assign y9322 = n29875 ;
  assign y9323 = ~n29876 ;
  assign y9324 = ~n29877 ;
  assign y9325 = n29879 ;
  assign y9326 = n29881 ;
  assign y9327 = ~n29882 ;
  assign y9328 = n29885 ;
  assign y9329 = ~n29890 ;
  assign y9330 = n29892 ;
  assign y9331 = n29894 ;
  assign y9332 = n29897 ;
  assign y9333 = ~n29899 ;
  assign y9334 = n29904 ;
  assign y9335 = n29906 ;
  assign y9336 = ~n29909 ;
  assign y9337 = ~n29911 ;
  assign y9338 = ~1'b0 ;
  assign y9339 = n29913 ;
  assign y9340 = ~1'b0 ;
  assign y9341 = ~1'b0 ;
  assign y9342 = ~n29915 ;
  assign y9343 = n29916 ;
  assign y9344 = n29918 ;
  assign y9345 = n29919 ;
  assign y9346 = n29921 ;
  assign y9347 = ~n13523 ;
  assign y9348 = ~n29926 ;
  assign y9349 = n29928 ;
  assign y9350 = n29932 ;
  assign y9351 = ~1'b0 ;
  assign y9352 = n29934 ;
  assign y9353 = n29938 ;
  assign y9354 = n29940 ;
  assign y9355 = ~n29942 ;
  assign y9356 = n29943 ;
  assign y9357 = ~n29944 ;
  assign y9358 = ~n29946 ;
  assign y9359 = ~1'b0 ;
  assign y9360 = ~1'b0 ;
  assign y9361 = n29947 ;
  assign y9362 = n29948 ;
  assign y9363 = ~n29952 ;
  assign y9364 = n29955 ;
  assign y9365 = n29956 ;
  assign y9366 = ~n29957 ;
  assign y9367 = n29960 ;
  assign y9368 = ~1'b0 ;
  assign y9369 = ~n29962 ;
  assign y9370 = ~1'b0 ;
  assign y9371 = ~n29964 ;
  assign y9372 = n29967 ;
  assign y9373 = n29970 ;
  assign y9374 = ~n29972 ;
  assign y9375 = ~n29974 ;
  assign y9376 = ~n29980 ;
  assign y9377 = n29981 ;
  assign y9378 = n29984 ;
  assign y9379 = ~n29988 ;
  assign y9380 = n29992 ;
  assign y9381 = n29994 ;
  assign y9382 = n29995 ;
  assign y9383 = n29996 ;
  assign y9384 = ~n29999 ;
  assign y9385 = ~n30004 ;
  assign y9386 = ~n30007 ;
  assign y9387 = ~n30009 ;
  assign y9388 = ~n30016 ;
  assign y9389 = n30020 ;
  assign y9390 = ~n30022 ;
  assign y9391 = ~1'b0 ;
  assign y9392 = ~n30025 ;
  assign y9393 = ~n30028 ;
  assign y9394 = ~n30032 ;
  assign y9395 = n30038 ;
  assign y9396 = ~n30039 ;
  assign y9397 = n30040 ;
  assign y9398 = n30042 ;
  assign y9399 = ~1'b0 ;
  assign y9400 = n30044 ;
  assign y9401 = n30045 ;
  assign y9402 = ~n30046 ;
  assign y9403 = n30051 ;
  assign y9404 = n30052 ;
  assign y9405 = ~n30053 ;
  assign y9406 = ~n30055 ;
  assign y9407 = ~n30063 ;
  assign y9408 = n30064 ;
  assign y9409 = n30066 ;
  assign y9410 = n30068 ;
  assign y9411 = ~1'b0 ;
  assign y9412 = n30071 ;
  assign y9413 = ~n30072 ;
  assign y9414 = ~n30073 ;
  assign y9415 = ~n30075 ;
  assign y9416 = ~n30079 ;
  assign y9417 = ~n30080 ;
  assign y9418 = n30082 ;
  assign y9419 = ~n30084 ;
  assign y9420 = ~n30087 ;
  assign y9421 = n30089 ;
  assign y9422 = ~n30091 ;
  assign y9423 = ~1'b0 ;
  assign y9424 = n30092 ;
  assign y9425 = ~n30094 ;
  assign y9426 = n30099 ;
  assign y9427 = n30100 ;
  assign y9428 = ~n30101 ;
  assign y9429 = n30105 ;
  assign y9430 = ~n30106 ;
  assign y9431 = ~n30108 ;
  assign y9432 = ~n30110 ;
  assign y9433 = ~n30114 ;
  assign y9434 = n30117 ;
  assign y9435 = n30118 ;
  assign y9436 = ~n30120 ;
  assign y9437 = n30128 ;
  assign y9438 = n30131 ;
  assign y9439 = n30132 ;
  assign y9440 = n30133 ;
  assign y9441 = ~1'b0 ;
  assign y9442 = n30135 ;
  assign y9443 = n30137 ;
  assign y9444 = ~1'b0 ;
  assign y9445 = ~n30138 ;
  assign y9446 = n30139 ;
  assign y9447 = ~n30141 ;
  assign y9448 = ~n30143 ;
  assign y9449 = ~n30150 ;
  assign y9450 = ~n30152 ;
  assign y9451 = n30155 ;
  assign y9452 = ~1'b0 ;
  assign y9453 = ~n30159 ;
  assign y9454 = n30161 ;
  assign y9455 = ~n30166 ;
  assign y9456 = n30167 ;
  assign y9457 = n30171 ;
  assign y9458 = n30172 ;
  assign y9459 = ~n30174 ;
  assign y9460 = n30175 ;
  assign y9461 = ~n30177 ;
  assign y9462 = ~n30180 ;
  assign y9463 = ~n30182 ;
  assign y9464 = ~1'b0 ;
  assign y9465 = ~n30185 ;
  assign y9466 = ~n30186 ;
  assign y9467 = n30187 ;
  assign y9468 = ~n30188 ;
  assign y9469 = ~1'b0 ;
  assign y9470 = ~n30190 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = n30196 ;
  assign y9473 = ~n30197 ;
  assign y9474 = ~n30199 ;
  assign y9475 = n30203 ;
  assign y9476 = ~n30207 ;
  assign y9477 = n30211 ;
  assign y9478 = ~n27969 ;
  assign y9479 = ~n30212 ;
  assign y9480 = ~1'b0 ;
  assign y9481 = ~n30214 ;
  assign y9482 = ~n30216 ;
  assign y9483 = ~1'b0 ;
  assign y9484 = ~n30217 ;
  assign y9485 = ~n30220 ;
  assign y9486 = n30222 ;
  assign y9487 = ~n30225 ;
  assign y9488 = n30228 ;
  assign y9489 = ~n30229 ;
  assign y9490 = n30233 ;
  assign y9491 = n30235 ;
  assign y9492 = n30236 ;
  assign y9493 = n30241 ;
  assign y9494 = ~n30242 ;
  assign y9495 = n30243 ;
  assign y9496 = n30248 ;
  assign y9497 = n30249 ;
  assign y9498 = ~n30251 ;
  assign y9499 = ~n30252 ;
  assign y9500 = ~n30257 ;
  assign y9501 = ~n30259 ;
  assign y9502 = ~n30261 ;
  assign y9503 = n30263 ;
  assign y9504 = ~n30265 ;
  assign y9505 = n30266 ;
  assign y9506 = n30267 ;
  assign y9507 = n30268 ;
  assign y9508 = ~n30271 ;
  assign y9509 = ~n30277 ;
  assign y9510 = n30279 ;
  assign y9511 = ~n30281 ;
  assign y9512 = n30283 ;
  assign y9513 = ~1'b0 ;
  assign y9514 = n30285 ;
  assign y9515 = ~n30287 ;
  assign y9516 = n30288 ;
  assign y9517 = ~n30289 ;
  assign y9518 = ~n30290 ;
  assign y9519 = n30292 ;
  assign y9520 = ~n30294 ;
  assign y9521 = ~n30296 ;
  assign y9522 = n30298 ;
  assign y9523 = ~1'b0 ;
  assign y9524 = ~1'b0 ;
  assign y9525 = ~n30302 ;
  assign y9526 = ~n30303 ;
  assign y9527 = n30305 ;
  assign y9528 = n30306 ;
  assign y9529 = ~n30307 ;
  assign y9530 = n30310 ;
  assign y9531 = ~n30313 ;
  assign y9532 = n30314 ;
  assign y9533 = n9251 ;
  assign y9534 = ~n30318 ;
  assign y9535 = n30320 ;
  assign y9536 = n30324 ;
  assign y9537 = ~n30325 ;
  assign y9538 = ~n30328 ;
  assign y9539 = n30331 ;
  assign y9540 = ~n30332 ;
  assign y9541 = n30333 ;
  assign y9542 = n30338 ;
  assign y9543 = ~n30339 ;
  assign y9544 = ~n30344 ;
  assign y9545 = n30347 ;
  assign y9546 = ~1'b0 ;
  assign y9547 = ~n30350 ;
  assign y9548 = ~n30353 ;
  assign y9549 = n30354 ;
  assign y9550 = ~n30355 ;
  assign y9551 = ~n30360 ;
  assign y9552 = ~n30361 ;
  assign y9553 = ~n30363 ;
  assign y9554 = ~n30366 ;
  assign y9555 = ~1'b0 ;
  assign y9556 = n30368 ;
  assign y9557 = ~n30370 ;
  assign y9558 = ~1'b0 ;
  assign y9559 = ~n30371 ;
  assign y9560 = ~n30373 ;
  assign y9561 = ~n30377 ;
  assign y9562 = n30383 ;
  assign y9563 = ~n30385 ;
  assign y9564 = ~n28002 ;
  assign y9565 = n30387 ;
  assign y9566 = ~1'b0 ;
  assign y9567 = ~n30389 ;
  assign y9568 = n30395 ;
  assign y9569 = ~n30396 ;
  assign y9570 = n30398 ;
  assign y9571 = n30399 ;
  assign y9572 = ~n30400 ;
  assign y9573 = n30403 ;
  assign y9574 = n30409 ;
  assign y9575 = n30413 ;
  assign y9576 = n30416 ;
  assign y9577 = n30418 ;
  assign y9578 = ~1'b0 ;
  assign y9579 = ~n30421 ;
  assign y9580 = ~n30425 ;
  assign y9581 = n30426 ;
  assign y9582 = n30429 ;
  assign y9583 = n30433 ;
  assign y9584 = ~n30436 ;
  assign y9585 = n30440 ;
  assign y9586 = ~n30444 ;
  assign y9587 = ~n30449 ;
  assign y9588 = ~n30451 ;
  assign y9589 = ~n30456 ;
  assign y9590 = ~n30463 ;
  assign y9591 = ~n30466 ;
  assign y9592 = ~n30468 ;
  assign y9593 = n30469 ;
  assign y9594 = ~n30476 ;
  assign y9595 = n30480 ;
  assign y9596 = ~n30484 ;
  assign y9597 = ~n30487 ;
  assign y9598 = ~n30491 ;
  assign y9599 = ~n30492 ;
  assign y9600 = ~n30494 ;
  assign y9601 = n30497 ;
  assign y9602 = ~n30499 ;
  assign y9603 = n24379 ;
  assign y9604 = n7412 ;
  assign y9605 = ~n30500 ;
  assign y9606 = n30503 ;
  assign y9607 = ~n30506 ;
  assign y9608 = n30509 ;
  assign y9609 = ~n30510 ;
  assign y9610 = n30511 ;
  assign y9611 = n30514 ;
  assign y9612 = n30517 ;
  assign y9613 = n30521 ;
  assign y9614 = n30526 ;
  assign y9615 = ~n30534 ;
  assign y9616 = ~n30536 ;
  assign y9617 = n30537 ;
  assign y9618 = ~n30538 ;
  assign y9619 = ~n30539 ;
  assign y9620 = n30540 ;
  assign y9621 = ~n30542 ;
  assign y9622 = ~n30544 ;
  assign y9623 = ~n30551 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = n30552 ;
  assign y9626 = n30555 ;
  assign y9627 = n30559 ;
  assign y9628 = ~n30561 ;
  assign y9629 = ~n30562 ;
  assign y9630 = ~n30569 ;
  assign y9631 = ~n30574 ;
  assign y9632 = ~n30576 ;
  assign y9633 = ~n30578 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = ~1'b0 ;
  assign y9636 = n30579 ;
  assign y9637 = ~n30581 ;
  assign y9638 = n30582 ;
  assign y9639 = n30585 ;
  assign y9640 = n30586 ;
  assign y9641 = n30588 ;
  assign y9642 = ~n30589 ;
  assign y9643 = n30591 ;
  assign y9644 = ~1'b0 ;
  assign y9645 = ~n30593 ;
  assign y9646 = ~1'b0 ;
  assign y9647 = n30601 ;
  assign y9648 = ~n30603 ;
  assign y9649 = ~n30608 ;
  assign y9650 = ~n30609 ;
  assign y9651 = n30610 ;
  assign y9652 = n30614 ;
  assign y9653 = n30617 ;
  assign y9654 = n30619 ;
  assign y9655 = ~n30621 ;
  assign y9656 = n30626 ;
  assign y9657 = n30632 ;
  assign y9658 = n30633 ;
  assign y9659 = n30634 ;
  assign y9660 = ~n30635 ;
  assign y9661 = n10118 ;
  assign y9662 = n30636 ;
  assign y9663 = n30637 ;
  assign y9664 = n30639 ;
  assign y9665 = ~1'b0 ;
  assign y9666 = n30641 ;
  assign y9667 = ~1'b0 ;
  assign y9668 = ~n30643 ;
  assign y9669 = ~n30645 ;
  assign y9670 = n30647 ;
  assign y9671 = n30655 ;
  assign y9672 = n30656 ;
  assign y9673 = ~n30661 ;
  assign y9674 = ~n30664 ;
  assign y9675 = n30665 ;
  assign y9676 = n30669 ;
  assign y9677 = ~n30671 ;
  assign y9678 = ~1'b0 ;
  assign y9679 = n30675 ;
  assign y9680 = n30676 ;
  assign y9681 = n30677 ;
  assign y9682 = n30678 ;
  assign y9683 = n30679 ;
  assign y9684 = ~n30681 ;
  assign y9685 = n30683 ;
  assign y9686 = ~n30685 ;
  assign y9687 = ~n30687 ;
  assign y9688 = ~1'b0 ;
  assign y9689 = ~1'b0 ;
  assign y9690 = ~n30689 ;
  assign y9691 = n30690 ;
  assign y9692 = n30691 ;
  assign y9693 = ~n30692 ;
  assign y9694 = ~n30697 ;
  assign y9695 = n30700 ;
  assign y9696 = n30702 ;
  assign y9697 = ~n30703 ;
  assign y9698 = n30706 ;
  assign y9699 = n30707 ;
  assign y9700 = ~n30710 ;
  assign y9701 = ~n30711 ;
  assign y9702 = ~n30714 ;
  assign y9703 = ~n30715 ;
  assign y9704 = n30716 ;
  assign y9705 = n30718 ;
  assign y9706 = n30719 ;
  assign y9707 = n30720 ;
  assign y9708 = n30721 ;
  assign y9709 = ~1'b0 ;
  assign y9710 = ~n30723 ;
  assign y9711 = ~n30727 ;
  assign y9712 = ~n30729 ;
  assign y9713 = ~n30734 ;
  assign y9714 = ~n30737 ;
  assign y9715 = n30740 ;
  assign y9716 = ~n30743 ;
  assign y9717 = n30745 ;
  assign y9718 = ~n30749 ;
  assign y9719 = n30753 ;
  assign y9720 = n30755 ;
  assign y9721 = n30759 ;
  assign y9722 = ~n30762 ;
  assign y9723 = n30767 ;
  assign y9724 = n30776 ;
  assign y9725 = ~n30780 ;
  assign y9726 = ~n30781 ;
  assign y9727 = ~n30792 ;
  assign y9728 = ~1'b0 ;
  assign y9729 = n30793 ;
  assign y9730 = ~n30795 ;
  assign y9731 = ~n30797 ;
  assign y9732 = ~n30798 ;
  assign y9733 = n30799 ;
  assign y9734 = n30800 ;
  assign y9735 = n30801 ;
  assign y9736 = n30806 ;
  assign y9737 = ~n30809 ;
  assign y9738 = ~n30811 ;
  assign y9739 = ~1'b0 ;
  assign y9740 = n30814 ;
  assign y9741 = ~n30817 ;
  assign y9742 = n30819 ;
  assign y9743 = ~n30821 ;
  assign y9744 = n30825 ;
  assign y9745 = ~n30828 ;
  assign y9746 = ~n30832 ;
  assign y9747 = ~n30833 ;
  assign y9748 = n17519 ;
  assign y9749 = ~1'b0 ;
  assign y9750 = n30837 ;
  assign y9751 = ~n30839 ;
  assign y9752 = ~n30841 ;
  assign y9753 = n30845 ;
  assign y9754 = n30846 ;
  assign y9755 = ~n30849 ;
  assign y9756 = ~n30851 ;
  assign y9757 = ~n30855 ;
  assign y9758 = n30858 ;
  assign y9759 = n30860 ;
  assign y9760 = ~1'b0 ;
  assign y9761 = ~n30862 ;
  assign y9762 = ~n30864 ;
  assign y9763 = n30867 ;
  assign y9764 = n30868 ;
  assign y9765 = n30871 ;
  assign y9766 = n30873 ;
  assign y9767 = ~1'b0 ;
  assign y9768 = ~1'b0 ;
  assign y9769 = n30878 ;
  assign y9770 = ~1'b0 ;
  assign y9771 = n30879 ;
  assign y9772 = ~n30880 ;
  assign y9773 = ~n30885 ;
  assign y9774 = n30886 ;
  assign y9775 = ~n30889 ;
  assign y9776 = n30890 ;
  assign y9777 = ~n30892 ;
  assign y9778 = ~n30894 ;
  assign y9779 = ~1'b0 ;
  assign y9780 = n30895 ;
  assign y9781 = ~n30898 ;
  assign y9782 = n30899 ;
  assign y9783 = ~n30903 ;
  assign y9784 = n30907 ;
  assign y9785 = n30910 ;
  assign y9786 = n30911 ;
  assign y9787 = n30912 ;
  assign y9788 = ~n30914 ;
  assign y9789 = n30918 ;
  assign y9790 = ~1'b0 ;
  assign y9791 = ~n30920 ;
  assign y9792 = ~1'b0 ;
  assign y9793 = n30921 ;
  assign y9794 = n30923 ;
  assign y9795 = ~x9 ;
  assign y9796 = ~n30928 ;
  assign y9797 = ~n30930 ;
  assign y9798 = n30931 ;
  assign y9799 = n30932 ;
  assign y9800 = n30933 ;
  assign y9801 = n30935 ;
  assign y9802 = n30937 ;
  assign y9803 = ~1'b0 ;
  assign y9804 = ~n30939 ;
  assign y9805 = n30940 ;
  assign y9806 = ~n30941 ;
  assign y9807 = ~n30942 ;
  assign y9808 = ~n30943 ;
  assign y9809 = ~n30944 ;
  assign y9810 = n30947 ;
  assign y9811 = ~1'b0 ;
  assign y9812 = ~n30948 ;
  assign y9813 = ~1'b0 ;
  assign y9814 = n30949 ;
  assign y9815 = ~n30953 ;
  assign y9816 = ~n30957 ;
  assign y9817 = n30958 ;
  assign y9818 = n30959 ;
  assign y9819 = n30961 ;
  assign y9820 = n30962 ;
  assign y9821 = ~n30964 ;
  assign y9822 = ~1'b0 ;
  assign y9823 = n30966 ;
  assign y9824 = n30970 ;
  assign y9825 = ~n30973 ;
  assign y9826 = n30982 ;
  assign y9827 = n30983 ;
  assign y9828 = n30985 ;
  assign y9829 = ~n30986 ;
  assign y9830 = n30989 ;
  assign y9831 = ~n30994 ;
  assign y9832 = ~n30997 ;
  assign y9833 = n30999 ;
  assign y9834 = n31003 ;
  assign y9835 = ~n31004 ;
  assign y9836 = n31005 ;
  assign y9837 = n31010 ;
  assign y9838 = ~n31012 ;
  assign y9839 = n31014 ;
  assign y9840 = n31017 ;
  assign y9841 = n31019 ;
  assign y9842 = ~1'b0 ;
  assign y9843 = n31022 ;
  assign y9844 = ~n31024 ;
  assign y9845 = ~n31025 ;
  assign y9846 = n31026 ;
  assign y9847 = ~n31031 ;
  assign y9848 = n31035 ;
  assign y9849 = n31036 ;
  assign y9850 = n31037 ;
  assign y9851 = ~n31039 ;
  assign y9852 = n18263 ;
  assign y9853 = ~n31042 ;
  assign y9854 = ~1'b0 ;
  assign y9855 = n31044 ;
  assign y9856 = ~n31045 ;
  assign y9857 = n31047 ;
  assign y9858 = n31052 ;
  assign y9859 = ~n31053 ;
  assign y9860 = ~n31055 ;
  assign y9861 = ~n31056 ;
  assign y9862 = ~n31058 ;
  assign y9863 = ~n31060 ;
  assign y9864 = ~1'b0 ;
  assign y9865 = ~n31062 ;
  assign y9866 = n31064 ;
  assign y9867 = ~n31068 ;
  assign y9868 = n31070 ;
  assign y9869 = n31073 ;
  assign y9870 = n31082 ;
  assign y9871 = n31087 ;
  assign y9872 = ~1'b0 ;
  assign y9873 = n31090 ;
  assign y9874 = ~n31094 ;
  assign y9875 = ~1'b0 ;
  assign y9876 = ~n31096 ;
  assign y9877 = ~n31098 ;
  assign y9878 = n31100 ;
  assign y9879 = n31110 ;
  assign y9880 = ~n31111 ;
  assign y9881 = n31112 ;
  assign y9882 = n31113 ;
  assign y9883 = ~n31119 ;
  assign y9884 = ~n31121 ;
  assign y9885 = ~1'b0 ;
  assign y9886 = n31123 ;
  assign y9887 = ~1'b0 ;
  assign y9888 = n3821 ;
  assign y9889 = n31124 ;
  assign y9890 = ~n31125 ;
  assign y9891 = ~n31127 ;
  assign y9892 = ~n31128 ;
  assign y9893 = n31130 ;
  assign y9894 = n31131 ;
  assign y9895 = n31132 ;
  assign y9896 = ~1'b0 ;
  assign y9897 = n31134 ;
  assign y9898 = ~1'b0 ;
  assign y9899 = ~n31135 ;
  assign y9900 = ~n31137 ;
  assign y9901 = ~n31138 ;
  assign y9902 = n31141 ;
  assign y9903 = n31142 ;
  assign y9904 = n31144 ;
  assign y9905 = ~n31147 ;
  assign y9906 = ~1'b0 ;
  assign y9907 = ~1'b0 ;
  assign y9908 = n31149 ;
  assign y9909 = n31152 ;
  assign y9910 = n31157 ;
  assign y9911 = n31158 ;
  assign y9912 = n31159 ;
  assign y9913 = ~n31162 ;
  assign y9914 = n31163 ;
  assign y9915 = n31168 ;
  assign y9916 = ~n31169 ;
  assign y9917 = ~1'b0 ;
  assign y9918 = ~1'b0 ;
  assign y9919 = n31170 ;
  assign y9920 = n31171 ;
  assign y9921 = n31175 ;
  assign y9922 = n31176 ;
  assign y9923 = ~n31177 ;
  assign y9924 = ~n31180 ;
  assign y9925 = n31183 ;
  assign y9926 = ~n31185 ;
  assign y9927 = ~n31188 ;
  assign y9928 = ~1'b0 ;
  assign y9929 = ~n31190 ;
  assign y9930 = n14060 ;
  assign y9931 = n31193 ;
  assign y9932 = n31195 ;
  assign y9933 = ~n31197 ;
  assign y9934 = ~n31198 ;
  assign y9935 = ~n31199 ;
  assign y9936 = n31200 ;
  assign y9937 = n31203 ;
  assign y9938 = ~n31205 ;
  assign y9939 = n31207 ;
  assign y9940 = n31209 ;
  assign y9941 = ~n31213 ;
  assign y9942 = n31219 ;
  assign y9943 = ~n31223 ;
  assign y9944 = ~n31226 ;
  assign y9945 = ~n31228 ;
  assign y9946 = ~n31230 ;
  assign y9947 = ~n31231 ;
  assign y9948 = ~1'b0 ;
  assign y9949 = ~n31236 ;
  assign y9950 = ~1'b0 ;
  assign y9951 = ~1'b0 ;
  assign y9952 = n31240 ;
  assign y9953 = ~n31243 ;
  assign y9954 = n31247 ;
  assign y9955 = n31248 ;
  assign y9956 = n31253 ;
  assign y9957 = ~n31254 ;
  assign y9958 = ~n31259 ;
  assign y9959 = n31261 ;
  assign y9960 = n31263 ;
  assign y9961 = ~n31266 ;
  assign y9962 = n31270 ;
  assign y9963 = n31271 ;
  assign y9964 = ~n31274 ;
  assign y9965 = n31278 ;
  assign y9966 = n31279 ;
  assign y9967 = n31281 ;
  assign y9968 = ~n31290 ;
  assign y9969 = ~1'b0 ;
  assign y9970 = ~n31292 ;
  assign y9971 = n31293 ;
  assign y9972 = n31300 ;
  assign y9973 = n31303 ;
  assign y9974 = n31306 ;
  assign y9975 = ~n31307 ;
  assign y9976 = ~n31311 ;
  assign y9977 = n31312 ;
  assign y9978 = ~n31313 ;
  assign y9979 = n31318 ;
  assign y9980 = ~n31324 ;
  assign y9981 = n31326 ;
  assign y9982 = ~1'b0 ;
  assign y9983 = n31328 ;
  assign y9984 = n31330 ;
  assign y9985 = n31332 ;
  assign y9986 = n31336 ;
  assign y9987 = ~n31340 ;
  assign y9988 = n31341 ;
  assign y9989 = ~n31343 ;
  assign y9990 = n31346 ;
  assign y9991 = n31349 ;
  assign y9992 = ~1'b0 ;
  assign y9993 = n31351 ;
  assign y9994 = ~1'b0 ;
  assign y9995 = ~n31352 ;
  assign y9996 = n31355 ;
  assign y9997 = n31362 ;
  assign y9998 = n31363 ;
  assign y9999 = ~n31364 ;
  assign y10000 = ~n31366 ;
  assign y10001 = n31367 ;
  assign y10002 = ~n31373 ;
  assign y10003 = n31377 ;
  assign y10004 = ~n31379 ;
  assign y10005 = ~1'b0 ;
  assign y10006 = ~n31380 ;
  assign y10007 = n31385 ;
  assign y10008 = ~n31387 ;
  assign y10009 = n31388 ;
  assign y10010 = ~n31389 ;
  assign y10011 = ~n31390 ;
  assign y10012 = ~n31392 ;
  assign y10013 = ~n31396 ;
  assign y10014 = ~n31397 ;
  assign y10015 = ~n31400 ;
  assign y10016 = n31402 ;
  assign y10017 = ~n31403 ;
  assign y10018 = n31405 ;
  assign y10019 = ~n31407 ;
  assign y10020 = ~n31408 ;
  assign y10021 = n31411 ;
  assign y10022 = ~n31412 ;
  assign y10023 = n31414 ;
  assign y10024 = ~1'b0 ;
  assign y10025 = ~n31416 ;
  assign y10026 = ~n31419 ;
  assign y10027 = ~n31424 ;
  assign y10028 = ~n31430 ;
  assign y10029 = n31431 ;
  assign y10030 = ~n31433 ;
  assign y10031 = n31434 ;
  assign y10032 = n31435 ;
  assign y10033 = n31443 ;
  assign y10034 = ~n31444 ;
  assign y10035 = ~n31447 ;
  assign y10036 = n31450 ;
  assign y10037 = n31452 ;
  assign y10038 = n31453 ;
  assign y10039 = n31454 ;
  assign y10040 = ~n31455 ;
  assign y10041 = n31459 ;
  assign y10042 = n31465 ;
  assign y10043 = ~n31467 ;
  assign y10044 = ~n31470 ;
  assign y10045 = ~n31472 ;
  assign y10046 = n31476 ;
  assign y10047 = n31478 ;
  assign y10048 = ~1'b0 ;
  assign y10049 = ~n31480 ;
  assign y10050 = ~n31484 ;
  assign y10051 = n31486 ;
  assign y10052 = n31489 ;
  assign y10053 = n31490 ;
  assign y10054 = ~n31491 ;
  assign y10055 = ~n31496 ;
  assign y10056 = ~1'b0 ;
  assign y10057 = ~1'b0 ;
  assign y10058 = ~1'b0 ;
  assign y10059 = n31498 ;
  assign y10060 = n31500 ;
  assign y10061 = ~n31503 ;
  assign y10062 = ~n31504 ;
  assign y10063 = n31506 ;
  assign y10064 = n31507 ;
  assign y10065 = ~n31508 ;
  assign y10066 = ~n31510 ;
  assign y10067 = ~n31512 ;
  assign y10068 = ~n31523 ;
  assign y10069 = ~1'b0 ;
  assign y10070 = n31524 ;
  assign y10071 = ~n31531 ;
  assign y10072 = ~n31532 ;
  assign y10073 = n31533 ;
  assign y10074 = ~n31534 ;
  assign y10075 = n31535 ;
  assign y10076 = ~n31536 ;
  assign y10077 = n31539 ;
  assign y10078 = n31550 ;
  assign y10079 = ~n31554 ;
  assign y10080 = ~1'b0 ;
  assign y10081 = n31558 ;
  assign y10082 = ~n31560 ;
  assign y10083 = n31561 ;
  assign y10084 = n31562 ;
  assign y10085 = n31564 ;
  assign y10086 = ~n31566 ;
  assign y10087 = n31567 ;
  assign y10088 = n31569 ;
  assign y10089 = n31570 ;
  assign y10090 = n31577 ;
  assign y10091 = ~n31579 ;
  assign y10092 = n31585 ;
  assign y10093 = ~n31586 ;
  assign y10094 = ~n31590 ;
  assign y10095 = n31592 ;
  assign y10096 = ~n31594 ;
  assign y10097 = n31595 ;
  assign y10098 = n31597 ;
  assign y10099 = n31599 ;
  assign y10100 = ~n31606 ;
  assign y10101 = ~n31609 ;
  assign y10102 = ~n31611 ;
  assign y10103 = ~n31612 ;
  assign y10104 = ~n31613 ;
  assign y10105 = ~n31614 ;
  assign y10106 = ~n31616 ;
  assign y10107 = ~n31617 ;
  assign y10108 = n31620 ;
  assign y10109 = n31621 ;
  assign y10110 = ~n31624 ;
  assign y10111 = n31626 ;
  assign y10112 = ~1'b0 ;
  assign y10113 = ~1'b0 ;
  assign y10114 = n31627 ;
  assign y10115 = n31631 ;
  assign y10116 = n31633 ;
  assign y10117 = n31634 ;
  assign y10118 = ~n31638 ;
  assign y10119 = ~n31641 ;
  assign y10120 = ~n31645 ;
  assign y10121 = ~n31648 ;
  assign y10122 = ~n31650 ;
  assign y10123 = n31652 ;
  assign y10124 = n31655 ;
  assign y10125 = ~n31656 ;
  assign y10126 = n31661 ;
  assign y10127 = ~n31664 ;
  assign y10128 = n31665 ;
  assign y10129 = n31666 ;
  assign y10130 = ~n31667 ;
  assign y10131 = ~n31669 ;
  assign y10132 = n31671 ;
  assign y10133 = ~1'b0 ;
  assign y10134 = n31672 ;
  assign y10135 = n31674 ;
  assign y10136 = ~n31675 ;
  assign y10137 = ~n31677 ;
  assign y10138 = ~n31678 ;
  assign y10139 = n31679 ;
  assign y10140 = n31683 ;
  assign y10141 = ~n31684 ;
  assign y10142 = ~n31687 ;
  assign y10143 = n31688 ;
  assign y10144 = ~1'b0 ;
  assign y10145 = n31691 ;
  assign y10146 = ~n31693 ;
  assign y10147 = ~n31698 ;
  assign y10148 = ~n31700 ;
  assign y10149 = n31702 ;
  assign y10150 = ~n31703 ;
  assign y10151 = ~n31708 ;
  assign y10152 = ~n31709 ;
  assign y10153 = ~n31711 ;
  assign y10154 = ~n31712 ;
  assign y10155 = ~1'b0 ;
  assign y10156 = ~n31714 ;
  assign y10157 = ~n31715 ;
  assign y10158 = ~n31717 ;
  assign y10159 = n31723 ;
  assign y10160 = n31725 ;
  assign y10161 = n31730 ;
  assign y10162 = ~n31733 ;
  assign y10163 = n31738 ;
  assign y10164 = ~n31739 ;
  assign y10165 = n31743 ;
  assign y10166 = 1'b0 ;
  assign y10167 = ~n31745 ;
  assign y10168 = ~1'b0 ;
  assign y10169 = n31750 ;
  assign y10170 = n31751 ;
  assign y10171 = ~n31756 ;
  assign y10172 = ~n31757 ;
  assign y10173 = n31758 ;
  assign y10174 = ~n31761 ;
  assign y10175 = ~n31762 ;
  assign y10176 = n31764 ;
  assign y10177 = ~1'b0 ;
  assign y10178 = n31765 ;
  assign y10179 = ~n31766 ;
  assign y10180 = n31767 ;
  assign y10181 = n31771 ;
  assign y10182 = n31776 ;
  assign y10183 = n31781 ;
  assign y10184 = n31785 ;
  assign y10185 = ~n31786 ;
  assign y10186 = n31790 ;
  assign y10187 = ~n31791 ;
  assign y10188 = ~n31793 ;
  assign y10189 = ~n31795 ;
  assign y10190 = ~1'b0 ;
  assign y10191 = ~n31797 ;
  assign y10192 = ~1'b0 ;
  assign y10193 = n31799 ;
  assign y10194 = ~n31803 ;
  assign y10195 = n31805 ;
  assign y10196 = ~n31808 ;
  assign y10197 = ~n31809 ;
  assign y10198 = n31815 ;
  assign y10199 = n31818 ;
  assign y10200 = ~n31821 ;
  assign y10201 = ~1'b0 ;
  assign y10202 = n31822 ;
  assign y10203 = n31825 ;
  assign y10204 = n31826 ;
  assign y10205 = n31827 ;
  assign y10206 = ~n31828 ;
  assign y10207 = ~n31829 ;
  assign y10208 = n31830 ;
  assign y10209 = n31832 ;
  assign y10210 = ~1'b0 ;
  assign y10211 = n31834 ;
  assign y10212 = ~n31836 ;
  assign y10213 = ~n31837 ;
  assign y10214 = ~n31840 ;
  assign y10215 = n31841 ;
  assign y10216 = ~n31849 ;
  assign y10217 = n10845 ;
  assign y10218 = ~n31851 ;
  assign y10219 = n31855 ;
  assign y10220 = ~n31856 ;
  assign y10221 = ~n31858 ;
  assign y10222 = ~n31863 ;
  assign y10223 = ~n31866 ;
  assign y10224 = n31867 ;
  assign y10225 = n31868 ;
  assign y10226 = n31871 ;
  assign y10227 = ~n31873 ;
  assign y10228 = n31874 ;
  assign y10229 = n31879 ;
  assign y10230 = ~n31880 ;
  assign y10231 = n31882 ;
  assign y10232 = n31884 ;
  assign y10233 = n31886 ;
  assign y10234 = n31891 ;
  assign y10235 = n31892 ;
  assign y10236 = n31895 ;
  assign y10237 = n31896 ;
  assign y10238 = ~n31899 ;
  assign y10239 = ~n31903 ;
  assign y10240 = n31904 ;
  assign y10241 = ~n31905 ;
  assign y10242 = n31907 ;
  assign y10243 = ~n798 ;
  assign y10244 = ~1'b0 ;
  assign y10245 = ~n31908 ;
  assign y10246 = ~n31911 ;
  assign y10247 = n31912 ;
  assign y10248 = n31915 ;
  assign y10249 = n31917 ;
  assign y10250 = n31921 ;
  assign y10251 = n31922 ;
  assign y10252 = ~1'b0 ;
  assign y10253 = ~1'b0 ;
  assign y10254 = n31924 ;
  assign y10255 = n31935 ;
  assign y10256 = n31938 ;
  assign y10257 = ~n31941 ;
  assign y10258 = ~n31944 ;
  assign y10259 = n31950 ;
  assign y10260 = n31952 ;
  assign y10261 = n31953 ;
  assign y10262 = ~n31963 ;
  assign y10263 = ~1'b0 ;
  assign y10264 = ~n31966 ;
  assign y10265 = n31968 ;
  assign y10266 = ~n31970 ;
  assign y10267 = ~n31973 ;
  assign y10268 = ~n31975 ;
  assign y10269 = ~n31977 ;
  assign y10270 = ~n31982 ;
  assign y10271 = ~n31987 ;
  assign y10272 = ~n31989 ;
  assign y10273 = n31992 ;
  assign y10274 = ~1'b0 ;
  assign y10275 = ~n31993 ;
  assign y10276 = ~n10402 ;
  assign y10277 = ~n31995 ;
  assign y10278 = ~n31999 ;
  assign y10279 = n32001 ;
  assign y10280 = ~n32006 ;
  assign y10281 = n32007 ;
  assign y10282 = n32008 ;
  assign y10283 = ~n32015 ;
  assign y10284 = n32021 ;
  assign y10285 = ~n32023 ;
  assign y10286 = ~1'b0 ;
  assign y10287 = ~n32024 ;
  assign y10288 = n32025 ;
  assign y10289 = n24756 ;
  assign y10290 = n32027 ;
  assign y10291 = n32028 ;
  assign y10292 = ~n32031 ;
  assign y10293 = ~n32032 ;
  assign y10294 = ~n32035 ;
  assign y10295 = n32037 ;
  assign y10296 = ~n32039 ;
  assign y10297 = ~n32041 ;
  assign y10298 = ~n32042 ;
  assign y10299 = ~n32044 ;
  assign y10300 = ~n32048 ;
  assign y10301 = ~n32049 ;
  assign y10302 = n32052 ;
  assign y10303 = n32057 ;
  assign y10304 = ~n32058 ;
  assign y10305 = ~1'b0 ;
  assign y10306 = ~n32060 ;
  assign y10307 = ~n32062 ;
  assign y10308 = ~1'b0 ;
  assign y10309 = ~n32065 ;
  assign y10310 = n32067 ;
  assign y10311 = n32068 ;
  assign y10312 = n32070 ;
  assign y10313 = ~n32075 ;
  assign y10314 = n32079 ;
  assign y10315 = n32081 ;
  assign y10316 = n32083 ;
  assign y10317 = ~n32084 ;
  assign y10318 = ~1'b0 ;
  assign y10319 = n32088 ;
endmodule
