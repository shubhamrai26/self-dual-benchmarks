module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 , y8929 , y8930 , y8931 , y8932 , y8933 , y8934 , y8935 , y8936 , y8937 , y8938 , y8939 , y8940 , y8941 , y8942 , y8943 , y8944 , y8945 , y8946 , y8947 , y8948 , y8949 , y8950 , y8951 , y8952 , y8953 , y8954 , y8955 , y8956 , y8957 , y8958 , y8959 , y8960 , y8961 , y8962 , y8963 , y8964 , y8965 , y8966 , y8967 , y8968 , y8969 , y8970 , y8971 , y8972 , y8973 , y8974 , y8975 , y8976 , y8977 , y8978 , y8979 , y8980 , y8981 , y8982 , y8983 , y8984 , y8985 , y8986 , y8987 , y8988 , y8989 , y8990 , y8991 , y8992 , y8993 , y8994 , y8995 , y8996 , y8997 , y8998 , y8999 , y9000 , y9001 , y9002 , y9003 , y9004 , y9005 , y9006 , y9007 , y9008 , y9009 , y9010 , y9011 , y9012 , y9013 , y9014 , y9015 , y9016 , y9017 , y9018 , y9019 , y9020 , y9021 , y9022 , y9023 , y9024 , y9025 , y9026 , y9027 , y9028 , y9029 , y9030 , y9031 , y9032 , y9033 , y9034 , y9035 , y9036 , y9037 , y9038 , y9039 , y9040 , y9041 , y9042 , y9043 , y9044 , y9045 , y9046 , y9047 , y9048 , y9049 , y9050 , y9051 , y9052 , y9053 , y9054 , y9055 , y9056 , y9057 , y9058 , y9059 , y9060 , y9061 , y9062 , y9063 , y9064 , y9065 , y9066 , y9067 , y9068 , y9069 , y9070 , y9071 , y9072 , y9073 , y9074 , y9075 , y9076 , y9077 , y9078 , y9079 , y9080 , y9081 , y9082 , y9083 , y9084 , y9085 , y9086 , y9087 , y9088 , y9089 , y9090 , y9091 , y9092 , y9093 , y9094 , y9095 , y9096 , y9097 , y9098 , y9099 , y9100 , y9101 , y9102 , y9103 , y9104 , y9105 , y9106 , y9107 , y9108 , y9109 , y9110 , y9111 , y9112 , y9113 , y9114 , y9115 , y9116 , y9117 , y9118 , y9119 , y9120 , y9121 , y9122 , y9123 , y9124 , y9125 , y9126 , y9127 , y9128 , y9129 , y9130 , y9131 , y9132 , y9133 , y9134 , y9135 , y9136 , y9137 , y9138 , y9139 , y9140 , y9141 , y9142 , y9143 , y9144 , y9145 , y9146 , y9147 , y9148 , y9149 , y9150 , y9151 , y9152 , y9153 , y9154 , y9155 , y9156 , y9157 , y9158 , y9159 , y9160 , y9161 , y9162 , y9163 , y9164 , y9165 , y9166 , y9167 , y9168 , y9169 , y9170 , y9171 , y9172 , y9173 , y9174 , y9175 , y9176 , y9177 , y9178 , y9179 , y9180 , y9181 , y9182 , y9183 , y9184 , y9185 , y9186 , y9187 , y9188 , y9189 , y9190 , y9191 , y9192 , y9193 , y9194 , y9195 , y9196 , y9197 , y9198 , y9199 , y9200 , y9201 , y9202 , y9203 , y9204 , y9205 , y9206 , y9207 , y9208 , y9209 , y9210 , y9211 , y9212 , y9213 , y9214 , y9215 , y9216 , y9217 , y9218 , y9219 , y9220 , y9221 , y9222 , y9223 , y9224 , y9225 , y9226 , y9227 , y9228 , y9229 , y9230 , y9231 , y9232 , y9233 , y9234 , y9235 , y9236 , y9237 , y9238 , y9239 , y9240 , y9241 , y9242 , y9243 , y9244 , y9245 , y9246 , y9247 , y9248 , y9249 , y9250 , y9251 , y9252 , y9253 , y9254 , y9255 , y9256 , y9257 , y9258 , y9259 , y9260 , y9261 , y9262 , y9263 , y9264 , y9265 , y9266 , y9267 , y9268 , y9269 , y9270 , y9271 , y9272 , y9273 , y9274 , y9275 , y9276 , y9277 , y9278 , y9279 , y9280 , y9281 , y9282 , y9283 , y9284 , y9285 , y9286 , y9287 , y9288 , y9289 , y9290 , y9291 , y9292 , y9293 , y9294 , y9295 , y9296 , y9297 , y9298 , y9299 , y9300 , y9301 , y9302 , y9303 , y9304 , y9305 , y9306 , y9307 , y9308 , y9309 , y9310 , y9311 , y9312 , y9313 , y9314 , y9315 , y9316 , y9317 , y9318 , y9319 , y9320 , y9321 , y9322 , y9323 , y9324 , y9325 , y9326 , y9327 , y9328 , y9329 , y9330 , y9331 , y9332 , y9333 , y9334 , y9335 , y9336 , y9337 , y9338 , y9339 , y9340 , y9341 , y9342 , y9343 , y9344 , y9345 , y9346 , y9347 , y9348 , y9349 , y9350 , y9351 , y9352 , y9353 , y9354 , y9355 , y9356 , y9357 , y9358 , y9359 , y9360 , y9361 , y9362 , y9363 , y9364 , y9365 , y9366 , y9367 , y9368 , y9369 , y9370 , y9371 , y9372 , y9373 , y9374 , y9375 , y9376 , y9377 , y9378 , y9379 , y9380 , y9381 , y9382 , y9383 , y9384 , y9385 , y9386 , y9387 , y9388 , y9389 , y9390 , y9391 , y9392 , y9393 , y9394 , y9395 , y9396 , y9397 , y9398 , y9399 , y9400 , y9401 , y9402 , y9403 , y9404 , y9405 , y9406 , y9407 , y9408 , y9409 , y9410 , y9411 , y9412 , y9413 , y9414 , y9415 , y9416 , y9417 , y9418 , y9419 , y9420 , y9421 , y9422 , y9423 , y9424 , y9425 , y9426 , y9427 , y9428 , y9429 , y9430 , y9431 , y9432 , y9433 , y9434 , y9435 , y9436 , y9437 , y9438 , y9439 , y9440 , y9441 , y9442 , y9443 , y9444 , y9445 , y9446 , y9447 , y9448 , y9449 , y9450 , y9451 , y9452 , y9453 , y9454 , y9455 , y9456 , y9457 , y9458 , y9459 , y9460 , y9461 , y9462 , y9463 , y9464 , y9465 , y9466 , y9467 , y9468 , y9469 , y9470 , y9471 , y9472 , y9473 , y9474 , y9475 , y9476 , y9477 , y9478 , y9479 , y9480 , y9481 , y9482 , y9483 , y9484 , y9485 , y9486 , y9487 , y9488 , y9489 , y9490 , y9491 , y9492 , y9493 , y9494 , y9495 , y9496 , y9497 , y9498 , y9499 , y9500 , y9501 , y9502 , y9503 , y9504 , y9505 , y9506 , y9507 , y9508 , y9509 , y9510 , y9511 , y9512 , y9513 , y9514 , y9515 , y9516 , y9517 , y9518 , y9519 , y9520 , y9521 , y9522 , y9523 , y9524 , y9525 , y9526 , y9527 , y9528 , y9529 , y9530 , y9531 , y9532 , y9533 , y9534 , y9535 , y9536 , y9537 , y9538 , y9539 , y9540 , y9541 , y9542 , y9543 , y9544 , y9545 , y9546 , y9547 , y9548 , y9549 , y9550 , y9551 , y9552 , y9553 , y9554 , y9555 , y9556 , y9557 , y9558 , y9559 , y9560 , y9561 , y9562 , y9563 , y9564 , y9565 , y9566 , y9567 , y9568 , y9569 , y9570 , y9571 , y9572 , y9573 , y9574 , y9575 , y9576 , y9577 , y9578 , y9579 , y9580 , y9581 , y9582 , y9583 , y9584 , y9585 , y9586 , y9587 , y9588 , y9589 , y9590 , y9591 , y9592 , y9593 , y9594 , y9595 , y9596 , y9597 , y9598 , y9599 , y9600 , y9601 , y9602 , y9603 , y9604 , y9605 , y9606 , y9607 , y9608 , y9609 , y9610 , y9611 , y9612 , y9613 , y9614 , y9615 , y9616 , y9617 , y9618 , y9619 , y9620 , y9621 , y9622 , y9623 , y9624 , y9625 , y9626 , y9627 , y9628 , y9629 , y9630 , y9631 , y9632 , y9633 , y9634 , y9635 , y9636 , y9637 , y9638 , y9639 , y9640 , y9641 , y9642 , y9643 , y9644 , y9645 , y9646 , y9647 , y9648 , y9649 , y9650 , y9651 , y9652 , y9653 , y9654 , y9655 , y9656 , y9657 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 ;
  assign n129 = ( ~x39 & x48 ) | ( ~x39 & x109 ) | ( x48 & x109 ) ;
  assign n130 = n129 ^ x124 ^ x43 ;
  assign n131 = n130 ^ x116 ^ x68 ;
  assign n132 = x71 & x75 ;
  assign n133 = n132 ^ x59 ^ 1'b0 ;
  assign n134 = x32 ^ x6 ^ 1'b0 ;
  assign n135 = ~n133 & n134 ;
  assign n136 = n135 ^ x4 ^ x0 ;
  assign n137 = x115 & x116 ;
  assign n138 = n137 ^ x123 ^ 1'b0 ;
  assign n139 = x52 ^ x14 ^ x7 ;
  assign n141 = ( x31 & x37 ) | ( x31 & ~x60 ) | ( x37 & ~x60 ) ;
  assign n142 = ( x14 & x108 ) | ( x14 & ~n141 ) | ( x108 & ~n141 ) ;
  assign n140 = ( x27 & x57 ) | ( x27 & ~x63 ) | ( x57 & ~x63 ) ;
  assign n143 = n142 ^ n140 ^ x110 ;
  assign n144 = x58 ^ x32 ^ 1'b0 ;
  assign n145 = x123 ^ x122 ^ 1'b0 ;
  assign n146 = x67 & ~n145 ;
  assign n147 = ( ~x75 & x76 ) | ( ~x75 & n146 ) | ( x76 & n146 ) ;
  assign n148 = ( ~x67 & x73 ) | ( ~x67 & x127 ) | ( x73 & x127 ) ;
  assign n149 = n148 ^ n131 ^ x125 ;
  assign n150 = ( x63 & x82 ) | ( x63 & n149 ) | ( x82 & n149 ) ;
  assign n151 = x100 & x114 ;
  assign n152 = ~x15 & n151 ;
  assign n153 = ( x1 & x115 ) | ( x1 & ~n141 ) | ( x115 & ~n141 ) ;
  assign n154 = x111 ^ x71 ^ x47 ;
  assign n155 = n154 ^ x109 ^ x49 ;
  assign n156 = x73 & x114 ;
  assign n157 = ~n155 & n156 ;
  assign n158 = x117 ^ x40 ^ x10 ;
  assign n159 = ( ~x70 & x120 ) | ( ~x70 & n158 ) | ( x120 & n158 ) ;
  assign n160 = ( x4 & ~x52 ) | ( x4 & n159 ) | ( ~x52 & n159 ) ;
  assign n161 = ( x10 & ~x112 ) | ( x10 & n160 ) | ( ~x112 & n160 ) ;
  assign n162 = ( x96 & n157 ) | ( x96 & n161 ) | ( n157 & n161 ) ;
  assign n172 = ( x18 & x67 ) | ( x18 & ~x99 ) | ( x67 & ~x99 ) ;
  assign n173 = n172 ^ x123 ^ x47 ;
  assign n169 = x65 ^ x37 ^ 1'b0 ;
  assign n170 = x51 & n169 ;
  assign n171 = ( x13 & ~n129 ) | ( x13 & n170 ) | ( ~n129 & n170 ) ;
  assign n167 = ( x49 & x71 ) | ( x49 & ~x73 ) | ( x71 & ~x73 ) ;
  assign n163 = ( x49 & ~x78 ) | ( x49 & x117 ) | ( ~x78 & x117 ) ;
  assign n164 = ( ~x31 & x63 ) | ( ~x31 & n163 ) | ( x63 & n163 ) ;
  assign n165 = n164 ^ x107 ^ x88 ;
  assign n166 = ( x24 & ~x86 ) | ( x24 & n165 ) | ( ~x86 & n165 ) ;
  assign n168 = n167 ^ n166 ^ x21 ;
  assign n174 = n173 ^ n171 ^ n168 ;
  assign n175 = x89 ^ x84 ^ x0 ;
  assign n176 = n175 ^ n165 ^ x66 ;
  assign n177 = x28 & ~x33 ;
  assign n178 = ( n170 & n176 ) | ( n170 & n177 ) | ( n176 & n177 ) ;
  assign n179 = ( x25 & ~x55 ) | ( x25 & n166 ) | ( ~x55 & n166 ) ;
  assign n180 = ( ~x81 & n163 ) | ( ~x81 & n175 ) | ( n163 & n175 ) ;
  assign n181 = n180 ^ n154 ^ x127 ;
  assign n189 = ( ~x3 & x31 ) | ( ~x3 & x103 ) | ( x31 & x103 ) ;
  assign n182 = ( x73 & ~x94 ) | ( x73 & n159 ) | ( ~x94 & n159 ) ;
  assign n183 = ( ~x10 & x99 ) | ( ~x10 & x105 ) | ( x99 & x105 ) ;
  assign n184 = n183 ^ x32 ^ x24 ;
  assign n185 = ( x11 & ~n133 ) | ( x11 & n184 ) | ( ~n133 & n184 ) ;
  assign n186 = ( ~x47 & x115 ) | ( ~x47 & n185 ) | ( x115 & n185 ) ;
  assign n187 = n186 ^ x112 ^ x84 ;
  assign n188 = ( n168 & n182 ) | ( n168 & n187 ) | ( n182 & n187 ) ;
  assign n190 = n189 ^ n188 ^ 1'b0 ;
  assign n191 = n181 | n190 ;
  assign n192 = ( x39 & ~x46 ) | ( x39 & x108 ) | ( ~x46 & x108 ) ;
  assign n193 = ( ~x35 & x74 ) | ( ~x35 & n192 ) | ( x74 & n192 ) ;
  assign n194 = ( x40 & x84 ) | ( x40 & n154 ) | ( x84 & n154 ) ;
  assign n195 = n194 ^ n163 ^ x90 ;
  assign n196 = x124 ^ x115 ^ x19 ;
  assign n197 = ( ~n135 & n145 ) | ( ~n135 & n196 ) | ( n145 & n196 ) ;
  assign n198 = ( x17 & n184 ) | ( x17 & n197 ) | ( n184 & n197 ) ;
  assign n199 = ( n193 & n195 ) | ( n193 & n198 ) | ( n195 & n198 ) ;
  assign n200 = ( x23 & ~x94 ) | ( x23 & n173 ) | ( ~x94 & n173 ) ;
  assign n201 = n200 ^ x55 ^ x35 ;
  assign n202 = ( x100 & x111 ) | ( x100 & ~x115 ) | ( x111 & ~x115 ) ;
  assign n203 = x41 & ~n176 ;
  assign n204 = ~x102 & n203 ;
  assign n205 = n202 & n204 ;
  assign n217 = x93 & ~n165 ;
  assign n218 = n217 ^ n145 ^ 1'b0 ;
  assign n216 = x77 & ~x120 ;
  assign n214 = x91 ^ x30 ^ x24 ;
  assign n207 = x118 ^ x43 ^ x21 ;
  assign n208 = n133 | n207 ;
  assign n209 = x125 ^ x106 ^ x61 ;
  assign n210 = x73 & ~n209 ;
  assign n211 = n210 ^ x44 ^ 1'b0 ;
  assign n212 = n211 ^ n166 ^ x94 ;
  assign n213 = ( x50 & ~n208 ) | ( x50 & n212 ) | ( ~n208 & n212 ) ;
  assign n206 = x76 & n145 ;
  assign n215 = n214 ^ n213 ^ n206 ;
  assign n219 = n218 ^ n216 ^ n215 ;
  assign n220 = x33 ^ x24 ^ x20 ;
  assign n221 = x85 & ~n220 ;
  assign n222 = n221 ^ x122 ^ 1'b0 ;
  assign n225 = x71 & x115 ;
  assign n226 = n225 ^ x46 ^ 1'b0 ;
  assign n223 = x83 ^ x46 ^ x9 ;
  assign n224 = n223 ^ x106 ^ 1'b0 ;
  assign n227 = n226 ^ n224 ^ 1'b0 ;
  assign n228 = ~n222 & n227 ;
  assign n234 = ( x48 & ~x64 ) | ( x48 & n129 ) | ( ~x64 & n129 ) ;
  assign n231 = x79 ^ x7 ^ 1'b0 ;
  assign n229 = ( x91 & ~x114 ) | ( x91 & n158 ) | ( ~x114 & n158 ) ;
  assign n230 = x60 & ~n229 ;
  assign n232 = n231 ^ n230 ^ 1'b0 ;
  assign n233 = n232 ^ x76 ^ x69 ;
  assign n235 = n234 ^ n233 ^ x36 ;
  assign n236 = x120 ^ x109 ^ x66 ;
  assign n237 = ( ~x11 & x39 ) | ( ~x11 & x126 ) | ( x39 & x126 ) ;
  assign n238 = ( ~x40 & n236 ) | ( ~x40 & n237 ) | ( n236 & n237 ) ;
  assign n239 = n182 ^ x61 ^ x56 ;
  assign n240 = ( x30 & x100 ) | ( x30 & ~n239 ) | ( x100 & ~n239 ) ;
  assign n241 = n136 ^ x79 ^ 1'b0 ;
  assign n242 = n240 & ~n241 ;
  assign n243 = ( x119 & n180 ) | ( x119 & ~n231 ) | ( n180 & ~n231 ) ;
  assign n244 = x106 ^ x99 ^ x53 ;
  assign n245 = x119 ^ x21 ^ x5 ;
  assign n246 = ( x78 & ~x114 ) | ( x78 & n245 ) | ( ~x114 & n245 ) ;
  assign n247 = ( x81 & n244 ) | ( x81 & ~n246 ) | ( n244 & ~n246 ) ;
  assign n248 = ( ~n136 & n243 ) | ( ~n136 & n247 ) | ( n243 & n247 ) ;
  assign n252 = n145 ^ x36 ^ x14 ;
  assign n253 = n252 ^ x47 ^ x27 ;
  assign n249 = n154 ^ x114 ^ x34 ;
  assign n250 = ( n167 & n181 ) | ( n167 & n249 ) | ( n181 & n249 ) ;
  assign n251 = n250 ^ x17 ^ 1'b0 ;
  assign n254 = n253 ^ n251 ^ n201 ;
  assign n255 = n254 ^ x125 ^ x96 ;
  assign n256 = x77 & x110 ;
  assign n257 = ( n146 & ~n231 ) | ( n146 & n256 ) | ( ~n231 & n256 ) ;
  assign n258 = n257 ^ n184 ^ n164 ;
  assign n259 = x98 ^ x18 ^ 1'b0 ;
  assign n260 = ~n160 & n259 ;
  assign n261 = ( ~n154 & n258 ) | ( ~n154 & n260 ) | ( n258 & n260 ) ;
  assign n262 = x43 & ~n218 ;
  assign n263 = n262 ^ x109 ^ 1'b0 ;
  assign n264 = ( ~x19 & x37 ) | ( ~x19 & n136 ) | ( x37 & n136 ) ;
  assign n265 = ( x72 & ~x91 ) | ( x72 & n264 ) | ( ~x91 & n264 ) ;
  assign n266 = n263 | n265 ;
  assign n267 = x20 & x99 ;
  assign n268 = n267 ^ x76 ^ 1'b0 ;
  assign n269 = n237 ^ n129 ^ 1'b0 ;
  assign n270 = x45 & n269 ;
  assign n271 = x48 & n270 ;
  assign n272 = n271 ^ n146 ^ 1'b0 ;
  assign n273 = ( ~n171 & n220 ) | ( ~n171 & n272 ) | ( n220 & n272 ) ;
  assign n274 = n257 | n273 ;
  assign n275 = n268 & ~n274 ;
  assign n276 = ( x36 & ~x45 ) | ( x36 & x114 ) | ( ~x45 & x114 ) ;
  assign n277 = ( n139 & n189 ) | ( n139 & n276 ) | ( n189 & n276 ) ;
  assign n278 = ( ~n165 & n275 ) | ( ~n165 & n277 ) | ( n275 & n277 ) ;
  assign n279 = ( x36 & x39 ) | ( x36 & n157 ) | ( x39 & n157 ) ;
  assign n280 = ( ~x17 & x70 ) | ( ~x17 & n279 ) | ( x70 & n279 ) ;
  assign n281 = n155 ^ x57 ^ 1'b0 ;
  assign n282 = n281 ^ n248 ^ n158 ;
  assign n283 = ( ~x23 & x57 ) | ( ~x23 & x112 ) | ( x57 & x112 ) ;
  assign n284 = n283 ^ n265 ^ n130 ;
  assign n285 = ( x117 & n249 ) | ( x117 & n284 ) | ( n249 & n284 ) ;
  assign n286 = x84 & x122 ;
  assign n287 = n286 ^ n236 ^ 1'b0 ;
  assign n288 = n287 ^ n129 ^ 1'b0 ;
  assign n289 = n285 & n288 ;
  assign n290 = x83 ^ x78 ^ x64 ;
  assign n291 = n290 ^ x118 ^ 1'b0 ;
  assign n292 = n291 ^ x116 ^ x101 ;
  assign n293 = x109 & n180 ;
  assign n294 = ( x99 & n168 ) | ( x99 & ~n293 ) | ( n168 & ~n293 ) ;
  assign n301 = n141 ^ x63 ^ x21 ;
  assign n295 = n206 ^ n180 ^ x10 ;
  assign n296 = ( ~n147 & n268 ) | ( ~n147 & n295 ) | ( n268 & n295 ) ;
  assign n297 = x111 & ~n154 ;
  assign n298 = ~n256 & n297 ;
  assign n299 = n298 ^ n196 ^ n143 ;
  assign n300 = n296 & n299 ;
  assign n302 = n301 ^ n300 ^ 1'b0 ;
  assign n303 = n302 ^ n146 ^ 1'b0 ;
  assign n304 = x21 & ~n303 ;
  assign n305 = n182 ^ x126 ^ x93 ;
  assign n306 = ( x58 & ~n240 ) | ( x58 & n305 ) | ( ~n240 & n305 ) ;
  assign n311 = x87 ^ x21 ^ 1'b0 ;
  assign n312 = x95 & n311 ;
  assign n308 = n149 & ~n176 ;
  assign n307 = x86 & x124 ;
  assign n309 = n308 ^ n307 ^ 1'b0 ;
  assign n310 = ( ~x60 & x117 ) | ( ~x60 & n309 ) | ( x117 & n309 ) ;
  assign n313 = n312 ^ n310 ^ 1'b0 ;
  assign n314 = n306 & ~n313 ;
  assign n317 = n301 ^ n193 ^ x82 ;
  assign n318 = x66 & n317 ;
  assign n315 = ( x0 & ~x43 ) | ( x0 & n296 ) | ( ~x43 & n296 ) ;
  assign n316 = ~n232 & n315 ;
  assign n319 = n318 ^ n316 ^ 1'b0 ;
  assign n320 = n289 ^ n238 ^ n218 ;
  assign n321 = n290 ^ n261 ^ x76 ;
  assign n322 = n265 ^ n222 ^ 1'b0 ;
  assign n323 = x127 & n322 ;
  assign n324 = x79 & n323 ;
  assign n325 = ~n321 & n324 ;
  assign n327 = x121 ^ x72 ^ x31 ;
  assign n328 = x105 ^ x17 ^ 1'b0 ;
  assign n329 = x34 & n328 ;
  assign n330 = n329 ^ x35 ^ 1'b0 ;
  assign n331 = x39 & n330 ;
  assign n332 = ( ~x11 & n164 ) | ( ~x11 & n331 ) | ( n164 & n331 ) ;
  assign n333 = ( ~x16 & n327 ) | ( ~x16 & n332 ) | ( n327 & n332 ) ;
  assign n326 = ( x3 & x87 ) | ( x3 & n152 ) | ( x87 & n152 ) ;
  assign n334 = n333 ^ n326 ^ n162 ;
  assign n336 = n175 ^ x119 ^ x61 ;
  assign n335 = ( ~x58 & x109 ) | ( ~x58 & n171 ) | ( x109 & n171 ) ;
  assign n337 = n336 ^ n335 ^ x87 ;
  assign n338 = n209 ^ x91 ^ x20 ;
  assign n339 = n338 ^ n293 ^ n292 ;
  assign n340 = x125 ^ x122 ^ x20 ;
  assign n341 = ~n224 & n340 ;
  assign n342 = x103 ^ x58 ^ x48 ;
  assign n343 = ( ~n291 & n336 ) | ( ~n291 & n342 ) | ( n336 & n342 ) ;
  assign n344 = n343 ^ n166 ^ x81 ;
  assign n345 = n344 ^ n199 ^ n177 ;
  assign n346 = ( x2 & ~n341 ) | ( x2 & n345 ) | ( ~n341 & n345 ) ;
  assign n347 = n170 ^ x124 ^ x68 ;
  assign n348 = ( n200 & ~n213 ) | ( n200 & n296 ) | ( ~n213 & n296 ) ;
  assign n349 = n348 ^ x95 ^ x45 ;
  assign n350 = ( ~x3 & x115 ) | ( ~x3 & x117 ) | ( x115 & x117 ) ;
  assign n351 = ( n153 & n185 ) | ( n153 & ~n350 ) | ( n185 & ~n350 ) ;
  assign n352 = n243 ^ x17 ^ 1'b0 ;
  assign n353 = ( ~n240 & n351 ) | ( ~n240 & n352 ) | ( n351 & n352 ) ;
  assign n354 = ( n347 & n349 ) | ( n347 & n353 ) | ( n349 & n353 ) ;
  assign n365 = x23 & x127 ;
  assign n366 = n365 ^ x29 ^ 1'b0 ;
  assign n367 = n366 ^ n291 ^ n228 ;
  assign n361 = n149 ^ x95 ^ 1'b0 ;
  assign n362 = x108 & ~n361 ;
  assign n363 = ( n158 & ~n201 ) | ( n158 & n362 ) | ( ~n201 & n362 ) ;
  assign n359 = ( x49 & x81 ) | ( x49 & n207 ) | ( x81 & n207 ) ;
  assign n360 = ~x74 & n359 ;
  assign n355 = x73 ^ x19 ^ x7 ;
  assign n356 = n355 ^ n194 ^ n142 ;
  assign n357 = ( n165 & n234 ) | ( n165 & ~n356 ) | ( n234 & ~n356 ) ;
  assign n358 = ( n184 & n232 ) | ( n184 & ~n357 ) | ( n232 & ~n357 ) ;
  assign n364 = n363 ^ n360 ^ n358 ;
  assign n368 = n367 ^ n364 ^ x100 ;
  assign n373 = x58 ^ x14 ^ x4 ;
  assign n374 = n373 ^ n173 ^ x8 ;
  assign n371 = x8 & ~n139 ;
  assign n372 = n371 ^ n189 ^ 1'b0 ;
  assign n369 = n209 ^ x101 ^ x76 ;
  assign n370 = n369 ^ n358 ^ n246 ;
  assign n375 = n374 ^ n372 ^ n370 ;
  assign n382 = x110 ^ x83 ^ x8 ;
  assign n383 = n382 ^ x41 ^ x17 ;
  assign n384 = n383 ^ n329 ^ n327 ;
  assign n380 = n129 ^ x124 ^ x89 ;
  assign n376 = n243 ^ x120 ^ 1'b0 ;
  assign n377 = n376 ^ x91 ^ 1'b0 ;
  assign n378 = ~n180 & n377 ;
  assign n379 = ~x90 & n378 ;
  assign n381 = n380 ^ n379 ^ x79 ;
  assign n385 = n384 ^ n381 ^ 1'b0 ;
  assign n386 = ( n154 & n234 ) | ( n154 & ~n385 ) | ( n234 & ~n385 ) ;
  assign n393 = ( x73 & ~x101 ) | ( x73 & n265 ) | ( ~x101 & n265 ) ;
  assign n394 = ( x90 & n228 ) | ( x90 & n393 ) | ( n228 & n393 ) ;
  assign n391 = n133 ^ x50 ^ x18 ;
  assign n390 = ( x30 & x71 ) | ( x30 & ~x119 ) | ( x71 & ~x119 ) ;
  assign n387 = x114 ^ x79 ^ x29 ;
  assign n388 = n387 ^ n380 ^ x18 ;
  assign n389 = ( x71 & ~n248 ) | ( x71 & n388 ) | ( ~n248 & n388 ) ;
  assign n392 = n391 ^ n390 ^ n389 ;
  assign n395 = n394 ^ n392 ^ n144 ;
  assign n396 = ( x6 & ~x58 ) | ( x6 & n341 ) | ( ~x58 & n341 ) ;
  assign n397 = ( x112 & n325 ) | ( x112 & n396 ) | ( n325 & n396 ) ;
  assign n402 = n152 ^ x79 ^ x20 ;
  assign n403 = n402 ^ n276 ^ 1'b0 ;
  assign n404 = n349 & n403 ;
  assign n405 = n191 ^ x109 ^ 1'b0 ;
  assign n406 = n404 & ~n405 ;
  assign n400 = n130 ^ x82 ^ x1 ;
  assign n401 = n299 & ~n400 ;
  assign n398 = ( x87 & ~x119 ) | ( x87 & n283 ) | ( ~x119 & n283 ) ;
  assign n399 = n398 ^ n320 ^ n145 ;
  assign n407 = n406 ^ n401 ^ n399 ;
  assign n408 = ( x70 & ~x98 ) | ( x70 & n309 ) | ( ~x98 & n309 ) ;
  assign n409 = ( n294 & n397 ) | ( n294 & ~n408 ) | ( n397 & ~n408 ) ;
  assign n410 = n213 ^ x40 ^ 1'b0 ;
  assign n411 = x119 ^ x115 ^ x38 ;
  assign n412 = n411 ^ n180 ^ x17 ;
  assign n413 = ( n216 & ~n301 ) | ( n216 & n412 ) | ( ~n301 & n412 ) ;
  assign n414 = ( ~x52 & n168 ) | ( ~x52 & n413 ) | ( n168 & n413 ) ;
  assign n417 = x87 ^ x47 ^ x24 ;
  assign n415 = x58 & ~n207 ;
  assign n416 = n415 ^ x7 ^ 1'b0 ;
  assign n418 = n417 ^ n416 ^ x61 ;
  assign n420 = x7 & ~n185 ;
  assign n419 = ( x120 & n178 ) | ( x120 & ~n326 ) | ( n178 & ~n326 ) ;
  assign n421 = n420 ^ n419 ^ n384 ;
  assign n422 = n226 ^ x118 ^ x90 ;
  assign n423 = ( x82 & n299 ) | ( x82 & ~n422 ) | ( n299 & ~n422 ) ;
  assign n424 = ( x18 & n162 ) | ( x18 & n195 ) | ( n162 & n195 ) ;
  assign n425 = n424 ^ n250 ^ x95 ;
  assign n426 = ( ~x57 & n423 ) | ( ~x57 & n425 ) | ( n423 & n425 ) ;
  assign n427 = ( x58 & ~n188 ) | ( x58 & n236 ) | ( ~n188 & n236 ) ;
  assign n428 = n427 ^ x96 ^ 1'b0 ;
  assign n433 = n143 ^ x26 ^ 1'b0 ;
  assign n434 = n298 | n433 ;
  assign n429 = ( ~x29 & x43 ) | ( ~x29 & x50 ) | ( x43 & x50 ) ;
  assign n430 = n429 ^ n305 ^ x101 ;
  assign n431 = n430 ^ n187 ^ 1'b0 ;
  assign n432 = n293 & n431 ;
  assign n435 = n434 ^ n432 ^ 1'b0 ;
  assign n436 = ( x127 & n428 ) | ( x127 & n435 ) | ( n428 & n435 ) ;
  assign n437 = n436 ^ n424 ^ 1'b0 ;
  assign n438 = ( x35 & n187 ) | ( x35 & ~n220 ) | ( n187 & ~n220 ) ;
  assign n439 = n438 ^ n147 ^ 1'b0 ;
  assign n440 = ( n421 & n437 ) | ( n421 & ~n439 ) | ( n437 & ~n439 ) ;
  assign n441 = n362 ^ x78 ^ x28 ;
  assign n443 = x27 & x123 ;
  assign n444 = n443 ^ x41 ^ 1'b0 ;
  assign n442 = n377 ^ n369 ^ n352 ;
  assign n445 = n444 ^ n442 ^ n168 ;
  assign n446 = x0 & n445 ;
  assign n447 = n367 & n446 ;
  assign n448 = ( n228 & n441 ) | ( n228 & ~n447 ) | ( n441 & ~n447 ) ;
  assign n449 = x29 ^ x13 ^ x5 ;
  assign n450 = ( ~x42 & x73 ) | ( ~x42 & n141 ) | ( x73 & n141 ) ;
  assign n451 = n450 ^ n408 ^ n291 ;
  assign n452 = n451 ^ n213 ^ 1'b0 ;
  assign n453 = ( n150 & n161 ) | ( n150 & ~n257 ) | ( n161 & ~n257 ) ;
  assign n454 = n453 ^ n312 ^ n232 ;
  assign n455 = n454 ^ n240 ^ 1'b0 ;
  assign n456 = x120 & n455 ;
  assign n457 = ( ~n449 & n452 ) | ( ~n449 & n456 ) | ( n452 & n456 ) ;
  assign n458 = ( x104 & n194 ) | ( x104 & ~n457 ) | ( n194 & ~n457 ) ;
  assign n459 = ( ~n358 & n374 ) | ( ~n358 & n458 ) | ( n374 & n458 ) ;
  assign n460 = n277 & ~n417 ;
  assign n461 = ( x58 & n206 ) | ( x58 & ~n460 ) | ( n206 & ~n460 ) ;
  assign n462 = n461 ^ n383 ^ 1'b0 ;
  assign n463 = n462 ^ x15 ^ 1'b0 ;
  assign n464 = ~n246 & n463 ;
  assign n465 = n205 | n461 ;
  assign n466 = n253 ^ n178 ^ x111 ;
  assign n467 = x94 & n466 ;
  assign n468 = n447 & n467 ;
  assign n471 = x100 ^ x52 ^ x19 ;
  assign n472 = n471 ^ n200 ^ x109 ;
  assign n469 = n237 ^ x86 ^ x56 ;
  assign n470 = n469 ^ x48 ^ 1'b0 ;
  assign n473 = n472 ^ n470 ^ n375 ;
  assign n481 = x98 & ~n449 ;
  assign n482 = n481 ^ n331 ^ 1'b0 ;
  assign n480 = ( ~n223 & n265 ) | ( ~n223 & n273 ) | ( n265 & n273 ) ;
  assign n477 = n299 ^ n181 ^ 1'b0 ;
  assign n478 = n477 ^ n240 ^ n140 ;
  assign n479 = n478 ^ n292 ^ 1'b0 ;
  assign n483 = n482 ^ n480 ^ n479 ;
  assign n474 = n373 ^ n340 ^ n194 ;
  assign n475 = ( ~x15 & n228 ) | ( ~x15 & n362 ) | ( n228 & n362 ) ;
  assign n476 = ( ~n391 & n474 ) | ( ~n391 & n475 ) | ( n474 & n475 ) ;
  assign n484 = n483 ^ n476 ^ n139 ;
  assign n485 = x59 & x105 ;
  assign n486 = ~x12 & n485 ;
  assign n487 = n486 ^ n369 ^ n138 ;
  assign n488 = ( n473 & n484 ) | ( n473 & n487 ) | ( n484 & n487 ) ;
  assign n489 = n301 ^ n205 ^ n201 ;
  assign n490 = n340 ^ x99 ^ 1'b0 ;
  assign n491 = x63 & ~n490 ;
  assign n492 = ( n223 & n408 ) | ( n223 & n491 ) | ( n408 & n491 ) ;
  assign n493 = ( x52 & n489 ) | ( x52 & n492 ) | ( n489 & n492 ) ;
  assign n498 = x125 ^ x124 ^ x96 ;
  assign n494 = x10 & x17 ;
  assign n495 = ~x16 & n494 ;
  assign n496 = ( x16 & n452 ) | ( x16 & ~n495 ) | ( n452 & ~n495 ) ;
  assign n497 = ( ~n435 & n439 ) | ( ~n435 & n496 ) | ( n439 & n496 ) ;
  assign n499 = n498 ^ n497 ^ n179 ;
  assign n500 = ( ~n264 & n493 ) | ( ~n264 & n499 ) | ( n493 & n499 ) ;
  assign n501 = ( n279 & ~n391 ) | ( n279 & n439 ) | ( ~n391 & n439 ) ;
  assign n502 = n209 ^ x119 ^ x94 ;
  assign n503 = ( x94 & ~n356 ) | ( x94 & n502 ) | ( ~n356 & n502 ) ;
  assign n504 = ~n178 & n503 ;
  assign n505 = n504 ^ n402 ^ 1'b0 ;
  assign n506 = n229 ^ n138 ^ 1'b0 ;
  assign n507 = ( x86 & n417 ) | ( x86 & ~n506 ) | ( n417 & ~n506 ) ;
  assign n508 = n507 ^ n238 ^ x91 ;
  assign n509 = n223 ^ x55 ^ x5 ;
  assign n510 = ( x62 & ~x78 ) | ( x62 & n509 ) | ( ~x78 & n509 ) ;
  assign n512 = x39 & ~n181 ;
  assign n511 = ( x78 & x104 ) | ( x78 & ~n194 ) | ( x104 & ~n194 ) ;
  assign n513 = n512 ^ n511 ^ n345 ;
  assign n514 = ( n195 & n510 ) | ( n195 & ~n513 ) | ( n510 & ~n513 ) ;
  assign n515 = ( x51 & n181 ) | ( x51 & n514 ) | ( n181 & n514 ) ;
  assign n516 = ( x26 & n424 ) | ( x26 & ~n477 ) | ( n424 & ~n477 ) ;
  assign n518 = n183 ^ x31 ^ 1'b0 ;
  assign n519 = n140 & n518 ;
  assign n517 = n359 ^ n202 ^ x54 ;
  assign n520 = n519 ^ n517 ^ x18 ;
  assign n521 = ( n202 & ~n516 ) | ( n202 & n520 ) | ( ~n516 & n520 ) ;
  assign n542 = x124 & ~n298 ;
  assign n543 = n542 ^ x41 ^ 1'b0 ;
  assign n544 = n270 & n391 ;
  assign n545 = n543 & n544 ;
  assign n546 = ( x77 & n199 ) | ( x77 & ~n545 ) | ( n199 & ~n545 ) ;
  assign n547 = n546 ^ n254 ^ n160 ;
  assign n537 = n291 ^ n253 ^ 1'b0 ;
  assign n538 = n220 | n537 ;
  assign n534 = ( ~n161 & n228 ) | ( ~n161 & n379 ) | ( n228 & n379 ) ;
  assign n535 = ( x97 & n283 ) | ( x97 & ~n534 ) | ( n283 & ~n534 ) ;
  assign n536 = n535 ^ x61 ^ x21 ;
  assign n531 = n164 & n331 ;
  assign n532 = n531 ^ x35 ^ 1'b0 ;
  assign n533 = n532 ^ n260 ^ n246 ;
  assign n539 = n538 ^ n536 ^ n533 ;
  assign n540 = n129 & n539 ;
  assign n541 = ~x104 & n540 ;
  assign n529 = n391 ^ n325 ^ x41 ;
  assign n524 = ( x42 & ~x64 ) | ( x42 & x96 ) | ( ~x64 & x96 ) ;
  assign n522 = x9 & x98 ;
  assign n523 = n522 ^ x111 ^ 1'b0 ;
  assign n525 = n524 ^ n523 ^ x15 ;
  assign n526 = ( ~x57 & n408 ) | ( ~x57 & n525 ) | ( n408 & n525 ) ;
  assign n527 = n167 ^ x103 ^ 1'b0 ;
  assign n528 = ( n495 & ~n526 ) | ( n495 & n527 ) | ( ~n526 & n527 ) ;
  assign n530 = n529 ^ n528 ^ n420 ;
  assign n548 = n547 ^ n541 ^ n530 ;
  assign n549 = ( n158 & ~n521 ) | ( n158 & n548 ) | ( ~n521 & n548 ) ;
  assign n561 = n404 ^ n231 ^ n196 ;
  assign n552 = ~n180 & n329 ;
  assign n553 = n552 ^ x96 ^ 1'b0 ;
  assign n550 = x99 ^ x48 ^ x40 ;
  assign n551 = n550 ^ n253 ^ n214 ;
  assign n554 = n553 ^ n551 ^ x121 ;
  assign n555 = ~n180 & n317 ;
  assign n556 = n554 & n555 ;
  assign n557 = n523 ^ n253 ^ x12 ;
  assign n558 = n557 ^ n349 ^ n133 ;
  assign n559 = n558 ^ n460 ^ n131 ;
  assign n560 = ( n459 & n556 ) | ( n459 & ~n559 ) | ( n556 & ~n559 ) ;
  assign n562 = n561 ^ n560 ^ x101 ;
  assign n563 = ( n181 & n273 ) | ( n181 & ~n301 ) | ( n273 & ~n301 ) ;
  assign n564 = n563 ^ n558 ^ n363 ;
  assign n565 = ( x108 & ~n344 ) | ( x108 & n564 ) | ( ~n344 & n564 ) ;
  assign n567 = n402 ^ n201 ^ 1'b0 ;
  assign n566 = n232 ^ n155 ^ 1'b0 ;
  assign n568 = n567 ^ n566 ^ n483 ;
  assign n569 = n346 ^ n309 ^ 1'b0 ;
  assign n570 = ( ~x113 & n475 ) | ( ~x113 & n569 ) | ( n475 & n569 ) ;
  assign n571 = ~n568 & n570 ;
  assign n572 = n565 & n571 ;
  assign n578 = n393 ^ n258 ^ n152 ;
  assign n573 = ( x35 & n155 ) | ( x35 & n373 ) | ( n155 & n373 ) ;
  assign n574 = n573 ^ x59 ^ x25 ;
  assign n575 = ( x110 & ~n495 ) | ( x110 & n574 ) | ( ~n495 & n574 ) ;
  assign n576 = n279 ^ n172 ^ x22 ;
  assign n577 = ( ~n388 & n575 ) | ( ~n388 & n576 ) | ( n575 & n576 ) ;
  assign n579 = n578 ^ n577 ^ n359 ;
  assign n580 = n343 ^ n301 ^ n212 ;
  assign n581 = ~x30 & x55 ;
  assign n582 = n581 ^ n139 ^ 1'b0 ;
  assign n583 = n159 ^ x125 ^ x79 ;
  assign n584 = n215 ^ n195 ^ x18 ;
  assign n585 = n583 & ~n584 ;
  assign n586 = n429 ^ n213 ^ n168 ;
  assign n587 = n586 ^ n367 ^ 1'b0 ;
  assign n588 = ~n585 & n587 ;
  assign n589 = ( x72 & n582 ) | ( x72 & ~n588 ) | ( n582 & ~n588 ) ;
  assign n591 = ( n166 & ~n240 ) | ( n166 & n296 ) | ( ~n240 & n296 ) ;
  assign n592 = ( x68 & n175 ) | ( x68 & n253 ) | ( n175 & n253 ) ;
  assign n593 = ( ~x96 & n298 ) | ( ~x96 & n592 ) | ( n298 & n592 ) ;
  assign n594 = n591 | n593 ;
  assign n595 = n486 & ~n594 ;
  assign n590 = ~x58 & n242 ;
  assign n596 = n595 ^ n590 ^ n348 ;
  assign n597 = n596 ^ n292 ^ x120 ;
  assign n598 = ( n580 & n589 ) | ( n580 & n597 ) | ( n589 & n597 ) ;
  assign n599 = n536 ^ n454 ^ x95 ;
  assign n600 = n344 ^ x115 ^ 1'b0 ;
  assign n601 = ~n177 & n600 ;
  assign n602 = n129 & n261 ;
  assign n603 = ~n240 & n602 ;
  assign n604 = n601 & ~n603 ;
  assign n605 = ~x97 & n604 ;
  assign n610 = n340 ^ n214 ^ x35 ;
  assign n611 = ( ~n231 & n506 ) | ( ~n231 & n610 ) | ( n506 & n610 ) ;
  assign n606 = n175 | n420 ;
  assign n607 = n382 & ~n606 ;
  assign n608 = x60 & ~n252 ;
  assign n609 = n607 & n608 ;
  assign n612 = n611 ^ n609 ^ n291 ;
  assign n614 = x58 & n434 ;
  assign n613 = ~x127 & n399 ;
  assign n615 = n614 ^ n613 ^ 1'b0 ;
  assign n616 = n183 & n615 ;
  assign n617 = n612 & n616 ;
  assign n618 = n617 ^ n583 ^ 1'b0 ;
  assign n635 = ( n167 & ~n402 ) | ( n167 & n507 ) | ( ~n402 & n507 ) ;
  assign n630 = n277 ^ n270 ^ 1'b0 ;
  assign n631 = n256 & n630 ;
  assign n632 = ~n309 & n631 ;
  assign n633 = ~n349 & n632 ;
  assign n628 = n236 ^ n196 ^ x113 ;
  assign n625 = x17 & n167 ;
  assign n626 = n625 ^ x79 ^ 1'b0 ;
  assign n627 = n626 ^ n380 ^ n250 ;
  assign n622 = x88 & n186 ;
  assign n623 = ~n185 & n622 ;
  assign n624 = ( ~n160 & n372 ) | ( ~n160 & n623 ) | ( n372 & n623 ) ;
  assign n629 = n628 ^ n627 ^ n624 ;
  assign n619 = ( x22 & x86 ) | ( x22 & ~n292 ) | ( x86 & ~n292 ) ;
  assign n620 = n460 ^ n425 ^ n232 ;
  assign n621 = ( n439 & ~n619 ) | ( n439 & n620 ) | ( ~n619 & n620 ) ;
  assign n634 = n633 ^ n629 ^ n621 ;
  assign n636 = n635 ^ n634 ^ x55 ;
  assign n637 = n301 ^ n185 ^ x112 ;
  assign n638 = ( x7 & n167 ) | ( x7 & ~n637 ) | ( n167 & ~n637 ) ;
  assign n639 = n638 ^ n377 ^ n216 ;
  assign n640 = ( n153 & ~n281 ) | ( n153 & n382 ) | ( ~n281 & n382 ) ;
  assign n641 = n640 ^ n329 ^ x26 ;
  assign n642 = n641 ^ n534 ^ n276 ;
  assign n643 = ( ~n347 & n639 ) | ( ~n347 & n642 ) | ( n639 & n642 ) ;
  assign n644 = n323 | n623 ;
  assign n645 = ( x11 & x22 ) | ( x11 & ~n249 ) | ( x22 & ~n249 ) ;
  assign n646 = ( n258 & n644 ) | ( n258 & ~n645 ) | ( n644 & ~n645 ) ;
  assign n647 = n573 ^ n336 ^ x109 ;
  assign n657 = n249 | n563 ;
  assign n654 = n543 ^ x67 ^ 1'b0 ;
  assign n653 = ( x115 & ~n350 ) | ( x115 & n573 ) | ( ~n350 & n573 ) ;
  assign n655 = n654 ^ n653 ^ n291 ;
  assign n648 = ( x1 & x84 ) | ( x1 & ~n491 ) | ( x84 & ~n491 ) ;
  assign n649 = ( x43 & x55 ) | ( x43 & ~n648 ) | ( x55 & ~n648 ) ;
  assign n650 = n525 & n649 ;
  assign n651 = n650 ^ n399 ^ 1'b0 ;
  assign n652 = n651 ^ x48 ^ 1'b0 ;
  assign n656 = n655 ^ n652 ^ n648 ;
  assign n658 = n657 ^ n656 ^ n547 ;
  assign n659 = ( x76 & n647 ) | ( x76 & ~n658 ) | ( n647 & ~n658 ) ;
  assign n660 = x52 & n323 ;
  assign n661 = n660 ^ x72 ^ 1'b0 ;
  assign n662 = n661 ^ x83 ^ x31 ;
  assign n663 = n314 ^ n244 ^ 1'b0 ;
  assign n664 = n629 & ~n663 ;
  assign n665 = n224 & n664 ;
  assign n675 = n543 ^ n374 ^ n295 ;
  assign n676 = ( ~n309 & n393 ) | ( ~n309 & n675 ) | ( n393 & n675 ) ;
  assign n677 = n676 ^ x15 ^ x1 ;
  assign n667 = n146 ^ x65 ^ x7 ;
  assign n668 = ( x33 & x103 ) | ( x33 & ~x112 ) | ( x103 & ~x112 ) ;
  assign n669 = n668 ^ n191 ^ x87 ;
  assign n670 = ~n543 & n669 ;
  assign n671 = ( x101 & n667 ) | ( x101 & ~n670 ) | ( n667 & ~n670 ) ;
  assign n666 = x14 & ~n162 ;
  assign n672 = n671 ^ n666 ^ 1'b0 ;
  assign n673 = ( x58 & n382 ) | ( x58 & ~n672 ) | ( n382 & ~n672 ) ;
  assign n674 = n673 ^ n345 ^ n247 ;
  assign n678 = n677 ^ n674 ^ n309 ;
  assign n679 = n206 ^ n140 ^ 1'b0 ;
  assign n680 = n670 & n679 ;
  assign n681 = ( n545 & n662 ) | ( n545 & ~n680 ) | ( n662 & ~n680 ) ;
  assign n682 = x41 & x88 ;
  assign n683 = n682 ^ x75 ^ 1'b0 ;
  assign n684 = n279 & ~n683 ;
  assign n685 = n684 ^ x58 ^ 1'b0 ;
  assign n686 = n685 ^ n363 ^ x32 ;
  assign n687 = n436 | n686 ;
  assign n688 = n348 & ~n687 ;
  assign n689 = ( x30 & n503 ) | ( x30 & n688 ) | ( n503 & n688 ) ;
  assign n690 = n601 & n689 ;
  assign n691 = n690 ^ n520 ^ 1'b0 ;
  assign n692 = ( x4 & n166 ) | ( x4 & ~n691 ) | ( n166 & ~n691 ) ;
  assign n693 = n628 ^ n543 ^ n257 ;
  assign n694 = n301 | n693 ;
  assign n695 = n175 ^ x62 ^ x50 ;
  assign n703 = x48 & n400 ;
  assign n704 = ~x113 & n703 ;
  assign n705 = ( x101 & ~n139 ) | ( x101 & n704 ) | ( ~n139 & n704 ) ;
  assign n706 = n705 ^ n278 ^ x95 ;
  assign n699 = ( n197 & n213 ) | ( n197 & ~n422 ) | ( n213 & ~n422 ) ;
  assign n700 = n581 | n699 ;
  assign n701 = n700 ^ x98 ^ 1'b0 ;
  assign n702 = ( n264 & ~n465 ) | ( n264 & n701 ) | ( ~n465 & n701 ) ;
  assign n707 = n706 ^ n702 ^ n473 ;
  assign n696 = x107 ^ x10 ^ 1'b0 ;
  assign n697 = n317 & n352 ;
  assign n698 = ( ~x63 & n696 ) | ( ~x63 & n697 ) | ( n696 & n697 ) ;
  assign n708 = n707 ^ n698 ^ n406 ;
  assign n709 = ( ~x68 & n206 ) | ( ~x68 & n427 ) | ( n206 & n427 ) ;
  assign n710 = ( n214 & n428 ) | ( n214 & n709 ) | ( n428 & n709 ) ;
  assign n711 = n710 ^ n143 ^ x35 ;
  assign n712 = ( x21 & x108 ) | ( x21 & n543 ) | ( x108 & n543 ) ;
  assign n713 = n669 ^ n273 ^ x98 ;
  assign n714 = n713 ^ n154 ^ 1'b0 ;
  assign n718 = n428 & n631 ;
  assign n715 = n183 ^ x64 ^ 1'b0 ;
  assign n716 = ~n218 & n715 ;
  assign n717 = ( ~n200 & n444 ) | ( ~n200 & n716 ) | ( n444 & n716 ) ;
  assign n719 = n718 ^ n717 ^ x13 ;
  assign n720 = n524 ^ n305 ^ n223 ;
  assign n722 = x86 ^ x79 ^ x7 ;
  assign n723 = ( n306 & ~n491 ) | ( n306 & n722 ) | ( ~n491 & n722 ) ;
  assign n724 = ( n153 & ~n704 ) | ( n153 & n723 ) | ( ~n704 & n723 ) ;
  assign n721 = ( n136 & n219 ) | ( n136 & ~n517 ) | ( n219 & ~n517 ) ;
  assign n725 = n724 ^ n721 ^ 1'b0 ;
  assign n733 = ( x46 & n309 ) | ( x46 & ~n438 ) | ( n309 & ~n438 ) ;
  assign n731 = x5 & x101 ;
  assign n732 = ( x37 & x125 ) | ( x37 & ~n731 ) | ( x125 & ~n731 ) ;
  assign n734 = n733 ^ n732 ^ x88 ;
  assign n726 = n233 & n317 ;
  assign n727 = n498 & n726 ;
  assign n728 = n727 ^ n669 ^ x13 ;
  assign n729 = ( x80 & n320 ) | ( x80 & n627 ) | ( n320 & n627 ) ;
  assign n730 = ( n569 & ~n728 ) | ( n569 & n729 ) | ( ~n728 & n729 ) ;
  assign n735 = n734 ^ n730 ^ n301 ;
  assign n736 = ( x41 & ~n173 ) | ( x41 & n735 ) | ( ~n173 & n735 ) ;
  assign n737 = ( ~n720 & n725 ) | ( ~n720 & n736 ) | ( n725 & n736 ) ;
  assign n745 = x75 & ~x109 ;
  assign n738 = ( x17 & ~x99 ) | ( x17 & n327 ) | ( ~x99 & n327 ) ;
  assign n739 = n738 ^ n495 ^ n477 ;
  assign n740 = ( ~x33 & x61 ) | ( ~x33 & x100 ) | ( x61 & x100 ) ;
  assign n741 = n637 & n740 ;
  assign n742 = ~x25 & n741 ;
  assign n743 = ( n360 & n438 ) | ( n360 & ~n742 ) | ( n438 & ~n742 ) ;
  assign n744 = n739 & n743 ;
  assign n746 = n745 ^ n744 ^ 1'b0 ;
  assign n747 = n224 | n359 ;
  assign n748 = ( x45 & n251 ) | ( x45 & n747 ) | ( n251 & n747 ) ;
  assign n749 = n748 ^ n590 ^ n557 ;
  assign n751 = n510 ^ n253 ^ x117 ;
  assign n750 = n295 ^ n294 ^ 1'b0 ;
  assign n752 = n751 ^ n750 ^ n525 ;
  assign n753 = ( n746 & n749 ) | ( n746 & ~n752 ) | ( n749 & ~n752 ) ;
  assign n754 = n579 ^ n437 ^ 1'b0 ;
  assign n755 = n754 ^ n220 ^ 1'b0 ;
  assign n756 = n448 & n755 ;
  assign n757 = n325 ^ n263 ^ 1'b0 ;
  assign n758 = n457 & n757 ;
  assign n759 = n758 ^ n667 ^ n423 ;
  assign n760 = n759 ^ n758 ^ x100 ;
  assign n761 = ( n314 & n693 ) | ( n314 & ~n760 ) | ( n693 & ~n760 ) ;
  assign n762 = ( ~x67 & n140 ) | ( ~x67 & n242 ) | ( n140 & n242 ) ;
  assign n763 = x28 & n762 ;
  assign n764 = ( ~x53 & n529 ) | ( ~x53 & n763 ) | ( n529 & n763 ) ;
  assign n765 = n764 ^ n342 ^ x80 ;
  assign n769 = ~x55 & x58 ;
  assign n767 = ( x60 & ~n201 ) | ( x60 & n480 ) | ( ~n201 & n480 ) ;
  assign n768 = ( ~n188 & n410 ) | ( ~n188 & n767 ) | ( n410 & n767 ) ;
  assign n766 = n642 ^ n181 ^ 1'b0 ;
  assign n770 = n769 ^ n768 ^ n766 ;
  assign n772 = n595 ^ n376 ^ n236 ;
  assign n771 = n489 ^ n411 ^ n148 ;
  assign n773 = n772 ^ n771 ^ 1'b0 ;
  assign n774 = ( n235 & n429 ) | ( n235 & ~n441 ) | ( n429 & ~n441 ) ;
  assign n775 = n774 ^ n740 ^ x7 ;
  assign n776 = ( n209 & ~n393 ) | ( n209 & n649 ) | ( ~n393 & n649 ) ;
  assign n777 = n776 ^ n305 ^ 1'b0 ;
  assign n778 = n777 ^ n654 ^ 1'b0 ;
  assign n779 = n517 ^ n223 ^ 1'b0 ;
  assign n780 = ~n532 & n779 ;
  assign n781 = n491 ^ n424 ^ 1'b0 ;
  assign n785 = n469 ^ x33 ^ 1'b0 ;
  assign n786 = n219 | n785 ;
  assign n782 = ( x38 & ~x78 ) | ( x38 & n149 ) | ( ~x78 & n149 ) ;
  assign n783 = n782 ^ n780 ^ x50 ;
  assign n784 = ( x82 & ~n749 ) | ( x82 & n783 ) | ( ~n749 & n783 ) ;
  assign n787 = n786 ^ n784 ^ n497 ;
  assign n788 = ( n780 & n781 ) | ( n780 & ~n787 ) | ( n781 & ~n787 ) ;
  assign n790 = n573 ^ x120 ^ x110 ;
  assign n789 = n366 | n545 ;
  assign n791 = n790 ^ n789 ^ 1'b0 ;
  assign n792 = x72 & ~n769 ;
  assign n793 = ~x78 & n792 ;
  assign n794 = ( ~n276 & n502 ) | ( ~n276 & n533 ) | ( n502 & n533 ) ;
  assign n795 = n794 ^ n380 ^ 1'b0 ;
  assign n796 = ( n505 & n793 ) | ( n505 & n795 ) | ( n793 & n795 ) ;
  assign n797 = ( x66 & ~n791 ) | ( x66 & n796 ) | ( ~n791 & n796 ) ;
  assign n798 = n565 ^ n373 ^ x83 ;
  assign n799 = n798 ^ n232 ^ x82 ;
  assign n800 = n799 ^ x73 ^ x27 ;
  assign n801 = n698 ^ n669 ^ n497 ;
  assign n802 = n369 & n516 ;
  assign n803 = n802 ^ n651 ^ 1'b0 ;
  assign n804 = n803 ^ n620 ^ 1'b0 ;
  assign n805 = ( x52 & n449 ) | ( x52 & n627 ) | ( n449 & n627 ) ;
  assign n806 = n251 ^ x83 ^ x14 ;
  assign n807 = n776 ^ x95 ^ 1'b0 ;
  assign n808 = x101 & n807 ;
  assign n809 = n808 ^ n491 ^ 1'b0 ;
  assign n810 = n809 ^ n727 ^ x126 ;
  assign n815 = n429 ^ n355 ^ x29 ;
  assign n811 = ( x80 & ~n383 ) | ( x80 & n408 ) | ( ~n383 & n408 ) ;
  assign n812 = n281 & ~n417 ;
  assign n813 = n812 ^ x105 ^ 1'b0 ;
  assign n814 = ( n133 & ~n811 ) | ( n133 & n813 ) | ( ~n811 & n813 ) ;
  assign n816 = n815 ^ n814 ^ n649 ;
  assign n817 = ( n360 & ~n613 ) | ( n360 & n816 ) | ( ~n613 & n816 ) ;
  assign n832 = n495 ^ n425 ^ n285 ;
  assign n830 = ~x62 & n312 ;
  assign n829 = ( x34 & x93 ) | ( x34 & n434 ) | ( x93 & n434 ) ;
  assign n818 = ( x126 & ~x127 ) | ( x126 & n285 ) | ( ~x127 & n285 ) ;
  assign n819 = n818 ^ n642 ^ n323 ;
  assign n820 = ( x47 & n411 ) | ( x47 & ~n451 ) | ( n411 & ~n451 ) ;
  assign n821 = x37 & n820 ;
  assign n822 = n821 ^ n174 ^ 1'b0 ;
  assign n825 = ( x12 & ~x61 ) | ( x12 & n268 ) | ( ~x61 & n268 ) ;
  assign n823 = n777 ^ n243 ^ 1'b0 ;
  assign n824 = x44 & ~n823 ;
  assign n826 = n825 ^ n824 ^ 1'b0 ;
  assign n827 = ( x54 & n822 ) | ( x54 & n826 ) | ( n822 & n826 ) ;
  assign n828 = n819 & ~n827 ;
  assign n831 = n830 ^ n829 ^ n828 ;
  assign n833 = n832 ^ n831 ^ x74 ;
  assign n834 = ( x71 & n523 ) | ( x71 & n667 ) | ( n523 & n667 ) ;
  assign n835 = n834 ^ n541 ^ n393 ;
  assign n836 = n318 & n731 ;
  assign n837 = n836 ^ n638 ^ 1'b0 ;
  assign n838 = ( n596 & n598 ) | ( n596 & n837 ) | ( n598 & n837 ) ;
  assign n839 = n642 | n838 ;
  assign n840 = n648 | n839 ;
  assign n841 = n776 ^ n577 ^ n356 ;
  assign n842 = n841 ^ n317 ^ n196 ;
  assign n843 = ~n232 & n740 ;
  assign n844 = n843 ^ n412 ^ 1'b0 ;
  assign n845 = n409 & n844 ;
  assign n846 = n212 & n845 ;
  assign n848 = x73 & n362 ;
  assign n849 = n848 ^ x2 ^ 1'b0 ;
  assign n850 = ( ~x25 & n488 ) | ( ~x25 & n728 ) | ( n488 & n728 ) ;
  assign n851 = ( n637 & ~n849 ) | ( n637 & n850 ) | ( ~n849 & n850 ) ;
  assign n847 = n336 & ~n389 ;
  assign n852 = n851 ^ n847 ^ 1'b0 ;
  assign n853 = n852 ^ n610 ^ 1'b0 ;
  assign n854 = ~n846 & n853 ;
  assign n855 = ( x111 & n354 ) | ( x111 & n591 ) | ( n354 & n591 ) ;
  assign n856 = n849 ^ n786 ^ n216 ;
  assign n857 = ( n187 & ~n855 ) | ( n187 & n856 ) | ( ~n855 & n856 ) ;
  assign n860 = n404 ^ n278 ^ n256 ;
  assign n861 = n780 & n860 ;
  assign n858 = ( x27 & n257 ) | ( x27 & n546 ) | ( n257 & n546 ) ;
  assign n859 = ( x71 & ~n783 ) | ( x71 & n858 ) | ( ~n783 & n858 ) ;
  assign n862 = n861 ^ n859 ^ n530 ;
  assign n863 = n676 ^ n430 ^ 1'b0 ;
  assign n864 = ( x76 & n290 ) | ( x76 & n787 ) | ( n290 & n787 ) ;
  assign n865 = n596 ^ n472 ^ x96 ;
  assign n866 = n865 ^ n176 ^ 1'b0 ;
  assign n867 = x38 & ~n866 ;
  assign n868 = n867 ^ n428 ^ n184 ;
  assign n869 = ( x73 & ~n161 ) | ( x73 & n341 ) | ( ~n161 & n341 ) ;
  assign n870 = n425 ^ n235 ^ 1'b0 ;
  assign n871 = n218 | n870 ;
  assign n872 = ( n643 & ~n869 ) | ( n643 & n871 ) | ( ~n869 & n871 ) ;
  assign n874 = n237 & ~n722 ;
  assign n875 = n874 ^ x8 ^ 1'b0 ;
  assign n873 = x80 | n412 ;
  assign n876 = n875 ^ n873 ^ 1'b0 ;
  assign n877 = n506 ^ x85 ^ x4 ;
  assign n878 = n424 ^ x14 ^ 1'b0 ;
  assign n879 = ( n407 & n877 ) | ( n407 & n878 ) | ( n877 & n878 ) ;
  assign n880 = ( n432 & n475 ) | ( n432 & n723 ) | ( n475 & n723 ) ;
  assign n881 = n633 ^ n155 ^ x15 ;
  assign n882 = n192 & n551 ;
  assign n883 = ( n880 & ~n881 ) | ( n880 & n882 ) | ( ~n881 & n882 ) ;
  assign n885 = ( n148 & ~n383 ) | ( n148 & n558 ) | ( ~n383 & n558 ) ;
  assign n886 = n885 ^ n381 ^ 1'b0 ;
  assign n884 = n401 | n647 ;
  assign n887 = n886 ^ n884 ^ 1'b0 ;
  assign n889 = n623 ^ n212 ^ 1'b0 ;
  assign n888 = n668 ^ n634 ^ n306 ;
  assign n890 = n889 ^ n888 ^ n838 ;
  assign n891 = ( n362 & n738 ) | ( n362 & n890 ) | ( n738 & n890 ) ;
  assign n892 = n809 ^ n762 ^ n550 ;
  assign n893 = ( n411 & n488 ) | ( n411 & n892 ) | ( n488 & n892 ) ;
  assign n894 = ( ~x20 & x61 ) | ( ~x20 & x122 ) | ( x61 & x122 ) ;
  assign n895 = x96 ^ x3 ^ 1'b0 ;
  assign n896 = ~n162 & n895 ;
  assign n897 = n896 ^ n648 ^ 1'b0 ;
  assign n898 = n894 & n897 ;
  assign n899 = ( n250 & n855 ) | ( n250 & ~n898 ) | ( n855 & ~n898 ) ;
  assign n900 = ( ~n174 & n548 ) | ( ~n174 & n661 ) | ( n548 & n661 ) ;
  assign n901 = ( n294 & n899 ) | ( n294 & n900 ) | ( n899 & n900 ) ;
  assign n902 = n593 ^ n465 ^ x120 ;
  assign n903 = n902 ^ n811 ^ n189 ;
  assign n904 = n903 ^ n852 ^ 1'b0 ;
  assign n905 = n669 & ~n904 ;
  assign n906 = n905 ^ n368 ^ 1'b0 ;
  assign n907 = x74 & x110 ;
  assign n908 = n907 ^ n482 ^ 1'b0 ;
  assign n909 = ( n283 & n623 ) | ( n283 & ~n908 ) | ( n623 & ~n908 ) ;
  assign n910 = n576 ^ n558 ^ 1'b0 ;
  assign n911 = n339 | n910 ;
  assign n912 = ( x21 & n363 ) | ( x21 & ~n528 ) | ( n363 & ~n528 ) ;
  assign n913 = ( n829 & ~n911 ) | ( n829 & n912 ) | ( ~n911 & n912 ) ;
  assign n914 = ( n256 & ~n273 ) | ( n256 & n393 ) | ( ~n273 & n393 ) ;
  assign n915 = n400 ^ n258 ^ 1'b0 ;
  assign n916 = ( n721 & n914 ) | ( n721 & n915 ) | ( n914 & n915 ) ;
  assign n917 = ( ~n268 & n355 ) | ( ~n268 & n593 ) | ( n355 & n593 ) ;
  assign n929 = n877 ^ n716 ^ n445 ;
  assign n921 = n229 ^ n160 ^ x96 ;
  assign n922 = n573 ^ n502 ^ n400 ;
  assign n923 = n922 ^ n251 ^ n231 ;
  assign n924 = ( n541 & n590 ) | ( n541 & ~n923 ) | ( n590 & ~n923 ) ;
  assign n925 = ( n493 & n921 ) | ( n493 & ~n924 ) | ( n921 & ~n924 ) ;
  assign n918 = n165 ^ n130 ^ 1'b0 ;
  assign n919 = ( n160 & n407 ) | ( n160 & n918 ) | ( n407 & n918 ) ;
  assign n920 = n919 ^ n710 ^ 1'b0 ;
  assign n926 = n925 ^ n920 ^ n266 ;
  assign n927 = n183 & n926 ;
  assign n928 = ~n908 & n927 ;
  assign n930 = n929 ^ n928 ^ n440 ;
  assign n931 = ( ~x127 & n452 ) | ( ~x127 & n512 ) | ( n452 & n512 ) ;
  assign n932 = ( x94 & n158 ) | ( x94 & n931 ) | ( n158 & n931 ) ;
  assign n933 = ( ~x94 & n465 ) | ( ~x94 & n880 ) | ( n465 & n880 ) ;
  assign n934 = ( x4 & n160 ) | ( x4 & n933 ) | ( n160 & n933 ) ;
  assign n935 = n165 ^ x44 ^ x10 ;
  assign n936 = ( x29 & n543 ) | ( x29 & n644 ) | ( n543 & n644 ) ;
  assign n937 = ( x101 & n935 ) | ( x101 & ~n936 ) | ( n935 & ~n936 ) ;
  assign n938 = x8 & n937 ;
  assign n939 = n938 ^ n331 ^ 1'b0 ;
  assign n940 = ( x14 & ~n934 ) | ( x14 & n939 ) | ( ~n934 & n939 ) ;
  assign n943 = ( n545 & ~n693 ) | ( n545 & n747 ) | ( ~n693 & n747 ) ;
  assign n944 = n943 ^ n704 ^ n496 ;
  assign n941 = n525 ^ n239 ^ x78 ;
  assign n942 = x75 & ~n941 ;
  assign n945 = n944 ^ n942 ^ 1'b0 ;
  assign n946 = ( x61 & ~n423 ) | ( x61 & n945 ) | ( ~n423 & n945 ) ;
  assign n947 = n291 ^ x68 ^ 1'b0 ;
  assign n948 = n946 & n947 ;
  assign n949 = n588 ^ n388 ^ n281 ;
  assign n950 = n471 | n636 ;
  assign n951 = n950 ^ n298 ^ 1'b0 ;
  assign n952 = n951 ^ n335 ^ n233 ;
  assign n953 = ( n135 & n155 ) | ( n135 & ~n171 ) | ( n155 & ~n171 ) ;
  assign n954 = n858 ^ n677 ^ 1'b0 ;
  assign n955 = n627 ^ x94 ^ x77 ;
  assign n956 = n955 ^ n412 ^ n258 ;
  assign n957 = n894 & ~n956 ;
  assign n958 = n954 & n957 ;
  assign n959 = ( x13 & n261 ) | ( x13 & ~n867 ) | ( n261 & ~n867 ) ;
  assign n960 = ( ~n545 & n958 ) | ( ~n545 & n959 ) | ( n958 & n959 ) ;
  assign n961 = n261 & ~n425 ;
  assign n962 = x95 ^ x77 ^ 1'b0 ;
  assign n963 = n962 ^ n716 ^ n380 ;
  assign n964 = ( n196 & ~n453 ) | ( n196 & n962 ) | ( ~n453 & n962 ) ;
  assign n965 = n418 ^ n374 ^ 1'b0 ;
  assign n966 = ~n340 & n965 ;
  assign n967 = n966 ^ n329 ^ 1'b0 ;
  assign n968 = ~n964 & n967 ;
  assign n969 = ( n961 & n963 ) | ( n961 & ~n968 ) | ( n963 & ~n968 ) ;
  assign n970 = n969 ^ n793 ^ n768 ;
  assign n971 = n426 & ~n970 ;
  assign n972 = n971 ^ n248 ^ 1'b0 ;
  assign n973 = ~n180 & n314 ;
  assign n974 = n972 & n973 ;
  assign n987 = n347 ^ n183 ^ x7 ;
  assign n988 = n987 ^ n825 ^ n396 ;
  assign n989 = n988 ^ n491 ^ n149 ;
  assign n981 = n583 ^ n272 ^ x62 ;
  assign n982 = n475 & ~n981 ;
  assign n983 = n982 ^ n543 ^ 1'b0 ;
  assign n984 = n344 & n983 ;
  assign n979 = n574 ^ n323 ^ 1'b0 ;
  assign n980 = x65 & ~n979 ;
  assign n985 = n984 ^ n980 ^ n464 ;
  assign n975 = x37 & n239 ;
  assign n976 = ( x91 & n237 ) | ( x91 & ~n423 ) | ( n237 & ~n423 ) ;
  assign n977 = ( x89 & x123 ) | ( x89 & ~n976 ) | ( x123 & ~n976 ) ;
  assign n978 = ( n947 & n975 ) | ( n947 & ~n977 ) | ( n975 & ~n977 ) ;
  assign n986 = n985 ^ n978 ^ n354 ;
  assign n990 = n989 ^ n986 ^ n861 ;
  assign n994 = ( x29 & ~x35 ) | ( x29 & n449 ) | ( ~x35 & n449 ) ;
  assign n991 = n424 ^ n289 ^ n237 ;
  assign n992 = ( ~n383 & n411 ) | ( ~n383 & n991 ) | ( n411 & n991 ) ;
  assign n993 = n992 ^ n729 ^ n157 ;
  assign n995 = n994 ^ n993 ^ n653 ;
  assign n996 = n995 ^ n978 ^ 1'b0 ;
  assign n997 = n996 ^ n582 ^ n384 ;
  assign n998 = ( n257 & n317 ) | ( n257 & n486 ) | ( n317 & n486 ) ;
  assign n999 = ( x58 & ~n284 ) | ( x58 & n998 ) | ( ~n284 & n998 ) ;
  assign n1000 = ( x0 & n209 ) | ( x0 & n783 ) | ( n209 & n783 ) ;
  assign n1001 = ( ~n302 & n999 ) | ( ~n302 & n1000 ) | ( n999 & n1000 ) ;
  assign n1002 = n1001 ^ n793 ^ 1'b0 ;
  assign n1003 = n404 & ~n1002 ;
  assign n1005 = ( n189 & n502 ) | ( n189 & n628 ) | ( n502 & n628 ) ;
  assign n1006 = ( n319 & ~n721 ) | ( n319 & n1005 ) | ( ~n721 & n1005 ) ;
  assign n1004 = ( n447 & n536 ) | ( n447 & n570 ) | ( n536 & n570 ) ;
  assign n1007 = n1006 ^ n1004 ^ n526 ;
  assign n1010 = n921 ^ n919 ^ x70 ;
  assign n1008 = ( n482 & n664 ) | ( n482 & ~n823 ) | ( n664 & ~n823 ) ;
  assign n1009 = n1008 ^ n728 ^ n648 ;
  assign n1011 = n1010 ^ n1009 ^ n634 ;
  assign n1012 = n981 ^ n380 ^ n294 ;
  assign n1013 = ~n573 & n592 ;
  assign n1014 = n629 ^ n176 ^ 1'b0 ;
  assign n1015 = ( ~n400 & n521 ) | ( ~n400 & n1014 ) | ( n521 & n1014 ) ;
  assign n1016 = ( n716 & ~n1013 ) | ( n716 & n1015 ) | ( ~n1013 & n1015 ) ;
  assign n1017 = ( n233 & n1012 ) | ( n233 & n1016 ) | ( n1012 & n1016 ) ;
  assign n1018 = ( n376 & n511 ) | ( n376 & ~n1017 ) | ( n511 & ~n1017 ) ;
  assign n1022 = n249 ^ n207 ^ x2 ;
  assign n1023 = n1022 ^ n635 ^ 1'b0 ;
  assign n1024 = n130 | n1023 ;
  assign n1020 = n613 ^ n343 ^ x85 ;
  assign n1021 = ( n413 & n875 ) | ( n413 & n1020 ) | ( n875 & n1020 ) ;
  assign n1019 = n725 ^ n367 ^ n338 ;
  assign n1025 = n1024 ^ n1021 ^ n1019 ;
  assign n1029 = x78 & ~n347 ;
  assign n1030 = n1029 ^ n545 ^ 1'b0 ;
  assign n1027 = x108 | n187 ;
  assign n1026 = n784 ^ n173 ^ x10 ;
  assign n1028 = n1027 ^ n1026 ^ 1'b0 ;
  assign n1031 = n1030 ^ n1028 ^ n796 ;
  assign n1032 = n983 ^ n372 ^ n131 ;
  assign n1033 = n442 & n1032 ;
  assign n1034 = n1033 ^ n645 ^ 1'b0 ;
  assign n1035 = n1034 ^ n639 ^ 1'b0 ;
  assign n1037 = ( n138 & ~n342 ) | ( n138 & n733 ) | ( ~n342 & n733 ) ;
  assign n1036 = n669 ^ n343 ^ n287 ;
  assign n1038 = n1037 ^ n1036 ^ n229 ;
  assign n1039 = ~n975 & n1038 ;
  assign n1041 = n430 & ~n523 ;
  assign n1040 = n325 ^ x87 ^ 1'b0 ;
  assign n1042 = n1041 ^ n1040 ^ n1000 ;
  assign n1048 = n999 ^ n199 ^ x89 ;
  assign n1047 = n935 ^ n198 ^ x17 ;
  assign n1045 = ( x86 & n373 ) | ( x86 & n450 ) | ( n373 & n450 ) ;
  assign n1043 = n226 ^ x52 ^ 1'b0 ;
  assign n1044 = n195 | n1043 ;
  assign n1046 = n1045 ^ n1044 ^ x116 ;
  assign n1049 = n1048 ^ n1047 ^ n1046 ;
  assign n1050 = n686 ^ n657 ^ n584 ;
  assign n1051 = n1050 ^ n188 ^ n148 ;
  assign n1052 = ( n605 & n1049 ) | ( n605 & ~n1051 ) | ( n1049 & ~n1051 ) ;
  assign n1053 = ( n368 & n1012 ) | ( n368 & n1052 ) | ( n1012 & n1052 ) ;
  assign n1055 = x62 & n144 ;
  assign n1054 = ( x38 & n654 ) | ( x38 & ~n995 ) | ( n654 & ~n995 ) ;
  assign n1056 = n1055 ^ n1054 ^ n145 ;
  assign n1057 = ( n167 & n298 ) | ( n167 & n696 ) | ( n298 & n696 ) ;
  assign n1058 = n1057 ^ n312 ^ 1'b0 ;
  assign n1059 = n592 ^ n223 ^ n133 ;
  assign n1060 = x61 & x108 ;
  assign n1061 = n1060 ^ n409 ^ 1'b0 ;
  assign n1062 = n1061 ^ x123 ^ x77 ;
  assign n1063 = ( x28 & n772 ) | ( x28 & ~n1062 ) | ( n772 & ~n1062 ) ;
  assign n1064 = ( ~n736 & n760 ) | ( ~n736 & n1063 ) | ( n760 & n1063 ) ;
  assign n1065 = n236 | n623 ;
  assign n1066 = n1065 ^ n480 ^ n188 ;
  assign n1067 = x118 & n1066 ;
  assign n1068 = n159 & n1067 ;
  assign n1070 = n215 & ~n782 ;
  assign n1071 = ~n406 & n1070 ;
  assign n1072 = ( ~n885 & n991 ) | ( ~n885 & n1071 ) | ( n991 & n1071 ) ;
  assign n1069 = ( x16 & ~x67 ) | ( x16 & n180 ) | ( ~x67 & n180 ) ;
  assign n1073 = n1072 ^ n1069 ^ x45 ;
  assign n1074 = n961 ^ n329 ^ 1'b0 ;
  assign n1075 = n1073 | n1074 ;
  assign n1076 = ( n426 & n505 ) | ( n426 & n1075 ) | ( n505 & n1075 ) ;
  assign n1077 = ( n717 & n810 ) | ( n717 & ~n908 ) | ( n810 & ~n908 ) ;
  assign n1078 = ( x22 & n1076 ) | ( x22 & ~n1077 ) | ( n1076 & ~n1077 ) ;
  assign n1082 = n577 & ~n626 ;
  assign n1083 = ~n732 & n1082 ;
  assign n1084 = ( n762 & ~n981 ) | ( n762 & n1083 ) | ( ~n981 & n1083 ) ;
  assign n1079 = n985 ^ n266 ^ x120 ;
  assign n1080 = n1079 ^ n828 ^ n466 ;
  assign n1081 = n1080 ^ n1032 ^ n302 ;
  assign n1085 = n1084 ^ n1081 ^ 1'b0 ;
  assign n1086 = ~n1078 & n1085 ;
  assign n1087 = ( n145 & n276 ) | ( n145 & ~n356 ) | ( n276 & ~n356 ) ;
  assign n1088 = ~n964 & n1087 ;
  assign n1097 = n244 | n292 ;
  assign n1098 = n386 & n1097 ;
  assign n1099 = n187 | n1098 ;
  assign n1100 = n1099 ^ n159 ^ 1'b0 ;
  assign n1089 = n554 ^ n407 ^ x73 ;
  assign n1090 = n815 & ~n1037 ;
  assign n1091 = n1090 ^ x51 ^ 1'b0 ;
  assign n1092 = n1091 ^ n899 ^ n661 ;
  assign n1093 = n209 ^ n149 ^ x8 ;
  assign n1094 = n1092 & n1093 ;
  assign n1095 = n1094 ^ n164 ^ 1'b0 ;
  assign n1096 = n1089 & ~n1095 ;
  assign n1101 = n1100 ^ n1096 ^ 1'b0 ;
  assign n1102 = n811 ^ n753 ^ n252 ;
  assign n1103 = ( x17 & n754 ) | ( x17 & n770 ) | ( n754 & n770 ) ;
  assign n1104 = ( n620 & n987 ) | ( n620 & ~n1103 ) | ( n987 & ~n1103 ) ;
  assign n1105 = ( ~n740 & n1102 ) | ( ~n740 & n1104 ) | ( n1102 & n1104 ) ;
  assign n1106 = n1105 ^ x57 ^ 1'b0 ;
  assign n1107 = n1101 & ~n1106 ;
  assign n1108 = n245 ^ n233 ^ 1'b0 ;
  assign n1109 = ( n256 & n1091 ) | ( n256 & ~n1108 ) | ( n1091 & ~n1108 ) ;
  assign n1110 = ~n961 & n1109 ;
  assign n1111 = n384 & ~n814 ;
  assign n1112 = ~n299 & n1111 ;
  assign n1113 = n237 ^ x87 ^ x17 ;
  assign n1114 = n1113 ^ x89 ^ 1'b0 ;
  assign n1115 = n621 | n651 ;
  assign n1133 = ( n352 & ~n478 ) | ( n352 & n716 ) | ( ~n478 & n716 ) ;
  assign n1132 = x20 & n495 ;
  assign n1134 = n1133 ^ n1132 ^ n649 ;
  assign n1116 = x20 | n492 ;
  assign n1117 = ( ~n149 & n499 ) | ( ~n149 & n1116 ) | ( n499 & n1116 ) ;
  assign n1118 = n335 & n1117 ;
  assign n1119 = n675 & n1118 ;
  assign n1120 = n1119 ^ n750 ^ n339 ;
  assign n1121 = n614 ^ n605 ^ n184 ;
  assign n1122 = ( ~n941 & n1120 ) | ( ~n941 & n1121 ) | ( n1120 & n1121 ) ;
  assign n1123 = ( x93 & n798 ) | ( x93 & ~n1122 ) | ( n798 & ~n1122 ) ;
  assign n1124 = n735 ^ n139 ^ x119 ;
  assign n1125 = n188 ^ x120 ^ x94 ;
  assign n1126 = ( n461 & n603 ) | ( n461 & ~n878 ) | ( n603 & ~n878 ) ;
  assign n1127 = ( x70 & n327 ) | ( x70 & n391 ) | ( n327 & n391 ) ;
  assign n1128 = ~n1126 & n1127 ;
  assign n1129 = ~n1125 & n1128 ;
  assign n1130 = n1124 | n1129 ;
  assign n1131 = n1123 & ~n1130 ;
  assign n1135 = n1134 ^ n1131 ^ n610 ;
  assign n1138 = n553 ^ n382 ^ x9 ;
  assign n1139 = ( n844 & n961 ) | ( n844 & ~n1138 ) | ( n961 & ~n1138 ) ;
  assign n1140 = ~n320 & n1139 ;
  assign n1141 = ~n377 & n1140 ;
  assign n1142 = ( ~n486 & n653 ) | ( ~n486 & n1141 ) | ( n653 & n1141 ) ;
  assign n1136 = n583 ^ x32 ^ x7 ;
  assign n1137 = n503 & n1136 ;
  assign n1143 = n1142 ^ n1137 ^ 1'b0 ;
  assign n1144 = ( n582 & n819 ) | ( n582 & n1143 ) | ( n819 & n1143 ) ;
  assign n1145 = n1110 ^ n1041 ^ n142 ;
  assign n1152 = n495 ^ n183 ^ x3 ;
  assign n1153 = n1152 ^ n936 ^ n626 ;
  assign n1154 = n505 ^ n471 ^ n292 ;
  assign n1155 = n285 & n693 ;
  assign n1156 = n1155 ^ n484 ^ 1'b0 ;
  assign n1157 = n1154 | n1156 ;
  assign n1158 = n1153 | n1157 ;
  assign n1148 = ( n142 & n145 ) | ( n142 & ~n237 ) | ( n145 & ~n237 ) ;
  assign n1149 = n631 ^ n533 ^ n475 ;
  assign n1150 = ( n837 & n1139 ) | ( n837 & ~n1149 ) | ( n1139 & ~n1149 ) ;
  assign n1151 = ( n391 & n1148 ) | ( n391 & n1150 ) | ( n1148 & n1150 ) ;
  assign n1146 = ( ~n434 & n655 ) | ( ~n434 & n722 ) | ( n655 & n722 ) ;
  assign n1147 = n1146 ^ n993 ^ x70 ;
  assign n1159 = n1158 ^ n1151 ^ n1147 ;
  assign n1160 = n1159 ^ n916 ^ n730 ;
  assign n1179 = ( ~n164 & n457 ) | ( ~n164 & n861 ) | ( n457 & n861 ) ;
  assign n1180 = n1179 ^ n437 ^ 1'b0 ;
  assign n1177 = ~n585 & n903 ;
  assign n1178 = ~n198 & n1177 ;
  assign n1175 = n556 ^ n258 ^ n191 ;
  assign n1169 = ( n238 & ~n382 ) | ( n238 & n588 ) | ( ~n382 & n588 ) ;
  assign n1170 = ( ~x93 & n554 ) | ( ~x93 & n1169 ) | ( n554 & n1169 ) ;
  assign n1171 = ( ~n145 & n360 ) | ( ~n145 & n575 ) | ( n360 & n575 ) ;
  assign n1172 = n1171 ^ n832 ^ n780 ;
  assign n1173 = x5 & n1172 ;
  assign n1174 = n1170 & n1173 ;
  assign n1165 = ( ~x71 & n506 ) | ( ~x71 & n535 ) | ( n506 & n535 ) ;
  assign n1163 = ( n351 & n860 ) | ( n351 & n1005 ) | ( n860 & n1005 ) ;
  assign n1164 = ( ~n298 & n1013 ) | ( ~n298 & n1163 ) | ( n1013 & n1163 ) ;
  assign n1166 = n1165 ^ n1164 ^ n610 ;
  assign n1167 = ( n815 & ~n1122 ) | ( n815 & n1166 ) | ( ~n1122 & n1166 ) ;
  assign n1161 = n470 ^ n229 ^ 1'b0 ;
  assign n1162 = n780 & n1161 ;
  assign n1168 = n1167 ^ n1162 ^ 1'b0 ;
  assign n1176 = n1175 ^ n1174 ^ n1168 ;
  assign n1181 = n1180 ^ n1178 ^ n1176 ;
  assign n1182 = n575 ^ n167 ^ x94 ;
  assign n1183 = n1182 ^ n722 ^ 1'b0 ;
  assign n1184 = ( x43 & n418 ) | ( x43 & n658 ) | ( n418 & n658 ) ;
  assign n1185 = n441 ^ n379 ^ 1'b0 ;
  assign n1186 = n1184 & n1185 ;
  assign n1187 = ( n211 & n1183 ) | ( n211 & n1186 ) | ( n1183 & n1186 ) ;
  assign n1188 = n728 ^ n441 ^ 1'b0 ;
  assign n1189 = n1188 ^ n1186 ^ n364 ;
  assign n1190 = n786 ^ x127 ^ 1'b0 ;
  assign n1191 = n491 & ~n1190 ;
  assign n1192 = ~n1133 & n1191 ;
  assign n1193 = n483 & n1192 ;
  assign n1194 = n1193 ^ n397 ^ x44 ;
  assign n1195 = n1194 ^ n165 ^ 1'b0 ;
  assign n1196 = n308 ^ x126 ^ 1'b0 ;
  assign n1197 = ~n181 & n1196 ;
  assign n1198 = ~n677 & n1197 ;
  assign n1199 = n1198 ^ x55 ^ 1'b0 ;
  assign n1200 = n750 & ~n1199 ;
  assign n1201 = n1200 ^ n628 ^ 1'b0 ;
  assign n1202 = n616 & n667 ;
  assign n1203 = n1202 ^ n722 ^ 1'b0 ;
  assign n1204 = ~n434 & n896 ;
  assign n1205 = n1204 ^ n395 ^ 1'b0 ;
  assign n1206 = ( n427 & ~n1203 ) | ( n427 & n1205 ) | ( ~n1203 & n1205 ) ;
  assign n1207 = ( n335 & n1201 ) | ( n335 & n1206 ) | ( n1201 & n1206 ) ;
  assign n1214 = n447 ^ n305 ^ x116 ;
  assign n1210 = n476 ^ x74 ^ x61 ;
  assign n1211 = ( ~n129 & n310 ) | ( ~n129 & n1210 ) | ( n310 & n1210 ) ;
  assign n1212 = n1211 ^ n791 ^ 1'b0 ;
  assign n1208 = n331 & n653 ;
  assign n1209 = n1208 ^ n1193 ^ 1'b0 ;
  assign n1213 = n1212 ^ n1209 ^ n1151 ;
  assign n1215 = n1214 ^ n1213 ^ n285 ;
  assign n1216 = n668 ^ n339 ^ n248 ;
  assign n1217 = n1216 ^ n923 ^ n871 ;
  assign n1218 = n1217 ^ n893 ^ n795 ;
  assign n1219 = n945 ^ n711 ^ n192 ;
  assign n1220 = ~n402 & n820 ;
  assign n1221 = n1220 ^ n1024 ^ 1'b0 ;
  assign n1222 = n547 & n1221 ;
  assign n1223 = n242 & n281 ;
  assign n1224 = n1223 ^ n418 ^ 1'b0 ;
  assign n1225 = n1224 ^ n408 ^ n318 ;
  assign n1226 = n834 ^ n575 ^ x33 ;
  assign n1227 = ( n497 & n921 ) | ( n497 & n1226 ) | ( n921 & n1226 ) ;
  assign n1228 = ( n381 & n1225 ) | ( n381 & ~n1227 ) | ( n1225 & ~n1227 ) ;
  assign n1229 = n962 & n1152 ;
  assign n1230 = x108 & n348 ;
  assign n1231 = n198 ^ x94 ^ 1'b0 ;
  assign n1232 = n384 ^ n198 ^ 1'b0 ;
  assign n1233 = ( n712 & n1231 ) | ( n712 & n1232 ) | ( n1231 & n1232 ) ;
  assign n1234 = n1233 ^ n694 ^ 1'b0 ;
  assign n1235 = n1234 ^ n721 ^ n229 ;
  assign n1236 = n260 & ~n1235 ;
  assign n1237 = ~n620 & n1236 ;
  assign n1241 = n681 ^ n461 ^ n189 ;
  assign n1238 = n592 ^ x40 ^ 1'b0 ;
  assign n1239 = n457 & n1238 ;
  assign n1240 = n289 & n1239 ;
  assign n1242 = n1241 ^ n1240 ^ 1'b0 ;
  assign n1243 = ( n503 & ~n1075 ) | ( n503 & n1242 ) | ( ~n1075 & n1242 ) ;
  assign n1244 = n652 ^ n647 ^ n397 ;
  assign n1245 = x110 & ~n1244 ;
  assign n1246 = n661 ^ n509 ^ x6 ;
  assign n1247 = ( x93 & n142 ) | ( x93 & ~n1246 ) | ( n142 & ~n1246 ) ;
  assign n1248 = n1247 ^ n818 ^ n404 ;
  assign n1249 = n1248 ^ n620 ^ 1'b0 ;
  assign n1250 = ( n244 & n1247 ) | ( n244 & n1249 ) | ( n1247 & n1249 ) ;
  assign n1251 = n818 ^ n391 ^ n370 ;
  assign n1252 = ( n220 & n456 ) | ( n220 & n1251 ) | ( n456 & n1251 ) ;
  assign n1253 = ( n831 & ~n881 ) | ( n831 & n1252 ) | ( ~n881 & n1252 ) ;
  assign n1254 = n1253 ^ n393 ^ n215 ;
  assign n1255 = ( x4 & ~n419 ) | ( x4 & n1124 ) | ( ~n419 & n1124 ) ;
  assign n1256 = n820 ^ x41 ^ 1'b0 ;
  assign n1257 = x119 & n1256 ;
  assign n1258 = ~x33 & n1257 ;
  assign n1259 = n1258 ^ n525 ^ n289 ;
  assign n1260 = n272 & n1259 ;
  assign n1261 = n1009 & n1260 ;
  assign n1262 = n1261 ^ n533 ^ 1'b0 ;
  assign n1266 = ( ~x13 & n129 ) | ( ~x13 & n247 ) | ( n129 & n247 ) ;
  assign n1263 = n774 ^ n398 ^ x49 ;
  assign n1264 = ~n730 & n798 ;
  assign n1265 = n1263 | n1264 ;
  assign n1267 = n1266 ^ n1265 ^ n891 ;
  assign n1268 = ( n1255 & n1262 ) | ( n1255 & n1267 ) | ( n1262 & n1267 ) ;
  assign n1270 = n1183 ^ n257 ^ x47 ;
  assign n1269 = n404 ^ x59 ^ x22 ;
  assign n1271 = n1270 ^ n1269 ^ x49 ;
  assign n1272 = n568 ^ n257 ^ x41 ;
  assign n1273 = n402 ^ n193 ^ x16 ;
  assign n1274 = ( x125 & ~n344 ) | ( x125 & n607 ) | ( ~n344 & n607 ) ;
  assign n1275 = n438 ^ n159 ^ x99 ;
  assign n1276 = ( n441 & ~n1274 ) | ( n441 & n1275 ) | ( ~n1274 & n1275 ) ;
  assign n1277 = n1276 ^ n658 ^ x52 ;
  assign n1278 = ( n1272 & n1273 ) | ( n1272 & ~n1277 ) | ( n1273 & ~n1277 ) ;
  assign n1279 = ( n135 & n325 ) | ( n135 & ~n923 ) | ( n325 & ~n923 ) ;
  assign n1280 = n1279 ^ n511 ^ n294 ;
  assign n1281 = n828 ^ n597 ^ 1'b0 ;
  assign n1282 = n1281 ^ n426 ^ 1'b0 ;
  assign n1283 = ( n434 & ~n1280 ) | ( n434 & n1282 ) | ( ~n1280 & n1282 ) ;
  assign n1284 = ( ~n772 & n852 ) | ( ~n772 & n1083 ) | ( n852 & n1083 ) ;
  assign n1285 = ( n420 & n568 ) | ( n420 & ~n1133 ) | ( n568 & ~n1133 ) ;
  assign n1286 = n1285 ^ n570 ^ n193 ;
  assign n1287 = ( n503 & ~n524 ) | ( n503 & n1159 ) | ( ~n524 & n1159 ) ;
  assign n1288 = n635 ^ n566 ^ 1'b0 ;
  assign n1289 = n1288 ^ n1063 ^ n235 ;
  assign n1290 = ( n1286 & ~n1287 ) | ( n1286 & n1289 ) | ( ~n1287 & n1289 ) ;
  assign n1292 = n472 ^ n408 ^ x109 ;
  assign n1296 = ( n701 & n820 ) | ( n701 & n1292 ) | ( n820 & n1292 ) ;
  assign n1291 = n509 ^ n242 ^ n234 ;
  assign n1293 = n149 | n1292 ;
  assign n1294 = n601 | n1293 ;
  assign n1295 = ( n665 & n1291 ) | ( n665 & n1294 ) | ( n1291 & n1294 ) ;
  assign n1297 = n1296 ^ n1295 ^ 1'b0 ;
  assign n1298 = n402 & ~n1297 ;
  assign n1299 = ~n1241 & n1298 ;
  assign n1300 = n1299 ^ n554 ^ 1'b0 ;
  assign n1308 = ( n226 & n476 ) | ( n226 & ~n799 ) | ( n476 & ~n799 ) ;
  assign n1304 = ( n541 & n975 ) | ( n541 & ~n1126 ) | ( n975 & ~n1126 ) ;
  assign n1305 = n358 | n1304 ;
  assign n1306 = ( ~x91 & x114 ) | ( ~x91 & n1305 ) | ( x114 & n1305 ) ;
  assign n1307 = ( ~n709 & n1291 ) | ( ~n709 & n1306 ) | ( n1291 & n1306 ) ;
  assign n1301 = n671 ^ n165 ^ 1'b0 ;
  assign n1302 = n209 | n1301 ;
  assign n1303 = n738 & ~n1302 ;
  assign n1309 = n1308 ^ n1307 ^ n1303 ;
  assign n1310 = ( n168 & ~n457 ) | ( n168 & n491 ) | ( ~n457 & n491 ) ;
  assign n1311 = x57 & n644 ;
  assign n1312 = n1311 ^ n131 ^ 1'b0 ;
  assign n1313 = ( n279 & n340 ) | ( n279 & ~n1312 ) | ( n340 & ~n1312 ) ;
  assign n1314 = ( n388 & ~n570 ) | ( n388 & n1313 ) | ( ~n570 & n1313 ) ;
  assign n1315 = ( n317 & ~n1310 ) | ( n317 & n1314 ) | ( ~n1310 & n1314 ) ;
  assign n1316 = n961 ^ n846 ^ x79 ;
  assign n1317 = n618 | n1316 ;
  assign n1320 = ( ~x33 & n406 ) | ( ~x33 & n513 ) | ( n406 & n513 ) ;
  assign n1318 = n837 ^ n512 ^ n401 ;
  assign n1319 = n1318 ^ n863 ^ n354 ;
  assign n1321 = n1320 ^ n1319 ^ 1'b0 ;
  assign n1322 = n1317 | n1321 ;
  assign n1323 = n264 | n1154 ;
  assign n1324 = n1323 ^ n1171 ^ 1'b0 ;
  assign n1325 = ( ~n855 & n1019 ) | ( ~n855 & n1324 ) | ( n1019 & n1324 ) ;
  assign n1326 = n1008 ^ n284 ^ 1'b0 ;
  assign n1327 = ( ~n482 & n698 ) | ( ~n482 & n1326 ) | ( n698 & n1326 ) ;
  assign n1328 = ( n206 & ~n1146 ) | ( n206 & n1327 ) | ( ~n1146 & n1327 ) ;
  assign n1337 = ( x23 & x81 ) | ( x23 & ~x109 ) | ( x81 & ~x109 ) ;
  assign n1329 = ~n223 & n1036 ;
  assign n1332 = n341 & n422 ;
  assign n1333 = n1332 ^ n584 ^ n557 ;
  assign n1334 = x119 & n1333 ;
  assign n1330 = n496 & ~n769 ;
  assign n1331 = ~n141 & n1330 ;
  assign n1335 = n1334 ^ n1331 ^ 1'b0 ;
  assign n1336 = ( n783 & ~n1329 ) | ( n783 & n1335 ) | ( ~n1329 & n1335 ) ;
  assign n1338 = n1337 ^ n1336 ^ 1'b0 ;
  assign n1339 = n1196 ^ n611 ^ x44 ;
  assign n1340 = n1170 | n1339 ;
  assign n1341 = n277 & n1340 ;
  assign n1342 = n1341 ^ n1273 ^ 1'b0 ;
  assign n1343 = ( x38 & ~n460 ) | ( x38 & n590 ) | ( ~n460 & n590 ) ;
  assign n1344 = n814 ^ n642 ^ n353 ;
  assign n1345 = n1161 ^ n425 ^ 1'b0 ;
  assign n1346 = n1344 & n1345 ;
  assign n1347 = ( n392 & n722 ) | ( n392 & n1346 ) | ( n722 & n1346 ) ;
  assign n1348 = n1347 ^ n1344 ^ n999 ;
  assign n1349 = ( ~n352 & n901 ) | ( ~n352 & n1348 ) | ( n901 & n1348 ) ;
  assign n1350 = n484 ^ n305 ^ n285 ;
  assign n1351 = ( x83 & n761 ) | ( x83 & n1350 ) | ( n761 & n1350 ) ;
  assign n1352 = x91 | n551 ;
  assign n1353 = n1332 ^ n444 ^ 1'b0 ;
  assign n1354 = n502 & n1353 ;
  assign n1355 = ~n341 & n707 ;
  assign n1356 = ~n936 & n1355 ;
  assign n1357 = n1025 ^ n1014 ^ n985 ;
  assign n1358 = n735 | n1357 ;
  assign n1359 = n1356 & ~n1358 ;
  assign n1360 = ( n1207 & ~n1354 ) | ( n1207 & n1359 ) | ( ~n1354 & n1359 ) ;
  assign n1361 = ( ~n1351 & n1352 ) | ( ~n1351 & n1360 ) | ( n1352 & n1360 ) ;
  assign n1362 = n1091 ^ n251 ^ x5 ;
  assign n1363 = n1292 ^ n466 ^ 1'b0 ;
  assign n1364 = ~n287 & n375 ;
  assign n1365 = ( n355 & ~n1363 ) | ( n355 & n1364 ) | ( ~n1363 & n1364 ) ;
  assign n1366 = ~n563 & n620 ;
  assign n1367 = n1366 ^ n468 ^ 1'b0 ;
  assign n1368 = n131 & ~n1102 ;
  assign n1369 = ( n1365 & n1367 ) | ( n1365 & ~n1368 ) | ( n1367 & ~n1368 ) ;
  assign n1372 = n197 ^ n168 ^ n165 ;
  assign n1373 = n1372 ^ n370 ^ x102 ;
  assign n1370 = ~n177 & n656 ;
  assign n1371 = n1370 ^ x7 ^ 1'b0 ;
  assign n1374 = n1373 ^ n1371 ^ n202 ;
  assign n1375 = ( x113 & ~n727 ) | ( x113 & n1374 ) | ( ~n727 & n1374 ) ;
  assign n1376 = ~n238 & n1375 ;
  assign n1377 = n1369 & n1376 ;
  assign n1378 = ( n1219 & n1362 ) | ( n1219 & n1377 ) | ( n1362 & n1377 ) ;
  assign n1380 = ( n200 & ~n214 ) | ( n200 & n696 ) | ( ~n214 & n696 ) ;
  assign n1381 = ( x124 & n842 ) | ( x124 & ~n1380 ) | ( n842 & ~n1380 ) ;
  assign n1379 = n1183 ^ n1104 ^ n1077 ;
  assign n1382 = n1381 ^ n1379 ^ n1015 ;
  assign n1383 = ~x127 & n521 ;
  assign n1384 = n1383 ^ n1112 ^ n859 ;
  assign n1385 = n369 & n1384 ;
  assign n1386 = n473 & ~n754 ;
  assign n1387 = n1231 ^ n974 ^ n162 ;
  assign n1392 = x29 & n222 ;
  assign n1393 = ( n182 & n514 ) | ( n182 & n1392 ) | ( n514 & n1392 ) ;
  assign n1389 = x19 & n440 ;
  assign n1390 = n1389 ^ x69 ^ 1'b0 ;
  assign n1391 = ( n810 & ~n1037 ) | ( n810 & n1390 ) | ( ~n1037 & n1390 ) ;
  assign n1388 = ( x46 & ~x74 ) | ( x46 & n599 ) | ( ~x74 & n599 ) ;
  assign n1394 = n1393 ^ n1391 ^ n1388 ;
  assign n1395 = n417 ^ n411 ^ x31 ;
  assign n1396 = ( n457 & ~n727 ) | ( n457 & n1395 ) | ( ~n727 & n1395 ) ;
  assign n1397 = n1396 ^ n1287 ^ 1'b0 ;
  assign n1398 = n525 ^ n513 ^ n424 ;
  assign n1399 = n1398 ^ n1313 ^ 1'b0 ;
  assign n1400 = n448 ^ n237 ^ 1'b0 ;
  assign n1401 = n1400 ^ n319 ^ 1'b0 ;
  assign n1402 = ( n323 & n1014 ) | ( n323 & ~n1065 ) | ( n1014 & ~n1065 ) ;
  assign n1403 = ~n157 & n1402 ;
  assign n1404 = x42 & ~n408 ;
  assign n1405 = n1404 ^ x0 ^ 1'b0 ;
  assign n1406 = n1405 ^ n987 ^ 1'b0 ;
  assign n1407 = ( ~n1078 & n1403 ) | ( ~n1078 & n1406 ) | ( n1403 & n1406 ) ;
  assign n1408 = n1401 & n1407 ;
  assign n1409 = ~n1399 & n1408 ;
  assign n1412 = n769 ^ n727 ^ x97 ;
  assign n1411 = ( n990 & n1071 ) | ( n990 & n1077 ) | ( n1071 & n1077 ) ;
  assign n1410 = ( x75 & n201 ) | ( x75 & n900 ) | ( n201 & n900 ) ;
  assign n1413 = n1412 ^ n1411 ^ n1410 ;
  assign n1414 = n1413 ^ n814 ^ n388 ;
  assign n1415 = ( n191 & ~n449 ) | ( n191 & n780 ) | ( ~n449 & n780 ) ;
  assign n1416 = n1050 ^ n1036 ^ 1'b0 ;
  assign n1417 = x26 & n188 ;
  assign n1418 = x97 & n428 ;
  assign n1419 = ( ~n157 & n1417 ) | ( ~n157 & n1418 ) | ( n1417 & n1418 ) ;
  assign n1420 = n1419 ^ n748 ^ n559 ;
  assign n1421 = ( ~n155 & n181 ) | ( ~n155 & n1022 ) | ( n181 & n1022 ) ;
  assign n1422 = n436 ^ x102 ^ 1'b0 ;
  assign n1423 = ( n539 & n1421 ) | ( n539 & ~n1422 ) | ( n1421 & ~n1422 ) ;
  assign n1424 = n1423 ^ n233 ^ 1'b0 ;
  assign n1425 = ( n885 & n1244 ) | ( n885 & n1424 ) | ( n1244 & n1424 ) ;
  assign n1426 = n1420 & n1425 ;
  assign n1427 = ~n1416 & n1426 ;
  assign n1428 = n257 & ~n1427 ;
  assign n1429 = n628 ^ n553 ^ 1'b0 ;
  assign n1430 = n186 & n1429 ;
  assign n1431 = n1430 ^ n849 ^ 1'b0 ;
  assign n1432 = n379 | n1431 ;
  assign n1433 = n1432 ^ n1076 ^ 1'b0 ;
  assign n1434 = ( n655 & ~n1055 ) | ( n655 & n1433 ) | ( ~n1055 & n1433 ) ;
  assign n1435 = n1428 & n1434 ;
  assign n1447 = n482 ^ n254 ^ n133 ;
  assign n1443 = x105 & ~n214 ;
  assign n1444 = n1443 ^ n173 ^ 1'b0 ;
  assign n1445 = n1444 ^ n575 ^ 1'b0 ;
  assign n1436 = n514 ^ x112 ^ x107 ;
  assign n1437 = ( x76 & n994 ) | ( x76 & n1436 ) | ( n994 & n1436 ) ;
  assign n1438 = n1437 ^ n675 ^ n582 ;
  assign n1439 = n239 & ~n340 ;
  assign n1440 = n507 & n1439 ;
  assign n1441 = n1440 ^ n1147 ^ n374 ;
  assign n1442 = n1438 & n1441 ;
  assign n1446 = n1445 ^ n1442 ^ 1'b0 ;
  assign n1448 = n1447 ^ n1446 ^ x26 ;
  assign n1452 = n1291 ^ n738 ^ 1'b0 ;
  assign n1453 = n1452 ^ n1154 ^ n776 ;
  assign n1449 = n457 ^ n320 ^ n168 ;
  assign n1450 = x44 & ~n838 ;
  assign n1451 = ~n1449 & n1450 ;
  assign n1454 = n1453 ^ n1451 ^ 1'b0 ;
  assign n1455 = x81 & ~n1454 ;
  assign n1456 = n1455 ^ n873 ^ n506 ;
  assign n1457 = ( ~n775 & n1265 ) | ( ~n775 & n1456 ) | ( n1265 & n1456 ) ;
  assign n1458 = n585 ^ n432 ^ n353 ;
  assign n1459 = n947 ^ n354 ^ 1'b0 ;
  assign n1460 = n215 & n1459 ;
  assign n1461 = n434 | n1418 ;
  assign n1462 = n1461 ^ n1055 ^ 1'b0 ;
  assign n1463 = n688 | n1462 ;
  assign n1464 = n1463 ^ n783 ^ n384 ;
  assign n1465 = ( n1011 & n1460 ) | ( n1011 & ~n1464 ) | ( n1460 & ~n1464 ) ;
  assign n1466 = n1465 ^ n547 ^ n153 ;
  assign n1467 = ( n912 & n953 ) | ( n912 & n1257 ) | ( n953 & n1257 ) ;
  assign n1468 = n582 & n968 ;
  assign n1469 = ~n356 & n1468 ;
  assign n1470 = n1469 ^ n302 ^ 1'b0 ;
  assign n1471 = ( n285 & n1467 ) | ( n285 & n1470 ) | ( n1467 & n1470 ) ;
  assign n1472 = n312 ^ n305 ^ x99 ;
  assign n1473 = n1472 ^ n312 ^ 1'b0 ;
  assign n1474 = ( n511 & n809 ) | ( n511 & n1372 ) | ( n809 & n1372 ) ;
  assign n1475 = ( n1149 & n1473 ) | ( n1149 & n1474 ) | ( n1473 & n1474 ) ;
  assign n1476 = ( x108 & n786 ) | ( x108 & n902 ) | ( n786 & n902 ) ;
  assign n1477 = n1476 ^ n1242 ^ n815 ;
  assign n1480 = ( ~n149 & n172 ) | ( ~n149 & n1417 ) | ( n172 & n1417 ) ;
  assign n1478 = n406 ^ n402 ^ n167 ;
  assign n1479 = ( n148 & ~n150 ) | ( n148 & n1478 ) | ( ~n150 & n1478 ) ;
  assign n1481 = n1480 ^ n1479 ^ n798 ;
  assign n1482 = n1481 ^ n778 ^ 1'b0 ;
  assign n1483 = n748 ^ n379 ^ x43 ;
  assign n1484 = ( x78 & n145 ) | ( x78 & n146 ) | ( n145 & n146 ) ;
  assign n1485 = ( n294 & ~n677 ) | ( n294 & n1484 ) | ( ~n677 & n1484 ) ;
  assign n1486 = n809 & n1485 ;
  assign n1487 = n1486 ^ n150 ^ 1'b0 ;
  assign n1488 = n937 ^ n672 ^ n551 ;
  assign n1489 = n1487 | n1488 ;
  assign n1490 = n1483 | n1489 ;
  assign n1491 = n1490 ^ n386 ^ n141 ;
  assign n1492 = n1491 ^ n1123 ^ n239 ;
  assign n1493 = n811 ^ x79 ^ x41 ;
  assign n1494 = ( ~n616 & n1102 ) | ( ~n616 & n1463 ) | ( n1102 & n1463 ) ;
  assign n1502 = ( x30 & n428 ) | ( x30 & ~n458 ) | ( n428 & ~n458 ) ;
  assign n1503 = ( x60 & n530 ) | ( x60 & n1502 ) | ( n530 & n1502 ) ;
  assign n1504 = n1503 ^ n1257 ^ n318 ;
  assign n1499 = n497 ^ n406 ^ n329 ;
  assign n1500 = n389 | n1499 ;
  assign n1501 = n1500 ^ n366 ^ 1'b0 ;
  assign n1496 = ( n159 & ~n341 ) | ( n159 & n865 ) | ( ~n341 & n865 ) ;
  assign n1497 = n1496 ^ n1055 ^ n402 ;
  assign n1495 = ( x93 & n536 ) | ( x93 & ~n1154 ) | ( n536 & ~n1154 ) ;
  assign n1498 = n1497 ^ n1495 ^ x103 ;
  assign n1505 = n1504 ^ n1501 ^ n1498 ;
  assign n1506 = n1110 & ~n1505 ;
  assign n1507 = n397 & n1506 ;
  assign n1508 = ( n1493 & n1494 ) | ( n1493 & ~n1507 ) | ( n1494 & ~n1507 ) ;
  assign n1509 = n714 & n937 ;
  assign n1510 = ~n573 & n1509 ;
  assign n1511 = n1510 ^ n1218 ^ n1001 ;
  assign n1522 = x85 & ~n252 ;
  assign n1523 = n1522 ^ n573 ^ 1'b0 ;
  assign n1524 = n1523 ^ n1125 ^ 1'b0 ;
  assign n1525 = n975 & ~n1524 ;
  assign n1526 = ( n401 & n478 ) | ( n401 & ~n1525 ) | ( n478 & ~n1525 ) ;
  assign n1512 = n416 | n786 ;
  assign n1513 = n1512 ^ n635 ^ 1'b0 ;
  assign n1517 = n528 ^ n513 ^ n339 ;
  assign n1514 = x13 & ~n652 ;
  assign n1515 = n291 & n1514 ;
  assign n1516 = ( n177 & ~n1080 ) | ( n177 & n1515 ) | ( ~n1080 & n1515 ) ;
  assign n1518 = n1517 ^ n1516 ^ n1051 ;
  assign n1519 = n1518 ^ n998 ^ n333 ;
  assign n1520 = ( ~n654 & n968 ) | ( ~n654 & n1519 ) | ( n968 & n1519 ) ;
  assign n1521 = ( n470 & ~n1513 ) | ( n470 & n1520 ) | ( ~n1513 & n1520 ) ;
  assign n1527 = n1526 ^ n1521 ^ n1364 ;
  assign n1529 = n239 & ~n626 ;
  assign n1530 = n1529 ^ n281 ^ 1'b0 ;
  assign n1528 = n1041 ^ n717 ^ 1'b0 ;
  assign n1531 = n1530 ^ n1528 ^ n1474 ;
  assign n1536 = n707 ^ x47 ^ 1'b0 ;
  assign n1532 = n674 & n858 ;
  assign n1533 = ~n242 & n1532 ;
  assign n1534 = n1501 ^ n207 ^ 1'b0 ;
  assign n1535 = ( ~n533 & n1533 ) | ( ~n533 & n1534 ) | ( n1533 & n1534 ) ;
  assign n1537 = n1536 ^ n1535 ^ n688 ;
  assign n1538 = n334 ^ n264 ^ x88 ;
  assign n1539 = n1538 ^ n578 ^ n479 ;
  assign n1540 = n1539 ^ x126 ^ 1'b0 ;
  assign n1541 = ~n538 & n1540 ;
  assign n1551 = ( n675 & n851 ) | ( n675 & n1444 ) | ( n851 & n1444 ) ;
  assign n1542 = n586 | n825 ;
  assign n1543 = n1463 ^ n590 ^ 1'b0 ;
  assign n1544 = n1542 | n1543 ;
  assign n1545 = ( x60 & n1400 ) | ( x60 & n1544 ) | ( n1400 & n1544 ) ;
  assign n1548 = n595 & ~n1013 ;
  assign n1546 = ( n465 & n610 ) | ( n465 & ~n831 ) | ( n610 & ~n831 ) ;
  assign n1547 = x28 & n1546 ;
  assign n1549 = n1548 ^ n1547 ^ 1'b0 ;
  assign n1550 = ( n1137 & ~n1545 ) | ( n1137 & n1549 ) | ( ~n1545 & n1549 ) ;
  assign n1552 = n1551 ^ n1550 ^ n673 ;
  assign n1575 = ( n133 & ~n363 ) | ( n133 & n628 ) | ( ~n363 & n628 ) ;
  assign n1571 = x20 & ~n1061 ;
  assign n1572 = n1571 ^ n147 ^ 1'b0 ;
  assign n1565 = ( n143 & ~n233 ) | ( n143 & n332 ) | ( ~n233 & n332 ) ;
  assign n1566 = n1050 | n1565 ;
  assign n1567 = n799 & ~n1566 ;
  assign n1568 = ( x99 & n309 ) | ( x99 & ~n464 ) | ( n309 & ~n464 ) ;
  assign n1569 = n1568 ^ n1183 ^ x92 ;
  assign n1570 = ( n398 & n1567 ) | ( n398 & n1569 ) | ( n1567 & n1569 ) ;
  assign n1573 = n1572 ^ n1570 ^ n1530 ;
  assign n1574 = n1573 ^ n1211 ^ 1'b0 ;
  assign n1562 = n1116 ^ n367 ^ n220 ;
  assign n1558 = x46 & n296 ;
  assign n1559 = n1373 ^ n1012 ^ n362 ;
  assign n1560 = ( ~n851 & n1558 ) | ( ~n851 & n1559 ) | ( n1558 & n1559 ) ;
  assign n1556 = n776 ^ n454 ^ 1'b0 ;
  assign n1557 = n256 & n1556 ;
  assign n1561 = n1560 ^ n1557 ^ n1116 ;
  assign n1555 = ( n279 & n609 ) | ( n279 & ~n1383 ) | ( n609 & ~n1383 ) ;
  assign n1563 = n1562 ^ n1561 ^ n1555 ;
  assign n1553 = n664 & ~n1421 ;
  assign n1554 = n1553 ^ n352 ^ 1'b0 ;
  assign n1564 = n1563 ^ n1554 ^ 1'b0 ;
  assign n1576 = n1575 ^ n1574 ^ n1564 ;
  assign n1577 = n172 & n272 ;
  assign n1578 = n1577 ^ n935 ^ n320 ;
  assign n1579 = n1578 ^ n1395 ^ n959 ;
  assign n1580 = ( n176 & n280 ) | ( n176 & ~n393 ) | ( n280 & ~n393 ) ;
  assign n1581 = ( x47 & n768 ) | ( x47 & ~n1580 ) | ( n768 & ~n1580 ) ;
  assign n1582 = ( ~n1216 & n1453 ) | ( ~n1216 & n1581 ) | ( n1453 & n1581 ) ;
  assign n1588 = n568 ^ x58 ^ 1'b0 ;
  assign n1583 = n1137 ^ n1050 ^ 1'b0 ;
  assign n1584 = n139 | n165 ;
  assign n1585 = ( n308 & n1014 ) | ( n308 & ~n1584 ) | ( n1014 & ~n1584 ) ;
  assign n1586 = n1585 ^ n1503 ^ n401 ;
  assign n1587 = ( n1039 & ~n1583 ) | ( n1039 & n1586 ) | ( ~n1583 & n1586 ) ;
  assign n1589 = n1588 ^ n1587 ^ n605 ;
  assign n1590 = n1485 & n1589 ;
  assign n1591 = n1590 ^ n236 ^ 1'b0 ;
  assign n1594 = x30 & ~n465 ;
  assign n1595 = n186 & ~n1594 ;
  assign n1596 = n1544 & n1595 ;
  assign n1599 = n235 ^ n164 ^ 1'b0 ;
  assign n1600 = n541 | n1599 ;
  assign n1597 = n1405 ^ n655 ^ n621 ;
  assign n1598 = ( n447 & ~n697 ) | ( n447 & n1597 ) | ( ~n697 & n1597 ) ;
  assign n1601 = n1600 ^ n1598 ^ 1'b0 ;
  assign n1602 = ( n352 & n1596 ) | ( n352 & ~n1601 ) | ( n1596 & ~n1601 ) ;
  assign n1603 = n1602 ^ n1425 ^ n1181 ;
  assign n1592 = n777 ^ n460 ^ x37 ;
  assign n1593 = ( x125 & n675 ) | ( x125 & ~n1592 ) | ( n675 & ~n1592 ) ;
  assign n1604 = n1603 ^ n1593 ^ n526 ;
  assign n1605 = n187 | n1390 ;
  assign n1606 = n725 & ~n1605 ;
  assign n1607 = n1138 ^ n837 ^ n458 ;
  assign n1610 = ( n131 & ~n377 ) | ( n131 & n649 ) | ( ~n377 & n649 ) ;
  assign n1608 = n564 ^ n184 ^ 1'b0 ;
  assign n1609 = ~n1440 & n1608 ;
  assign n1611 = n1610 ^ n1609 ^ n827 ;
  assign n1612 = n1365 ^ n1280 ^ n368 ;
  assign n1613 = n838 ^ n669 ^ 1'b0 ;
  assign n1614 = n1612 | n1613 ;
  assign n1615 = n1212 ^ n383 ^ 1'b0 ;
  assign n1616 = n808 ^ n129 ^ 1'b0 ;
  assign n1617 = ~n181 & n1616 ;
  assign n1618 = ( n201 & n1424 ) | ( n201 & ~n1617 ) | ( n1424 & ~n1617 ) ;
  assign n1619 = n1618 ^ n935 ^ 1'b0 ;
  assign n1620 = n1615 | n1619 ;
  assign n1621 = ( ~n393 & n1614 ) | ( ~n393 & n1620 ) | ( n1614 & n1620 ) ;
  assign n1622 = n1167 & ~n1621 ;
  assign n1623 = n1611 & n1622 ;
  assign n1624 = n1006 & ~n1623 ;
  assign n1625 = n1607 & n1624 ;
  assign n1639 = ( n236 & n677 ) | ( n236 & ~n786 ) | ( n677 & ~n786 ) ;
  assign n1626 = ( n213 & n377 ) | ( n213 & ~n677 ) | ( n377 & ~n677 ) ;
  assign n1627 = ( ~x6 & n672 ) | ( ~x6 & n1626 ) | ( n672 & n1626 ) ;
  assign n1632 = ( n191 & n677 ) | ( n191 & n1163 ) | ( n677 & n1163 ) ;
  assign n1630 = ( ~n419 & n580 ) | ( ~n419 & n1332 ) | ( n580 & n1332 ) ;
  assign n1631 = n693 | n1630 ;
  assign n1628 = ( n209 & ~n557 ) | ( n209 & n673 ) | ( ~n557 & n673 ) ;
  assign n1629 = n1628 ^ n1626 ^ n141 ;
  assign n1633 = n1632 ^ n1631 ^ n1629 ;
  assign n1634 = ( n451 & n577 ) | ( n451 & ~n718 ) | ( n577 & ~n718 ) ;
  assign n1635 = ( n793 & ~n956 ) | ( n793 & n1634 ) | ( ~n956 & n1634 ) ;
  assign n1636 = ( n968 & n980 ) | ( n968 & ~n1635 ) | ( n980 & ~n1635 ) ;
  assign n1637 = ( n1627 & ~n1633 ) | ( n1627 & n1636 ) | ( ~n1633 & n1636 ) ;
  assign n1638 = n1637 ^ n407 ^ 1'b0 ;
  assign n1640 = n1639 ^ n1638 ^ 1'b0 ;
  assign n1641 = x99 & ~n1640 ;
  assign n1642 = ~n634 & n780 ;
  assign n1643 = n749 ^ n142 ^ 1'b0 ;
  assign n1644 = n1642 & ~n1643 ;
  assign n1645 = n1480 ^ n750 ^ n408 ;
  assign n1646 = ~n1504 & n1645 ;
  assign n1647 = ~n908 & n1646 ;
  assign n1648 = n1647 ^ n1642 ^ n1570 ;
  assign n1662 = n577 ^ n564 ^ x99 ;
  assign n1663 = ~n620 & n1662 ;
  assign n1664 = n1663 ^ n1463 ^ n834 ;
  assign n1649 = n659 ^ n519 ^ n239 ;
  assign n1651 = ~n187 & n620 ;
  assign n1652 = ~n820 & n1651 ;
  assign n1653 = ( n383 & n871 ) | ( n383 & ~n1652 ) | ( n871 & ~n1652 ) ;
  assign n1654 = n1653 ^ n998 ^ n765 ;
  assign n1655 = ( ~x58 & n559 ) | ( ~x58 & n1654 ) | ( n559 & n1654 ) ;
  assign n1650 = ~n538 & n1127 ;
  assign n1656 = n1655 ^ n1650 ^ 1'b0 ;
  assign n1657 = n484 ^ x16 ^ 1'b0 ;
  assign n1658 = n984 ^ n685 ^ n426 ;
  assign n1659 = ( n304 & n429 ) | ( n304 & ~n1658 ) | ( n429 & ~n1658 ) ;
  assign n1660 = ( n841 & ~n1657 ) | ( n841 & n1659 ) | ( ~n1657 & n1659 ) ;
  assign n1661 = ( ~n1649 & n1656 ) | ( ~n1649 & n1660 ) | ( n1656 & n1660 ) ;
  assign n1665 = n1664 ^ n1661 ^ x15 ;
  assign n1666 = x47 & n1351 ;
  assign n1667 = ~n888 & n1666 ;
  assign n1668 = n1667 ^ n1574 ^ n1147 ;
  assign n1669 = x121 & n162 ;
  assign n1670 = ( n1526 & n1668 ) | ( n1526 & ~n1669 ) | ( n1668 & ~n1669 ) ;
  assign n1671 = n693 & ~n1075 ;
  assign n1672 = n1671 ^ n1407 ^ 1'b0 ;
  assign n1673 = ~n243 & n459 ;
  assign n1674 = n1673 ^ n1020 ^ 1'b0 ;
  assign n1675 = n635 & ~n1674 ;
  assign n1678 = ( n205 & n637 ) | ( n205 & ~n947 ) | ( n637 & ~n947 ) ;
  assign n1679 = n1678 ^ n414 ^ n317 ;
  assign n1676 = x110 & ~n349 ;
  assign n1677 = n1676 ^ n391 ^ 1'b0 ;
  assign n1680 = n1679 ^ n1677 ^ n564 ;
  assign n1681 = ~n436 & n1521 ;
  assign n1682 = n1681 ^ n194 ^ 1'b0 ;
  assign n1686 = ( ~n244 & n1068 ) | ( ~n244 & n1300 ) | ( n1068 & n1300 ) ;
  assign n1683 = n1004 ^ x103 ^ 1'b0 ;
  assign n1684 = n746 & ~n1683 ;
  assign n1685 = n1684 ^ n1053 ^ n179 ;
  assign n1687 = n1686 ^ n1685 ^ n868 ;
  assign n1688 = n1658 ^ n243 ^ 1'b0 ;
  assign n1689 = n1688 ^ n1631 ^ n1003 ;
  assign n1690 = n1689 ^ n1557 ^ 1'b0 ;
  assign n1691 = n1658 ^ n1515 ^ 1'b0 ;
  assign n1692 = n1126 ^ n130 ^ 1'b0 ;
  assign n1693 = ~n1691 & n1692 ;
  assign n1694 = ( x122 & ~n170 ) | ( x122 & n611 ) | ( ~n170 & n611 ) ;
  assign n1695 = n1636 ^ n731 ^ n681 ;
  assign n1697 = n1105 ^ x22 ^ 1'b0 ;
  assign n1698 = ( x1 & x91 ) | ( x1 & n1697 ) | ( x91 & n1697 ) ;
  assign n1699 = n1698 ^ n1367 ^ n1282 ;
  assign n1696 = n168 & n1041 ;
  assign n1700 = n1699 ^ n1696 ^ 1'b0 ;
  assign n1701 = n1700 ^ n507 ^ x42 ;
  assign n1705 = n1642 ^ n882 ^ n363 ;
  assign n1703 = n1191 ^ x121 ^ x107 ;
  assign n1704 = n1703 ^ n627 ^ n575 ;
  assign n1702 = n1016 ^ n815 ^ x117 ;
  assign n1706 = n1705 ^ n1704 ^ n1702 ;
  assign n1707 = n1706 ^ n1530 ^ n745 ;
  assign n1708 = n1061 ^ n429 ^ 1'b0 ;
  assign n1709 = ( n276 & n1083 ) | ( n276 & n1339 ) | ( n1083 & n1339 ) ;
  assign n1710 = ( n628 & n669 ) | ( n628 & n1709 ) | ( n669 & n1709 ) ;
  assign n1711 = n1710 ^ n445 ^ 1'b0 ;
  assign n1712 = n1484 ^ n841 ^ n339 ;
  assign n1713 = n341 & ~n1712 ;
  assign n1716 = n707 ^ n561 ^ n242 ;
  assign n1717 = n1716 ^ n1518 ^ n948 ;
  assign n1714 = n667 ^ n228 ^ 1'b0 ;
  assign n1715 = ~n1292 & n1714 ;
  assign n1718 = n1717 ^ n1715 ^ n706 ;
  assign n1719 = ( ~n1149 & n1713 ) | ( ~n1149 & n1718 ) | ( n1713 & n1718 ) ;
  assign n1728 = n669 ^ n564 ^ n372 ;
  assign n1726 = n1373 ^ n1191 ^ x55 ;
  assign n1727 = ( ~n851 & n1198 ) | ( ~n851 & n1726 ) | ( n1198 & n1726 ) ;
  assign n1721 = n376 ^ n187 ^ n167 ;
  assign n1722 = n458 & n1721 ;
  assign n1723 = n849 & n1722 ;
  assign n1724 = n1723 ^ n1642 ^ 1'b0 ;
  assign n1720 = n1001 & n1580 ;
  assign n1725 = n1724 ^ n1720 ^ 1'b0 ;
  assign n1729 = n1728 ^ n1727 ^ n1725 ;
  assign n1730 = n743 ^ n738 ^ n240 ;
  assign n1731 = ( n1215 & n1313 ) | ( n1215 & ~n1730 ) | ( n1313 & ~n1730 ) ;
  assign n1732 = n1125 ^ n672 ^ 1'b0 ;
  assign n1733 = ~n138 & n1615 ;
  assign n1734 = n411 ^ n357 ^ n213 ;
  assign n1735 = ( ~n1523 & n1557 ) | ( ~n1523 & n1734 ) | ( n1557 & n1734 ) ;
  assign n1736 = n643 & ~n983 ;
  assign n1737 = n829 & n1596 ;
  assign n1748 = ( n176 & n195 ) | ( n176 & n317 ) | ( n195 & n317 ) ;
  assign n1749 = n1748 ^ n1332 ^ n484 ;
  assign n1745 = ( ~x59 & n429 ) | ( ~x59 & n991 ) | ( n429 & n991 ) ;
  assign n1746 = ~n397 & n1745 ;
  assign n1747 = n1746 ^ n206 ^ 1'b0 ;
  assign n1750 = n1749 ^ n1747 ^ n186 ;
  assign n1738 = n419 & n1610 ;
  assign n1739 = n1738 ^ n667 ^ 1'b0 ;
  assign n1740 = n376 & ~n1739 ;
  assign n1741 = ( n477 & ~n486 ) | ( n477 & n1211 ) | ( ~n486 & n1211 ) ;
  assign n1742 = n1741 ^ n553 ^ n362 ;
  assign n1743 = ( n197 & n1740 ) | ( n197 & n1742 ) | ( n1740 & n1742 ) ;
  assign n1744 = n1743 ^ n232 ^ n193 ;
  assign n1751 = n1750 ^ n1744 ^ n1727 ;
  assign n1752 = n567 & ~n590 ;
  assign n1753 = n1752 ^ n391 ^ n152 ;
  assign n1754 = ~n767 & n1753 ;
  assign n1755 = ~n1346 & n1754 ;
  assign n1756 = n1755 ^ n1738 ^ x0 ;
  assign n1757 = ( ~n1214 & n1632 ) | ( ~n1214 & n1756 ) | ( n1632 & n1756 ) ;
  assign n1758 = n214 | n928 ;
  assign n1759 = n260 | n1758 ;
  assign n1764 = n818 ^ n337 ^ 1'b0 ;
  assign n1765 = n231 & ~n1764 ;
  assign n1766 = n1765 ^ n1291 ^ n214 ;
  assign n1760 = ( x116 & n277 ) | ( x116 & n686 ) | ( n277 & n686 ) ;
  assign n1761 = ( n252 & n1161 ) | ( n252 & ~n1653 ) | ( n1161 & ~n1653 ) ;
  assign n1762 = n1760 & ~n1761 ;
  assign n1763 = ~x66 & n1762 ;
  assign n1767 = n1766 ^ n1763 ^ 1'b0 ;
  assign n1778 = n868 ^ n158 ^ x30 ;
  assign n1776 = ( n507 & n601 ) | ( n507 & n1273 ) | ( n601 & n1273 ) ;
  assign n1777 = ( n527 & n1538 ) | ( n527 & n1776 ) | ( n1538 & n1776 ) ;
  assign n1768 = n984 ^ n880 ^ n471 ;
  assign n1769 = n976 ^ x124 ^ 1'b0 ;
  assign n1770 = n945 & n1769 ;
  assign n1771 = n1216 ^ n163 ^ 1'b0 ;
  assign n1772 = ~n470 & n1771 ;
  assign n1773 = ( n1041 & n1545 ) | ( n1041 & ~n1632 ) | ( n1545 & ~n1632 ) ;
  assign n1774 = ( n1761 & n1772 ) | ( n1761 & ~n1773 ) | ( n1772 & ~n1773 ) ;
  assign n1775 = ( n1768 & n1770 ) | ( n1768 & ~n1774 ) | ( n1770 & ~n1774 ) ;
  assign n1779 = n1778 ^ n1777 ^ n1775 ;
  assign n1780 = n1089 ^ n586 ^ x37 ;
  assign n1781 = n541 ^ n242 ^ n139 ;
  assign n1782 = n1476 ^ n451 ^ x99 ;
  assign n1783 = ( n1780 & n1781 ) | ( n1780 & n1782 ) | ( n1781 & n1782 ) ;
  assign n1788 = n345 ^ n157 ^ x44 ;
  assign n1787 = ( n372 & n570 ) | ( n372 & ~n1480 ) | ( n570 & ~n1480 ) ;
  assign n1789 = n1788 ^ n1787 ^ n1645 ;
  assign n1784 = ~x68 & n926 ;
  assign n1785 = n1784 ^ n1352 ^ 1'b0 ;
  assign n1786 = n1592 | n1785 ;
  assign n1790 = n1789 ^ n1786 ^ n1723 ;
  assign n1791 = n1790 ^ n970 ^ n829 ;
  assign n1792 = ( n459 & ~n934 ) | ( n459 & n1022 ) | ( ~n934 & n1022 ) ;
  assign n1793 = ~n257 & n1792 ;
  assign n1794 = n1793 ^ x122 ^ 1'b0 ;
  assign n1796 = n1292 ^ n707 ^ 1'b0 ;
  assign n1795 = n368 & ~n754 ;
  assign n1797 = n1796 ^ n1795 ^ 1'b0 ;
  assign n1798 = n1286 ^ n678 ^ 1'b0 ;
  assign n1800 = ( ~x94 & x99 ) | ( ~x94 & n472 ) | ( x99 & n472 ) ;
  assign n1799 = n1430 ^ n1022 ^ n735 ;
  assign n1801 = n1800 ^ n1799 ^ n512 ;
  assign n1802 = ( ~x113 & n1089 ) | ( ~x113 & n1801 ) | ( n1089 & n1801 ) ;
  assign n1803 = n1798 & ~n1802 ;
  assign n1804 = n1259 ^ n882 ^ n453 ;
  assign n1805 = ( ~n323 & n857 ) | ( ~n323 & n877 ) | ( n857 & n877 ) ;
  assign n1806 = ( n488 & n1577 ) | ( n488 & n1805 ) | ( n1577 & n1805 ) ;
  assign n1807 = n908 ^ n517 ^ x48 ;
  assign n1808 = n429 & n623 ;
  assign n1809 = n693 & ~n1808 ;
  assign n1810 = ~x54 & n1809 ;
  assign n1811 = n852 | n1810 ;
  assign n1812 = n500 & ~n1811 ;
  assign n1813 = ( n877 & n1658 ) | ( n877 & n1812 ) | ( n1658 & n1812 ) ;
  assign n1814 = ( n335 & n445 ) | ( n335 & n1813 ) | ( n445 & n1813 ) ;
  assign n1815 = n1807 & n1814 ;
  assign n1816 = n1815 ^ n1684 ^ 1'b0 ;
  assign n1817 = n849 | n1816 ;
  assign n1818 = n1806 & ~n1817 ;
  assign n1819 = n823 | n1818 ;
  assign n1820 = n1804 | n1819 ;
  assign n1829 = n1117 | n1324 ;
  assign n1824 = n141 & ~n161 ;
  assign n1825 = ~x14 & n1824 ;
  assign n1826 = ( x106 & n816 ) | ( x106 & ~n1721 ) | ( n816 & ~n1721 ) ;
  assign n1827 = ( n264 & n567 ) | ( n264 & n819 ) | ( n567 & n819 ) ;
  assign n1828 = ( n1825 & ~n1826 ) | ( n1825 & n1827 ) | ( ~n1826 & n1827 ) ;
  assign n1822 = n1211 ^ x57 ^ 1'b0 ;
  assign n1821 = ( x59 & n428 ) | ( x59 & n987 ) | ( n428 & n987 ) ;
  assign n1823 = n1822 ^ n1821 ^ n483 ;
  assign n1830 = n1829 ^ n1828 ^ n1823 ;
  assign n1834 = n1032 ^ n830 ^ 1'b0 ;
  assign n1835 = n1063 ^ n977 ^ n931 ;
  assign n1836 = ~n498 & n1835 ;
  assign n1837 = ( n293 & n1834 ) | ( n293 & ~n1836 ) | ( n1834 & ~n1836 ) ;
  assign n1838 = n804 & n1837 ;
  assign n1831 = ( n771 & n1480 ) | ( n771 & n1612 ) | ( n1480 & n1612 ) ;
  assign n1832 = n1831 ^ n285 ^ 1'b0 ;
  assign n1833 = n390 & ~n1832 ;
  assign n1839 = n1838 ^ n1833 ^ 1'b0 ;
  assign n1840 = n212 | n1839 ;
  assign n1841 = ( n196 & ~n1830 ) | ( n196 & n1840 ) | ( ~n1830 & n1840 ) ;
  assign n1842 = n680 ^ n198 ^ x71 ;
  assign n1843 = n1659 & n1842 ;
  assign n1844 = ~n1546 & n1843 ;
  assign n1846 = n1020 & n1745 ;
  assign n1847 = n1822 & n1846 ;
  assign n1845 = ~n652 & n873 ;
  assign n1848 = n1847 ^ n1845 ^ 1'b0 ;
  assign n1849 = n1848 ^ n653 ^ n314 ;
  assign n1850 = ( n933 & n1216 ) | ( n933 & n1849 ) | ( n1216 & n1849 ) ;
  assign n1865 = n638 ^ n264 ^ n247 ;
  assign n1859 = n728 & ~n1743 ;
  assign n1860 = ~n346 & n1859 ;
  assign n1861 = ( ~n469 & n1198 ) | ( ~n469 & n1860 ) | ( n1198 & n1860 ) ;
  assign n1862 = n302 & ~n398 ;
  assign n1863 = n1862 ^ n856 ^ n543 ;
  assign n1864 = ( n1166 & n1861 ) | ( n1166 & n1863 ) | ( n1861 & n1863 ) ;
  assign n1857 = ( x127 & n336 ) | ( x127 & n1308 ) | ( n336 & n1308 ) ;
  assign n1855 = n614 ^ n411 ^ n295 ;
  assign n1856 = n1855 ^ n1493 ^ x100 ;
  assign n1851 = n465 & ~n759 ;
  assign n1852 = n1851 ^ n639 ^ 1'b0 ;
  assign n1853 = n1852 ^ n1635 ^ n379 ;
  assign n1854 = ( n471 & n1161 ) | ( n471 & n1853 ) | ( n1161 & n1853 ) ;
  assign n1858 = n1857 ^ n1856 ^ n1854 ;
  assign n1866 = n1865 ^ n1864 ^ n1858 ;
  assign n1869 = ( n566 & n899 ) | ( n566 & n1164 ) | ( n899 & n1164 ) ;
  assign n1867 = ( x127 & n559 ) | ( x127 & n1334 ) | ( n559 & n1334 ) ;
  assign n1868 = ( n1499 & n1539 ) | ( n1499 & ~n1867 ) | ( n1539 & ~n1867 ) ;
  assign n1870 = n1869 ^ n1868 ^ n1797 ;
  assign n1871 = ( ~n165 & n219 ) | ( ~n165 & n841 ) | ( n219 & n841 ) ;
  assign n1872 = n742 & n1536 ;
  assign n1873 = ( n528 & n768 ) | ( n528 & n1872 ) | ( n768 & n1872 ) ;
  assign n1874 = n1161 ^ n669 ^ 1'b0 ;
  assign n1875 = n1822 ^ n947 ^ n569 ;
  assign n1876 = ( n671 & ~n728 ) | ( n671 & n1875 ) | ( ~n728 & n1875 ) ;
  assign n1877 = n1863 | n1876 ;
  assign n1878 = n1874 | n1877 ;
  assign n1879 = ~n978 & n1878 ;
  assign n1896 = n731 ^ n441 ^ n130 ;
  assign n1894 = n698 ^ n457 ^ x104 ;
  assign n1895 = n1894 ^ n223 ^ 1'b0 ;
  assign n1897 = n1896 ^ n1895 ^ n1172 ;
  assign n1891 = n362 & n1066 ;
  assign n1892 = n1891 ^ x18 ^ 1'b0 ;
  assign n1890 = n609 ^ n578 ^ x21 ;
  assign n1893 = n1892 ^ n1890 ^ n714 ;
  assign n1886 = n623 ^ x116 ^ x115 ;
  assign n1887 = ~n1726 & n1886 ;
  assign n1888 = n1887 ^ n1463 ^ x49 ;
  assign n1880 = n994 ^ n578 ^ n407 ;
  assign n1881 = n958 ^ n357 ^ 1'b0 ;
  assign n1882 = n1880 & n1881 ;
  assign n1883 = n846 ^ n445 ^ n208 ;
  assign n1884 = ( n472 & n1882 ) | ( n472 & n1883 ) | ( n1882 & n1883 ) ;
  assign n1885 = n341 | n1884 ;
  assign n1889 = n1888 ^ n1885 ^ 1'b0 ;
  assign n1898 = n1897 ^ n1893 ^ n1889 ;
  assign n1899 = x124 & ~n309 ;
  assign n1900 = n1899 ^ n160 ^ 1'b0 ;
  assign n1901 = n1898 | n1900 ;
  assign n1910 = ( x124 & n554 ) | ( x124 & n1087 ) | ( n554 & n1087 ) ;
  assign n1911 = ( n306 & n1149 ) | ( n306 & ~n1910 ) | ( n1149 & ~n1910 ) ;
  assign n1912 = n1911 ^ n1864 ^ n1231 ;
  assign n1904 = n867 ^ x94 ^ x53 ;
  assign n1905 = n1904 ^ n964 ^ 1'b0 ;
  assign n1906 = n426 & n1905 ;
  assign n1907 = n1906 ^ n294 ^ n256 ;
  assign n1908 = ( n1027 & n1441 ) | ( n1027 & ~n1907 ) | ( n1441 & ~n1907 ) ;
  assign n1902 = n468 ^ n445 ^ n138 ;
  assign n1903 = n1902 ^ n1174 ^ n661 ;
  assign n1909 = n1908 ^ n1903 ^ n589 ;
  assign n1913 = n1912 ^ n1909 ^ n776 ;
  assign n1914 = n1324 ^ n326 ^ 1'b0 ;
  assign n1915 = n346 & ~n1869 ;
  assign n1916 = n1914 & n1915 ;
  assign n1920 = ( n1182 & n1749 ) | ( n1182 & n1880 ) | ( n1749 & n1880 ) ;
  assign n1921 = ( n810 & n1530 ) | ( n810 & n1920 ) | ( n1530 & n1920 ) ;
  assign n1917 = ( ~n251 & n649 ) | ( ~n251 & n1863 ) | ( n649 & n1863 ) ;
  assign n1918 = ( n1095 & ~n1612 ) | ( n1095 & n1917 ) | ( ~n1612 & n1917 ) ;
  assign n1919 = n1918 ^ n1633 ^ n357 ;
  assign n1922 = n1921 ^ n1919 ^ 1'b0 ;
  assign n1925 = n1717 ^ n719 ^ n185 ;
  assign n1923 = n1346 ^ n782 ^ x22 ;
  assign n1924 = n1923 ^ n435 ^ n427 ;
  assign n1926 = n1925 ^ n1924 ^ n1079 ;
  assign n1927 = ( n197 & ~n273 ) | ( n197 & n1179 ) | ( ~n273 & n1179 ) ;
  assign n1928 = ( ~n379 & n1558 ) | ( ~n379 & n1927 ) | ( n1558 & n1927 ) ;
  assign n1929 = n1928 ^ n1108 ^ n183 ;
  assign n1930 = ( ~n197 & n778 ) | ( ~n197 & n1929 ) | ( n778 & n1929 ) ;
  assign n1931 = n1205 ^ n581 ^ 1'b0 ;
  assign n1932 = n438 & ~n1931 ;
  assign n1933 = ( n251 & ~n497 ) | ( n251 & n1932 ) | ( ~n497 & n1932 ) ;
  assign n1934 = n500 & n1032 ;
  assign n1935 = ~n676 & n783 ;
  assign n1936 = ~n1484 & n1935 ;
  assign n1937 = n464 ^ n281 ^ 1'b0 ;
  assign n1938 = ( n1302 & n1936 ) | ( n1302 & n1937 ) | ( n1936 & n1937 ) ;
  assign n1939 = n470 & ~n738 ;
  assign n1940 = n1455 & n1939 ;
  assign n1941 = ( n1114 & n1938 ) | ( n1114 & ~n1940 ) | ( n1938 & ~n1940 ) ;
  assign n1942 = n1941 ^ n898 ^ n444 ;
  assign n1943 = n1942 ^ n1022 ^ 1'b0 ;
  assign n1944 = n1934 & ~n1943 ;
  assign n1945 = n140 & n749 ;
  assign n1946 = ~n364 & n1945 ;
  assign n1947 = n456 & ~n1946 ;
  assign n1948 = ~n864 & n1947 ;
  assign n1950 = ( n213 & ~n222 ) | ( n213 & n627 ) | ( ~n222 & n627 ) ;
  assign n1949 = n1131 ^ n689 ^ n353 ;
  assign n1951 = n1950 ^ n1949 ^ 1'b0 ;
  assign n1952 = n1787 | n1951 ;
  assign n1953 = n1027 ^ n1020 ^ 1'b0 ;
  assign n1954 = n354 | n1953 ;
  assign n1955 = x121 ^ x104 ^ 1'b0 ;
  assign n1956 = ( ~n424 & n1954 ) | ( ~n424 & n1955 ) | ( n1954 & n1955 ) ;
  assign n1960 = n318 | n921 ;
  assign n1957 = ( n202 & n216 ) | ( n202 & ~n419 ) | ( n216 & ~n419 ) ;
  assign n1958 = ( n689 & n1037 ) | ( n689 & n1957 ) | ( n1037 & n1957 ) ;
  assign n1959 = n1958 ^ n1071 ^ n528 ;
  assign n1961 = n1960 ^ n1959 ^ 1'b0 ;
  assign n1962 = ( n470 & n1017 ) | ( n470 & n1961 ) | ( n1017 & n1961 ) ;
  assign n1963 = n1848 ^ n881 ^ 1'b0 ;
  assign n1964 = n1780 & n1963 ;
  assign n1965 = ( x4 & n1122 ) | ( x4 & ~n1964 ) | ( n1122 & ~n1964 ) ;
  assign n1966 = ( n245 & n1198 ) | ( n245 & ~n1327 ) | ( n1198 & ~n1327 ) ;
  assign n1967 = ( n1962 & n1965 ) | ( n1962 & n1966 ) | ( n1965 & n1966 ) ;
  assign n1968 = ( n1952 & n1956 ) | ( n1952 & ~n1967 ) | ( n1956 & ~n1967 ) ;
  assign n1969 = ( n591 & ~n742 ) | ( n591 & n820 ) | ( ~n742 & n820 ) ;
  assign n1970 = n1161 ^ x43 ^ 1'b0 ;
  assign n1971 = ( ~n1055 & n1969 ) | ( ~n1055 & n1970 ) | ( n1969 & n1970 ) ;
  assign n1972 = ( x84 & n1016 ) | ( x84 & ~n1496 ) | ( n1016 & ~n1496 ) ;
  assign n1973 = n1972 ^ n1862 ^ n545 ;
  assign n1974 = ( n624 & n1971 ) | ( n624 & ~n1973 ) | ( n1971 & ~n1973 ) ;
  assign n1975 = n762 & n1974 ;
  assign n1976 = n498 & n1975 ;
  assign n1977 = n915 & ~n1976 ;
  assign n1978 = n1760 ^ n1493 ^ n573 ;
  assign n1979 = ( n372 & n404 ) | ( n372 & ~n1978 ) | ( n404 & ~n1978 ) ;
  assign n1983 = ( x37 & n293 ) | ( x37 & n1050 ) | ( n293 & n1050 ) ;
  assign n1980 = ( x40 & ~n270 ) | ( x40 & n296 ) | ( ~n270 & n296 ) ;
  assign n1981 = ( x82 & n258 ) | ( x82 & ~n1120 ) | ( n258 & ~n1120 ) ;
  assign n1982 = ( n1446 & n1980 ) | ( n1446 & n1981 ) | ( n1980 & n1981 ) ;
  assign n1984 = n1983 ^ n1982 ^ n1541 ;
  assign n1985 = ( x13 & n1222 ) | ( x13 & n1984 ) | ( n1222 & n1984 ) ;
  assign n1991 = n505 & n1536 ;
  assign n1988 = ( n627 & n1138 ) | ( n627 & n1161 ) | ( n1138 & n1161 ) ;
  assign n1986 = n1617 ^ n528 ^ 1'b0 ;
  assign n1987 = n399 & n1986 ;
  assign n1989 = n1988 ^ n1987 ^ 1'b0 ;
  assign n1990 = n211 | n1989 ;
  assign n1992 = n1991 ^ n1990 ^ 1'b0 ;
  assign n1994 = n1577 ^ n573 ^ n196 ;
  assign n1993 = x60 & ~n733 ;
  assign n1995 = n1994 ^ n1993 ^ 1'b0 ;
  assign n1996 = n1995 ^ n1214 ^ n596 ;
  assign n1997 = n1996 ^ n1869 ^ n1810 ;
  assign n1998 = n964 ^ n759 ^ n249 ;
  assign n1999 = n1998 ^ n728 ^ 1'b0 ;
  assign n2006 = n533 | n1493 ;
  assign n2000 = ( ~x3 & x45 ) | ( ~x3 & x95 ) | ( x45 & x95 ) ;
  assign n2001 = ~n388 & n528 ;
  assign n2002 = ~n819 & n2001 ;
  assign n2003 = n163 & ~n2002 ;
  assign n2004 = n2003 ^ n1211 ^ 1'b0 ;
  assign n2005 = n2000 & n2004 ;
  assign n2007 = n2006 ^ n2005 ^ 1'b0 ;
  assign n2010 = ( n140 & n166 ) | ( n140 & n218 ) | ( n166 & n218 ) ;
  assign n2011 = ( n247 & n1743 ) | ( n247 & n2010 ) | ( n1743 & n2010 ) ;
  assign n2008 = n388 ^ n140 ^ x58 ;
  assign n2009 = n2008 ^ n1280 ^ n532 ;
  assign n2012 = n2011 ^ n2009 ^ n401 ;
  assign n2013 = n2012 ^ n1531 ^ n329 ;
  assign n2015 = n878 ^ n810 ^ 1'b0 ;
  assign n2016 = n1084 ^ n499 ^ n464 ;
  assign n2017 = ( n975 & n2015 ) | ( n975 & ~n2016 ) | ( n2015 & ~n2016 ) ;
  assign n2018 = n2017 ^ n1874 ^ 1'b0 ;
  assign n2014 = n287 & n306 ;
  assign n2019 = n2018 ^ n2014 ^ 1'b0 ;
  assign n2022 = ( n153 & n1612 ) | ( n153 & ~n1855 ) | ( n1612 & ~n1855 ) ;
  assign n2020 = ( x51 & n168 ) | ( x51 & ~n765 ) | ( n168 & ~n765 ) ;
  assign n2021 = n2020 ^ n454 ^ x8 ;
  assign n2023 = n2022 ^ n2021 ^ 1'b0 ;
  assign n2024 = n1412 ^ x102 ^ 1'b0 ;
  assign n2025 = ( ~n1272 & n1517 ) | ( ~n1272 & n1741 ) | ( n1517 & n1741 ) ;
  assign n2026 = ( ~n142 & n1420 ) | ( ~n142 & n2025 ) | ( n1420 & n2025 ) ;
  assign n2027 = n2024 & n2026 ;
  assign n2028 = n778 ^ n704 ^ 1'b0 ;
  assign n2029 = n1575 & ~n2028 ;
  assign n2030 = n2029 ^ n2000 ^ n1072 ;
  assign n2038 = n944 ^ n706 ^ 1'b0 ;
  assign n2031 = n209 & n1195 ;
  assign n2032 = n2031 ^ x8 ^ 1'b0 ;
  assign n2033 = n1801 ^ n750 ^ x93 ;
  assign n2034 = ~n1805 & n2033 ;
  assign n2035 = n1890 & ~n2034 ;
  assign n2036 = n2035 ^ n1383 ^ 1'b0 ;
  assign n2037 = ( n2012 & ~n2032 ) | ( n2012 & n2036 ) | ( ~n2032 & n2036 ) ;
  assign n2039 = n2038 ^ n2037 ^ n719 ;
  assign n2040 = n1034 ^ n823 ^ 1'b0 ;
  assign n2041 = n2000 ^ n1678 ^ n686 ;
  assign n2042 = n2041 ^ n1336 ^ n539 ;
  assign n2043 = ( ~n1294 & n2040 ) | ( ~n1294 & n2042 ) | ( n2040 & n2042 ) ;
  assign n2044 = n1880 ^ n599 ^ 1'b0 ;
  assign n2045 = ( n701 & n2043 ) | ( n701 & n2044 ) | ( n2043 & n2044 ) ;
  assign n2046 = ( n658 & n1041 ) | ( n658 & ~n1906 ) | ( n1041 & ~n1906 ) ;
  assign n2047 = ( n436 & n1743 ) | ( n436 & n2046 ) | ( n1743 & n2046 ) ;
  assign n2048 = n370 | n1044 ;
  assign n2049 = n1768 | n2048 ;
  assign n2050 = n1288 ^ n337 ^ n170 ;
  assign n2051 = ( n1181 & n2049 ) | ( n1181 & ~n2050 ) | ( n2049 & ~n2050 ) ;
  assign n2052 = n863 & ~n2051 ;
  assign n2053 = n2047 & n2052 ;
  assign n2054 = n315 ^ n235 ^ 1'b0 ;
  assign n2055 = n2054 ^ n1038 ^ x110 ;
  assign n2056 = n2055 ^ n1936 ^ n756 ;
  assign n2057 = ~n972 & n2056 ;
  assign n2058 = ~n1210 & n2057 ;
  assign n2059 = n731 & n1772 ;
  assign n2060 = ~n453 & n2059 ;
  assign n2061 = ( n1246 & ~n1247 ) | ( n1246 & n2060 ) | ( ~n1247 & n2060 ) ;
  assign n2062 = n688 ^ n272 ^ x95 ;
  assign n2063 = ~n1265 & n2062 ;
  assign n2064 = ~n1351 & n2063 ;
  assign n2065 = ( n270 & n2061 ) | ( n270 & ~n2064 ) | ( n2061 & ~n2064 ) ;
  assign n2066 = n1801 ^ n678 ^ 1'b0 ;
  assign n2067 = n2066 ^ n560 ^ 1'b0 ;
  assign n2068 = ~n1212 & n2067 ;
  assign n2069 = ( n977 & ~n985 ) | ( n977 & n1523 ) | ( ~n985 & n1523 ) ;
  assign n2070 = n2069 ^ n1875 ^ n612 ;
  assign n2071 = ( n2065 & ~n2068 ) | ( n2065 & n2070 ) | ( ~n2068 & n2070 ) ;
  assign n2074 = ( n211 & ~n232 ) | ( n211 & n386 ) | ( ~n232 & n386 ) ;
  assign n2072 = n1405 ^ n609 ^ 1'b0 ;
  assign n2073 = x25 & n2072 ;
  assign n2075 = n2074 ^ n2073 ^ n1515 ;
  assign n2076 = ( n553 & ~n1510 ) | ( n553 & n1664 ) | ( ~n1510 & n1664 ) ;
  assign n2077 = ( ~n1030 & n1562 ) | ( ~n1030 & n2076 ) | ( n1562 & n2076 ) ;
  assign n2078 = n2077 ^ n1038 ^ n623 ;
  assign n2079 = ( ~n413 & n745 ) | ( ~n413 & n1022 ) | ( n745 & n1022 ) ;
  assign n2080 = ~n1562 & n2079 ;
  assign n2081 = n2078 & n2080 ;
  assign n2082 = n735 & n1880 ;
  assign n2083 = ~n381 & n2082 ;
  assign n2086 = n676 ^ n591 ^ n202 ;
  assign n2084 = ( n675 & n834 ) | ( n675 & ~n1865 ) | ( n834 & ~n1865 ) ;
  assign n2085 = ( n312 & n654 ) | ( n312 & n2084 ) | ( n654 & n2084 ) ;
  assign n2087 = n2086 ^ n2085 ^ 1'b0 ;
  assign n2089 = ( n158 & ~n310 ) | ( n158 & n422 ) | ( ~n310 & n422 ) ;
  assign n2088 = ( x83 & n720 ) | ( x83 & ~n896 ) | ( n720 & ~n896 ) ;
  assign n2090 = n2089 ^ n2088 ^ n1451 ;
  assign n2091 = ( n645 & n729 ) | ( n645 & ~n915 ) | ( n729 & ~n915 ) ;
  assign n2092 = ( n279 & n1575 ) | ( n279 & ~n1896 ) | ( n1575 & ~n1896 ) ;
  assign n2093 = n576 & n2092 ;
  assign n2094 = n1485 & ~n2093 ;
  assign n2095 = ( n229 & ~n417 ) | ( n229 & n2094 ) | ( ~n417 & n2094 ) ;
  assign n2096 = n2095 ^ n833 ^ n337 ;
  assign n2097 = n1391 & n2096 ;
  assign n2098 = ~n2091 & n2097 ;
  assign n2099 = n2090 & ~n2098 ;
  assign n2100 = n2087 & n2099 ;
  assign n2101 = n1334 ^ n354 ^ 1'b0 ;
  assign n2102 = n1304 ^ n1071 ^ n851 ;
  assign n2103 = n2101 & n2102 ;
  assign n2104 = ( x120 & n728 ) | ( x120 & n2103 ) | ( n728 & n2103 ) ;
  assign n2105 = n2002 ^ n932 ^ 1'b0 ;
  assign n2106 = n1048 ^ n846 ^ n457 ;
  assign n2107 = ( n710 & n2105 ) | ( n710 & ~n2106 ) | ( n2105 & ~n2106 ) ;
  assign n2108 = n2107 ^ n545 ^ n470 ;
  assign n2109 = n478 & n2108 ;
  assign n2110 = ~n1887 & n2109 ;
  assign n2112 = ( n1284 & n1390 ) | ( n1284 & n1982 ) | ( n1390 & n1982 ) ;
  assign n2111 = n1515 | n1731 ;
  assign n2113 = n2112 ^ n2111 ^ 1'b0 ;
  assign n2122 = n556 | n1483 ;
  assign n2123 = ( n173 & ~n637 ) | ( n173 & n2122 ) | ( ~n637 & n2122 ) ;
  assign n2119 = ( ~x74 & n461 ) | ( ~x74 & n1422 ) | ( n461 & n1422 ) ;
  assign n2114 = ( ~x64 & n400 ) | ( ~x64 & n533 ) | ( n400 & n533 ) ;
  assign n2115 = ( x104 & n258 ) | ( x104 & n1314 ) | ( n258 & n1314 ) ;
  assign n2116 = x90 & ~n1217 ;
  assign n2117 = ( n1194 & ~n2115 ) | ( n1194 & n2116 ) | ( ~n2115 & n2116 ) ;
  assign n2118 = ~n2114 & n2117 ;
  assign n2120 = n2119 ^ n2118 ^ n989 ;
  assign n2121 = ( n129 & n251 ) | ( n129 & n2120 ) | ( n251 & n2120 ) ;
  assign n2124 = n2123 ^ n2121 ^ n654 ;
  assign n2140 = n1163 ^ n865 ^ n194 ;
  assign n2141 = n406 & n465 ;
  assign n2142 = n2140 & n2141 ;
  assign n2126 = n509 & ~n860 ;
  assign n2127 = n2126 ^ n1292 ^ 1'b0 ;
  assign n2128 = ( x80 & x108 ) | ( x80 & ~n2127 ) | ( x108 & ~n2127 ) ;
  assign n2129 = ( ~n205 & n628 ) | ( ~n205 & n2128 ) | ( n628 & n2128 ) ;
  assign n2130 = n911 & ~n1523 ;
  assign n2131 = n2090 ^ n667 ^ n474 ;
  assign n2132 = n805 ^ n636 ^ 1'b0 ;
  assign n2133 = n597 ^ n579 ^ 1'b0 ;
  assign n2134 = ~n2132 & n2133 ;
  assign n2135 = ( x39 & n1198 ) | ( x39 & n2134 ) | ( n1198 & n2134 ) ;
  assign n2136 = ( n1961 & ~n2131 ) | ( n1961 & n2135 ) | ( ~n2131 & n2135 ) ;
  assign n2137 = ( n2128 & n2130 ) | ( n2128 & n2136 ) | ( n2130 & n2136 ) ;
  assign n2138 = ( n980 & n2129 ) | ( n980 & ~n2137 ) | ( n2129 & ~n2137 ) ;
  assign n2125 = n629 & n714 ;
  assign n2139 = n2138 ^ n2125 ^ 1'b0 ;
  assign n2143 = n2142 ^ n2139 ^ 1'b0 ;
  assign n2144 = ( n149 & n528 ) | ( n149 & n856 ) | ( n528 & n856 ) ;
  assign n2145 = ( n372 & ~n1134 ) | ( n372 & n1380 ) | ( ~n1134 & n1380 ) ;
  assign n2146 = n612 | n964 ;
  assign n2147 = ~n1320 & n2146 ;
  assign n2148 = n1337 & ~n2147 ;
  assign n2149 = n2148 ^ n538 ^ 1'b0 ;
  assign n2150 = ( ~n1496 & n1941 ) | ( ~n1496 & n2149 ) | ( n1941 & n2149 ) ;
  assign n2151 = ( n1567 & n2145 ) | ( n1567 & n2150 ) | ( n2145 & n2150 ) ;
  assign n2152 = ( ~n172 & n2144 ) | ( ~n172 & n2151 ) | ( n2144 & n2151 ) ;
  assign n2153 = n933 ^ n756 ^ 1'b0 ;
  assign n2154 = ( n992 & ~n1810 ) | ( n992 & n1818 ) | ( ~n1810 & n1818 ) ;
  assign n2155 = n638 & n1066 ;
  assign n2156 = n2155 ^ n1662 ^ 1'b0 ;
  assign n2157 = n2156 ^ n832 ^ n780 ;
  assign n2158 = ( n281 & n1402 ) | ( n281 & ~n2157 ) | ( n1402 & ~n2157 ) ;
  assign n2159 = n2158 ^ n129 ^ 1'b0 ;
  assign n2160 = n272 & n2159 ;
  assign n2161 = n941 ^ n312 ^ n220 ;
  assign n2162 = n868 | n2161 ;
  assign n2163 = n2162 ^ n810 ^ 1'b0 ;
  assign n2164 = ( ~x8 & n2160 ) | ( ~x8 & n2163 ) | ( n2160 & n2163 ) ;
  assign n2165 = n1897 ^ n1895 ^ n243 ;
  assign n2166 = ~n188 & n2165 ;
  assign n2167 = ~n131 & n2166 ;
  assign n2168 = ( n674 & ~n2140 ) | ( n674 & n2167 ) | ( ~n2140 & n2167 ) ;
  assign n2169 = n1142 ^ n460 ^ 1'b0 ;
  assign n2176 = n1065 ^ n955 ^ 1'b0 ;
  assign n2177 = x108 & ~n2176 ;
  assign n2175 = n1371 ^ n1310 ^ n272 ;
  assign n2170 = n1294 ^ n896 ^ n474 ;
  assign n2171 = ( ~n191 & n197 ) | ( ~n191 & n1083 ) | ( n197 & n1083 ) ;
  assign n2172 = n573 ^ n421 ^ n389 ;
  assign n2173 = ( n761 & n1972 ) | ( n761 & n2172 ) | ( n1972 & n2172 ) ;
  assign n2174 = ( ~n2170 & n2171 ) | ( ~n2170 & n2173 ) | ( n2171 & n2173 ) ;
  assign n2178 = n2177 ^ n2175 ^ n2174 ;
  assign n2179 = ( n1036 & n2042 ) | ( n1036 & n2178 ) | ( n2042 & n2178 ) ;
  assign n2180 = n980 ^ x127 ^ 1'b0 ;
  assign n2181 = ~n149 & n2180 ;
  assign n2182 = ( ~n457 & n1718 ) | ( ~n457 & n2181 ) | ( n1718 & n2181 ) ;
  assign n2190 = n681 ^ n422 ^ n397 ;
  assign n2184 = ~n341 & n649 ;
  assign n2185 = n2184 ^ n388 ^ 1'b0 ;
  assign n2186 = ( n1065 & n1483 ) | ( n1065 & n1787 ) | ( n1483 & n1787 ) ;
  assign n2187 = n1175 ^ n364 ^ 1'b0 ;
  assign n2188 = n1047 & ~n2187 ;
  assign n2189 = ( n2185 & n2186 ) | ( n2185 & n2188 ) | ( n2186 & n2188 ) ;
  assign n2183 = n951 ^ n364 ^ 1'b0 ;
  assign n2191 = n2190 ^ n2189 ^ n2183 ;
  assign n2192 = n477 ^ x13 ^ 1'b0 ;
  assign n2193 = n863 & ~n2192 ;
  assign n2194 = x55 & n2193 ;
  assign n2195 = n2191 & n2194 ;
  assign n2196 = ( n966 & ~n1417 ) | ( n966 & n1424 ) | ( ~n1417 & n1424 ) ;
  assign n2197 = n2196 ^ n398 ^ 1'b0 ;
  assign n2198 = n505 | n2197 ;
  assign n2199 = n165 | n1196 ;
  assign n2200 = n2199 ^ n936 ^ 1'b0 ;
  assign n2201 = ( ~n1052 & n1287 ) | ( ~n1052 & n2200 ) | ( n1287 & n2200 ) ;
  assign n2202 = ( ~n237 & n2023 ) | ( ~n237 & n2201 ) | ( n2023 & n2201 ) ;
  assign n2203 = n245 & ~n1141 ;
  assign n2204 = n2203 ^ n706 ^ n427 ;
  assign n2205 = ( n805 & n1703 ) | ( n805 & ~n2204 ) | ( n1703 & ~n2204 ) ;
  assign n2206 = n1249 ^ n1049 ^ n788 ;
  assign n2207 = n1391 & n1684 ;
  assign n2208 = ( n496 & n2206 ) | ( n496 & ~n2207 ) | ( n2206 & ~n2207 ) ;
  assign n2215 = n803 ^ n281 ^ n191 ;
  assign n2216 = n2215 ^ n585 ^ n158 ;
  assign n2217 = n772 ^ n266 ^ n239 ;
  assign n2218 = n2217 ^ n1642 ^ n215 ;
  assign n2219 = n2218 ^ n1813 ^ 1'b0 ;
  assign n2220 = n2216 | n2219 ;
  assign n2221 = n502 & n1001 ;
  assign n2222 = n2221 ^ n1772 ^ 1'b0 ;
  assign n2223 = n2220 | n2222 ;
  assign n2224 = n1207 | n2223 ;
  assign n2212 = ( n146 & n279 ) | ( n146 & n996 ) | ( n279 & n996 ) ;
  assign n2209 = n1363 ^ n1244 ^ n231 ;
  assign n2210 = ~x91 & n2209 ;
  assign n2211 = n2210 ^ n1069 ^ n658 ;
  assign n2213 = n2212 ^ n2211 ^ 1'b0 ;
  assign n2214 = n1328 | n2213 ;
  assign n2225 = n2224 ^ n2214 ^ 1'b0 ;
  assign n2229 = ( x13 & n1401 ) | ( x13 & n1755 ) | ( n1401 & n1755 ) ;
  assign n2226 = ( x9 & ~n1015 ) | ( x9 & n1588 ) | ( ~n1015 & n1588 ) ;
  assign n2227 = n2226 ^ x103 ^ 1'b0 ;
  assign n2228 = ~n1491 & n2227 ;
  assign n2230 = n2229 ^ n2228 ^ n1276 ;
  assign n2233 = ( n480 & n728 ) | ( n480 & n1488 ) | ( n728 & n1488 ) ;
  assign n2234 = n2233 ^ n1048 ^ 1'b0 ;
  assign n2231 = ( ~n388 & n390 ) | ( ~n388 & n790 ) | ( n390 & n790 ) ;
  assign n2232 = n2231 ^ n1479 ^ n198 ;
  assign n2235 = n2234 ^ n2232 ^ n577 ;
  assign n2236 = ( ~n479 & n1052 ) | ( ~n479 & n2235 ) | ( n1052 & n2235 ) ;
  assign n2237 = ( ~x2 & x62 ) | ( ~x2 & n1012 ) | ( x62 & n1012 ) ;
  assign n2238 = ( ~n2056 & n2069 ) | ( ~n2056 & n2237 ) | ( n2069 & n2237 ) ;
  assign n2239 = n1127 ^ n809 ^ n224 ;
  assign n2240 = n570 ^ n473 ^ n421 ;
  assign n2241 = n362 & ~n404 ;
  assign n2242 = n1280 ^ n818 ^ n416 ;
  assign n2243 = n840 & ~n2242 ;
  assign n2244 = n1860 & n2243 ;
  assign n2245 = ( n708 & n1515 ) | ( n708 & ~n2244 ) | ( n1515 & ~n2244 ) ;
  assign n2246 = n2245 ^ n914 ^ 1'b0 ;
  assign n2247 = ~n1611 & n2246 ;
  assign n2248 = n2241 & n2247 ;
  assign n2249 = ( n421 & n805 ) | ( n421 & ~n2248 ) | ( n805 & ~n2248 ) ;
  assign n2250 = n1142 & ~n2033 ;
  assign n2251 = n1179 & n2250 ;
  assign n2252 = n2251 ^ n765 ^ 1'b0 ;
  assign n2256 = n1044 ^ n963 ^ n301 ;
  assign n2255 = n867 ^ n809 ^ n263 ;
  assign n2257 = n2256 ^ n2255 ^ x67 ;
  assign n2253 = n1465 & ~n1667 ;
  assign n2254 = ~n1658 & n2253 ;
  assign n2258 = n2257 ^ n2254 ^ n1702 ;
  assign n2259 = n1149 ^ n1005 ^ x64 ;
  assign n2260 = ( x9 & ~n1787 ) | ( x9 & n2259 ) | ( ~n1787 & n2259 ) ;
  assign n2261 = n2260 ^ n1808 ^ 1'b0 ;
  assign n2262 = n462 & ~n2261 ;
  assign n2263 = n2262 ^ n335 ^ 1'b0 ;
  assign n2264 = ~n2258 & n2263 ;
  assign n2265 = n1006 ^ n383 ^ x109 ;
  assign n2269 = ( ~x97 & n858 ) | ( ~x97 & n1005 ) | ( n858 & n1005 ) ;
  assign n2270 = n2269 ^ n750 ^ n621 ;
  assign n2267 = n1452 ^ n892 ^ 1'b0 ;
  assign n2266 = n863 & ~n1331 ;
  assign n2268 = n2267 ^ n2266 ^ 1'b0 ;
  assign n2271 = n2270 ^ n2268 ^ x91 ;
  assign n2272 = ( n893 & n2265 ) | ( n893 & n2271 ) | ( n2265 & n2271 ) ;
  assign n2273 = ( ~n220 & n435 ) | ( ~n220 & n1073 ) | ( n435 & n1073 ) ;
  assign n2274 = ( n686 & ~n1365 ) | ( n686 & n2273 ) | ( ~n1365 & n2273 ) ;
  assign n2275 = n880 ^ n397 ^ n251 ;
  assign n2276 = ( x17 & ~n1789 ) | ( x17 & n2275 ) | ( ~n1789 & n2275 ) ;
  assign n2277 = n198 & n1480 ;
  assign n2278 = n2277 ^ n1689 ^ 1'b0 ;
  assign n2279 = n2276 & ~n2278 ;
  assign n2280 = n2183 ^ n752 ^ 1'b0 ;
  assign n2281 = ( n226 & n1000 ) | ( n226 & ~n2280 ) | ( n1000 & ~n2280 ) ;
  assign n2282 = n2279 & n2281 ;
  assign n2283 = n2274 & n2282 ;
  assign n2284 = ~n334 & n731 ;
  assign n2285 = n2283 & n2284 ;
  assign n2286 = n1703 ^ n1013 ^ n425 ;
  assign n2287 = n2286 ^ n916 ^ x105 ;
  assign n2291 = n2251 ^ n597 ^ n301 ;
  assign n2292 = n662 ^ n442 ^ n247 ;
  assign n2293 = ( ~n223 & n2291 ) | ( ~n223 & n2292 ) | ( n2291 & n2292 ) ;
  assign n2288 = n1798 & n2131 ;
  assign n2289 = n1481 & n2288 ;
  assign n2290 = n1955 & ~n2289 ;
  assign n2294 = n2293 ^ n2290 ^ 1'b0 ;
  assign n2295 = n2294 ^ n1932 ^ x113 ;
  assign n2296 = n2287 | n2295 ;
  assign n2298 = n295 & n983 ;
  assign n2299 = ~n809 & n2298 ;
  assign n2297 = n293 ^ n256 ^ 1'b0 ;
  assign n2300 = n2299 ^ n2297 ^ n1611 ;
  assign n2301 = n564 | n1481 ;
  assign n2302 = n2301 ^ n1705 ^ 1'b0 ;
  assign n2303 = n2302 ^ n1878 ^ n1831 ;
  assign n2304 = n448 & n2303 ;
  assign n2305 = n896 ^ n158 ^ 1'b0 ;
  assign n2306 = ( ~n877 & n996 ) | ( ~n877 & n2305 ) | ( n996 & n2305 ) ;
  assign n2309 = n1312 ^ n1165 ^ n538 ;
  assign n2310 = n2309 ^ n305 ^ n135 ;
  assign n2307 = n1536 ^ n1104 ^ n224 ;
  assign n2308 = n429 & n2307 ;
  assign n2311 = n2310 ^ n2308 ^ 1'b0 ;
  assign n2312 = n2311 ^ n2156 ^ n456 ;
  assign n2313 = n1258 ^ n546 ^ n526 ;
  assign n2314 = n1064 | n2313 ;
  assign n2315 = n1022 & ~n2314 ;
  assign n2316 = ~n716 & n2315 ;
  assign n2317 = n224 ^ x17 ^ 1'b0 ;
  assign n2318 = n2317 ^ n1523 ^ x93 ;
  assign n2319 = n358 | n2318 ;
  assign n2320 = n2319 ^ n1676 ^ 1'b0 ;
  assign n2321 = n649 & ~n2320 ;
  assign n2322 = n2321 ^ n591 ^ 1'b0 ;
  assign n2323 = ( n473 & n588 ) | ( n473 & ~n2009 ) | ( n588 & ~n2009 ) ;
  assign n2324 = n2323 ^ n1959 ^ 1'b0 ;
  assign n2325 = ~n2220 & n2324 ;
  assign n2326 = ( n1842 & n1990 ) | ( n1842 & n2325 ) | ( n1990 & n2325 ) ;
  assign n2327 = ( x56 & n1014 ) | ( x56 & n1837 ) | ( n1014 & n1837 ) ;
  assign n2328 = ( ~x106 & n454 ) | ( ~x106 & n1226 ) | ( n454 & n1226 ) ;
  assign n2329 = n710 ^ n228 ^ 1'b0 ;
  assign n2330 = ~n1216 & n1337 ;
  assign n2331 = ( ~n1264 & n2329 ) | ( ~n1264 & n2330 ) | ( n2329 & n2330 ) ;
  assign n2332 = n2328 | n2331 ;
  assign n2333 = n2332 ^ n382 ^ 1'b0 ;
  assign n2334 = n2327 & n2333 ;
  assign n2335 = ( ~n192 & n342 ) | ( ~n192 & n1046 ) | ( n342 & n1046 ) ;
  assign n2336 = n2335 ^ n678 ^ x43 ;
  assign n2337 = n449 | n1396 ;
  assign n2338 = ( n358 & n1127 ) | ( n358 & ~n1569 ) | ( n1127 & ~n1569 ) ;
  assign n2339 = n2338 ^ n321 ^ 1'b0 ;
  assign n2340 = x107 & ~n2339 ;
  assign n2341 = ( ~n194 & n343 ) | ( ~n194 & n869 ) | ( n343 & n869 ) ;
  assign n2342 = ( n358 & ~n1768 ) | ( n358 & n2341 ) | ( ~n1768 & n2341 ) ;
  assign n2343 = n1259 ^ x81 ^ 1'b0 ;
  assign n2344 = ( n1496 & n2342 ) | ( n1496 & n2343 ) | ( n2342 & n2343 ) ;
  assign n2345 = n2344 ^ n2105 ^ n1542 ;
  assign n2346 = n2345 ^ n1789 ^ 1'b0 ;
  assign n2347 = x96 & n1907 ;
  assign n2348 = n2347 ^ n149 ^ 1'b0 ;
  assign n2349 = n1338 & ~n2348 ;
  assign n2350 = ~n832 & n2349 ;
  assign n2351 = ( ~x21 & n419 ) | ( ~x21 & n2000 ) | ( n419 & n2000 ) ;
  assign n2352 = n2351 ^ n2206 ^ n1247 ;
  assign n2353 = ( ~n1481 & n1699 ) | ( ~n1481 & n2352 ) | ( n1699 & n2352 ) ;
  assign n2354 = ( n570 & ~n1065 ) | ( n570 & n1574 ) | ( ~n1065 & n1574 ) ;
  assign n2364 = n1867 ^ n1034 ^ n914 ;
  assign n2355 = n1156 ^ n1100 ^ x14 ;
  assign n2356 = n913 | n2355 ;
  assign n2357 = n506 & ~n1015 ;
  assign n2358 = n2357 ^ n595 ^ 1'b0 ;
  assign n2359 = n2358 ^ n1886 ^ 1'b0 ;
  assign n2360 = n1969 & n2359 ;
  assign n2361 = n2360 ^ n711 ^ n667 ;
  assign n2362 = n2361 ^ n1193 ^ 1'b0 ;
  assign n2363 = n2356 | n2362 ;
  assign n2365 = n2364 ^ n2363 ^ n469 ;
  assign n2378 = n1483 ^ n1139 ^ 1'b0 ;
  assign n2376 = n476 | n2305 ;
  assign n2377 = ( x85 & n1789 ) | ( x85 & ~n2376 ) | ( n1789 & ~n2376 ) ;
  assign n2366 = n1076 ^ n825 ^ 1'b0 ;
  assign n2367 = n991 & n2366 ;
  assign n2372 = n528 ^ x67 ^ x16 ;
  assign n2373 = n2372 ^ n1852 ^ n314 ;
  assign n2369 = n390 & n1231 ;
  assign n2370 = n758 & n2369 ;
  assign n2371 = ~n2145 & n2370 ;
  assign n2368 = n1575 ^ n1446 ^ 1'b0 ;
  assign n2374 = n2373 ^ n2371 ^ n2368 ;
  assign n2375 = ( ~n683 & n2367 ) | ( ~n683 & n2374 ) | ( n2367 & n2374 ) ;
  assign n2379 = n2378 ^ n2377 ^ n2375 ;
  assign n2380 = ( n1668 & n2365 ) | ( n1668 & n2379 ) | ( n2365 & n2379 ) ;
  assign n2381 = n2380 ^ n677 ^ x90 ;
  assign n2382 = n728 & ~n1440 ;
  assign n2383 = ~n983 & n2382 ;
  assign n2384 = ( ~n507 & n576 ) | ( ~n507 & n945 ) | ( n576 & n945 ) ;
  assign n2385 = n2384 ^ n515 ^ 1'b0 ;
  assign n2386 = n2385 ^ n184 ^ 1'b0 ;
  assign n2387 = n2386 ^ n567 ^ x87 ;
  assign n2388 = ~n1564 & n2387 ;
  assign n2389 = ( n1528 & ~n2045 ) | ( n1528 & n2388 ) | ( ~n2045 & n2388 ) ;
  assign n2393 = ( x79 & n369 ) | ( x79 & n1787 ) | ( n369 & n1787 ) ;
  assign n2394 = n2393 ^ n793 ^ x106 ;
  assign n2395 = ( ~x68 & n934 ) | ( ~x68 & n2394 ) | ( n934 & n2394 ) ;
  assign n2396 = n2395 ^ n497 ^ x33 ;
  assign n2397 = n917 & ~n2396 ;
  assign n2391 = ~n636 & n1304 ;
  assign n2392 = n2391 ^ n1028 ^ n992 ;
  assign n2390 = ( n442 & ~n748 ) | ( n442 & n1656 ) | ( ~n748 & n1656 ) ;
  assign n2398 = n2397 ^ n2392 ^ n2390 ;
  assign n2399 = n566 ^ n135 ^ 1'b0 ;
  assign n2400 = n302 & ~n2399 ;
  assign n2401 = n1004 ^ n486 ^ 1'b0 ;
  assign n2402 = n2400 & n2401 ;
  assign n2403 = ( ~n189 & n1008 ) | ( ~n189 & n2402 ) | ( n1008 & n2402 ) ;
  assign n2404 = n315 & ~n1319 ;
  assign n2405 = n2404 ^ n1753 ^ 1'b0 ;
  assign n2406 = n2405 ^ n348 ^ n240 ;
  assign n2407 = n1013 | n2406 ;
  assign n2408 = n2403 | n2407 ;
  assign n2414 = ( n579 & n920 ) | ( n579 & n1148 ) | ( n920 & n1148 ) ;
  assign n2409 = ( n1122 & n1780 ) | ( n1122 & n1828 ) | ( n1780 & n1828 ) ;
  assign n2410 = ~n574 & n2409 ;
  assign n2411 = ~x62 & n2410 ;
  assign n2412 = x94 & n2411 ;
  assign n2413 = n2412 ^ n1406 ^ n705 ;
  assign n2415 = n2414 ^ n2413 ^ x66 ;
  assign n2416 = n881 & ~n1421 ;
  assign n2417 = ~n460 & n2416 ;
  assign n2418 = n2417 ^ n2289 ^ n1120 ;
  assign n2419 = n1012 ^ n516 ^ 1'b0 ;
  assign n2420 = n2419 ^ n452 ^ 1'b0 ;
  assign n2421 = ( ~n969 & n2418 ) | ( ~n969 & n2420 ) | ( n2418 & n2420 ) ;
  assign n2422 = n933 ^ n662 ^ n162 ;
  assign n2423 = n155 & n2422 ;
  assign n2424 = n2423 ^ n1178 ^ 1'b0 ;
  assign n2425 = n1592 ^ n1347 ^ n409 ;
  assign n2426 = ( ~n1792 & n2424 ) | ( ~n1792 & n2425 ) | ( n2424 & n2425 ) ;
  assign n2427 = x33 & ~n252 ;
  assign n2428 = n2182 ^ n1568 ^ 1'b0 ;
  assign n2429 = ( n2426 & ~n2427 ) | ( n2426 & n2428 ) | ( ~n2427 & n2428 ) ;
  assign n2430 = n2185 ^ n441 ^ x118 ;
  assign n2431 = ( n329 & ~n2069 ) | ( n329 & n2430 ) | ( ~n2069 & n2430 ) ;
  assign n2432 = n1541 ^ n787 ^ n425 ;
  assign n2433 = n2432 ^ n2039 ^ n418 ;
  assign n2438 = ( n258 & n699 ) | ( n258 & n1865 ) | ( n699 & n1865 ) ;
  assign n2434 = ( ~x28 & n452 ) | ( ~x28 & n2079 ) | ( n452 & n2079 ) ;
  assign n2435 = n2434 ^ n1641 ^ n289 ;
  assign n2436 = n978 ^ n702 ^ 1'b0 ;
  assign n2437 = ( ~n664 & n2435 ) | ( ~n664 & n2436 ) | ( n2435 & n2436 ) ;
  assign n2439 = n2438 ^ n2437 ^ n2161 ;
  assign n2440 = n1876 ^ n1729 ^ n1660 ;
  assign n2441 = ( n814 & n1153 ) | ( n814 & ~n1380 ) | ( n1153 & ~n1380 ) ;
  assign n2442 = ( ~n1490 & n2062 ) | ( ~n1490 & n2441 ) | ( n2062 & n2441 ) ;
  assign n2443 = n2442 ^ n1343 ^ n233 ;
  assign n2444 = n1759 ^ n1272 ^ x5 ;
  assign n2445 = ( ~n1909 & n2443 ) | ( ~n1909 & n2444 ) | ( n2443 & n2444 ) ;
  assign n2446 = ( n732 & n2440 ) | ( n732 & n2445 ) | ( n2440 & n2445 ) ;
  assign n2447 = n1183 ^ n811 ^ x90 ;
  assign n2448 = ( ~x114 & n377 ) | ( ~x114 & n2447 ) | ( n377 & n2447 ) ;
  assign n2449 = ( n1045 & ~n1664 ) | ( n1045 & n2448 ) | ( ~n1664 & n2448 ) ;
  assign n2450 = n1638 ^ n1158 ^ x60 ;
  assign n2451 = n1292 ^ n553 ^ 1'b0 ;
  assign n2452 = n285 & n2451 ;
  assign n2453 = ( n143 & n502 ) | ( n143 & ~n2452 ) | ( n502 & ~n2452 ) ;
  assign n2454 = n2453 ^ n1075 ^ 1'b0 ;
  assign n2455 = n2450 & n2454 ;
  assign n2456 = ( x58 & n838 ) | ( x58 & ~n1336 ) | ( n838 & ~n1336 ) ;
  assign n2457 = ( ~n1949 & n2455 ) | ( ~n1949 & n2456 ) | ( n2455 & n2456 ) ;
  assign n2469 = n952 | n1691 ;
  assign n2470 = n2469 ^ n1610 ^ n263 ;
  assign n2458 = n987 ^ n656 ^ 1'b0 ;
  assign n2459 = n748 ^ n199 ^ x124 ;
  assign n2460 = n277 & n2459 ;
  assign n2461 = ~n873 & n2460 ;
  assign n2462 = n627 | n2461 ;
  assign n2463 = n2462 ^ n850 ^ 1'b0 ;
  assign n2464 = n2463 ^ n2146 ^ n905 ;
  assign n2465 = ( ~n1137 & n1612 ) | ( ~n1137 & n2464 ) | ( n1612 & n2464 ) ;
  assign n2466 = n1983 & n2411 ;
  assign n2467 = n2465 & n2466 ;
  assign n2468 = ~n2458 & n2467 ;
  assign n2471 = n2470 ^ n2468 ^ n961 ;
  assign n2472 = n394 & n452 ;
  assign n2478 = ( n476 & n565 ) | ( n476 & n668 ) | ( n565 & n668 ) ;
  assign n2473 = ( n502 & ~n898 ) | ( n502 & n1314 ) | ( ~n898 & n1314 ) ;
  assign n2474 = n1587 | n2473 ;
  assign n2475 = n2297 | n2474 ;
  assign n2476 = ~n1212 & n2475 ;
  assign n2477 = ( n414 & n2066 ) | ( n414 & ~n2476 ) | ( n2066 & ~n2476 ) ;
  assign n2479 = n2478 ^ n2477 ^ n503 ;
  assign n2480 = ( ~n888 & n1186 ) | ( ~n888 & n2438 ) | ( n1186 & n2438 ) ;
  assign n2481 = n2480 ^ n1995 ^ n1535 ;
  assign n2482 = ( n198 & n2379 ) | ( n198 & ~n2481 ) | ( n2379 & ~n2481 ) ;
  assign n2483 = n758 | n1049 ;
  assign n2484 = ( n424 & n1755 ) | ( n424 & n2483 ) | ( n1755 & n2483 ) ;
  assign n2485 = n442 ^ n258 ^ n160 ;
  assign n2486 = ( n1276 & n2412 ) | ( n1276 & ~n2485 ) | ( n2412 & ~n2485 ) ;
  assign n2487 = n2406 ^ n1723 ^ 1'b0 ;
  assign n2488 = ( ~n513 & n673 ) | ( ~n513 & n2487 ) | ( n673 & n2487 ) ;
  assign n2493 = n464 ^ n440 ^ n147 ;
  assign n2491 = n468 | n1533 ;
  assign n2492 = n2491 ^ n657 ^ 1'b0 ;
  assign n2494 = n2493 ^ n2492 ^ n191 ;
  assign n2489 = ( x52 & n925 ) | ( x52 & n1179 ) | ( n925 & n1179 ) ;
  assign n2490 = n808 & ~n2489 ;
  assign n2495 = n2494 ^ n2490 ^ 1'b0 ;
  assign n2499 = ( ~n293 & n459 ) | ( ~n293 & n878 ) | ( n459 & n878 ) ;
  assign n2500 = ~n1904 & n2499 ;
  assign n2501 = n2500 ^ n354 ^ 1'b0 ;
  assign n2502 = ( ~n685 & n951 ) | ( ~n685 & n1052 ) | ( n951 & n1052 ) ;
  assign n2503 = n1251 & ~n2502 ;
  assign n2504 = n2503 ^ n1825 ^ 1'b0 ;
  assign n2505 = n429 & n2504 ;
  assign n2506 = n1988 & n2505 ;
  assign n2507 = ( n1829 & ~n2501 ) | ( n1829 & n2506 ) | ( ~n2501 & n2506 ) ;
  assign n2496 = n1728 ^ n1568 ^ n158 ;
  assign n2497 = ( n1091 & ~n1703 ) | ( n1091 & n2496 ) | ( ~n1703 & n2496 ) ;
  assign n2498 = n399 & n2497 ;
  assign n2508 = n2507 ^ n2498 ^ 1'b0 ;
  assign n2509 = ~n1745 & n2508 ;
  assign n2510 = ( ~x120 & n399 ) | ( ~x120 & n1400 ) | ( n399 & n1400 ) ;
  assign n2511 = n2129 ^ n949 ^ x21 ;
  assign n2512 = ( n1010 & n2510 ) | ( n1010 & n2511 ) | ( n2510 & n2511 ) ;
  assign n2513 = n2458 ^ n2452 ^ n905 ;
  assign n2514 = n2512 | n2513 ;
  assign n2515 = n2509 & ~n2514 ;
  assign n2516 = ( n2488 & n2495 ) | ( n2488 & ~n2515 ) | ( n2495 & ~n2515 ) ;
  assign n2517 = n1380 & n2516 ;
  assign n2518 = x39 & n819 ;
  assign n2519 = ~n141 & n2518 ;
  assign n2520 = x45 & ~n500 ;
  assign n2521 = n2309 & n2520 ;
  assign n2522 = n2521 ^ x103 ^ 1'b0 ;
  assign n2523 = x1 & ~n2522 ;
  assign n2524 = n1398 ^ n981 ^ n206 ;
  assign n2525 = n2524 ^ n565 ^ 1'b0 ;
  assign n2526 = ( ~n653 & n2523 ) | ( ~n653 & n2525 ) | ( n2523 & n2525 ) ;
  assign n2527 = n186 | n256 ;
  assign n2528 = ( n837 & n862 ) | ( n837 & n2527 ) | ( n862 & n2527 ) ;
  assign n2529 = ~n454 & n1452 ;
  assign n2530 = ( x119 & n424 ) | ( x119 & n2529 ) | ( n424 & n2529 ) ;
  assign n2531 = ( ~x9 & x58 ) | ( ~x9 & n484 ) | ( x58 & n484 ) ;
  assign n2532 = n869 ^ n598 ^ n182 ;
  assign n2533 = ( n2530 & n2531 ) | ( n2530 & ~n2532 ) | ( n2531 & ~n2532 ) ;
  assign n2534 = n2528 & ~n2533 ;
  assign n2535 = ( n2519 & n2526 ) | ( n2519 & n2534 ) | ( n2526 & n2534 ) ;
  assign n2536 = n2430 ^ n575 ^ 1'b0 ;
  assign n2537 = ( n219 & ~n1290 ) | ( n219 & n1516 ) | ( ~n1290 & n1516 ) ;
  assign n2538 = ( x14 & n264 ) | ( x14 & ~n668 ) | ( n264 & ~n668 ) ;
  assign n2539 = n2538 ^ n1391 ^ n189 ;
  assign n2540 = ~n940 & n2539 ;
  assign n2548 = ( n590 & n816 ) | ( n590 & ~n1852 ) | ( n816 & ~n1852 ) ;
  assign n2549 = n1294 ^ n581 ^ n160 ;
  assign n2550 = ( n698 & n2548 ) | ( n698 & n2549 ) | ( n2548 & n2549 ) ;
  assign n2551 = n2550 ^ n2089 ^ n1808 ;
  assign n2542 = ( x42 & n228 ) | ( x42 & n998 ) | ( n228 & n998 ) ;
  assign n2543 = ~n1237 & n2542 ;
  assign n2544 = n1418 & n2543 ;
  assign n2545 = n2544 ^ n556 ^ 1'b0 ;
  assign n2541 = ~n1327 & n1659 ;
  assign n2546 = n2545 ^ n2541 ^ 1'b0 ;
  assign n2547 = n2546 ^ n909 ^ 1'b0 ;
  assign n2552 = n2551 ^ n2547 ^ 1'b0 ;
  assign n2554 = n1617 ^ n524 ^ 1'b0 ;
  assign n2553 = n153 & ~n915 ;
  assign n2555 = n2554 ^ n2553 ^ 1'b0 ;
  assign n2556 = ( x33 & ~n319 ) | ( x33 & n2275 ) | ( ~n319 & n2275 ) ;
  assign n2557 = n1958 ^ n1781 ^ n1050 ;
  assign n2558 = ( x59 & ~n2556 ) | ( x59 & n2557 ) | ( ~n2556 & n2557 ) ;
  assign n2559 = ( n2549 & ~n2555 ) | ( n2549 & n2558 ) | ( ~n2555 & n2558 ) ;
  assign n2560 = ( ~n2540 & n2552 ) | ( ~n2540 & n2559 ) | ( n2552 & n2559 ) ;
  assign n2561 = n2560 ^ n1780 ^ n1580 ;
  assign n2562 = n1807 ^ n1073 ^ n879 ;
  assign n2563 = n2562 ^ n1036 ^ 1'b0 ;
  assign n2568 = n2232 ^ n543 ^ x123 ;
  assign n2564 = n1407 ^ n851 ^ 1'b0 ;
  assign n2565 = n289 & n2564 ;
  assign n2566 = ( n940 & n1383 ) | ( n940 & ~n2565 ) | ( n1383 & ~n2565 ) ;
  assign n2567 = n1541 & ~n2566 ;
  assign n2569 = n2568 ^ n2567 ^ 1'b0 ;
  assign n2570 = ( x74 & ~n2563 ) | ( x74 & n2569 ) | ( ~n2563 & n2569 ) ;
  assign n2571 = n2302 ^ n1200 ^ n212 ;
  assign n2572 = n786 & ~n2571 ;
  assign n2573 = ( ~x16 & x102 ) | ( ~x16 & n1995 ) | ( x102 & n1995 ) ;
  assign n2574 = x21 & ~n2573 ;
  assign n2575 = ( n427 & n688 ) | ( n427 & n868 ) | ( n688 & n868 ) ;
  assign n2576 = n992 ^ n396 ^ 1'b0 ;
  assign n2577 = n2576 ^ n937 ^ n609 ;
  assign n2578 = ~x5 & n2577 ;
  assign n2579 = n2578 ^ n1918 ^ 1'b0 ;
  assign n2580 = ~n173 & n1288 ;
  assign n2581 = ~n758 & n2580 ;
  assign n2582 = n2581 ^ n242 ^ 1'b0 ;
  assign n2583 = n1149 & ~n2582 ;
  assign n2584 = ( n2313 & ~n2579 ) | ( n2313 & n2583 ) | ( ~n2579 & n2583 ) ;
  assign n2585 = n2304 ^ n2218 ^ n1266 ;
  assign n2586 = n790 ^ n597 ^ 1'b0 ;
  assign n2587 = n2586 ^ n1087 ^ x3 ;
  assign n2588 = n2587 ^ n624 ^ 1'b0 ;
  assign n2593 = n1291 ^ n980 ^ n814 ;
  assign n2589 = ( n735 & n1493 ) | ( n735 & n1752 ) | ( n1493 & n1752 ) ;
  assign n2590 = n2589 ^ x90 ^ 1'b0 ;
  assign n2591 = n510 & n2590 ;
  assign n2592 = n2591 ^ n2573 ^ n1552 ;
  assign n2594 = n2593 ^ n2592 ^ n1587 ;
  assign n2595 = ( x92 & n881 ) | ( x92 & ~n945 ) | ( n881 & ~n945 ) ;
  assign n2596 = n2275 ^ n1560 ^ 1'b0 ;
  assign n2597 = n1867 & n2596 ;
  assign n2598 = n1836 & n2597 ;
  assign n2599 = ( n346 & ~n864 ) | ( n346 & n1487 ) | ( ~n864 & n1487 ) ;
  assign n2600 = n1842 & n2066 ;
  assign n2601 = n2599 & n2600 ;
  assign n2602 = ( n2595 & ~n2598 ) | ( n2595 & n2601 ) | ( ~n2598 & n2601 ) ;
  assign n2603 = ( n766 & ~n946 ) | ( n766 & n1560 ) | ( ~n946 & n1560 ) ;
  assign n2604 = ( n2343 & n2375 ) | ( n2343 & n2603 ) | ( n2375 & n2603 ) ;
  assign n2606 = ( n890 & n1437 ) | ( n890 & ~n1773 ) | ( n1437 & ~n1773 ) ;
  assign n2605 = ( x107 & n478 ) | ( x107 & ~n2297 ) | ( n478 & ~n2297 ) ;
  assign n2607 = n2606 ^ n2605 ^ n2515 ;
  assign n2608 = ( n1923 & n2604 ) | ( n1923 & ~n2607 ) | ( n2604 & ~n2607 ) ;
  assign n2612 = ( x97 & n526 ) | ( x97 & ~n1464 ) | ( n526 & ~n1464 ) ;
  assign n2609 = n2286 ^ n1375 ^ n1228 ;
  assign n2610 = n296 & ~n2609 ;
  assign n2611 = n1787 | n2610 ;
  assign n2613 = n2612 ^ n2611 ^ 1'b0 ;
  assign n2614 = n1992 ^ n1011 ^ 1'b0 ;
  assign n2615 = n1788 ^ n1705 ^ n858 ;
  assign n2616 = n2615 ^ n1855 ^ 1'b0 ;
  assign n2617 = n2614 | n2616 ;
  assign n2618 = n1354 ^ n984 ^ x69 ;
  assign n2619 = n539 ^ n315 ^ 1'b0 ;
  assign n2620 = ( ~n892 & n1584 ) | ( ~n892 & n2619 ) | ( n1584 & n2619 ) ;
  assign n2621 = ( n1462 & n2138 ) | ( n1462 & n2620 ) | ( n2138 & n2620 ) ;
  assign n2622 = ( n223 & ~n2618 ) | ( n223 & n2621 ) | ( ~n2618 & n2621 ) ;
  assign n2623 = n2501 ^ n223 ^ n146 ;
  assign n2624 = n2623 ^ n1853 ^ n1455 ;
  assign n2625 = ( ~n1888 & n2622 ) | ( ~n1888 & n2624 ) | ( n2622 & n2624 ) ;
  assign n2629 = ( n578 & n580 ) | ( n578 & ~n719 ) | ( n580 & ~n719 ) ;
  assign n2626 = ( n228 & n1688 ) | ( n228 & ~n2144 ) | ( n1688 & ~n2144 ) ;
  assign n2627 = n2626 ^ n793 ^ 1'b0 ;
  assign n2628 = ~n1563 & n2627 ;
  assign n2630 = n2629 ^ n2628 ^ n226 ;
  assign n2631 = n2630 ^ n2309 ^ n2089 ;
  assign n2632 = n2631 ^ n1102 ^ 1'b0 ;
  assign n2633 = ( n296 & n776 ) | ( n296 & ~n1572 ) | ( n776 & ~n1572 ) ;
  assign n2634 = n2633 ^ n1546 ^ 1'b0 ;
  assign n2635 = n2634 ^ n1836 ^ n146 ;
  assign n2636 = ( ~x53 & n314 ) | ( ~x53 & n1034 ) | ( n314 & n1034 ) ;
  assign n2637 = ( n447 & n2391 ) | ( n447 & ~n2636 ) | ( n2391 & ~n2636 ) ;
  assign n2638 = ~n2385 & n2637 ;
  assign n2639 = n2635 & n2638 ;
  assign n2640 = ( n239 & n280 ) | ( n239 & n388 ) | ( n280 & n388 ) ;
  assign n2641 = n1493 & ~n1575 ;
  assign n2642 = ~n2640 & n2641 ;
  assign n2643 = n1422 | n2642 ;
  assign n2644 = ( ~n1534 & n2639 ) | ( ~n1534 & n2643 ) | ( n2639 & n2643 ) ;
  assign n2645 = x16 & n1165 ;
  assign n2646 = n2645 ^ n2310 ^ 1'b0 ;
  assign n2647 = n2646 ^ n2388 ^ n249 ;
  assign n2648 = n1962 ^ n970 ^ n858 ;
  assign n2649 = n1954 ^ n717 ^ x42 ;
  assign n2650 = n958 | n1298 ;
  assign n2651 = n2650 ^ n2337 ^ n178 ;
  assign n2652 = ~n1243 & n2651 ;
  assign n2664 = n1372 ^ n565 ^ n165 ;
  assign n2665 = ( n301 & ~n326 ) | ( n301 & n2664 ) | ( ~n326 & n2664 ) ;
  assign n2666 = n2665 ^ n306 ^ 1'b0 ;
  assign n2667 = n2666 ^ n557 ^ n333 ;
  assign n2658 = ( ~n817 & n1056 ) | ( ~n817 & n1127 ) | ( n1056 & n1127 ) ;
  assign n2657 = x70 & ~n166 ;
  assign n2659 = n2658 ^ n2657 ^ 1'b0 ;
  assign n2660 = n2659 ^ n1066 ^ n820 ;
  assign n2661 = n2521 & ~n2660 ;
  assign n2662 = n2422 ^ n1135 ^ n206 ;
  assign n2663 = ( x65 & n2661 ) | ( x65 & n2662 ) | ( n2661 & n2662 ) ;
  assign n2655 = n1019 ^ x78 ^ 1'b0 ;
  assign n2653 = ( x92 & n515 ) | ( x92 & ~n1075 ) | ( n515 & ~n1075 ) ;
  assign n2654 = n2653 ^ n2512 ^ n1557 ;
  assign n2656 = n2655 ^ n2654 ^ n282 ;
  assign n2668 = n2667 ^ n2663 ^ n2656 ;
  assign n2669 = ~n216 & n731 ;
  assign n2670 = n2669 ^ x46 ^ 1'b0 ;
  assign n2671 = ( n2373 & ~n2571 ) | ( n2373 & n2670 ) | ( ~n2571 & n2670 ) ;
  assign n2676 = n1645 ^ n784 ^ n152 ;
  assign n2675 = n198 & ~n430 ;
  assign n2677 = n2676 ^ n2675 ^ 1'b0 ;
  assign n2673 = n1523 ^ n626 ^ n597 ;
  assign n2674 = ( n1607 & n2106 ) | ( n1607 & n2673 ) | ( n2106 & n2673 ) ;
  assign n2678 = n2677 ^ n2674 ^ x7 ;
  assign n2672 = n302 & ~n1542 ;
  assign n2679 = n2678 ^ n2672 ^ 1'b0 ;
  assign n2680 = n2076 ^ n351 ^ n175 ;
  assign n2681 = ( ~n1230 & n1776 ) | ( ~n1230 & n2090 ) | ( n1776 & n2090 ) ;
  assign n2682 = n2680 & n2681 ;
  assign n2683 = n2679 & n2682 ;
  assign n2684 = n2665 ^ n1367 ^ 1'b0 ;
  assign n2685 = n2226 & ~n2684 ;
  assign n2686 = ( n147 & n704 ) | ( n147 & n1957 ) | ( n704 & n1957 ) ;
  assign n2687 = ~n543 & n2686 ;
  assign n2688 = ( n838 & n2685 ) | ( n838 & ~n2687 ) | ( n2685 & ~n2687 ) ;
  assign n2690 = n1503 ^ n1126 ^ x120 ;
  assign n2689 = n164 & ~n450 ;
  assign n2691 = n2690 ^ n2689 ^ n1010 ;
  assign n2692 = ( n751 & n1702 ) | ( n751 & n2691 ) | ( n1702 & n2691 ) ;
  assign n2693 = n2688 & ~n2692 ;
  assign n2694 = n1748 & n2693 ;
  assign n2695 = n2683 | n2694 ;
  assign n2696 = ( n2124 & n2671 ) | ( n2124 & ~n2695 ) | ( n2671 & ~n2695 ) ;
  assign n2698 = ( x18 & n452 ) | ( x18 & n947 ) | ( n452 & n947 ) ;
  assign n2699 = n2698 ^ n1037 ^ n408 ;
  assign n2697 = n1781 ^ n1497 ^ n763 ;
  assign n2700 = n2699 ^ n2697 ^ n2144 ;
  assign n2701 = n1101 & ~n1820 ;
  assign n2702 = ( n827 & n911 ) | ( n827 & ~n1313 ) | ( n911 & ~n1313 ) ;
  assign n2703 = ( n1936 & n2229 ) | ( n1936 & n2702 ) | ( n2229 & n2702 ) ;
  assign n2704 = n2703 ^ n1585 ^ n1502 ;
  assign n2705 = ( n343 & n890 ) | ( n343 & n2704 ) | ( n890 & n2704 ) ;
  assign n2706 = ( x113 & ~n2248 ) | ( x113 & n2705 ) | ( ~n2248 & n2705 ) ;
  assign n2721 = ( ~x57 & n1855 ) | ( ~x57 & n2185 ) | ( n1855 & n2185 ) ;
  assign n2718 = n2438 ^ n1842 ^ n838 ;
  assign n2716 = n152 & n2576 ;
  assign n2715 = ( n981 & n1893 ) | ( n981 & n2132 ) | ( n1893 & n2132 ) ;
  assign n2717 = n2716 ^ n2715 ^ n364 ;
  assign n2719 = n2718 ^ n2717 ^ n583 ;
  assign n2720 = n2719 ^ n1847 ^ n1406 ;
  assign n2711 = ( x75 & ~n857 ) | ( x75 & n1510 ) | ( ~n857 & n1510 ) ;
  assign n2712 = ~n1080 & n1517 ;
  assign n2713 = ( n893 & n2612 ) | ( n893 & n2712 ) | ( n2612 & n2712 ) ;
  assign n2714 = ( n2493 & n2711 ) | ( n2493 & n2713 ) | ( n2711 & n2713 ) ;
  assign n2722 = n2721 ^ n2720 ^ n2714 ;
  assign n2707 = n2047 ^ x96 ^ 1'b0 ;
  assign n2708 = n474 | n2707 ;
  assign n2709 = n2708 ^ n762 ^ n582 ;
  assign n2710 = n2637 & n2709 ;
  assign n2723 = n2722 ^ n2710 ^ 1'b0 ;
  assign n2724 = ( ~n678 & n712 ) | ( ~n678 & n855 ) | ( n712 & n855 ) ;
  assign n2728 = n677 & ~n754 ;
  assign n2729 = n1852 ^ n497 ^ n340 ;
  assign n2730 = ( n138 & ~n771 ) | ( n138 & n1436 ) | ( ~n771 & n1436 ) ;
  assign n2731 = ( n775 & ~n2729 ) | ( n775 & n2730 ) | ( ~n2729 & n2730 ) ;
  assign n2732 = ( n1129 & ~n2728 ) | ( n1129 & n2731 ) | ( ~n2728 & n2731 ) ;
  assign n2726 = ( n401 & n705 ) | ( n401 & n1119 ) | ( n705 & n1119 ) ;
  assign n2725 = ( ~x22 & n1718 ) | ( ~x22 & n2670 ) | ( n1718 & n2670 ) ;
  assign n2727 = n2726 ^ n2725 ^ n1774 ;
  assign n2733 = n2732 ^ n2727 ^ n2199 ;
  assign n2734 = ( n986 & n2724 ) | ( n986 & n2733 ) | ( n2724 & n2733 ) ;
  assign n2735 = ( n2706 & n2723 ) | ( n2706 & ~n2734 ) | ( n2723 & ~n2734 ) ;
  assign n2736 = n1479 ^ n701 ^ 1'b0 ;
  assign n2737 = n911 | n2736 ;
  assign n2738 = ( n276 & n2530 ) | ( n276 & ~n2737 ) | ( n2530 & ~n2737 ) ;
  assign n2739 = ( n728 & n1266 ) | ( n728 & ~n2738 ) | ( n1266 & ~n2738 ) ;
  assign n2740 = ( n429 & n1618 ) | ( n429 & ~n2739 ) | ( n1618 & ~n2739 ) ;
  assign n2741 = n798 ^ n535 ^ 1'b0 ;
  assign n2742 = n2741 ^ n1857 ^ n937 ;
  assign n2743 = ( n2328 & n2544 ) | ( n2328 & n2742 ) | ( n2544 & n2742 ) ;
  assign n2744 = n931 & n1125 ;
  assign n2745 = ( n478 & ~n1077 ) | ( n478 & n2744 ) | ( ~n1077 & n2744 ) ;
  assign n2746 = n969 ^ n256 ^ 1'b0 ;
  assign n2747 = ( ~n1633 & n1849 ) | ( ~n1633 & n2746 ) | ( n1849 & n2746 ) ;
  assign n2748 = n1723 ^ n1654 ^ n1224 ;
  assign n2752 = ( n628 & n670 ) | ( n628 & n2523 ) | ( n670 & n2523 ) ;
  assign n2750 = n689 ^ n254 ^ n208 ;
  assign n2749 = n2160 ^ n1974 ^ n293 ;
  assign n2751 = n2750 ^ n2749 ^ x75 ;
  assign n2753 = n2752 ^ n2751 ^ n2058 ;
  assign n2754 = n2464 ^ n1021 ^ n187 ;
  assign n2755 = ( n956 & n1597 ) | ( n956 & ~n2754 ) | ( n1597 & ~n2754 ) ;
  assign n2758 = ( ~n869 & n1774 ) | ( ~n869 & n1995 ) | ( n1774 & n1995 ) ;
  assign n2759 = n2758 ^ n963 ^ n751 ;
  assign n2756 = n505 ^ n439 ^ x114 ;
  assign n2757 = n2756 ^ n1417 ^ x126 ;
  assign n2760 = n2759 ^ n2757 ^ n2200 ;
  assign n2769 = ( ~n828 & n941 ) | ( ~n828 & n1224 ) | ( n941 & n1224 ) ;
  assign n2770 = ( n627 & ~n1855 ) | ( n627 & n2769 ) | ( ~n1855 & n2769 ) ;
  assign n2761 = n483 ^ n226 ^ 1'b0 ;
  assign n2762 = n2761 ^ n862 ^ n516 ;
  assign n2763 = n306 & ~n1568 ;
  assign n2764 = n2763 ^ x76 ^ 1'b0 ;
  assign n2765 = n2762 | n2764 ;
  assign n2766 = n2765 ^ n737 ^ 1'b0 ;
  assign n2767 = n2766 ^ n2563 ^ n723 ;
  assign n2768 = n2713 & n2767 ;
  assign n2771 = n2770 ^ n2768 ^ 1'b0 ;
  assign n2772 = x58 & n392 ;
  assign n2773 = n2772 ^ n1116 ^ 1'b0 ;
  assign n2774 = ( ~n1677 & n2317 ) | ( ~n1677 & n2773 ) | ( n2317 & n2773 ) ;
  assign n2775 = ( n468 & n1559 ) | ( n468 & ~n2774 ) | ( n1559 & ~n2774 ) ;
  assign n2776 = ( n402 & ~n2372 ) | ( n402 & n2775 ) | ( ~n2372 & n2775 ) ;
  assign n2777 = n2776 ^ n1679 ^ x93 ;
  assign n2796 = n662 & n1030 ;
  assign n2797 = n2796 ^ n178 ^ 1'b0 ;
  assign n2798 = n2752 & n2797 ;
  assign n2799 = ~n282 & n2798 ;
  assign n2800 = ( ~n252 & n911 ) | ( ~n252 & n2799 ) | ( n911 & n2799 ) ;
  assign n2778 = ( ~x111 & n256 ) | ( ~x111 & n448 ) | ( n256 & n448 ) ;
  assign n2779 = ~n1703 & n1960 ;
  assign n2780 = n2779 ^ n382 ^ 1'b0 ;
  assign n2781 = ( n258 & n2778 ) | ( n258 & ~n2780 ) | ( n2778 & ~n2780 ) ;
  assign n2782 = ( ~n883 & n1076 ) | ( ~n883 & n1226 ) | ( n1076 & n1226 ) ;
  assign n2783 = n849 ^ x54 ^ 1'b0 ;
  assign n2784 = ( ~n451 & n1251 ) | ( ~n451 & n2783 ) | ( n1251 & n2783 ) ;
  assign n2785 = n2093 ^ n275 ^ 1'b0 ;
  assign n2786 = ~n675 & n2785 ;
  assign n2787 = ( n742 & n2784 ) | ( n742 & ~n2786 ) | ( n2784 & ~n2786 ) ;
  assign n2788 = ( n350 & ~n538 ) | ( n350 & n2787 ) | ( ~n538 & n2787 ) ;
  assign n2789 = n1523 ^ n720 ^ x95 ;
  assign n2790 = ( ~n1167 & n1296 ) | ( ~n1167 & n2789 ) | ( n1296 & n2789 ) ;
  assign n2791 = n654 & n2790 ;
  assign n2792 = ~n2310 & n2791 ;
  assign n2793 = n2792 ^ n2628 ^ n258 ;
  assign n2794 = ( n2782 & n2788 ) | ( n2782 & n2793 ) | ( n2788 & n2793 ) ;
  assign n2795 = ( n765 & n2781 ) | ( n765 & n2794 ) | ( n2781 & n2794 ) ;
  assign n2801 = n2800 ^ n2795 ^ n192 ;
  assign n2802 = ( n746 & n1154 ) | ( n746 & ~n2186 ) | ( n1154 & ~n2186 ) ;
  assign n2803 = n1120 | n2579 ;
  assign n2804 = ( n2120 & n2802 ) | ( n2120 & ~n2803 ) | ( n2802 & ~n2803 ) ;
  assign n2805 = n273 | n706 ;
  assign n2806 = n1604 & ~n2805 ;
  assign n2807 = n2200 | n2806 ;
  assign n2808 = n1112 & ~n2807 ;
  assign n2809 = ( n374 & ~n488 ) | ( n374 & n1740 ) | ( ~n488 & n1740 ) ;
  assign n2810 = n1016 ^ n709 ^ n385 ;
  assign n2811 = n249 & n2810 ;
  assign n2812 = n2811 ^ n2593 ^ 1'b0 ;
  assign n2813 = n2812 ^ n2228 ^ n2215 ;
  assign n2814 = n2813 ^ x91 ^ 1'b0 ;
  assign n2815 = n1594 | n2814 ;
  assign n2816 = ( n1932 & ~n2809 ) | ( n1932 & n2815 ) | ( ~n2809 & n2815 ) ;
  assign n2817 = n2816 ^ n1644 ^ 1'b0 ;
  assign n2818 = n510 & n2817 ;
  assign n2819 = ( ~n1520 & n2138 ) | ( ~n1520 & n2144 ) | ( n2138 & n2144 ) ;
  assign n2820 = x52 & ~n1510 ;
  assign n2821 = ( ~n822 & n885 ) | ( ~n822 & n2156 ) | ( n885 & n2156 ) ;
  assign n2822 = n2821 ^ n762 ^ n192 ;
  assign n2823 = n772 ^ n716 ^ 1'b0 ;
  assign n2824 = n2823 ^ n388 ^ 1'b0 ;
  assign n2825 = ~n2822 & n2824 ;
  assign n2826 = ( x25 & n2820 ) | ( x25 & ~n2825 ) | ( n2820 & ~n2825 ) ;
  assign n2827 = n2819 & n2826 ;
  assign n2828 = ( n583 & n1643 ) | ( n583 & ~n2827 ) | ( n1643 & ~n2827 ) ;
  assign n2829 = x37 & ~n1999 ;
  assign n2835 = n1822 ^ n1768 ^ 1'b0 ;
  assign n2833 = n536 ^ n272 ^ 1'b0 ;
  assign n2834 = n1283 & ~n2833 ;
  assign n2830 = n153 ^ x56 ^ x4 ;
  assign n2831 = n2830 ^ n1279 ^ n171 ;
  assign n2832 = n2521 & n2831 ;
  assign n2836 = n2835 ^ n2834 ^ n2832 ;
  assign n2843 = n209 ^ n152 ^ n149 ;
  assign n2844 = ( n438 & n1647 ) | ( n438 & ~n2843 ) | ( n1647 & ~n2843 ) ;
  assign n2845 = n2844 ^ n1949 ^ n1171 ;
  assign n2842 = n1981 ^ n272 ^ 1'b0 ;
  assign n2839 = n2036 ^ n1936 ^ n534 ;
  assign n2840 = ( n589 & ~n1314 ) | ( n589 & n2839 ) | ( ~n1314 & n2839 ) ;
  assign n2838 = n2435 ^ n1292 ^ n159 ;
  assign n2837 = n2797 ^ n1690 ^ n1441 ;
  assign n2841 = n2840 ^ n2838 ^ n2837 ;
  assign n2846 = n2845 ^ n2842 ^ n2841 ;
  assign n2847 = n639 | n2846 ;
  assign n2848 = n2769 ^ n257 ^ 1'b0 ;
  assign n2849 = x6 & ~n2848 ;
  assign n2850 = ( x26 & n1064 ) | ( x26 & ~n2849 ) | ( n1064 & ~n2849 ) ;
  assign n2851 = ( n234 & ~n256 ) | ( n234 & n841 ) | ( ~n256 & n841 ) ;
  assign n2852 = n2851 ^ n145 ^ 1'b0 ;
  assign n2855 = n1332 ^ n1045 ^ n445 ;
  assign n2853 = ( n226 & n495 ) | ( n226 & n561 ) | ( n495 & n561 ) ;
  assign n2854 = ( n1476 & ~n1485 ) | ( n1476 & n2853 ) | ( ~n1485 & n2853 ) ;
  assign n2856 = n2855 ^ n2854 ^ n645 ;
  assign n2857 = ~n2852 & n2856 ;
  assign n2859 = n2293 ^ n1072 ^ n174 ;
  assign n2858 = ( ~n823 & n890 ) | ( ~n823 & n1757 ) | ( n890 & n1757 ) ;
  assign n2860 = n2859 ^ n2858 ^ n1528 ;
  assign n2861 = ( n1036 & ~n2857 ) | ( n1036 & n2860 ) | ( ~n2857 & n2860 ) ;
  assign n2862 = ( n647 & n1789 ) | ( n647 & ~n2086 ) | ( n1789 & ~n2086 ) ;
  assign n2863 = n2862 ^ n1886 ^ 1'b0 ;
  assign n2864 = n2689 | n2863 ;
  assign n2865 = ~n1174 & n1664 ;
  assign n2866 = n1694 & n2865 ;
  assign n2867 = ~n421 & n1610 ;
  assign n2868 = n2867 ^ n159 ^ 1'b0 ;
  assign n2869 = n2868 ^ n285 ^ n268 ;
  assign n2870 = n1419 ^ x101 ^ 1'b0 ;
  assign n2871 = ~n849 & n2870 ;
  assign n2872 = ( n489 & n2869 ) | ( n489 & n2871 ) | ( n2869 & n2871 ) ;
  assign n2873 = ( n1577 & n2054 ) | ( n1577 & ~n2872 ) | ( n2054 & ~n2872 ) ;
  assign n2874 = ( n1369 & ~n2356 ) | ( n1369 & n2873 ) | ( ~n2356 & n2873 ) ;
  assign n2887 = n437 & n747 ;
  assign n2888 = n2887 ^ x92 ^ 1'b0 ;
  assign n2885 = ( n308 & ~n560 ) | ( n308 & n772 ) | ( ~n560 & n772 ) ;
  assign n2886 = ( n1054 & n1488 ) | ( n1054 & n2885 ) | ( n1488 & n2885 ) ;
  assign n2876 = ( n468 & ~n924 ) | ( n468 & n1010 ) | ( ~n924 & n1010 ) ;
  assign n2875 = ( n1097 & n1176 ) | ( n1097 & ~n1765 ) | ( n1176 & ~n1765 ) ;
  assign n2877 = n2876 ^ n2875 ^ n2082 ;
  assign n2881 = ( n347 & n380 ) | ( n347 & ~n769 ) | ( n380 & ~n769 ) ;
  assign n2880 = ( n724 & ~n1473 ) | ( n724 & n1712 ) | ( ~n1473 & n1712 ) ;
  assign n2882 = n2881 ^ n2880 ^ n1507 ;
  assign n2878 = n1847 ^ n1484 ^ n1152 ;
  assign n2879 = ( n1007 & n1550 ) | ( n1007 & n2878 ) | ( n1550 & n2878 ) ;
  assign n2883 = n2882 ^ n2879 ^ n1779 ;
  assign n2884 = ( n2234 & n2877 ) | ( n2234 & ~n2883 ) | ( n2877 & ~n2883 ) ;
  assign n2889 = n2888 ^ n2886 ^ n2884 ;
  assign n2890 = ( x63 & ~x74 ) | ( x63 & n200 ) | ( ~x74 & n200 ) ;
  assign n2891 = n2890 ^ n2529 ^ n1276 ;
  assign n2892 = n2891 ^ n1125 ^ n747 ;
  assign n2893 = ( ~n462 & n488 ) | ( ~n462 & n1392 ) | ( n488 & n1392 ) ;
  assign n2894 = n2892 & ~n2893 ;
  assign n2895 = n2894 ^ n1254 ^ 1'b0 ;
  assign n2896 = n1076 ^ n588 ^ 1'b0 ;
  assign n2897 = n601 ^ n417 ^ 1'b0 ;
  assign n2898 = n912 ^ n451 ^ x7 ;
  assign n2899 = n491 & ~n2898 ;
  assign n2900 = n2897 & n2899 ;
  assign n2901 = n1430 ^ n937 ^ x104 ;
  assign n2902 = n1491 ^ n512 ^ x31 ;
  assign n2903 = n2902 ^ n2573 ^ n386 ;
  assign n2904 = ( n567 & n2901 ) | ( n567 & n2903 ) | ( n2901 & n2903 ) ;
  assign n2905 = ( n1735 & n2186 ) | ( n1735 & ~n2904 ) | ( n2186 & ~n2904 ) ;
  assign n2906 = ( n1226 & ~n2900 ) | ( n1226 & n2905 ) | ( ~n2900 & n2905 ) ;
  assign n2907 = n2274 ^ n2220 ^ n969 ;
  assign n2908 = ~n1887 & n2907 ;
  assign n2909 = n239 & ~n2908 ;
  assign n2910 = n567 | n1936 ;
  assign n2911 = n2910 ^ n915 ^ 1'b0 ;
  assign n2912 = n2241 | n2911 ;
  assign n2913 = n1971 | n2912 ;
  assign n2914 = ( x93 & n1319 ) | ( x93 & ~n1697 ) | ( n1319 & ~n1697 ) ;
  assign n2915 = ( n996 & n1453 ) | ( n996 & ~n2914 ) | ( n1453 & ~n2914 ) ;
  assign n2916 = ( n698 & n833 ) | ( n698 & n1279 ) | ( n833 & n1279 ) ;
  assign n2917 = ~n367 & n2916 ;
  assign n2918 = ~n2040 & n2917 ;
  assign n2919 = ~n1405 & n1858 ;
  assign n2920 = n2918 & n2919 ;
  assign n2921 = n2800 ^ n1206 ^ n1080 ;
  assign n2923 = ( n457 & n514 ) | ( n457 & ~n541 ) | ( n514 & ~n541 ) ;
  assign n2924 = ( n275 & ~n1282 ) | ( n275 & n2923 ) | ( ~n1282 & n2923 ) ;
  assign n2925 = ( n422 & n588 ) | ( n422 & n2924 ) | ( n588 & n2924 ) ;
  assign n2922 = n2323 ^ n2129 ^ n1149 ;
  assign n2926 = n2925 ^ n2922 ^ n678 ;
  assign n2927 = ( n2341 & n2921 ) | ( n2341 & n2926 ) | ( n2921 & n2926 ) ;
  assign n2928 = n2927 ^ n1835 ^ n1447 ;
  assign n2929 = n1488 ^ n1273 ^ n445 ;
  assign n2931 = n850 ^ n562 ^ n238 ;
  assign n2930 = n534 & n1142 ;
  assign n2932 = n2931 ^ n2930 ^ n1545 ;
  assign n2933 = ( ~n272 & n894 ) | ( ~n272 & n2309 ) | ( n894 & n2309 ) ;
  assign n2934 = ( n689 & n2932 ) | ( n689 & n2933 ) | ( n2932 & n2933 ) ;
  assign n2935 = x80 & n364 ;
  assign n2936 = n2935 ^ n1523 ^ 1'b0 ;
  assign n2937 = ~n344 & n2936 ;
  assign n2938 = n2937 ^ n1749 ^ n1257 ;
  assign n2939 = n2938 ^ n1748 ^ 1'b0 ;
  assign n2940 = n1340 & n2939 ;
  assign n2941 = ( ~x125 & n512 ) | ( ~x125 & n610 ) | ( n512 & n610 ) ;
  assign n2942 = n1225 & ~n2941 ;
  assign n2943 = ~n2940 & n2942 ;
  assign n2944 = ( n2929 & n2934 ) | ( n2929 & ~n2943 ) | ( n2934 & ~n2943 ) ;
  assign n2945 = n2348 ^ n1753 ^ n248 ;
  assign n2946 = n1107 & ~n1113 ;
  assign n2947 = n2011 & n2946 ;
  assign n2948 = n2945 | n2947 ;
  assign n2949 = n450 & n1032 ;
  assign n2950 = ( n1526 & n2471 ) | ( n1526 & ~n2949 ) | ( n2471 & ~n2949 ) ;
  assign n2951 = n612 & n1159 ;
  assign n2952 = ~n1416 & n2951 ;
  assign n2954 = n2442 ^ n1168 ^ 1'b0 ;
  assign n2955 = ( ~n597 & n867 ) | ( ~n597 & n2954 ) | ( n867 & n2954 ) ;
  assign n2953 = ( ~n640 & n1828 ) | ( ~n640 & n2741 ) | ( n1828 & n2741 ) ;
  assign n2956 = n2955 ^ n2953 ^ n214 ;
  assign n2957 = ( ~n1292 & n2952 ) | ( ~n1292 & n2956 ) | ( n2952 & n2956 ) ;
  assign n2964 = ( n475 & n721 ) | ( n475 & n1101 ) | ( n721 & n1101 ) ;
  assign n2965 = n2964 ^ n2732 ^ n2038 ;
  assign n2958 = n1318 & n1695 ;
  assign n2960 = n736 ^ n258 ^ x78 ;
  assign n2959 = ( ~n295 & n507 ) | ( ~n295 & n2422 ) | ( n507 & n2422 ) ;
  assign n2961 = n2960 ^ n2959 ^ 1'b0 ;
  assign n2962 = n854 & ~n2961 ;
  assign n2963 = n2958 & n2962 ;
  assign n2966 = n2965 ^ n2963 ^ n1455 ;
  assign n2967 = n1704 ^ n1576 ^ n664 ;
  assign n2971 = x24 & n997 ;
  assign n2968 = ( n273 & n1487 ) | ( n273 & ~n2064 ) | ( n1487 & ~n2064 ) ;
  assign n2969 = n2968 ^ n2670 ^ n233 ;
  assign n2970 = n2969 ^ n1478 ^ n429 ;
  assign n2972 = n2971 ^ n2970 ^ n582 ;
  assign n2973 = n440 & n1936 ;
  assign n2974 = ( ~n886 & n1789 ) | ( ~n886 & n2973 ) | ( n1789 & n2973 ) ;
  assign n2975 = ~n469 & n728 ;
  assign n2976 = n2975 ^ n987 ^ 1'b0 ;
  assign n2977 = ( n1980 & n2974 ) | ( n1980 & ~n2976 ) | ( n2974 & ~n2976 ) ;
  assign n2978 = ( ~n133 & n1559 ) | ( ~n133 & n2977 ) | ( n1559 & n2977 ) ;
  assign n2981 = n2028 ^ n1211 ^ n858 ;
  assign n2982 = n2981 ^ n627 ^ n564 ;
  assign n2983 = ( ~n2043 & n2120 ) | ( ~n2043 & n2982 ) | ( n2120 & n2982 ) ;
  assign n2979 = n394 & ~n810 ;
  assign n2980 = ( n339 & n1061 ) | ( n339 & ~n2979 ) | ( n1061 & ~n2979 ) ;
  assign n2984 = n2983 ^ n2980 ^ n442 ;
  assign n2985 = n2800 ^ n2135 ^ n1554 ;
  assign n2986 = n2985 ^ n1421 ^ 1'b0 ;
  assign n2987 = n1492 | n2986 ;
  assign n2988 = ( ~n642 & n735 ) | ( ~n642 & n804 ) | ( n735 & n804 ) ;
  assign n2989 = n2988 ^ n2851 ^ 1'b0 ;
  assign n2990 = n2989 ^ n680 ^ 1'b0 ;
  assign n2991 = ( n369 & ~n1346 ) | ( n369 & n2990 ) | ( ~n1346 & n2990 ) ;
  assign n2992 = n1456 ^ n1374 ^ 1'b0 ;
  assign n2993 = ~n2216 & n2992 ;
  assign n2996 = ~n178 & n987 ;
  assign n2997 = n2996 ^ n141 ^ 1'b0 ;
  assign n2998 = ( n2135 & n2142 ) | ( n2135 & ~n2997 ) | ( n2142 & ~n2997 ) ;
  assign n2994 = n1362 & n1647 ;
  assign n2995 = ~n1660 & n2994 ;
  assign n2999 = n2998 ^ n2995 ^ 1'b0 ;
  assign n3003 = ( x90 & n375 ) | ( x90 & ~n1046 ) | ( n375 & ~n1046 ) ;
  assign n3000 = ( n310 & ~n814 ) | ( n310 & n2094 ) | ( ~n814 & n2094 ) ;
  assign n3001 = n3000 ^ n360 ^ 1'b0 ;
  assign n3002 = n1036 | n3001 ;
  assign n3004 = n3003 ^ n3002 ^ 1'b0 ;
  assign n3005 = n219 & ~n333 ;
  assign n3006 = n3005 ^ n2440 ^ n2038 ;
  assign n3007 = ( ~n676 & n767 ) | ( ~n676 & n2752 ) | ( n767 & n2752 ) ;
  assign n3008 = ( n421 & ~n2386 ) | ( n421 & n3007 ) | ( ~n2386 & n3007 ) ;
  assign n3009 = ( n890 & n1153 ) | ( n890 & ~n1373 ) | ( n1153 & ~n1373 ) ;
  assign n3010 = ( n1284 & ~n1542 ) | ( n1284 & n3009 ) | ( ~n1542 & n3009 ) ;
  assign n3011 = n3010 ^ n2555 ^ n999 ;
  assign n3013 = ( n651 & n896 ) | ( n651 & n1539 ) | ( n896 & n1539 ) ;
  assign n3012 = n530 | n2982 ;
  assign n3014 = n3013 ^ n3012 ^ n1015 ;
  assign n3015 = ( n253 & ~n773 ) | ( n253 & n1035 ) | ( ~n773 & n1035 ) ;
  assign n3016 = n3015 ^ n997 ^ 1'b0 ;
  assign n3017 = n1279 & n3016 ;
  assign n3018 = n3017 ^ n497 ^ 1'b0 ;
  assign n3019 = x27 & n511 ;
  assign n3020 = n822 & n3019 ;
  assign n3021 = n651 | n2966 ;
  assign n3022 = ( n224 & ~n3020 ) | ( n224 & n3021 ) | ( ~n3020 & n3021 ) ;
  assign n3023 = ( x79 & ~n448 ) | ( x79 & n924 ) | ( ~n448 & n924 ) ;
  assign n3024 = ( ~n1303 & n2504 ) | ( ~n1303 & n3023 ) | ( n2504 & n3023 ) ;
  assign n3025 = ( x11 & ~n1609 ) | ( x11 & n3024 ) | ( ~n1609 & n3024 ) ;
  assign n3026 = n2916 ^ n1239 ^ n1175 ;
  assign n3027 = n3026 ^ n2411 ^ 1'b0 ;
  assign n3028 = n3025 & ~n3027 ;
  assign n3029 = ~n1818 & n3028 ;
  assign n3030 = ~n1305 & n3029 ;
  assign n3031 = n3030 ^ n425 ^ n392 ;
  assign n3032 = ~n1428 & n3031 ;
  assign n3033 = n1853 ^ n771 ^ n497 ;
  assign n3034 = n1799 ^ n260 ^ 1'b0 ;
  assign n3035 = n3034 ^ n1676 ^ n1102 ;
  assign n3036 = ( ~n1823 & n3033 ) | ( ~n1823 & n3035 ) | ( n3033 & n3035 ) ;
  assign n3037 = n3036 ^ n1806 ^ n337 ;
  assign n3038 = ( n280 & n368 ) | ( n280 & ~n3037 ) | ( n368 & ~n3037 ) ;
  assign n3039 = ( ~x50 & n382 ) | ( ~x50 & n801 ) | ( n382 & n801 ) ;
  assign n3040 = ( n816 & n2140 ) | ( n816 & ~n2835 ) | ( n2140 & ~n2835 ) ;
  assign n3041 = ( n337 & ~n3039 ) | ( n337 & n3040 ) | ( ~n3039 & n3040 ) ;
  assign n3042 = n3041 ^ n202 ^ 1'b0 ;
  assign n3043 = ~n1933 & n3042 ;
  assign n3044 = n3043 ^ n425 ^ 1'b0 ;
  assign n3045 = ( n743 & n804 ) | ( n743 & n1421 ) | ( n804 & n1421 ) ;
  assign n3046 = ( n992 & n1835 ) | ( n992 & n2546 ) | ( n1835 & n2546 ) ;
  assign n3047 = n3045 | n3046 ;
  assign n3048 = ( n596 & n619 ) | ( n596 & ~n1344 ) | ( n619 & ~n1344 ) ;
  assign n3049 = n3048 ^ n1225 ^ x108 ;
  assign n3050 = n2842 ^ n353 ^ 1'b0 ;
  assign n3051 = ( ~n183 & n3049 ) | ( ~n183 & n3050 ) | ( n3049 & n3050 ) ;
  assign n3052 = n582 & n2706 ;
  assign n3053 = n1723 ^ n1504 ^ 1'b0 ;
  assign n3054 = ( n173 & n740 ) | ( n173 & n3053 ) | ( n740 & n3053 ) ;
  assign n3056 = ( n186 & n440 ) | ( n186 & ~n2218 ) | ( n440 & ~n2218 ) ;
  assign n3055 = n1193 | n1703 ;
  assign n3057 = n3056 ^ n3055 ^ 1'b0 ;
  assign n3058 = ( n516 & n735 ) | ( n516 & ~n3057 ) | ( n735 & ~n3057 ) ;
  assign n3059 = ( n573 & n1061 ) | ( n573 & n2483 ) | ( n1061 & n2483 ) ;
  assign n3060 = ( ~n2169 & n2922 ) | ( ~n2169 & n3059 ) | ( n2922 & n3059 ) ;
  assign n3061 = n1220 ^ n1080 ^ 1'b0 ;
  assign n3062 = n3061 ^ n2079 ^ n1747 ;
  assign n3063 = n1453 & ~n3062 ;
  assign n3069 = ( n1000 & n1488 ) | ( n1000 & n2034 ) | ( n1488 & n2034 ) ;
  assign n3068 = n1147 ^ n1119 ^ n704 ;
  assign n3070 = n3069 ^ n3068 ^ 1'b0 ;
  assign n3071 = n345 | n3070 ;
  assign n3072 = n1786 & ~n3071 ;
  assign n3064 = n1383 ^ n1050 ^ x50 ;
  assign n3065 = ~n1217 & n3064 ;
  assign n3066 = n3065 ^ n1852 ^ 1'b0 ;
  assign n3067 = ( x2 & x56 ) | ( x2 & ~n3066 ) | ( x56 & ~n3066 ) ;
  assign n3073 = n3072 ^ n3067 ^ n218 ;
  assign n3074 = ( n2507 & n3063 ) | ( n2507 & ~n3073 ) | ( n3063 & ~n3073 ) ;
  assign n3080 = n1883 ^ n1175 ^ x15 ;
  assign n3079 = n2646 ^ n1928 ^ n1611 ;
  assign n3081 = n3080 ^ n3079 ^ 1'b0 ;
  assign n3082 = ~n255 & n294 ;
  assign n3083 = n2140 ^ n718 ^ 1'b0 ;
  assign n3084 = n3082 & n3083 ;
  assign n3085 = ( x108 & n1114 ) | ( x108 & ~n3084 ) | ( n1114 & ~n3084 ) ;
  assign n3086 = n2047 ^ n989 ^ n919 ;
  assign n3087 = ( ~n774 & n3085 ) | ( ~n774 & n3086 ) | ( n3085 & n3086 ) ;
  assign n3088 = ( n1479 & n1928 ) | ( n1479 & n3087 ) | ( n1928 & n3087 ) ;
  assign n3089 = n3081 | n3088 ;
  assign n3077 = ( n720 & n791 ) | ( n720 & n1139 ) | ( n791 & n1139 ) ;
  assign n3075 = n2868 ^ n304 ^ x68 ;
  assign n3076 = n1731 | n3075 ;
  assign n3078 = n3077 ^ n3076 ^ 1'b0 ;
  assign n3090 = n3089 ^ n3078 ^ n2322 ;
  assign n3091 = n1343 ^ n1279 ^ 1'b0 ;
  assign n3094 = ( n309 & ~n2275 ) | ( n309 & n2533 ) | ( ~n2275 & n2533 ) ;
  assign n3095 = ( ~n287 & n317 ) | ( ~n287 & n3094 ) | ( n317 & n3094 ) ;
  assign n3096 = n714 ^ x10 ^ 1'b0 ;
  assign n3097 = ( ~n2576 & n3095 ) | ( ~n2576 & n3096 ) | ( n3095 & n3096 ) ;
  assign n3098 = ( n2171 & n2858 ) | ( n2171 & n3097 ) | ( n2858 & n3097 ) ;
  assign n3092 = n2174 ^ n567 ^ x12 ;
  assign n3093 = ( n580 & n1351 ) | ( n580 & ~n3092 ) | ( n1351 & ~n3092 ) ;
  assign n3099 = n3098 ^ n3093 ^ n508 ;
  assign n3102 = n1801 ^ n1510 ^ n1224 ;
  assign n3103 = n814 & n3102 ;
  assign n3100 = ( ~n1209 & n1270 ) | ( ~n1209 & n2787 ) | ( n1270 & n2787 ) ;
  assign n3101 = ( n1414 & n3086 ) | ( n1414 & ~n3100 ) | ( n3086 & ~n3100 ) ;
  assign n3104 = n3103 ^ n3101 ^ n580 ;
  assign n3110 = n557 & ~n2157 ;
  assign n3113 = n1752 ^ n656 ^ 1'b0 ;
  assign n3114 = n2554 & n3113 ;
  assign n3115 = n3114 ^ n1356 ^ 1'b0 ;
  assign n3111 = ( ~n1017 & n1388 ) | ( ~n1017 & n2717 ) | ( n1388 & n2717 ) ;
  assign n3112 = ( n2599 & n2716 ) | ( n2599 & ~n3111 ) | ( n2716 & ~n3111 ) ;
  assign n3116 = n3115 ^ n3112 ^ 1'b0 ;
  assign n3117 = ~n3110 & n3116 ;
  assign n3105 = n586 ^ n383 ^ n323 ;
  assign n3106 = n3105 ^ n2089 ^ n858 ;
  assign n3107 = n3106 ^ n1633 ^ 1'b0 ;
  assign n3108 = n2714 ^ n2240 ^ n163 ;
  assign n3109 = ( n347 & n3107 ) | ( n347 & n3108 ) | ( n3107 & n3108 ) ;
  assign n3118 = n3117 ^ n3109 ^ n430 ;
  assign n3126 = ( ~x13 & n426 ) | ( ~x13 & n1431 ) | ( n426 & n1431 ) ;
  assign n3125 = ~n579 & n1463 ;
  assign n3127 = n3126 ^ n3125 ^ 1'b0 ;
  assign n3124 = ( n464 & n1536 ) | ( n464 & n1545 ) | ( n1536 & n1545 ) ;
  assign n3128 = n3127 ^ n3124 ^ n1892 ;
  assign n3120 = ( x68 & n627 ) | ( x68 & n2458 ) | ( n627 & n2458 ) ;
  assign n3121 = ( n261 & n2506 ) | ( n261 & n3120 ) | ( n2506 & n3120 ) ;
  assign n3119 = ( n676 & ~n811 ) | ( n676 & n881 ) | ( ~n811 & n881 ) ;
  assign n3122 = n3121 ^ n3119 ^ n1581 ;
  assign n3123 = n1150 | n3122 ;
  assign n3129 = n3128 ^ n3123 ^ 1'b0 ;
  assign n3130 = ( x18 & n1567 ) | ( x18 & ~n2231 ) | ( n1567 & ~n2231 ) ;
  assign n3131 = ( n738 & n849 ) | ( n738 & ~n1773 ) | ( n849 & ~n1773 ) ;
  assign n3132 = n2129 & ~n3131 ;
  assign n3133 = n3132 ^ n3025 ^ 1'b0 ;
  assign n3134 = n3133 ^ n1575 ^ n1125 ;
  assign n3135 = ( ~x20 & x55 ) | ( ~x20 & x100 ) | ( x55 & x100 ) ;
  assign n3136 = ( ~x83 & n549 ) | ( ~x83 & n3135 ) | ( n549 & n3135 ) ;
  assign n3137 = ( n554 & n1827 ) | ( n554 & ~n2259 ) | ( n1827 & ~n2259 ) ;
  assign n3138 = ( ~n149 & n1981 ) | ( ~n149 & n2130 ) | ( n1981 & n2130 ) ;
  assign n3139 = ( n263 & n906 ) | ( n263 & n1705 ) | ( n906 & n1705 ) ;
  assign n3140 = n1789 | n3139 ;
  assign n3141 = ( ~n3137 & n3138 ) | ( ~n3137 & n3140 ) | ( n3138 & n3140 ) ;
  assign n3142 = ( x107 & n483 ) | ( x107 & ~n992 ) | ( n483 & ~n992 ) ;
  assign n3143 = ( n598 & n1093 ) | ( n598 & ~n3142 ) | ( n1093 & ~n3142 ) ;
  assign n3144 = ( n3136 & n3141 ) | ( n3136 & ~n3143 ) | ( n3141 & ~n3143 ) ;
  assign n3145 = ( n1095 & n1496 ) | ( n1095 & n3144 ) | ( n1496 & n3144 ) ;
  assign n3146 = n1908 ^ n1480 ^ n1420 ;
  assign n3147 = ( n806 & n1019 ) | ( n806 & ~n1594 ) | ( n1019 & ~n1594 ) ;
  assign n3148 = n3147 ^ n502 ^ 1'b0 ;
  assign n3149 = x44 & n3148 ;
  assign n3150 = n3146 & n3149 ;
  assign n3151 = n669 ^ n487 ^ 1'b0 ;
  assign n3152 = n2047 ^ n1775 ^ n1394 ;
  assign n3153 = ( ~n1163 & n3151 ) | ( ~n1163 & n3152 ) | ( n3151 & n3152 ) ;
  assign n3154 = ( n1195 & n2480 ) | ( n1195 & ~n2924 ) | ( n2480 & ~n2924 ) ;
  assign n3155 = n3154 ^ n2022 ^ n1844 ;
  assign n3156 = n1614 ^ n1107 ^ n915 ;
  assign n3157 = n3156 ^ n1292 ^ 1'b0 ;
  assign n3158 = ( ~n1800 & n3155 ) | ( ~n1800 & n3157 ) | ( n3155 & n3157 ) ;
  assign n3159 = n984 & n2706 ;
  assign n3160 = n3159 ^ n3086 ^ 1'b0 ;
  assign n3161 = ( n1774 & n2840 ) | ( n1774 & n3160 ) | ( n2840 & n3160 ) ;
  assign n3166 = n374 | n1148 ;
  assign n3167 = n3166 ^ n1300 ^ 1'b0 ;
  assign n3168 = n1413 & n3167 ;
  assign n3162 = ( ~x51 & n417 ) | ( ~x51 & n1557 ) | ( n417 & n1557 ) ;
  assign n3163 = x74 & ~n3162 ;
  assign n3164 = n3163 ^ n2640 ^ 1'b0 ;
  assign n3165 = n3164 ^ n1718 ^ n228 ;
  assign n3169 = n3168 ^ n3165 ^ 1'b0 ;
  assign n3170 = n3161 & n3169 ;
  assign n3171 = n2589 ^ n228 ^ n148 ;
  assign n3172 = ( n1076 & n2181 ) | ( n1076 & n3171 ) | ( n2181 & n3171 ) ;
  assign n3173 = n315 ^ x40 ^ x7 ;
  assign n3174 = n3173 ^ n3015 ^ n1551 ;
  assign n3175 = n321 | n3174 ;
  assign n3179 = ( x26 & ~n1049 ) | ( x26 & n2372 ) | ( ~n1049 & n2372 ) ;
  assign n3180 = ( ~n611 & n1196 ) | ( ~n611 & n1633 ) | ( n1196 & n1633 ) ;
  assign n3181 = ~n813 & n1419 ;
  assign n3182 = n3181 ^ n1182 ^ 1'b0 ;
  assign n3183 = n3182 ^ n447 ^ 1'b0 ;
  assign n3184 = n3180 & ~n3183 ;
  assign n3185 = ( n2374 & n3179 ) | ( n2374 & n3184 ) | ( n3179 & n3184 ) ;
  assign n3176 = n3013 ^ n1592 ^ n1356 ;
  assign n3177 = n1181 ^ n719 ^ 1'b0 ;
  assign n3178 = n3176 | n3177 ;
  assign n3186 = n3185 ^ n3178 ^ n3025 ;
  assign n3187 = ( n3172 & ~n3175 ) | ( n3172 & n3186 ) | ( ~n3175 & n3186 ) ;
  assign n3188 = ( n579 & n1248 ) | ( n579 & ~n2729 ) | ( n1248 & ~n2729 ) ;
  assign n3189 = n1383 & n3188 ;
  assign n3190 = n3189 ^ n3053 ^ x40 ;
  assign n3191 = ( n634 & ~n2572 ) | ( n634 & n3190 ) | ( ~n2572 & n3190 ) ;
  assign n3204 = n2531 ^ n344 ^ x93 ;
  assign n3194 = n2809 ^ x91 ^ 1'b0 ;
  assign n3195 = ~n2123 & n3194 ;
  assign n3193 = n613 ^ n595 ^ n425 ;
  assign n3192 = ( n1032 & n1117 ) | ( n1032 & n1264 ) | ( n1117 & n1264 ) ;
  assign n3196 = n3195 ^ n3193 ^ n3192 ;
  assign n3198 = ~n517 & n976 ;
  assign n3199 = n3198 ^ n783 ^ n582 ;
  assign n3200 = n3199 ^ n2555 ^ n756 ;
  assign n3197 = ( n1490 & n1798 ) | ( n1490 & n2222 ) | ( n1798 & n2222 ) ;
  assign n3201 = n3200 ^ n3197 ^ n661 ;
  assign n3202 = n3196 & ~n3201 ;
  assign n3203 = n417 & n3202 ;
  assign n3205 = n3204 ^ n3203 ^ n909 ;
  assign n3206 = n2923 ^ n1186 ^ n640 ;
  assign n3207 = n3206 ^ n1831 ^ 1'b0 ;
  assign n3208 = ( ~n572 & n2575 ) | ( ~n572 & n3207 ) | ( n2575 & n3207 ) ;
  assign n3209 = n3208 ^ n2631 ^ n1380 ;
  assign n3210 = ~n449 & n1504 ;
  assign n3212 = n1006 ^ n878 ^ n402 ;
  assign n3213 = ( n936 & ~n2089 ) | ( n936 & n3212 ) | ( ~n2089 & n3212 ) ;
  assign n3214 = n3213 ^ n1592 ^ n1136 ;
  assign n3211 = x38 & n2576 ;
  assign n3215 = n3214 ^ n3211 ^ 1'b0 ;
  assign n3216 = ( n2377 & n3210 ) | ( n2377 & n3215 ) | ( n3210 & n3215 ) ;
  assign n3230 = n731 ^ n588 ^ 1'b0 ;
  assign n3229 = n1226 ^ n692 ^ n176 ;
  assign n3231 = n3230 ^ n3229 ^ n678 ;
  assign n3217 = ( ~n197 & n676 ) | ( ~n197 & n838 ) | ( n676 & n838 ) ;
  assign n3218 = ( n215 & ~n281 ) | ( n215 & n977 ) | ( ~n281 & n977 ) ;
  assign n3222 = ( n480 & n560 ) | ( n480 & n579 ) | ( n560 & n579 ) ;
  assign n3223 = n2119 ^ n1853 ^ 1'b0 ;
  assign n3224 = n3222 | n3223 ;
  assign n3219 = ( ~n761 & n1449 ) | ( ~n761 & n1515 ) | ( n1449 & n1515 ) ;
  assign n3220 = n214 | n2292 ;
  assign n3221 = ( ~n2311 & n3219 ) | ( ~n2311 & n3220 ) | ( n3219 & n3220 ) ;
  assign n3225 = n3224 ^ n3221 ^ 1'b0 ;
  assign n3226 = n3225 ^ n1112 ^ n814 ;
  assign n3227 = n3226 ^ n787 ^ n178 ;
  assign n3228 = ( ~n3217 & n3218 ) | ( ~n3217 & n3227 ) | ( n3218 & n3227 ) ;
  assign n3232 = n3231 ^ n3228 ^ n1938 ;
  assign n3242 = n846 ^ n276 ^ x103 ;
  assign n3243 = n1135 ^ n672 ^ n601 ;
  assign n3244 = ( x26 & ~n3242 ) | ( x26 & n3243 ) | ( ~n3242 & n3243 ) ;
  assign n3239 = n1530 ^ x84 ^ 1'b0 ;
  assign n3240 = n1745 & ~n3239 ;
  assign n3237 = x36 | n1655 ;
  assign n3233 = ( x17 & n256 ) | ( x17 & ~n2750 ) | ( n256 & ~n2750 ) ;
  assign n3234 = n1822 | n3233 ;
  assign n3235 = n3234 ^ n2190 ^ 1'b0 ;
  assign n3236 = n3235 ^ n1561 ^ n331 ;
  assign n3238 = n3237 ^ n3236 ^ 1'b0 ;
  assign n3241 = n3240 ^ n3238 ^ n2523 ;
  assign n3245 = n3244 ^ n3241 ^ 1'b0 ;
  assign n3246 = n590 | n3245 ;
  assign n3247 = n1003 ^ n171 ^ 1'b0 ;
  assign n3248 = ( n398 & n985 ) | ( n398 & n2215 ) | ( n985 & n2215 ) ;
  assign n3249 = n3248 ^ n2873 ^ n1292 ;
  assign n3250 = n3249 ^ n184 ^ 1'b0 ;
  assign n3251 = ( n1394 & ~n1799 ) | ( n1394 & n2066 ) | ( ~n1799 & n2066 ) ;
  assign n3252 = n3251 ^ n2722 ^ n2561 ;
  assign n3253 = n370 & ~n1625 ;
  assign n3254 = n2630 ^ n1159 ^ n438 ;
  assign n3255 = ( ~x119 & n2151 ) | ( ~x119 & n3254 ) | ( n2151 & n3254 ) ;
  assign n3256 = n1019 ^ n1000 ^ x17 ;
  assign n3257 = ~n1407 & n3256 ;
  assign n3259 = ( ~n1329 & n2352 ) | ( ~n1329 & n3005 ) | ( n2352 & n3005 ) ;
  assign n3260 = ( n1266 & ~n2643 ) | ( n1266 & n3259 ) | ( ~n2643 & n3259 ) ;
  assign n3258 = n3094 ^ n974 ^ 1'b0 ;
  assign n3261 = n3260 ^ n3258 ^ n3165 ;
  assign n3262 = ~n3257 & n3261 ;
  assign n3263 = ( n599 & ~n1054 ) | ( n599 & n1887 ) | ( ~n1054 & n1887 ) ;
  assign n3264 = ( ~n912 & n1320 ) | ( ~n912 & n2839 ) | ( n1320 & n2839 ) ;
  assign n3265 = n1641 & n3264 ;
  assign n3266 = ~n1610 & n3265 ;
  assign n3267 = n2910 ^ n923 ^ n683 ;
  assign n3268 = n2685 ^ n833 ^ n655 ;
  assign n3269 = ( n1062 & n3267 ) | ( n1062 & ~n3268 ) | ( n3267 & ~n3268 ) ;
  assign n3270 = ( n3263 & n3266 ) | ( n3263 & ~n3269 ) | ( n3266 & ~n3269 ) ;
  assign n3271 = n3270 ^ n2232 ^ n477 ;
  assign n3272 = ( n466 & ~n637 ) | ( n466 & n1977 ) | ( ~n637 & n1977 ) ;
  assign n3273 = ( n655 & n1315 ) | ( n655 & ~n3272 ) | ( n1315 & ~n3272 ) ;
  assign n3274 = n3057 & n3273 ;
  assign n3275 = n3271 & n3274 ;
  assign n3276 = n2181 ^ n1895 ^ 1'b0 ;
  assign n3277 = ~n175 & n631 ;
  assign n3278 = ( n3011 & n3276 ) | ( n3011 & n3277 ) | ( n3276 & n3277 ) ;
  assign n3287 = ( ~n154 & n236 ) | ( ~n154 & n739 ) | ( n236 & n739 ) ;
  assign n3288 = ( n1542 & n1577 ) | ( n1542 & n3287 ) | ( n1577 & n3287 ) ;
  assign n3284 = n168 & n3135 ;
  assign n3285 = n1324 & n3284 ;
  assign n3286 = n3285 ^ n959 ^ n298 ;
  assign n3279 = n1910 ^ n780 ^ n406 ;
  assign n3280 = n2557 | n3279 ;
  assign n3281 = n568 & ~n3280 ;
  assign n3282 = n3281 ^ n2396 ^ 1'b0 ;
  assign n3283 = n903 & n3282 ;
  assign n3289 = n3288 ^ n3286 ^ n3283 ;
  assign n3290 = n2073 ^ n872 ^ x5 ;
  assign n3291 = ~n607 & n1239 ;
  assign n3292 = n3291 ^ n1660 ^ n1284 ;
  assign n3293 = n1800 ^ n1781 ^ n1284 ;
  assign n3294 = n3146 ^ n1210 ^ n1125 ;
  assign n3295 = ( n1231 & n3293 ) | ( n1231 & ~n3294 ) | ( n3293 & ~n3294 ) ;
  assign n3297 = n2916 ^ n2671 ^ n1271 ;
  assign n3296 = n2480 ^ n2392 ^ n2235 ;
  assign n3298 = n3297 ^ n3296 ^ 1'b0 ;
  assign n3299 = n238 | n3298 ;
  assign n3300 = n2666 ^ n2453 ^ 1'b0 ;
  assign n3301 = ~n627 & n3300 ;
  assign n3302 = n3301 ^ n421 ^ 1'b0 ;
  assign n3303 = n3302 ^ n2733 ^ n1876 ;
  assign n3311 = n2105 ^ n1781 ^ 1'b0 ;
  assign n3312 = n3040 ^ n2259 ^ 1'b0 ;
  assign n3313 = n3311 & ~n3312 ;
  assign n3309 = ( n575 & n860 ) | ( n575 & n1093 ) | ( n860 & n1093 ) ;
  assign n3308 = n1047 ^ n639 ^ n524 ;
  assign n3307 = ( n147 & n1497 ) | ( n147 & ~n2047 ) | ( n1497 & ~n2047 ) ;
  assign n3310 = n3309 ^ n3308 ^ n3307 ;
  assign n3304 = n1503 ^ n445 ^ n176 ;
  assign n3305 = n3304 ^ n3279 ^ n2285 ;
  assign n3306 = n1695 & n3305 ;
  assign n3314 = n3313 ^ n3310 ^ n3306 ;
  assign n3317 = n2531 ^ n1528 ^ n456 ;
  assign n3315 = ~n1230 & n2469 ;
  assign n3316 = n3315 ^ n2245 ^ n337 ;
  assign n3318 = n3317 ^ n3316 ^ n2827 ;
  assign n3319 = ( n740 & n1188 ) | ( n740 & n3318 ) | ( n1188 & n3318 ) ;
  assign n3320 = n3319 ^ n2198 ^ n236 ;
  assign n3321 = n586 | n3320 ;
  assign n3322 = ( x127 & ~n1480 ) | ( x127 & n2049 ) | ( ~n1480 & n2049 ) ;
  assign n3323 = n3322 ^ n1184 ^ n1100 ;
  assign n3324 = n1867 ^ x4 ^ 1'b0 ;
  assign n3326 = n944 | n1787 ;
  assign n3327 = n879 | n3326 ;
  assign n3325 = n2720 ^ n1939 ^ n239 ;
  assign n3328 = n3327 ^ n3325 ^ 1'b0 ;
  assign n3329 = ( n1864 & ~n2287 ) | ( n1864 & n2818 ) | ( ~n2287 & n2818 ) ;
  assign n3334 = n501 ^ n318 ^ x81 ;
  assign n3335 = n293 ^ x53 ^ x8 ;
  assign n3336 = n3335 ^ n1233 ^ 1'b0 ;
  assign n3337 = ( n769 & n3334 ) | ( n769 & n3336 ) | ( n3334 & n3336 ) ;
  assign n3338 = n2121 | n3337 ;
  assign n3339 = n3338 ^ n2237 ^ n675 ;
  assign n3330 = ( n1016 & n1788 ) | ( n1016 & n2851 ) | ( n1788 & n2851 ) ;
  assign n3331 = n2348 ^ n786 ^ n148 ;
  assign n3332 = n3331 ^ n1265 ^ 1'b0 ;
  assign n3333 = n3330 & n3332 ;
  assign n3340 = n3339 ^ n3333 ^ 1'b0 ;
  assign n3341 = ( ~n1704 & n1949 ) | ( ~n1704 & n3131 ) | ( n1949 & n3131 ) ;
  assign n3342 = n3341 ^ n2892 ^ n370 ;
  assign n3343 = x109 & ~n3342 ;
  assign n3344 = n3343 ^ n2229 ^ 1'b0 ;
  assign n3345 = n3344 ^ n826 ^ 1'b0 ;
  assign n3346 = ( ~n2464 & n3340 ) | ( ~n2464 & n3345 ) | ( n3340 & n3345 ) ;
  assign n3347 = n1032 & n2188 ;
  assign n3348 = n553 & n3347 ;
  assign n3349 = ~n607 & n1593 ;
  assign n3350 = ( n258 & n712 ) | ( n258 & ~n1030 ) | ( n712 & ~n1030 ) ;
  assign n3351 = n3350 ^ n1030 ^ 1'b0 ;
  assign n3352 = n2856 & n3351 ;
  assign n3353 = ~n689 & n2068 ;
  assign n3361 = n2844 ^ n2171 ^ n1611 ;
  assign n3360 = ( n298 & n462 ) | ( n298 & n2633 ) | ( n462 & n2633 ) ;
  assign n3354 = ( x7 & ~n1917 ) | ( x7 & n3121 ) | ( ~n1917 & n3121 ) ;
  assign n3355 = n683 | n3354 ;
  assign n3356 = ( ~n1332 & n2140 ) | ( ~n1332 & n3355 ) | ( n2140 & n3355 ) ;
  assign n3357 = n3356 ^ n2524 ^ n362 ;
  assign n3358 = n3357 ^ n609 ^ 1'b0 ;
  assign n3359 = n2789 & n3358 ;
  assign n3362 = n3361 ^ n3360 ^ n3359 ;
  assign n3363 = ( n315 & ~n538 ) | ( n315 & n1828 ) | ( ~n538 & n1828 ) ;
  assign n3364 = ( ~n764 & n1410 ) | ( ~n764 & n3363 ) | ( n1410 & n3363 ) ;
  assign n3376 = n805 ^ n404 ^ n309 ;
  assign n3377 = n806 | n3376 ;
  assign n3371 = ( n804 & n1129 ) | ( n804 & ~n1488 ) | ( n1129 & ~n1488 ) ;
  assign n3372 = n1544 ^ n906 ^ 1'b0 ;
  assign n3373 = ( n407 & ~n3371 ) | ( n407 & n3372 ) | ( ~n3371 & n3372 ) ;
  assign n3374 = ( ~n1000 & n1163 ) | ( ~n1000 & n2778 ) | ( n1163 & n2778 ) ;
  assign n3375 = ( n1920 & n3373 ) | ( n1920 & ~n3374 ) | ( n3373 & ~n3374 ) ;
  assign n3365 = x78 & n1214 ;
  assign n3366 = n991 ^ n963 ^ 1'b0 ;
  assign n3367 = n386 & n3366 ;
  assign n3368 = n3367 ^ n1153 ^ n993 ;
  assign n3369 = n3048 ^ n2744 ^ 1'b0 ;
  assign n3370 = ( n3365 & ~n3368 ) | ( n3365 & n3369 ) | ( ~n3368 & n3369 ) ;
  assign n3378 = n3377 ^ n3375 ^ n3370 ;
  assign n3379 = n1126 | n2033 ;
  assign n3383 = n417 | n2002 ;
  assign n3384 = n3383 ^ n649 ^ 1'b0 ;
  assign n3385 = ( n1637 & ~n2770 ) | ( n1637 & n3384 ) | ( ~n2770 & n3384 ) ;
  assign n3380 = n2279 ^ n184 ^ 1'b0 ;
  assign n3381 = n1051 | n3380 ;
  assign n3382 = n3381 ^ n2799 ^ 1'b0 ;
  assign n3386 = n3385 ^ n3382 ^ n908 ;
  assign n3387 = ( n2767 & n3379 ) | ( n2767 & n3386 ) | ( n3379 & n3386 ) ;
  assign n3396 = n2420 ^ n1938 ^ n991 ;
  assign n3394 = n1702 ^ n543 ^ 1'b0 ;
  assign n3395 = ~n209 & n3394 ;
  assign n3397 = n3396 ^ n3395 ^ n1398 ;
  assign n3388 = n969 | n1510 ;
  assign n3389 = n3388 ^ n1071 ^ 1'b0 ;
  assign n3390 = n3389 ^ n398 ^ 1'b0 ;
  assign n3391 = n1007 | n3390 ;
  assign n3392 = ( n1241 & n2064 ) | ( n1241 & ~n3391 ) | ( n2064 & ~n3391 ) ;
  assign n3393 = ~n413 & n3392 ;
  assign n3398 = n3397 ^ n3393 ^ 1'b0 ;
  assign n3399 = n182 | n626 ;
  assign n3400 = n3399 ^ n2626 ^ 1'b0 ;
  assign n3401 = n2907 ^ n595 ^ 1'b0 ;
  assign n3402 = n3400 | n3401 ;
  assign n3403 = n949 & ~n1261 ;
  assign n3404 = ~n1728 & n3403 ;
  assign n3405 = ~n1273 & n3404 ;
  assign n3406 = ( n240 & ~n2754 ) | ( n240 & n3023 ) | ( ~n2754 & n3023 ) ;
  assign n3408 = n1263 ^ n1180 ^ 1'b0 ;
  assign n3409 = n2049 & n3408 ;
  assign n3407 = ~n1263 & n2270 ;
  assign n3410 = n3409 ^ n3407 ^ 1'b0 ;
  assign n3411 = ~n3406 & n3410 ;
  assign n3412 = n3119 ^ n645 ^ 1'b0 ;
  assign n3413 = ~n1335 & n3412 ;
  assign n3414 = n1406 ^ n880 ^ 1'b0 ;
  assign n3415 = n528 & ~n3414 ;
  assign n3416 = ~n778 & n3415 ;
  assign n3417 = ( n246 & ~n616 ) | ( n246 & n3416 ) | ( ~n616 & n3416 ) ;
  assign n3418 = n3417 ^ n2568 ^ n1716 ;
  assign n3422 = ~n2047 & n2941 ;
  assign n3419 = ( n655 & ~n1493 ) | ( n655 & n2554 ) | ( ~n1493 & n2554 ) ;
  assign n3420 = n1938 ^ n1937 ^ n861 ;
  assign n3421 = n3419 & ~n3420 ;
  assign n3423 = n3422 ^ n3421 ^ 1'b0 ;
  assign n3424 = n2174 ^ n2028 ^ n451 ;
  assign n3425 = ( ~n394 & n591 ) | ( ~n394 & n1384 ) | ( n591 & n1384 ) ;
  assign n3426 = n2869 ^ n2459 ^ n892 ;
  assign n3427 = n194 | n3426 ;
  assign n3428 = ( n3316 & ~n3425 ) | ( n3316 & n3427 ) | ( ~n3425 & n3427 ) ;
  assign n3429 = x16 | n2287 ;
  assign n3430 = ( n944 & n1765 ) | ( n944 & n3429 ) | ( n1765 & n3429 ) ;
  assign n3431 = n2493 & n3430 ;
  assign n3432 = ~n3428 & n3431 ;
  assign n3433 = ( n748 & n3424 ) | ( n748 & n3432 ) | ( n3424 & n3432 ) ;
  assign n3434 = ( n597 & n3423 ) | ( n597 & n3433 ) | ( n3423 & n3433 ) ;
  assign n3437 = n2360 ^ n849 ^ n411 ;
  assign n3435 = ( x15 & n677 ) | ( x15 & ~n712 ) | ( n677 & ~n712 ) ;
  assign n3436 = n3435 ^ n3337 ^ 1'b0 ;
  assign n3438 = n3437 ^ n3436 ^ 1'b0 ;
  assign n3439 = n3434 & ~n3438 ;
  assign n3440 = n616 & ~n2704 ;
  assign n3441 = n3440 ^ n1476 ^ 1'b0 ;
  assign n3442 = ( n1806 & n3135 ) | ( n1806 & ~n3441 ) | ( n3135 & ~n3441 ) ;
  assign n3443 = n3442 ^ n2283 ^ n2268 ;
  assign n3451 = n3061 ^ n207 ^ n157 ;
  assign n3452 = ( ~n1661 & n3164 ) | ( ~n1661 & n3451 ) | ( n3164 & n3451 ) ;
  assign n3448 = n249 & n1403 ;
  assign n3449 = ~n1225 & n3448 ;
  assign n3450 = ( n2932 & n3120 ) | ( n2932 & n3449 ) | ( n3120 & n3449 ) ;
  assign n3444 = ( ~n1957 & n2478 ) | ( ~n1957 & n2619 ) | ( n2478 & n2619 ) ;
  assign n3445 = ( n620 & n2025 ) | ( n620 & n3444 ) | ( n2025 & n3444 ) ;
  assign n3446 = n1654 & n2810 ;
  assign n3447 = ~n3445 & n3446 ;
  assign n3453 = n3452 ^ n3450 ^ n3447 ;
  assign n3454 = n2685 ^ n2604 ^ n536 ;
  assign n3455 = n2422 ^ n1534 ^ n177 ;
  assign n3456 = n497 & n3455 ;
  assign n3457 = ~n3454 & n3456 ;
  assign n3458 = ~n420 & n1813 ;
  assign n3459 = n3458 ^ n2830 ^ n2086 ;
  assign n3460 = ( x109 & ~n2038 ) | ( x109 & n2554 ) | ( ~n2038 & n2554 ) ;
  assign n3461 = ( n3243 & ~n3337 ) | ( n3243 & n3460 ) | ( ~n3337 & n3460 ) ;
  assign n3462 = ~n882 & n3461 ;
  assign n3463 = ( n272 & n505 ) | ( n272 & n2477 ) | ( n505 & n2477 ) ;
  assign n3464 = n3463 ^ n2446 ^ n2053 ;
  assign n3465 = ~n176 & n349 ;
  assign n3466 = ~n1246 & n3465 ;
  assign n3467 = n1411 ^ n1281 ^ n842 ;
  assign n3468 = ( n208 & n716 ) | ( n208 & ~n2502 ) | ( n716 & ~n2502 ) ;
  assign n3469 = ( n3466 & n3467 ) | ( n3466 & ~n3468 ) | ( n3467 & ~n3468 ) ;
  assign n3472 = ( x98 & ~n1456 ) | ( x98 & n1518 ) | ( ~n1456 & n1518 ) ;
  assign n3470 = n1485 ^ n1108 ^ n413 ;
  assign n3471 = ( n187 & n2157 ) | ( n187 & n3470 ) | ( n2157 & n3470 ) ;
  assign n3473 = n3472 ^ n3471 ^ n2395 ;
  assign n3474 = ~n1254 & n3473 ;
  assign n3475 = n2033 & n3474 ;
  assign n3476 = x64 & n878 ;
  assign n3477 = n3476 ^ n263 ^ 1'b0 ;
  assign n3478 = ( ~n2201 & n3315 ) | ( ~n2201 & n3477 ) | ( n3315 & n3477 ) ;
  assign n3479 = n3153 | n3478 ;
  assign n3480 = ( n255 & n1351 ) | ( n255 & ~n2473 ) | ( n1351 & ~n2473 ) ;
  assign n3481 = n521 & ~n3480 ;
  assign n3491 = ( ~x119 & n2741 ) | ( ~x119 & n3374 ) | ( n2741 & n3374 ) ;
  assign n3492 = ( ~x36 & n1347 ) | ( ~x36 & n3491 ) | ( n1347 & n3491 ) ;
  assign n3482 = n2199 ^ n305 ^ 1'b0 ;
  assign n3483 = n3172 | n3482 ;
  assign n3484 = ( ~n1036 & n1210 ) | ( ~n1036 & n3483 ) | ( n1210 & n3483 ) ;
  assign n3485 = n668 ^ n554 ^ n391 ;
  assign n3486 = n3485 ^ n2718 ^ n2499 ;
  assign n3487 = ( n501 & n958 ) | ( n501 & n3486 ) | ( n958 & n3486 ) ;
  assign n3488 = n3487 ^ n1117 ^ n868 ;
  assign n3489 = n3488 ^ n3158 ^ 1'b0 ;
  assign n3490 = n3484 & ~n3489 ;
  assign n3493 = n3492 ^ n3490 ^ 1'b0 ;
  assign n3494 = n2183 & n3304 ;
  assign n3496 = ( n1024 & ~n1193 ) | ( n1024 & n1281 ) | ( ~n1193 & n1281 ) ;
  assign n3495 = ~n634 & n1268 ;
  assign n3497 = n3496 ^ n3495 ^ n1990 ;
  assign n3498 = n1481 & ~n1841 ;
  assign n3499 = n3172 ^ n2885 ^ n418 ;
  assign n3500 = ( n187 & n717 ) | ( n187 & ~n3499 ) | ( n717 & ~n3499 ) ;
  assign n3501 = n2635 | n3500 ;
  assign n3502 = n3498 & ~n3501 ;
  assign n3503 = ( n759 & n2456 ) | ( n759 & ~n3502 ) | ( n2456 & ~n3502 ) ;
  assign n3508 = n276 ^ x63 ^ 1'b0 ;
  assign n3504 = n293 & ~n921 ;
  assign n3505 = n3504 ^ x30 ^ 1'b0 ;
  assign n3506 = n1810 ^ n325 ^ 1'b0 ;
  assign n3507 = ~n3505 & n3506 ;
  assign n3509 = n3508 ^ n3507 ^ 1'b0 ;
  assign n3510 = n2475 ^ n1667 ^ n1423 ;
  assign n3511 = n3510 ^ n2542 ^ n1663 ;
  assign n3517 = x95 & n2676 ;
  assign n3518 = n1097 & n3517 ;
  assign n3512 = n2064 ^ n1141 ^ n216 ;
  assign n3513 = ( ~n1458 & n3112 ) | ( ~n1458 & n3512 ) | ( n3112 & n3512 ) ;
  assign n3514 = ~n1781 & n2425 ;
  assign n3515 = n1326 & n1752 ;
  assign n3516 = ( n3513 & n3514 ) | ( n3513 & n3515 ) | ( n3514 & n3515 ) ;
  assign n3519 = n3518 ^ n3516 ^ n2100 ;
  assign n3522 = n1904 ^ n786 ^ x48 ;
  assign n3520 = ( n425 & ~n1403 ) | ( n425 & n2851 ) | ( ~n1403 & n2851 ) ;
  assign n3521 = n3049 | n3520 ;
  assign n3523 = n3522 ^ n3521 ^ n1833 ;
  assign n3524 = ( n1606 & ~n2042 ) | ( n1606 & n3523 ) | ( ~n2042 & n3523 ) ;
  assign n3525 = n447 ^ n196 ^ 1'b0 ;
  assign n3526 = ( n597 & ~n1131 ) | ( n597 & n3525 ) | ( ~n1131 & n3525 ) ;
  assign n3527 = n3526 ^ n859 ^ 1'b0 ;
  assign n3528 = ~n290 & n3527 ;
  assign n3529 = ~n2639 & n3528 ;
  assign n3530 = ( n2007 & n3524 ) | ( n2007 & ~n3529 ) | ( n3524 & ~n3529 ) ;
  assign n3531 = ( x51 & ~n3070 ) | ( x51 & n3133 ) | ( ~n3070 & n3133 ) ;
  assign n3532 = n3531 ^ n3232 ^ 1'b0 ;
  assign n3535 = n1504 ^ n773 ^ n135 ;
  assign n3536 = n3535 ^ n1394 ^ n244 ;
  assign n3533 = n1600 ^ x85 ^ 1'b0 ;
  assign n3534 = n3266 | n3533 ;
  assign n3537 = n3536 ^ n3534 ^ n981 ;
  assign n3552 = ( ~n282 & n1289 ) | ( ~n282 & n2982 ) | ( n1289 & n2982 ) ;
  assign n3548 = n294 & ~n676 ;
  assign n3549 = n3548 ^ n1464 ^ 1'b0 ;
  assign n3538 = n1369 ^ n1014 ^ n745 ;
  assign n3539 = n815 ^ n161 ^ n153 ;
  assign n3540 = n1787 ^ n499 ^ n347 ;
  assign n3541 = n1374 ^ n956 ^ 1'b0 ;
  assign n3542 = ( n130 & n886 ) | ( n130 & n3541 ) | ( n886 & n3541 ) ;
  assign n3543 = ( n732 & ~n784 ) | ( n732 & n3542 ) | ( ~n784 & n3542 ) ;
  assign n3544 = n1669 & ~n3543 ;
  assign n3545 = ~n3540 & n3544 ;
  assign n3546 = ( ~n1490 & n3539 ) | ( ~n1490 & n3545 ) | ( n3539 & n3545 ) ;
  assign n3547 = ( n2189 & ~n3538 ) | ( n2189 & n3546 ) | ( ~n3538 & n3546 ) ;
  assign n3550 = n3549 ^ n3547 ^ n1343 ;
  assign n3551 = ( ~n1276 & n2733 ) | ( ~n1276 & n3550 ) | ( n2733 & n3550 ) ;
  assign n3553 = n3552 ^ n3551 ^ n1860 ;
  assign n3554 = ~n3537 & n3553 ;
  assign n3555 = ( n921 & n1422 ) | ( n921 & n1625 ) | ( n1422 & n1625 ) ;
  assign n3556 = n3555 ^ n3192 ^ 1'b0 ;
  assign n3557 = n2634 & ~n3556 ;
  assign n3558 = ( n1940 & n2340 ) | ( n1940 & ~n3515 ) | ( n2340 & ~n3515 ) ;
  assign n3560 = ( n239 & ~n1048 ) | ( n239 & n1274 ) | ( ~n1048 & n1274 ) ;
  assign n3561 = n3560 ^ n2242 ^ x46 ;
  assign n3562 = n3561 ^ n2674 ^ x52 ;
  assign n3559 = ( ~n688 & n1261 ) | ( ~n688 & n2465 ) | ( n1261 & n2465 ) ;
  assign n3563 = n3562 ^ n3559 ^ 1'b0 ;
  assign n3564 = ( n205 & ~n1747 ) | ( n205 & n3563 ) | ( ~n1747 & n3563 ) ;
  assign n3568 = n2329 ^ n1211 ^ n454 ;
  assign n3565 = x3 & n1577 ;
  assign n3566 = n579 & n3565 ;
  assign n3567 = n3566 ^ n3400 ^ n1733 ;
  assign n3569 = n3568 ^ n3567 ^ n1567 ;
  assign n3570 = n3564 & ~n3569 ;
  assign n3574 = n773 ^ n515 ^ n512 ;
  assign n3571 = n603 | n2737 ;
  assign n3572 = n1630 & ~n3571 ;
  assign n3573 = n3572 ^ n349 ^ x62 ;
  assign n3575 = n3574 ^ n3573 ^ 1'b0 ;
  assign n3576 = ~n1707 & n3575 ;
  assign n3577 = ~n691 & n3576 ;
  assign n3578 = ~n1643 & n3577 ;
  assign n3583 = n2417 ^ n1726 ^ n129 ;
  assign n3584 = n3583 ^ n3426 ^ 1'b0 ;
  assign n3579 = ( n881 & n1813 ) | ( n881 & n3062 ) | ( n1813 & n3062 ) ;
  assign n3580 = ~n3540 & n3579 ;
  assign n3581 = ( ~n1172 & n2754 ) | ( ~n1172 & n3580 ) | ( n2754 & n3580 ) ;
  assign n3582 = n3581 ^ n1643 ^ x48 ;
  assign n3585 = n3584 ^ n3582 ^ n2795 ;
  assign n3586 = ( n383 & n651 ) | ( n383 & ~n1829 ) | ( n651 & ~n1829 ) ;
  assign n3587 = ( n970 & n1163 ) | ( n970 & ~n3586 ) | ( n1163 & ~n3586 ) ;
  assign n3588 = ( n3578 & n3585 ) | ( n3578 & ~n3587 ) | ( n3585 & ~n3587 ) ;
  assign n3589 = n732 ^ n593 ^ n392 ;
  assign n3590 = n1814 ^ n1201 ^ n452 ;
  assign n3591 = ( ~n2744 & n3589 ) | ( ~n2744 & n3590 ) | ( n3589 & n3590 ) ;
  assign n3592 = n3561 ^ n2981 ^ n1362 ;
  assign n3593 = n3592 ^ n2020 ^ n1906 ;
  assign n3594 = ( n475 & ~n1205 ) | ( n475 & n3593 ) | ( ~n1205 & n3593 ) ;
  assign n3595 = ( x32 & n251 ) | ( x32 & n3594 ) | ( n251 & n3594 ) ;
  assign n3596 = n1902 ^ n1849 ^ n1042 ;
  assign n3597 = n3522 ^ n2136 ^ n247 ;
  assign n3598 = ~n3596 & n3597 ;
  assign n3599 = ~n3595 & n3598 ;
  assign n3601 = n3162 ^ n2982 ^ 1'b0 ;
  assign n3600 = n3315 ^ n1648 ^ n159 ;
  assign n3602 = n3601 ^ n3600 ^ 1'b0 ;
  assign n3607 = n1861 ^ n1270 ^ n417 ;
  assign n3603 = ( ~n914 & n1220 ) | ( ~n914 & n1477 ) | ( n1220 & n1477 ) ;
  assign n3604 = n3603 ^ n1749 ^ 1'b0 ;
  assign n3605 = n3604 ^ n1802 ^ n894 ;
  assign n3606 = n3605 ^ n1927 ^ 1'b0 ;
  assign n3608 = n3607 ^ n3606 ^ n3040 ;
  assign n3609 = n1894 ^ n447 ^ x113 ;
  assign n3610 = n3609 ^ n702 ^ n473 ;
  assign n3612 = ( ~n214 & n294 ) | ( ~n214 & n2274 ) | ( n294 & n2274 ) ;
  assign n3611 = n2408 & n3384 ;
  assign n3613 = n3612 ^ n3611 ^ 1'b0 ;
  assign n3614 = ( n2083 & n3610 ) | ( n2083 & ~n3613 ) | ( n3610 & ~n3613 ) ;
  assign n3615 = ( n2653 & n2909 ) | ( n2653 & n3614 ) | ( n2909 & n3614 ) ;
  assign n3624 = ( n355 & n692 ) | ( n355 & ~n1507 ) | ( n692 & ~n1507 ) ;
  assign n3621 = n2066 ^ n526 ^ n355 ;
  assign n3622 = n350 & ~n369 ;
  assign n3623 = ( n197 & n3621 ) | ( n197 & ~n3622 ) | ( n3621 & ~n3622 ) ;
  assign n3618 = n1519 ^ n1084 ^ n944 ;
  assign n3619 = ( n1027 & n3095 ) | ( n1027 & n3618 ) | ( n3095 & n3618 ) ;
  assign n3616 = n234 & ~n1332 ;
  assign n3617 = ( n1307 & ~n3215 ) | ( n1307 & n3616 ) | ( ~n3215 & n3616 ) ;
  assign n3620 = n3619 ^ n3617 ^ n2653 ;
  assign n3625 = n3624 ^ n3623 ^ n3620 ;
  assign n3626 = ~n363 & n1133 ;
  assign n3627 = ~n2620 & n3077 ;
  assign n3628 = n3432 & n3627 ;
  assign n3629 = ( ~n2777 & n3626 ) | ( ~n2777 & n3628 ) | ( n3626 & n3628 ) ;
  assign n3630 = n585 ^ x72 ^ 1'b0 ;
  assign n3631 = x86 & ~n3630 ;
  assign n3632 = n778 | n2557 ;
  assign n3633 = n3632 ^ n1336 ^ 1'b0 ;
  assign n3634 = ( n2488 & n3631 ) | ( n2488 & ~n3633 ) | ( n3631 & ~n3633 ) ;
  assign n3635 = n2235 ^ n1682 ^ n1286 ;
  assign n3636 = n2501 & ~n3635 ;
  assign n3637 = n3636 ^ n3535 ^ n2789 ;
  assign n3651 = ( n250 & n691 ) | ( n250 & n709 ) | ( n691 & n709 ) ;
  assign n3652 = n3651 ^ n1822 ^ n1365 ;
  assign n3653 = ( n601 & ~n2458 ) | ( n601 & n2762 ) | ( ~n2458 & n2762 ) ;
  assign n3654 = n1457 ^ n447 ^ 1'b0 ;
  assign n3655 = ( n3652 & n3653 ) | ( n3652 & n3654 ) | ( n3653 & n3654 ) ;
  assign n3646 = n3188 ^ n863 ^ 1'b0 ;
  assign n3647 = n875 | n3646 ;
  assign n3648 = n3647 ^ n1187 ^ 1'b0 ;
  assign n3649 = n2660 & n3648 ;
  assign n3650 = n3649 ^ n2809 ^ n1914 ;
  assign n3638 = n292 & n776 ;
  assign n3639 = n3638 ^ n1081 ^ 1'b0 ;
  assign n3640 = ( n908 & n2033 ) | ( n908 & n3639 ) | ( n2033 & n3639 ) ;
  assign n3641 = n3121 ^ n2545 ^ n2134 ;
  assign n3642 = ( ~n484 & n2132 ) | ( ~n484 & n2177 ) | ( n2132 & n2177 ) ;
  assign n3643 = n3642 ^ n2690 ^ n1455 ;
  assign n3644 = ( n3640 & n3641 ) | ( n3640 & ~n3643 ) | ( n3641 & ~n3643 ) ;
  assign n3645 = n3644 ^ x116 ^ x96 ;
  assign n3656 = n3655 ^ n3650 ^ n3645 ;
  assign n3657 = ( n513 & n852 ) | ( n513 & ~n2618 ) | ( n852 & ~n2618 ) ;
  assign n3658 = n997 & n3657 ;
  assign n3659 = n3658 ^ n3218 ^ 1'b0 ;
  assign n3660 = n1233 ^ n1217 ^ x55 ;
  assign n3661 = n3660 ^ n2526 ^ x115 ;
  assign n3662 = n3661 ^ n191 ^ 1'b0 ;
  assign n3663 = n3607 | n3662 ;
  assign n3664 = ( x27 & n565 ) | ( x27 & ~n1052 ) | ( n565 & ~n1052 ) ;
  assign n3665 = ( ~n1097 & n1908 ) | ( ~n1097 & n3664 ) | ( n1908 & n3664 ) ;
  assign n3666 = n1849 ^ n177 ^ x36 ;
  assign n3667 = n2554 ^ n767 ^ n441 ;
  assign n3668 = n3667 ^ n3081 ^ n1270 ;
  assign n3669 = n3668 ^ n3307 ^ n2670 ;
  assign n3670 = ( ~n3068 & n3666 ) | ( ~n3068 & n3669 ) | ( n3666 & n3669 ) ;
  assign n3671 = ( x42 & n3665 ) | ( x42 & n3670 ) | ( n3665 & n3670 ) ;
  assign n3672 = n2338 ^ n1294 ^ 1'b0 ;
  assign n3673 = n3671 & ~n3672 ;
  assign n3674 = ( n2082 & n2922 ) | ( n2082 & n3673 ) | ( n2922 & n3673 ) ;
  assign n3679 = n935 & n2844 ;
  assign n3680 = n3679 ^ n1914 ^ 1'b0 ;
  assign n3677 = ( n289 & ~n825 ) | ( n289 & n1596 ) | ( ~n825 & n1596 ) ;
  assign n3675 = n1280 | n2258 ;
  assign n3676 = n2851 | n3675 ;
  assign n3678 = n3677 ^ n3676 ^ n1865 ;
  assign n3681 = n3680 ^ n3678 ^ 1'b0 ;
  assign n3682 = n1897 | n3681 ;
  assign n3683 = ( n401 & ~n1055 ) | ( n401 & n2094 ) | ( ~n1055 & n2094 ) ;
  assign n3684 = ( n1287 & n2531 ) | ( n1287 & ~n2840 ) | ( n2531 & ~n2840 ) ;
  assign n3685 = n1493 & ~n3684 ;
  assign n3686 = ( n2413 & n3384 ) | ( n2413 & ~n3685 ) | ( n3384 & ~n3685 ) ;
  assign n3687 = ( n3040 & n3683 ) | ( n3040 & n3686 ) | ( n3683 & n3686 ) ;
  assign n3688 = n3621 ^ n2304 ^ 1'b0 ;
  assign n3689 = ( n1393 & n3687 ) | ( n1393 & n3688 ) | ( n3687 & n3688 ) ;
  assign n3697 = n2405 ^ n2046 ^ n620 ;
  assign n3698 = n1056 ^ n956 ^ 1'b0 ;
  assign n3699 = ~n2029 & n3698 ;
  assign n3700 = ( ~n778 & n3371 ) | ( ~n778 & n3699 ) | ( n3371 & n3699 ) ;
  assign n3701 = ( n2655 & n3697 ) | ( n2655 & n3700 ) | ( n3697 & n3700 ) ;
  assign n3690 = n2593 ^ n1867 ^ n794 ;
  assign n3693 = ~n1012 & n1340 ;
  assign n3694 = ( x115 & ~n277 ) | ( x115 & n3693 ) | ( ~n277 & n3693 ) ;
  assign n3691 = n1937 ^ n1304 ^ n447 ;
  assign n3692 = n1627 | n3691 ;
  assign n3695 = n3694 ^ n3692 ^ n1531 ;
  assign n3696 = ~n3690 & n3695 ;
  assign n3702 = n3701 ^ n3696 ^ n224 ;
  assign n3715 = n1072 | n1789 ;
  assign n3716 = n1226 & ~n3715 ;
  assign n3717 = n3716 ^ n129 ^ x31 ;
  assign n3718 = n1219 & n3717 ;
  assign n3719 = n3718 ^ n1210 ^ 1'b0 ;
  assign n3720 = n3719 ^ n3056 ^ n427 ;
  assign n3721 = n902 ^ n705 ^ 1'b0 ;
  assign n3722 = ( ~n1393 & n1902 ) | ( ~n1393 & n3721 ) | ( n1902 & n3721 ) ;
  assign n3723 = n3720 & n3722 ;
  assign n3724 = n1322 & n3723 ;
  assign n3703 = ( n291 & n583 ) | ( n291 & ~n827 ) | ( n583 & ~n827 ) ;
  assign n3704 = n3703 ^ n1705 ^ n1132 ;
  assign n3705 = n3704 ^ n956 ^ 1'b0 ;
  assign n3706 = n3705 ^ n2601 ^ n1725 ;
  assign n3707 = ( ~n419 & n1660 ) | ( ~n419 & n2513 ) | ( n1660 & n2513 ) ;
  assign n3708 = n3707 ^ n3573 ^ 1'b0 ;
  assign n3709 = n3160 | n3708 ;
  assign n3710 = ( n818 & n3706 ) | ( n818 & ~n3709 ) | ( n3706 & ~n3709 ) ;
  assign n3711 = ( x92 & n532 ) | ( x92 & ~n734 ) | ( n532 & ~n734 ) ;
  assign n3712 = n3711 ^ n2247 ^ n1704 ;
  assign n3713 = n3712 ^ n3085 ^ n1344 ;
  assign n3714 = ( n2182 & n3710 ) | ( n2182 & n3713 ) | ( n3710 & n3713 ) ;
  assign n3725 = n3724 ^ n3714 ^ 1'b0 ;
  assign n3726 = n3558 ^ n2688 ^ n368 ;
  assign n3727 = n349 & n1805 ;
  assign n3728 = n2034 ^ n777 ^ n261 ;
  assign n3729 = ( n1828 & ~n2342 ) | ( n1828 & n3728 ) | ( ~n2342 & n3728 ) ;
  assign n3730 = n916 | n2803 ;
  assign n3731 = n2497 | n3730 ;
  assign n3732 = ( n2079 & n2487 ) | ( n2079 & n3731 ) | ( n2487 & n3731 ) ;
  assign n3733 = ( n199 & ~n940 ) | ( n199 & n1727 ) | ( ~n940 & n1727 ) ;
  assign n3734 = n3733 ^ n483 ^ 1'b0 ;
  assign n3735 = n3734 ^ n2183 ^ n977 ;
  assign n3736 = ~n1342 & n2323 ;
  assign n3737 = n2670 ^ n2291 ^ n1025 ;
  assign n3738 = n3737 ^ n1743 ^ 1'b0 ;
  assign n3739 = n3152 & ~n3738 ;
  assign n3742 = n2711 ^ n1755 ^ n754 ;
  assign n3743 = n638 ^ n245 ^ 1'b0 ;
  assign n3744 = n3742 & ~n3743 ;
  assign n3740 = n2952 ^ n1179 ^ n641 ;
  assign n3741 = n3740 ^ n379 ^ 1'b0 ;
  assign n3745 = n3744 ^ n3741 ^ n903 ;
  assign n3746 = n810 ^ n432 ^ n163 ;
  assign n3747 = n3746 ^ n1066 ^ n929 ;
  assign n3748 = ( n1338 & n1826 ) | ( n1338 & ~n3747 ) | ( n1826 & ~n3747 ) ;
  assign n3749 = ~n791 & n3748 ;
  assign n3750 = n2885 & n3749 ;
  assign n3751 = n1261 | n1539 ;
  assign n3752 = n3751 ^ n3269 ^ n1242 ;
  assign n3753 = ( n458 & n3750 ) | ( n458 & ~n3752 ) | ( n3750 & ~n3752 ) ;
  assign n3754 = n2786 ^ n578 ^ x99 ;
  assign n3755 = n3754 ^ n1230 ^ n393 ;
  assign n3756 = n2840 ^ n389 ^ n239 ;
  assign n3757 = ( x2 & n2414 ) | ( x2 & n3756 ) | ( n2414 & n3756 ) ;
  assign n3758 = ( n751 & n3755 ) | ( n751 & n3757 ) | ( n3755 & n3757 ) ;
  assign n3759 = ( n2829 & n3270 ) | ( n2829 & n3702 ) | ( n3270 & n3702 ) ;
  assign n3760 = n3583 ^ n3338 ^ n696 ;
  assign n3761 = ( ~n290 & n1757 ) | ( ~n290 & n3760 ) | ( n1757 & n3760 ) ;
  assign n3762 = ( n139 & n194 ) | ( n139 & ~n1767 ) | ( n194 & ~n1767 ) ;
  assign n3763 = ( n935 & ~n3761 ) | ( n935 & n3762 ) | ( ~n3761 & n3762 ) ;
  assign n3764 = n304 & n558 ;
  assign n3765 = ~n141 & n3764 ;
  assign n3766 = n579 | n3062 ;
  assign n3767 = ( ~n3428 & n3765 ) | ( ~n3428 & n3766 ) | ( n3765 & n3766 ) ;
  assign n3768 = ( x31 & n1457 ) | ( x31 & ~n3767 ) | ( n1457 & ~n3767 ) ;
  assign n3769 = ( n266 & n2185 ) | ( n266 & ~n2206 ) | ( n2185 & ~n2206 ) ;
  assign n3770 = ~n1076 & n3769 ;
  assign n3771 = n672 & n3770 ;
  assign n3772 = n3771 ^ n2859 ^ n708 ;
  assign n3773 = n3101 ^ n1703 ^ n1241 ;
  assign n3774 = ( n2245 & n2874 ) | ( n2245 & n3773 ) | ( n2874 & n3773 ) ;
  assign n3776 = n2773 ^ n2245 ^ n1700 ;
  assign n3777 = ( ~n565 & n1052 ) | ( ~n565 & n1352 ) | ( n1052 & n1352 ) ;
  assign n3778 = ~n1805 & n3777 ;
  assign n3779 = n3778 ^ n454 ^ 1'b0 ;
  assign n3780 = ( ~n2964 & n3776 ) | ( ~n2964 & n3779 ) | ( n3776 & n3779 ) ;
  assign n3775 = ( n196 & n1265 ) | ( n196 & ~n2980 ) | ( n1265 & ~n2980 ) ;
  assign n3781 = n3780 ^ n3775 ^ n1589 ;
  assign n3797 = ( ~x27 & n2049 ) | ( ~x27 & n2355 ) | ( n2049 & n2355 ) ;
  assign n3798 = n3106 & ~n3797 ;
  assign n3795 = n2127 ^ n1580 ^ 1'b0 ;
  assign n3796 = n192 & n3795 ;
  assign n3799 = n3798 ^ n3796 ^ 1'b0 ;
  assign n3788 = n1987 & ~n2477 ;
  assign n3789 = n3733 & n3788 ;
  assign n3790 = n3384 ^ n1411 ^ n671 ;
  assign n3791 = n3790 ^ n2859 ^ n2177 ;
  assign n3792 = n1471 & n3791 ;
  assign n3793 = ~n1132 & n3792 ;
  assign n3794 = n3789 & n3793 ;
  assign n3784 = ( x3 & n546 ) | ( x3 & n1491 ) | ( n546 & n1491 ) ;
  assign n3783 = n607 | n702 ;
  assign n3785 = n3784 ^ n3783 ^ 1'b0 ;
  assign n3786 = n3785 ^ n2228 ^ n1865 ;
  assign n3782 = n3589 ^ n2241 ^ n756 ;
  assign n3787 = n3786 ^ n3782 ^ 1'b0 ;
  assign n3800 = n3799 ^ n3794 ^ n3787 ;
  assign n3801 = n1670 & ~n2529 ;
  assign n3802 = ( ~n2170 & n3013 ) | ( ~n2170 & n3801 ) | ( n3013 & n3801 ) ;
  assign n3803 = ( ~x68 & n207 ) | ( ~x68 & n1104 ) | ( n207 & n1104 ) ;
  assign n3804 = n3468 & ~n3803 ;
  assign n3805 = ( x115 & ~n1430 ) | ( x115 & n1712 ) | ( ~n1430 & n1712 ) ;
  assign n3806 = n2501 ^ n760 ^ n567 ;
  assign n3807 = n3806 ^ n3560 ^ n2241 ;
  assign n3808 = ( n2479 & ~n3805 ) | ( n2479 & n3807 ) | ( ~n3805 & n3807 ) ;
  assign n3809 = n1344 ^ n470 ^ 1'b0 ;
  assign n3810 = n1807 & ~n3809 ;
  assign n3811 = n3810 ^ n2129 ^ 1'b0 ;
  assign n3812 = n193 & n3811 ;
  assign n3813 = n3812 ^ n2661 ^ 1'b0 ;
  assign n3814 = n1474 & ~n3813 ;
  assign n3815 = ( n2034 & n2739 ) | ( n2034 & ~n3287 ) | ( n2739 & ~n3287 ) ;
  assign n3816 = ( n1103 & n1872 ) | ( n1103 & ~n2897 ) | ( n1872 & ~n2897 ) ;
  assign n3817 = n3816 ^ n1644 ^ n658 ;
  assign n3824 = n599 & n1557 ;
  assign n3825 = n2941 & n3824 ;
  assign n3826 = x39 & ~n3825 ;
  assign n3827 = ~n282 & n3826 ;
  assign n3822 = n497 & n1937 ;
  assign n3820 = ( n2269 & n2750 ) | ( n2269 & n2758 ) | ( n2750 & n2758 ) ;
  assign n3821 = ( ~n145 & n2021 ) | ( ~n145 & n3820 ) | ( n2021 & n3820 ) ;
  assign n3823 = n3822 ^ n3821 ^ n3165 ;
  assign n3828 = n3827 ^ n3823 ^ 1'b0 ;
  assign n3818 = n3056 ^ n1287 ^ n527 ;
  assign n3819 = x115 & ~n3818 ;
  assign n3829 = n3828 ^ n3819 ^ 1'b0 ;
  assign n3830 = ( n3815 & n3817 ) | ( n3815 & n3829 ) | ( n3817 & n3829 ) ;
  assign n3831 = n1655 ^ n712 ^ 1'b0 ;
  assign n3832 = ( n215 & n460 ) | ( n215 & n2200 ) | ( n460 & n2200 ) ;
  assign n3833 = ~n1656 & n3832 ;
  assign n3838 = n774 & ~n1561 ;
  assign n3835 = n999 ^ x112 ^ 1'b0 ;
  assign n3834 = n314 & n844 ;
  assign n3836 = n3835 ^ n3834 ^ 1'b0 ;
  assign n3837 = n3836 ^ n1715 ^ n733 ;
  assign n3839 = n3838 ^ n3837 ^ n2878 ;
  assign n3844 = ~n1093 & n1165 ;
  assign n3845 = ( x46 & ~n1416 ) | ( x46 & n3844 ) | ( ~n1416 & n3844 ) ;
  assign n3846 = ( ~n2872 & n2890 ) | ( ~n2872 & n3845 ) | ( n2890 & n3845 ) ;
  assign n3841 = n3505 ^ n1409 ^ n1189 ;
  assign n3842 = ( ~n3193 & n3487 ) | ( ~n3193 & n3841 ) | ( n3487 & n3841 ) ;
  assign n3840 = n2635 ^ n1055 ^ n827 ;
  assign n3843 = n3842 ^ n3840 ^ n2483 ;
  assign n3847 = n3846 ^ n3843 ^ n2529 ;
  assign n3848 = n3847 ^ n2365 ^ n1861 ;
  assign n3854 = ( n538 & n2086 ) | ( n538 & n3034 ) | ( n2086 & n3034 ) ;
  assign n3855 = n3854 ^ n2764 ^ n2445 ;
  assign n3849 = n2356 ^ n1405 ^ n1350 ;
  assign n3850 = n2131 & ~n2603 ;
  assign n3851 = n3850 ^ n1662 ^ 1'b0 ;
  assign n3852 = n3851 ^ n3697 ^ n1075 ;
  assign n3853 = ( ~n3653 & n3849 ) | ( ~n3653 & n3852 ) | ( n3849 & n3852 ) ;
  assign n3856 = n3855 ^ n3853 ^ n1690 ;
  assign n3857 = ( n1634 & ~n2346 ) | ( n1634 & n3856 ) | ( ~n2346 & n3856 ) ;
  assign n3858 = ( n673 & ~n959 ) | ( n673 & n1807 ) | ( ~n959 & n1807 ) ;
  assign n3859 = n250 & n961 ;
  assign n3860 = n3859 ^ n1228 ^ n629 ;
  assign n3861 = n3860 ^ n1633 ^ n1368 ;
  assign n3862 = ( n1191 & n3858 ) | ( n1191 & ~n3861 ) | ( n3858 & ~n3861 ) ;
  assign n3875 = ( n162 & n1633 ) | ( n162 & n1790 ) | ( n1633 & n1790 ) ;
  assign n3876 = n3875 ^ n969 ^ 1'b0 ;
  assign n3877 = ( n1884 & ~n2634 ) | ( n1884 & n3876 ) | ( ~n2634 & n3876 ) ;
  assign n3871 = ~n389 & n497 ;
  assign n3872 = ~x76 & n3871 ;
  assign n3873 = ( n1445 & n2778 ) | ( n1445 & n3872 ) | ( n2778 & n3872 ) ;
  assign n3874 = ~n1374 & n3873 ;
  assign n3878 = n3877 ^ n3874 ^ 1'b0 ;
  assign n3867 = ( n420 & ~n661 ) | ( n420 & n1277 ) | ( ~n661 & n1277 ) ;
  assign n3868 = n3867 ^ n1318 ^ n1229 ;
  assign n3863 = n724 ^ x3 ^ 1'b0 ;
  assign n3864 = n2727 ^ n892 ^ 1'b0 ;
  assign n3865 = n3863 & ~n3864 ;
  assign n3866 = n3865 ^ n2730 ^ n2689 ;
  assign n3869 = n3868 ^ n3866 ^ 1'b0 ;
  assign n3870 = n434 | n3869 ;
  assign n3879 = n3878 ^ n3870 ^ 1'b0 ;
  assign n3880 = ( ~n1207 & n2163 ) | ( ~n1207 & n3518 ) | ( n2163 & n3518 ) ;
  assign n3881 = n1424 | n3880 ;
  assign n3882 = n1723 ^ n730 ^ n364 ;
  assign n3883 = n3882 ^ n3166 ^ n2813 ;
  assign n3884 = ( ~n3331 & n3881 ) | ( ~n3331 & n3883 ) | ( n3881 & n3883 ) ;
  assign n3885 = n325 & ~n2206 ;
  assign n3886 = n2215 & n2325 ;
  assign n3887 = n588 & n3886 ;
  assign n3888 = n3887 ^ n949 ^ 1'b0 ;
  assign n3889 = ( n387 & ~n2114 ) | ( n387 & n3888 ) | ( ~n2114 & n3888 ) ;
  assign n3890 = ( n1335 & n2891 ) | ( n1335 & ~n3716 ) | ( n2891 & ~n3716 ) ;
  assign n3891 = n3242 ^ n2117 ^ 1'b0 ;
  assign n3892 = ~n2010 & n3891 ;
  assign n3893 = ( n1302 & n1421 ) | ( n1302 & n3892 ) | ( n1421 & n3892 ) ;
  assign n3894 = n1089 ^ n277 ^ 1'b0 ;
  assign n3895 = n1890 & n3894 ;
  assign n3896 = n3895 ^ n3586 ^ 1'b0 ;
  assign n3897 = ( n181 & n3574 ) | ( n181 & n3896 ) | ( n3574 & n3896 ) ;
  assign n3898 = n1498 & ~n3897 ;
  assign n3899 = ~n3138 & n3898 ;
  assign n3900 = n3899 ^ n2738 ^ n859 ;
  assign n3901 = ( ~n2994 & n3893 ) | ( ~n2994 & n3900 ) | ( n3893 & n3900 ) ;
  assign n3902 = n3901 ^ n2586 ^ 1'b0 ;
  assign n3903 = n3541 & n3902 ;
  assign n3904 = n3890 | n3903 ;
  assign n3905 = ( n144 & ~n409 ) | ( n144 & n3039 ) | ( ~n409 & n3039 ) ;
  assign n3906 = n772 | n3905 ;
  assign n3907 = n3906 ^ n2295 ^ 1'b0 ;
  assign n3908 = ( ~x66 & n1908 ) | ( ~x66 & n2103 ) | ( n1908 & n2103 ) ;
  assign n3909 = ( ~n3752 & n3907 ) | ( ~n3752 & n3908 ) | ( n3907 & n3908 ) ;
  assign n3910 = n1405 ^ n735 ^ n254 ;
  assign n3911 = ( ~n157 & n559 ) | ( ~n157 & n1924 ) | ( n559 & n1924 ) ;
  assign n3912 = ( n1102 & n2202 ) | ( n1102 & n3911 ) | ( n2202 & n3911 ) ;
  assign n3913 = ( n1400 & n3910 ) | ( n1400 & ~n3912 ) | ( n3910 & ~n3912 ) ;
  assign n3918 = n1756 ^ n1262 ^ n995 ;
  assign n3914 = n2927 ^ n2417 ^ 1'b0 ;
  assign n3915 = n2949 & ~n3914 ;
  assign n3916 = n3915 ^ n1071 ^ n1038 ;
  assign n3917 = n3916 ^ n3402 ^ n2228 ;
  assign n3919 = n3918 ^ n3917 ^ 1'b0 ;
  assign n3920 = n1823 ^ n1515 ^ x97 ;
  assign n3921 = n1244 ^ n497 ^ n160 ;
  assign n3922 = n3921 ^ n913 ^ 1'b0 ;
  assign n3923 = ~n3538 & n3922 ;
  assign n3924 = ( n3235 & n3920 ) | ( n3235 & n3923 ) | ( n3920 & n3923 ) ;
  assign n3938 = ( ~n896 & n977 ) | ( ~n896 & n1036 ) | ( n977 & n1036 ) ;
  assign n3925 = n1411 & n1546 ;
  assign n3926 = ~n1142 & n3925 ;
  assign n3927 = ( n2782 & n2880 ) | ( n2782 & n3168 ) | ( n2880 & n3168 ) ;
  assign n3928 = ( n462 & n1289 ) | ( n462 & n1309 ) | ( n1289 & n1309 ) ;
  assign n3929 = ( n732 & n3384 ) | ( n732 & ~n3928 ) | ( n3384 & ~n3928 ) ;
  assign n3930 = ~n159 & n3929 ;
  assign n3931 = n180 & n3930 ;
  assign n3932 = ( n1904 & n2228 ) | ( n1904 & n3931 ) | ( n2228 & n3931 ) ;
  assign n3933 = n3237 ^ n2952 ^ 1'b0 ;
  assign n3934 = n3933 ^ n1833 ^ 1'b0 ;
  assign n3935 = ( n3153 & ~n3932 ) | ( n3153 & n3934 ) | ( ~n3932 & n3934 ) ;
  assign n3936 = ( n2425 & ~n3927 ) | ( n2425 & n3935 ) | ( ~n3927 & n3935 ) ;
  assign n3937 = n3926 & ~n3936 ;
  assign n3939 = n3938 ^ n3937 ^ n2087 ;
  assign n3940 = ~n737 & n2810 ;
  assign n3941 = ( n1006 & n1057 ) | ( n1006 & ~n3940 ) | ( n1057 & ~n3940 ) ;
  assign n3942 = ( n1254 & ~n3308 ) | ( n1254 & n3941 ) | ( ~n3308 & n3941 ) ;
  assign n3943 = n1658 ^ n714 ^ x2 ;
  assign n3944 = n3943 ^ n3102 ^ n1142 ;
  assign n3945 = ~n2800 & n3944 ;
  assign n3946 = n3174 & n3945 ;
  assign n3947 = n2789 & ~n3946 ;
  assign n3948 = n3947 ^ n3417 ^ 1'b0 ;
  assign n3949 = n3948 ^ n2818 ^ n373 ;
  assign n3950 = ( n620 & ~n3942 ) | ( n620 & n3949 ) | ( ~n3942 & n3949 ) ;
  assign n3951 = n3950 ^ n1139 ^ 1'b0 ;
  assign n3955 = n3146 & ~n3603 ;
  assign n3956 = ~n646 & n3955 ;
  assign n3952 = n1790 ^ n705 ^ x77 ;
  assign n3953 = n1365 ^ n1332 ^ x4 ;
  assign n3954 = ( ~n813 & n3952 ) | ( ~n813 & n3953 ) | ( n3952 & n3953 ) ;
  assign n3957 = n3956 ^ n3954 ^ n1973 ;
  assign n3958 = n3957 ^ n2633 ^ n740 ;
  assign n3961 = n850 | n1373 ;
  assign n3962 = n3961 ^ n1412 ^ 1'b0 ;
  assign n3963 = n2925 & ~n3962 ;
  assign n3964 = ~n701 & n3963 ;
  assign n3959 = n2145 | n2891 ;
  assign n3960 = n1580 & n3959 ;
  assign n3965 = n3964 ^ n3960 ^ 1'b0 ;
  assign n3966 = ( n545 & n1447 ) | ( n545 & n3619 ) | ( n1447 & n3619 ) ;
  assign n3967 = n3966 ^ n1647 ^ n430 ;
  assign n3968 = ( n1121 & ~n1572 ) | ( n1121 & n3126 ) | ( ~n1572 & n3126 ) ;
  assign n3969 = ( n1331 & n3243 ) | ( n1331 & ~n3968 ) | ( n3243 & ~n3968 ) ;
  assign n3970 = ~n698 & n2341 ;
  assign n3971 = n3970 ^ n3171 ^ x89 ;
  assign n3972 = n2642 ^ n987 ^ n305 ;
  assign n3973 = ( n655 & ~n3971 ) | ( n655 & n3972 ) | ( ~n3971 & n3972 ) ;
  assign n3974 = n3973 ^ n3485 ^ n419 ;
  assign n3976 = n2665 ^ n1899 ^ n1340 ;
  assign n3975 = ( n182 & n2691 ) | ( n182 & n2728 ) | ( n2691 & n2728 ) ;
  assign n3977 = n3976 ^ n3975 ^ n2013 ;
  assign n3978 = ( n651 & n3349 ) | ( n651 & ~n3610 ) | ( n3349 & ~n3610 ) ;
  assign n3979 = n1131 ^ n739 ^ 1'b0 ;
  assign n3980 = ( ~n1490 & n1998 ) | ( ~n1490 & n2028 ) | ( n1998 & n2028 ) ;
  assign n3981 = n3980 ^ n155 ^ 1'b0 ;
  assign n3982 = n3981 ^ n2574 ^ n1327 ;
  assign n3983 = n2650 ^ n1675 ^ 1'b0 ;
  assign n3984 = ( ~x20 & n2686 ) | ( ~x20 & n3311 ) | ( n2686 & n3311 ) ;
  assign n3985 = ( n3882 & n3983 ) | ( n3882 & ~n3984 ) | ( n3983 & ~n3984 ) ;
  assign n3986 = ( n3979 & n3982 ) | ( n3979 & ~n3985 ) | ( n3982 & ~n3985 ) ;
  assign n3987 = n3477 ^ n1346 ^ x115 ;
  assign n3988 = ( ~n1538 & n2037 ) | ( ~n1538 & n3987 ) | ( n2037 & n3987 ) ;
  assign n3989 = n1927 ^ n358 ^ n338 ;
  assign n3990 = n3989 ^ n260 ^ 1'b0 ;
  assign n3991 = ( n3235 & n3331 ) | ( n3235 & n3990 ) | ( n3331 & n3990 ) ;
  assign n3992 = n3640 ^ n773 ^ n146 ;
  assign n3997 = n1348 ^ n867 ^ n636 ;
  assign n3998 = n1214 & n3997 ;
  assign n3993 = ( n618 & ~n2040 ) | ( n618 & n2188 ) | ( ~n2040 & n2188 ) ;
  assign n3994 = ~x43 & n858 ;
  assign n3995 = ( n1222 & n3993 ) | ( n1222 & n3994 ) | ( n3993 & n3994 ) ;
  assign n3996 = ( n1663 & n1971 ) | ( n1663 & n3995 ) | ( n1971 & n3995 ) ;
  assign n3999 = n3998 ^ n3996 ^ 1'b0 ;
  assign n4000 = n769 ^ n291 ^ 1'b0 ;
  assign n4001 = n4000 ^ n879 ^ n811 ;
  assign n4002 = ~n1424 & n3691 ;
  assign n4003 = n229 & n4002 ;
  assign n4004 = ( n3999 & ~n4001 ) | ( n3999 & n4003 ) | ( ~n4001 & n4003 ) ;
  assign n4013 = n1895 ^ n1549 ^ n1143 ;
  assign n4014 = ( n691 & ~n1295 ) | ( n691 & n4013 ) | ( ~n1295 & n4013 ) ;
  assign n4015 = ( n426 & ~n3798 ) | ( n426 & n4014 ) | ( ~n3798 & n4014 ) ;
  assign n4016 = n4015 ^ n3805 ^ 1'b0 ;
  assign n4005 = n1229 & n1520 ;
  assign n4006 = ~n1971 & n4005 ;
  assign n4007 = x55 & n426 ;
  assign n4008 = n4007 ^ n404 ^ 1'b0 ;
  assign n4009 = n4008 ^ n1729 ^ n509 ;
  assign n4010 = ( n247 & ~n4006 ) | ( n247 & n4009 ) | ( ~n4006 & n4009 ) ;
  assign n4011 = ( n1796 & n3933 ) | ( n1796 & n4010 ) | ( n3933 & n4010 ) ;
  assign n4012 = n469 | n4011 ;
  assign n4017 = n4016 ^ n4012 ^ n793 ;
  assign n4018 = ( n1888 & n2910 ) | ( n1888 & ~n3177 ) | ( n2910 & ~n3177 ) ;
  assign n4019 = ( n209 & n1391 ) | ( n209 & n1492 ) | ( n1391 & n1492 ) ;
  assign n4020 = ( n642 & n1600 ) | ( n642 & ~n3162 ) | ( n1600 & ~n3162 ) ;
  assign n4021 = n4020 ^ n767 ^ n293 ;
  assign n4022 = ~n238 & n1380 ;
  assign n4023 = n4022 ^ n2295 ^ n1644 ;
  assign n4024 = n3368 ^ n2902 ^ 1'b0 ;
  assign n4025 = n3613 ^ n421 ^ 1'b0 ;
  assign n4026 = n962 & n4025 ;
  assign n4027 = n4026 ^ n3128 ^ 1'b0 ;
  assign n4028 = ( n4023 & n4024 ) | ( n4023 & ~n4027 ) | ( n4024 & ~n4027 ) ;
  assign n4029 = n2129 ^ n1209 ^ 1'b0 ;
  assign n4030 = n4029 ^ n3225 ^ n1661 ;
  assign n4031 = n2076 ^ n1182 ^ n737 ;
  assign n4032 = n4031 ^ n3765 ^ n1292 ;
  assign n4033 = ~n3705 & n4032 ;
  assign n4034 = n4030 & n4033 ;
  assign n4039 = ~n1652 & n1890 ;
  assign n4040 = n4039 ^ n3603 ^ n2557 ;
  assign n4037 = n725 | n1072 ;
  assign n4036 = ( n2027 & n2569 ) | ( n2027 & ~n3953 ) | ( n2569 & ~n3953 ) ;
  assign n4035 = ( ~n1435 & n1880 ) | ( ~n1435 & n3093 ) | ( n1880 & n3093 ) ;
  assign n4038 = n4037 ^ n4036 ^ n4035 ;
  assign n4041 = n4040 ^ n4038 ^ n512 ;
  assign n4042 = n1716 ^ n864 ^ x45 ;
  assign n4043 = n762 ^ n654 ^ n349 ;
  assign n4044 = n4043 ^ n2328 ^ 1'b0 ;
  assign n4045 = n4044 ^ n491 ^ 1'b0 ;
  assign n4046 = n4045 ^ n733 ^ n558 ;
  assign n4047 = n497 & n4046 ;
  assign n4048 = ~n4042 & n4047 ;
  assign n4049 = ~n1365 & n3149 ;
  assign n4050 = ~n4012 & n4049 ;
  assign n4051 = n1534 ^ n799 ^ 1'b0 ;
  assign n4052 = n1068 | n4051 ;
  assign n4053 = ( ~x50 & x120 ) | ( ~x50 & n3025 ) | ( x120 & n3025 ) ;
  assign n4054 = ( ~n554 & n1892 ) | ( ~n554 & n2039 ) | ( n1892 & n2039 ) ;
  assign n4055 = ( n710 & n4053 ) | ( n710 & ~n4054 ) | ( n4053 & ~n4054 ) ;
  assign n4056 = n701 & ~n963 ;
  assign n4057 = n291 | n992 ;
  assign n4058 = ( n282 & ~n450 ) | ( n282 & n2397 ) | ( ~n450 & n2397 ) ;
  assign n4059 = ( n484 & ~n1279 ) | ( n484 & n4058 ) | ( ~n1279 & n4058 ) ;
  assign n4060 = ~n4057 & n4059 ;
  assign n4061 = ( n641 & ~n3385 ) | ( n641 & n3653 ) | ( ~n3385 & n3653 ) ;
  assign n4062 = ~n4060 & n4061 ;
  assign n4063 = n4056 & n4062 ;
  assign n4064 = n1138 ^ n901 ^ 1'b0 ;
  assign n4065 = ( n1009 & n3172 ) | ( n1009 & n4064 ) | ( n3172 & n4064 ) ;
  assign n4066 = ( n421 & ~n489 ) | ( n421 & n4065 ) | ( ~n489 & n4065 ) ;
  assign n4079 = ( n914 & n1960 ) | ( n914 & ~n2378 ) | ( n1960 & ~n2378 ) ;
  assign n4080 = ( n1980 & ~n3785 ) | ( n1980 & n4079 ) | ( ~n3785 & n4079 ) ;
  assign n4078 = n2242 ^ n514 ^ n432 ;
  assign n4081 = n4080 ^ n4078 ^ n3954 ;
  assign n4074 = n142 ^ x65 ^ 1'b0 ;
  assign n4075 = ~n1332 & n4074 ;
  assign n4076 = ( n1653 & ~n2094 ) | ( n1653 & n4075 ) | ( ~n2094 & n4075 ) ;
  assign n4071 = ( n1041 & ~n2420 ) | ( n1041 & n3867 ) | ( ~n2420 & n3867 ) ;
  assign n4072 = n4071 ^ n2658 ^ 1'b0 ;
  assign n4073 = n771 | n4072 ;
  assign n4067 = n3304 ^ n1107 ^ 1'b0 ;
  assign n4068 = n145 & n4067 ;
  assign n4069 = n4068 ^ n1400 ^ n416 ;
  assign n4070 = n4069 ^ n2532 ^ 1'b0 ;
  assign n4077 = n4076 ^ n4073 ^ n4070 ;
  assign n4082 = n4081 ^ n4077 ^ 1'b0 ;
  assign n4083 = n1826 & ~n4082 ;
  assign n4084 = n1436 & ~n2317 ;
  assign n4085 = ~n1430 & n4084 ;
  assign n4086 = ( n154 & ~n482 ) | ( n154 & n539 ) | ( ~n482 & n539 ) ;
  assign n4087 = n4086 ^ n3980 ^ 1'b0 ;
  assign n4088 = n4087 ^ n167 ^ 1'b0 ;
  assign n4089 = ( n4006 & ~n4085 ) | ( n4006 & n4088 ) | ( ~n4085 & n4088 ) ;
  assign n4090 = n4089 ^ n2151 ^ n385 ;
  assign n4091 = n3664 ^ n2783 ^ n1497 ;
  assign n4092 = n593 | n4091 ;
  assign n4093 = n1742 | n4092 ;
  assign n4094 = n4093 ^ n1336 ^ n539 ;
  assign n4095 = n752 & n4094 ;
  assign n4096 = ~n570 & n4095 ;
  assign n4097 = n2510 ^ n562 ^ 1'b0 ;
  assign n4098 = n4097 ^ n3592 ^ n2480 ;
  assign n4099 = n2506 ^ n198 ^ 1'b0 ;
  assign n4100 = ( ~n2932 & n3182 ) | ( ~n2932 & n4099 ) | ( n3182 & n4099 ) ;
  assign n4101 = n4100 ^ n3370 ^ n2574 ;
  assign n4102 = ( ~n4096 & n4098 ) | ( ~n4096 & n4101 ) | ( n4098 & n4101 ) ;
  assign n4103 = n951 ^ n254 ^ 1'b0 ;
  assign n4104 = n4102 & ~n4103 ;
  assign n4105 = n3106 ^ n2297 ^ n1241 ;
  assign n4106 = n4105 ^ n3761 ^ n3691 ;
  assign n4107 = n4068 ^ n3435 ^ n214 ;
  assign n4108 = n4107 ^ n2303 ^ 1'b0 ;
  assign n4109 = n4108 ^ n2073 ^ 1'b0 ;
  assign n4110 = n1349 | n4109 ;
  assign n4111 = ( ~n414 & n1826 ) | ( ~n414 & n2274 ) | ( n1826 & n2274 ) ;
  assign n4112 = ( ~n998 & n1996 ) | ( ~n998 & n2991 ) | ( n1996 & n2991 ) ;
  assign n4113 = ( n2854 & n3518 ) | ( n2854 & n4112 ) | ( n3518 & n4112 ) ;
  assign n4121 = n3968 ^ n2898 ^ n1088 ;
  assign n4122 = n4121 ^ n1606 ^ n524 ;
  assign n4123 = n2539 & ~n4122 ;
  assign n4114 = n1667 ^ n688 ^ n568 ;
  assign n4115 = ( n832 & ~n1994 ) | ( n832 & n4114 ) | ( ~n1994 & n4114 ) ;
  assign n4116 = ( n459 & n1587 ) | ( n459 & ~n2990 ) | ( n1587 & ~n2990 ) ;
  assign n4117 = n2764 ^ n2367 ^ 1'b0 ;
  assign n4118 = n1113 | n4117 ;
  assign n4119 = n4118 ^ n2189 ^ n256 ;
  assign n4120 = ( ~n4115 & n4116 ) | ( ~n4115 & n4119 ) | ( n4116 & n4119 ) ;
  assign n4124 = n4123 ^ n4120 ^ n131 ;
  assign n4125 = n1560 ^ n201 ^ 1'b0 ;
  assign n4126 = n3070 | n4125 ;
  assign n4127 = n519 | n4126 ;
  assign n4128 = n4127 ^ n1922 ^ n580 ;
  assign n4129 = ( ~n1335 & n1346 ) | ( ~n1335 & n3308 ) | ( n1346 & n3308 ) ;
  assign n4130 = ~n224 & n4129 ;
  assign n4131 = ~n4128 & n4130 ;
  assign n4132 = n2481 ^ n1340 ^ n1234 ;
  assign n4133 = n4132 ^ n3746 ^ n626 ;
  assign n4134 = ~n2603 & n3818 ;
  assign n4135 = n4133 & ~n4134 ;
  assign n4136 = n1391 | n4135 ;
  assign n4137 = ( n3114 & ~n4131 ) | ( n3114 & n4136 ) | ( ~n4131 & n4136 ) ;
  assign n4138 = n2185 ^ n653 ^ 1'b0 ;
  assign n4139 = ~n923 & n4138 ;
  assign n4140 = n3692 & n3744 ;
  assign n4141 = ~n4139 & n4140 ;
  assign n4142 = ( n549 & n2538 ) | ( n549 & ~n4141 ) | ( n2538 & ~n4141 ) ;
  assign n4143 = ( ~n4124 & n4137 ) | ( ~n4124 & n4142 ) | ( n4137 & n4142 ) ;
  assign n4144 = n2028 ^ x104 ^ x40 ;
  assign n4145 = n2788 & n4144 ;
  assign n4146 = n4145 ^ n2694 ^ 1'b0 ;
  assign n4147 = ( ~n235 & n1059 ) | ( ~n235 & n4146 ) | ( n1059 & n4146 ) ;
  assign n4148 = ( n906 & ~n2260 ) | ( n906 & n4115 ) | ( ~n2260 & n4115 ) ;
  assign n4149 = x11 & n4148 ;
  assign n4150 = n1800 & n4149 ;
  assign n4151 = n4150 ^ n1496 ^ n199 ;
  assign n4152 = n2235 & ~n3588 ;
  assign n4153 = n4152 ^ n1889 ^ 1'b0 ;
  assign n4154 = n3349 ^ n3311 ^ n804 ;
  assign n4155 = n4154 ^ n3182 ^ n1232 ;
  assign n4156 = x92 & n1647 ;
  assign n4157 = ~n285 & n2664 ;
  assign n4158 = ( n304 & ~n4156 ) | ( n304 & n4157 ) | ( ~n4156 & n4157 ) ;
  assign n4159 = n2286 & n4158 ;
  assign n4170 = ~n1409 & n3594 ;
  assign n4171 = ~x65 & n4170 ;
  assign n4168 = n3063 ^ n2066 ^ n591 ;
  assign n4160 = ( n235 & n397 ) | ( n235 & ~n1884 ) | ( n397 & ~n1884 ) ;
  assign n4161 = ( n255 & ~n1050 ) | ( n255 & n4160 ) | ( ~n1050 & n4160 ) ;
  assign n4162 = ~n509 & n2015 ;
  assign n4163 = ( n1016 & n3664 ) | ( n1016 & n4162 ) | ( n3664 & n4162 ) ;
  assign n4164 = n1550 ^ n790 ^ 1'b0 ;
  assign n4165 = n4163 & ~n4164 ;
  assign n4166 = ( n1536 & n3259 ) | ( n1536 & ~n4165 ) | ( n3259 & ~n4165 ) ;
  assign n4167 = ( n3562 & n4161 ) | ( n3562 & n4166 ) | ( n4161 & n4166 ) ;
  assign n4169 = n4168 ^ n4167 ^ n3193 ;
  assign n4172 = n4171 ^ n4169 ^ n474 ;
  assign n4176 = n2396 ^ n964 ^ n312 ;
  assign n4177 = n4176 ^ n1941 ^ 1'b0 ;
  assign n4178 = n4177 ^ n3593 ^ n2021 ;
  assign n4179 = n1848 & ~n4178 ;
  assign n4173 = n2557 ^ n1151 ^ n366 ;
  assign n4174 = ( n2094 & n3285 ) | ( n2094 & ~n4173 ) | ( n3285 & ~n4173 ) ;
  assign n4175 = ( ~n1126 & n3821 ) | ( ~n1126 & n4174 ) | ( n3821 & n4174 ) ;
  assign n4180 = n4179 ^ n4175 ^ n2539 ;
  assign n4181 = n2260 ^ n786 ^ 1'b0 ;
  assign n4182 = n1938 ^ n553 ^ 1'b0 ;
  assign n4183 = ~n4181 & n4182 ;
  assign n4184 = n3057 ^ n2204 ^ n1792 ;
  assign n4185 = ( n1286 & n4183 ) | ( n1286 & ~n4184 ) | ( n4183 & ~n4184 ) ;
  assign n4186 = ( n1027 & ~n2487 ) | ( n1027 & n4185 ) | ( ~n2487 & n4185 ) ;
  assign n4187 = ( n1229 & n1314 ) | ( n1229 & ~n2666 ) | ( n1314 & ~n2666 ) ;
  assign n4188 = n4187 ^ n628 ^ 1'b0 ;
  assign n4190 = ( x121 & n232 ) | ( x121 & n707 ) | ( n232 & n707 ) ;
  assign n4189 = n695 ^ n314 ^ 1'b0 ;
  assign n4191 = n4190 ^ n4189 ^ n187 ;
  assign n4192 = n4191 ^ n2083 ^ 1'b0 ;
  assign n4193 = n2421 & ~n4192 ;
  assign n4194 = ( n1664 & ~n2060 ) | ( n1664 & n3188 ) | ( ~n2060 & n3188 ) ;
  assign n4195 = ( n1856 & ~n1928 ) | ( n1856 & n4194 ) | ( ~n1928 & n4194 ) ;
  assign n4196 = n2429 ^ n1713 ^ n1200 ;
  assign n4198 = ~n1069 & n1281 ;
  assign n4199 = n2532 & n4198 ;
  assign n4200 = n4199 ^ n2174 ^ n920 ;
  assign n4201 = n4200 ^ n1960 ^ n1555 ;
  assign n4202 = n868 | n4201 ;
  assign n4197 = n1841 | n2760 ;
  assign n4203 = n4202 ^ n4197 ^ 1'b0 ;
  assign n4204 = ( n1312 & n4196 ) | ( n1312 & n4203 ) | ( n4196 & n4203 ) ;
  assign n4205 = ( ~n1188 & n4195 ) | ( ~n1188 & n4204 ) | ( n4195 & n4204 ) ;
  assign n4213 = ( ~n1546 & n1701 ) | ( ~n1546 & n2977 ) | ( n1701 & n2977 ) ;
  assign n4206 = n575 & ~n627 ;
  assign n4207 = n1295 & n4206 ;
  assign n4209 = n2557 ^ n2532 ^ 1'b0 ;
  assign n4210 = ~n2858 & n4209 ;
  assign n4208 = n2859 ^ n1721 ^ n1338 ;
  assign n4211 = n4210 ^ n4208 ^ n2360 ;
  assign n4212 = ~n4207 & n4211 ;
  assign n4214 = n4213 ^ n4212 ^ 1'b0 ;
  assign n4215 = n3881 ^ n2333 ^ 1'b0 ;
  assign n4216 = n2418 & n4215 ;
  assign n4217 = n1520 ^ n854 ^ n145 ;
  assign n4218 = n4217 ^ n1865 ^ n951 ;
  assign n4219 = n4218 ^ n1902 ^ 1'b0 ;
  assign n4220 = n1335 ^ n710 ^ 1'b0 ;
  assign n4221 = n2419 & ~n4220 ;
  assign n4222 = n1166 ^ n794 ^ n167 ;
  assign n4223 = n4222 ^ n1728 ^ n142 ;
  assign n4227 = ( n416 & n1588 ) | ( n416 & ~n3281 ) | ( n1588 & ~n3281 ) ;
  assign n4224 = x115 & n2420 ;
  assign n4225 = ( n2949 & n3680 ) | ( n2949 & n4224 ) | ( n3680 & n4224 ) ;
  assign n4226 = ~n2890 & n4225 ;
  assign n4228 = n4227 ^ n4226 ^ 1'b0 ;
  assign n4229 = n2179 ^ n1717 ^ 1'b0 ;
  assign n4230 = n4134 | n4229 ;
  assign n4231 = ( ~n850 & n1024 ) | ( ~n850 & n2666 ) | ( n1024 & n2666 ) ;
  assign n4232 = n4231 ^ n1156 ^ n458 ;
  assign n4233 = n1141 & n1159 ;
  assign n4234 = n4233 ^ n624 ^ x26 ;
  assign n4235 = n282 | n1615 ;
  assign n4236 = n4235 ^ n2435 ^ n1241 ;
  assign n4237 = n3953 | n4236 ;
  assign n4238 = n840 | n4237 ;
  assign n4239 = ( n4232 & n4234 ) | ( n4232 & n4238 ) | ( n4234 & n4238 ) ;
  assign n4240 = ( n793 & ~n1248 ) | ( n793 & n3102 ) | ( ~n1248 & n3102 ) ;
  assign n4241 = ( n170 & ~n1802 ) | ( n170 & n4240 ) | ( ~n1802 & n4240 ) ;
  assign n4242 = ( n1100 & n1383 ) | ( n1100 & ~n4241 ) | ( n1383 & ~n4241 ) ;
  assign n4246 = n1744 ^ n1615 ^ n343 ;
  assign n4247 = n1895 ^ n1531 ^ x43 ;
  assign n4248 = n3220 ^ n2023 ^ x13 ;
  assign n4249 = ( n4246 & n4247 ) | ( n4246 & ~n4248 ) | ( n4247 & ~n4248 ) ;
  assign n4250 = ~n2328 & n4249 ;
  assign n4251 = n334 & n4250 ;
  assign n4243 = ( n237 & n2843 ) | ( n237 & ~n3279 ) | ( n2843 & ~n3279 ) ;
  assign n4244 = ( ~n389 & n1485 ) | ( ~n389 & n2338 ) | ( n1485 & n2338 ) ;
  assign n4245 = n4243 & n4244 ;
  assign n4252 = n4251 ^ n4245 ^ 1'b0 ;
  assign n4254 = ( n226 & n480 ) | ( n226 & n1294 ) | ( n480 & n1294 ) ;
  assign n4253 = n1738 & n3547 ;
  assign n4255 = n4254 ^ n4253 ^ n3249 ;
  assign n4256 = n1124 | n3981 ;
  assign n4257 = n4256 ^ n1585 ^ 1'b0 ;
  assign n4258 = ( n816 & n1531 ) | ( n816 & ~n4257 ) | ( n1531 & ~n4257 ) ;
  assign n4259 = ( n2245 & ~n3559 ) | ( n2245 & n4168 ) | ( ~n3559 & n4168 ) ;
  assign n4263 = n3197 ^ n733 ^ n595 ;
  assign n4260 = ( n158 & n381 ) | ( n158 & ~n2274 ) | ( n381 & ~n2274 ) ;
  assign n4261 = ( n896 & n2220 ) | ( n896 & n4260 ) | ( n2220 & n4260 ) ;
  assign n4262 = n4261 ^ n2916 ^ n1899 ;
  assign n4264 = n4263 ^ n4262 ^ n1254 ;
  assign n4265 = n1401 & ~n2147 ;
  assign n4266 = ~n2065 & n4265 ;
  assign n4267 = n3508 ^ n1814 ^ n1203 ;
  assign n4268 = ( n1243 & n1946 ) | ( n1243 & ~n4267 ) | ( n1946 & ~n4267 ) ;
  assign n4269 = ( n2137 & n4266 ) | ( n2137 & n4268 ) | ( n4266 & n4268 ) ;
  assign n4272 = ( ~n207 & n1139 ) | ( ~n207 & n2890 ) | ( n1139 & n2890 ) ;
  assign n4270 = n517 & ~n1156 ;
  assign n4271 = n4270 ^ n2830 ^ n598 ;
  assign n4273 = n4272 ^ n4271 ^ n399 ;
  assign n4274 = n4078 ^ n1269 ^ 1'b0 ;
  assign n4275 = ~n2355 & n4274 ;
  assign n4279 = n2304 & n3973 ;
  assign n4280 = n2749 & n4279 ;
  assign n4276 = n1760 & ~n3652 ;
  assign n4277 = n1542 & n4276 ;
  assign n4278 = ( ~n2134 & n3467 ) | ( ~n2134 & n4277 ) | ( n3467 & n4277 ) ;
  assign n4281 = n4280 ^ n4278 ^ 1'b0 ;
  assign n4282 = n2189 | n2244 ;
  assign n4283 = n2963 ^ n1464 ^ n596 ;
  assign n4284 = n4283 ^ n2515 ^ n395 ;
  assign n4289 = n2945 ^ n1254 ^ 1'b0 ;
  assign n4290 = ( ~n940 & n3803 ) | ( ~n940 & n4289 ) | ( n3803 & n4289 ) ;
  assign n4285 = n317 & ~n525 ;
  assign n4286 = ( ~n423 & n1578 ) | ( ~n423 & n4285 ) | ( n1578 & n4285 ) ;
  assign n4287 = n501 & ~n4286 ;
  assign n4288 = ( n881 & n2202 ) | ( n881 & n4287 ) | ( n2202 & n4287 ) ;
  assign n4291 = n4290 ^ n4288 ^ n678 ;
  assign n4292 = ( n209 & n657 ) | ( n209 & ~n2276 ) | ( n657 & ~n2276 ) ;
  assign n4293 = n1789 | n4292 ;
  assign n4294 = n1627 & ~n4293 ;
  assign n4295 = ( n723 & n2725 ) | ( n723 & ~n4294 ) | ( n2725 & ~n4294 ) ;
  assign n4296 = ( n633 & n1744 ) | ( n633 & ~n3716 ) | ( n1744 & ~n3716 ) ;
  assign n4298 = ( x36 & x48 ) | ( x36 & n3779 ) | ( x48 & n3779 ) ;
  assign n4297 = n747 & ~n1552 ;
  assign n4299 = n4298 ^ n4297 ^ 1'b0 ;
  assign n4300 = ( n4295 & ~n4296 ) | ( n4295 & n4299 ) | ( ~n4296 & n4299 ) ;
  assign n4301 = ( n3016 & n3024 ) | ( n3016 & n4300 ) | ( n3024 & n4300 ) ;
  assign n4302 = ( n1188 & n2216 ) | ( n1188 & n2997 ) | ( n2216 & n2997 ) ;
  assign n4303 = n315 & n465 ;
  assign n4304 = n4303 ^ n2558 ^ n1171 ;
  assign n4305 = n678 & n3264 ;
  assign n4306 = n4305 ^ n3168 ^ 1'b0 ;
  assign n4307 = n3677 & ~n4306 ;
  assign n4308 = n4304 & n4307 ;
  assign n4309 = n4308 ^ n226 ^ 1'b0 ;
  assign n4310 = ( ~x39 & n4302 ) | ( ~x39 & n4309 ) | ( n4302 & n4309 ) ;
  assign n4311 = n4310 ^ n1171 ^ n829 ;
  assign n4312 = n937 & ~n985 ;
  assign n4313 = ~n426 & n4312 ;
  assign n4314 = n4313 ^ n2936 ^ 1'b0 ;
  assign n4315 = n2660 | n4314 ;
  assign n4316 = ( ~n2783 & n3229 ) | ( ~n2783 & n4315 ) | ( n3229 & n4315 ) ;
  assign n4321 = n2200 ^ n1510 ^ n232 ;
  assign n4322 = n4321 ^ n418 ^ x86 ;
  assign n4317 = n201 & ~n2666 ;
  assign n4318 = n1427 & n4317 ;
  assign n4319 = n1050 | n4318 ;
  assign n4320 = n4319 ^ n2819 ^ 1'b0 ;
  assign n4323 = n4322 ^ n4320 ^ 1'b0 ;
  assign n4324 = n928 ^ x83 ^ 1'b0 ;
  assign n4325 = n800 ^ n704 ^ 1'b0 ;
  assign n4326 = ( n2384 & n4324 ) | ( n2384 & ~n4325 ) | ( n4324 & ~n4325 ) ;
  assign n4327 = n4326 ^ n3478 ^ n1928 ;
  assign n4328 = ( n642 & n4323 ) | ( n642 & ~n4327 ) | ( n4323 & ~n4327 ) ;
  assign n4329 = n525 | n1272 ;
  assign n4330 = n255 | n4329 ;
  assign n4331 = n4267 ^ n3101 ^ n145 ;
  assign n4332 = n4331 ^ n1274 ^ 1'b0 ;
  assign n4338 = n977 & ~n3890 ;
  assign n4339 = ~n1917 & n4338 ;
  assign n4340 = ~n576 & n4339 ;
  assign n4335 = n1821 ^ n1225 ^ 1'b0 ;
  assign n4336 = ~n1193 & n4335 ;
  assign n4337 = ( n1901 & n3059 ) | ( n1901 & ~n4336 ) | ( n3059 & ~n4336 ) ;
  assign n4341 = n4340 ^ n4337 ^ n2989 ;
  assign n4333 = ( n1865 & n2850 ) | ( n1865 & n3407 ) | ( n2850 & n3407 ) ;
  assign n4334 = ( n1467 & ~n3395 ) | ( n1467 & n4333 ) | ( ~n3395 & n4333 ) ;
  assign n4342 = n4341 ^ n4334 ^ n3977 ;
  assign n4344 = n2251 ^ n1639 ^ n838 ;
  assign n4343 = n1924 & ~n3746 ;
  assign n4345 = n4344 ^ n4343 ^ 1'b0 ;
  assign n4349 = n567 & n1396 ;
  assign n4350 = n4349 ^ n1217 ^ 1'b0 ;
  assign n4351 = ( ~n2806 & n3316 ) | ( ~n2806 & n4350 ) | ( n3316 & n4350 ) ;
  assign n4352 = n1193 | n4351 ;
  assign n4346 = ~x108 & n2079 ;
  assign n4347 = n1218 | n4346 ;
  assign n4348 = n1193 & ~n4347 ;
  assign n4353 = n4352 ^ n4348 ^ 1'b0 ;
  assign n4354 = n1852 | n4353 ;
  assign n4356 = n3212 ^ n1580 ^ n828 ;
  assign n4357 = n2618 ^ n1174 ^ n1170 ;
  assign n4358 = n4357 ^ n3086 ^ n924 ;
  assign n4359 = ~n3546 & n4358 ;
  assign n4360 = n4356 & n4359 ;
  assign n4355 = n4202 ^ n2877 ^ n450 ;
  assign n4361 = n4360 ^ n4355 ^ n659 ;
  assign n4362 = n2006 ^ n899 ^ 1'b0 ;
  assign n4364 = n3875 ^ n3873 ^ n1910 ;
  assign n4363 = ( n1324 & n1496 ) | ( n1324 & n3336 ) | ( n1496 & n3336 ) ;
  assign n4365 = n4364 ^ n4363 ^ n207 ;
  assign n4366 = ( n2144 & ~n4362 ) | ( n2144 & n4365 ) | ( ~n4362 & n4365 ) ;
  assign n4367 = n4366 ^ n2464 ^ 1'b0 ;
  assign n4371 = n1974 ^ n1565 ^ n395 ;
  assign n4368 = n533 ^ n179 ^ x28 ;
  assign n4369 = n1707 ^ n1678 ^ 1'b0 ;
  assign n4370 = ( n1626 & n4368 ) | ( n1626 & n4369 ) | ( n4368 & n4369 ) ;
  assign n4372 = n4371 ^ n4370 ^ n523 ;
  assign n4373 = ( n1726 & ~n2861 ) | ( n1726 & n2871 ) | ( ~n2861 & n2871 ) ;
  assign n4380 = n477 | n1423 ;
  assign n4381 = n717 | n4380 ;
  assign n4382 = ( ~n150 & n3048 ) | ( ~n150 & n4381 ) | ( n3048 & n4381 ) ;
  assign n4383 = n818 & n4382 ;
  assign n4374 = n1787 ^ n867 ^ 1'b0 ;
  assign n4375 = n4374 ^ n3854 ^ x92 ;
  assign n4376 = n4375 ^ n3220 ^ n332 ;
  assign n4377 = ( n529 & n613 ) | ( n529 & n1568 ) | ( n613 & n1568 ) ;
  assign n4378 = ( n1502 & ~n1682 ) | ( n1502 & n4377 ) | ( ~n1682 & n4377 ) ;
  assign n4379 = ( ~n2115 & n4376 ) | ( ~n2115 & n4378 ) | ( n4376 & n4378 ) ;
  assign n4384 = n4383 ^ n4379 ^ n2830 ;
  assign n4385 = n4373 & ~n4384 ;
  assign n4386 = ~n4372 & n4385 ;
  assign n4387 = n2876 ^ n572 ^ 1'b0 ;
  assign n4388 = ( n801 & ~n1072 ) | ( n801 & n4387 ) | ( ~n1072 & n4387 ) ;
  assign n4389 = ( n1108 & n1218 ) | ( n1108 & ~n4099 ) | ( n1218 & ~n4099 ) ;
  assign n4391 = n2499 & n2650 ;
  assign n4392 = n2043 & n4391 ;
  assign n4390 = n3717 ^ n2094 ^ n250 ;
  assign n4393 = n4392 ^ n4390 ^ 1'b0 ;
  assign n4394 = ~n4389 & n4393 ;
  assign n4395 = n3868 ^ n3094 ^ n2193 ;
  assign n4396 = n1362 ^ n769 ^ n171 ;
  assign n4397 = n4396 ^ n1802 ^ 1'b0 ;
  assign n4398 = ~n974 & n4397 ;
  assign n4399 = ( n680 & n1849 ) | ( n680 & n4398 ) | ( n1849 & n4398 ) ;
  assign n4400 = ( n2363 & n2930 ) | ( n2363 & ~n4399 ) | ( n2930 & ~n4399 ) ;
  assign n4401 = ( n2427 & ~n2719 ) | ( n2427 & n4400 ) | ( ~n2719 & n4400 ) ;
  assign n4402 = n4395 & n4401 ;
  assign n4403 = n4402 ^ n2465 ^ 1'b0 ;
  assign n4404 = n4403 ^ n2453 ^ n408 ;
  assign n4405 = n869 & n4404 ;
  assign n4406 = n3120 ^ n2076 ^ n903 ;
  assign n4407 = x79 & n1637 ;
  assign n4408 = ( n1268 & n2598 ) | ( n1268 & ~n2910 ) | ( n2598 & ~n2910 ) ;
  assign n4409 = ( ~n891 & n4407 ) | ( ~n891 & n4408 ) | ( n4407 & n4408 ) ;
  assign n4410 = ( n1549 & n4406 ) | ( n1549 & n4409 ) | ( n4406 & n4409 ) ;
  assign n4413 = n1259 & ~n1733 ;
  assign n4411 = n368 & ~n1390 ;
  assign n4412 = n1966 & n4411 ;
  assign n4414 = n4413 ^ n4412 ^ n2440 ;
  assign n4415 = ( ~n1415 & n4410 ) | ( ~n1415 & n4414 ) | ( n4410 & n4414 ) ;
  assign n4424 = n2218 ^ x88 ^ x33 ;
  assign n4425 = n4424 ^ n689 ^ x74 ;
  assign n4420 = n1032 ^ n898 ^ 1'b0 ;
  assign n4416 = n911 ^ n178 ^ 1'b0 ;
  assign n4417 = n1493 & n4416 ;
  assign n4418 = ( n452 & ~n616 ) | ( n452 & n879 ) | ( ~n616 & n879 ) ;
  assign n4419 = n4417 | n4418 ;
  assign n4421 = n4420 ^ n4419 ^ n541 ;
  assign n4422 = n4421 ^ n3166 ^ n2463 ;
  assign n4423 = ( n1154 & ~n1992 ) | ( n1154 & n4422 ) | ( ~n1992 & n4422 ) ;
  assign n4426 = n4425 ^ n4423 ^ n1447 ;
  assign n4427 = n3849 & ~n4426 ;
  assign n4428 = n4427 ^ n1753 ^ 1'b0 ;
  assign n4429 = n1699 ^ n1690 ^ n1625 ;
  assign n4430 = n4295 & ~n4429 ;
  assign n4431 = n4428 | n4430 ;
  assign n4432 = n4431 ^ n4075 ^ 1'b0 ;
  assign n4433 = ( x124 & n442 ) | ( x124 & ~n1121 ) | ( n442 & ~n1121 ) ;
  assign n4434 = n4433 ^ n3591 ^ n915 ;
  assign n4436 = n400 & ~n1069 ;
  assign n4437 = n4436 ^ n200 ^ 1'b0 ;
  assign n4438 = n1387 & n4437 ;
  assign n4439 = n1049 & n4438 ;
  assign n4440 = n4439 ^ n3243 ^ n2270 ;
  assign n4435 = n3967 ^ n3149 ^ n1054 ;
  assign n4441 = n4440 ^ n4435 ^ x103 ;
  assign n4442 = ( n681 & n4434 ) | ( n681 & ~n4441 ) | ( n4434 & ~n4441 ) ;
  assign n4443 = n1849 & n3260 ;
  assign n4444 = ( ~n412 & n855 ) | ( ~n412 & n859 ) | ( n855 & n859 ) ;
  assign n4445 = ( n2157 & ~n2502 ) | ( n2157 & n2535 ) | ( ~n2502 & n2535 ) ;
  assign n4446 = ( n163 & ~n4444 ) | ( n163 & n4445 ) | ( ~n4444 & n4445 ) ;
  assign n4447 = n4009 ^ n2267 ^ n1274 ;
  assign n4448 = ( ~n1847 & n3081 ) | ( ~n1847 & n4447 ) | ( n3081 & n4447 ) ;
  assign n4449 = n2029 | n2782 ;
  assign n4450 = n4449 ^ n996 ^ 1'b0 ;
  assign n4451 = ( n896 & n1136 ) | ( n896 & n4407 ) | ( n1136 & n4407 ) ;
  assign n4452 = ( ~n623 & n722 ) | ( ~n623 & n1410 ) | ( n722 & n1410 ) ;
  assign n4453 = ( n2938 & ~n4161 ) | ( n2938 & n4452 ) | ( ~n4161 & n4452 ) ;
  assign n4454 = ~n1567 & n4453 ;
  assign n4455 = n4454 ^ n1687 ^ 1'b0 ;
  assign n4456 = ( n4450 & n4451 ) | ( n4450 & n4455 ) | ( n4451 & n4455 ) ;
  assign n4457 = n1250 & n4456 ;
  assign n4458 = ~n2358 & n4457 ;
  assign n4459 = n2974 ^ n746 ^ 1'b0 ;
  assign n4460 = ( n3157 & ~n4458 ) | ( n3157 & n4459 ) | ( ~n4458 & n4459 ) ;
  assign n4461 = ( n1076 & n2421 ) | ( n1076 & n4306 ) | ( n2421 & n4306 ) ;
  assign n4462 = x19 & n1580 ;
  assign n4463 = ~n3496 & n4462 ;
  assign n4464 = ~n940 & n2730 ;
  assign n4465 = n2251 & n4464 ;
  assign n4466 = ( n395 & n3858 ) | ( n395 & n4465 ) | ( n3858 & n4465 ) ;
  assign n4467 = n4466 ^ n1998 ^ 1'b0 ;
  assign n4468 = ~n4463 & n4467 ;
  assign n4469 = n4468 ^ n272 ^ 1'b0 ;
  assign n4470 = ( n2153 & n4461 ) | ( n2153 & ~n4469 ) | ( n4461 & ~n4469 ) ;
  assign n4471 = ( n398 & ~n1987 ) | ( n398 & n2849 ) | ( ~n1987 & n2849 ) ;
  assign n4472 = ( ~x111 & n1503 ) | ( ~x111 & n1647 ) | ( n1503 & n1647 ) ;
  assign n4473 = ( ~n2971 & n3195 ) | ( ~n2971 & n4472 ) | ( n3195 & n4472 ) ;
  assign n4474 = ( n249 & ~n860 ) | ( n249 & n4473 ) | ( ~n860 & n4473 ) ;
  assign n4475 = n4474 ^ n2677 ^ 1'b0 ;
  assign n4476 = n1582 & ~n4475 ;
  assign n4477 = n4476 ^ n3020 ^ n1617 ;
  assign n4478 = n4321 ^ n2990 ^ n798 ;
  assign n4479 = n4478 ^ n3302 ^ n1013 ;
  assign n4480 = ( n4471 & n4477 ) | ( n4471 & n4479 ) | ( n4477 & n4479 ) ;
  assign n4481 = n2070 & ~n2837 ;
  assign n4488 = ( ~n869 & n1022 ) | ( ~n869 & n1544 ) | ( n1022 & n1544 ) ;
  assign n4485 = ( n1887 & ~n2554 ) | ( n1887 & n3420 ) | ( ~n2554 & n3420 ) ;
  assign n4486 = n2106 ^ n1491 ^ n1269 ;
  assign n4487 = ( n427 & n4485 ) | ( n427 & n4486 ) | ( n4485 & n4486 ) ;
  assign n4482 = n3508 ^ n1680 ^ n411 ;
  assign n4483 = n1129 | n4482 ;
  assign n4484 = n2464 | n4483 ;
  assign n4489 = n4488 ^ n4487 ^ n4484 ;
  assign n4490 = ( n2874 & n4481 ) | ( n2874 & n4489 ) | ( n4481 & n4489 ) ;
  assign n4491 = n1212 & n2173 ;
  assign n4492 = n2745 | n4491 ;
  assign n4493 = n4492 ^ n3251 ^ 1'b0 ;
  assign n4494 = ( n373 & n725 ) | ( n373 & ~n1141 ) | ( n725 & ~n1141 ) ;
  assign n4495 = n276 & n4494 ;
  assign n4496 = n4495 ^ n1803 ^ 1'b0 ;
  assign n4497 = ( n2662 & ~n3039 ) | ( n2662 & n4389 ) | ( ~n3039 & n4389 ) ;
  assign n4498 = n1957 & ~n4497 ;
  assign n4499 = n4498 ^ n2836 ^ 1'b0 ;
  assign n4500 = n2674 & n4187 ;
  assign n4501 = ( n4496 & n4499 ) | ( n4496 & ~n4500 ) | ( n4499 & ~n4500 ) ;
  assign n4502 = n3746 ^ n1503 ^ n813 ;
  assign n4503 = n492 | n4502 ;
  assign n4504 = ( n1347 & ~n1544 ) | ( n1347 & n4503 ) | ( ~n1544 & n4503 ) ;
  assign n4505 = n3116 ^ n2786 ^ n1533 ;
  assign n4506 = n4505 ^ n3643 ^ n1672 ;
  assign n4512 = ~n436 & n4064 ;
  assign n4513 = n4512 ^ n1757 ^ 1'b0 ;
  assign n4509 = n2960 & ~n3342 ;
  assign n4510 = n4509 ^ n1517 ^ 1'b0 ;
  assign n4507 = n4292 ^ n3952 ^ 1'b0 ;
  assign n4508 = n4507 ^ n3164 ^ n550 ;
  assign n4511 = n4510 ^ n4508 ^ x50 ;
  assign n4514 = n4513 ^ n4511 ^ n4134 ;
  assign n4515 = n4514 ^ n2581 ^ 1'b0 ;
  assign n4516 = ( n1597 & ~n1708 ) | ( n1597 & n4515 ) | ( ~n1708 & n4515 ) ;
  assign n4518 = x49 & n3435 ;
  assign n4519 = n4518 ^ n199 ^ 1'b0 ;
  assign n4520 = n4519 ^ n2320 ^ n1972 ;
  assign n4517 = ~n2507 & n2584 ;
  assign n4521 = n4520 ^ n4517 ^ 1'b0 ;
  assign n4522 = ( n2560 & n3573 ) | ( n2560 & ~n3949 ) | ( n3573 & ~n3949 ) ;
  assign n4523 = n1171 | n3518 ;
  assign n4524 = n1390 & ~n4523 ;
  assign n4525 = n4524 ^ n3139 ^ 1'b0 ;
  assign n4526 = n3407 & n4525 ;
  assign n4527 = n4526 ^ n1743 ^ 1'b0 ;
  assign n4528 = n4527 ^ n3920 ^ n476 ;
  assign n4529 = ( ~n497 & n1318 ) | ( ~n497 & n2210 ) | ( n1318 & n2210 ) ;
  assign n4530 = n4529 ^ n1016 ^ n465 ;
  assign n4531 = n4530 ^ x85 ^ 1'b0 ;
  assign n4532 = x75 & n4531 ;
  assign n4533 = n4532 ^ n2750 ^ x103 ;
  assign n4534 = n4533 ^ n3642 ^ n3088 ;
  assign n4535 = ( ~n766 & n2450 ) | ( ~n766 & n4015 ) | ( n2450 & n4015 ) ;
  assign n4536 = n1629 ^ n1578 ^ n386 ;
  assign n4537 = n4536 ^ n2699 ^ 1'b0 ;
  assign n4538 = n4535 | n4537 ;
  assign n4539 = n1634 | n2507 ;
  assign n4540 = ( n934 & n2717 ) | ( n934 & ~n4539 ) | ( n2717 & ~n4539 ) ;
  assign n4541 = ( n143 & n912 ) | ( n143 & ~n2100 ) | ( n912 & ~n2100 ) ;
  assign n4542 = n2915 ^ n2047 ^ 1'b0 ;
  assign n4543 = ( n3145 & ~n4541 ) | ( n3145 & n4542 ) | ( ~n4541 & n4542 ) ;
  assign n4544 = n3790 ^ n2358 ^ n787 ;
  assign n4545 = n4544 ^ n2880 ^ 1'b0 ;
  assign n4546 = n4322 ^ n1998 ^ 1'b0 ;
  assign n4547 = n2732 ^ n885 ^ n293 ;
  assign n4548 = ( ~n902 & n4546 ) | ( ~n902 & n4547 ) | ( n4546 & n4547 ) ;
  assign n4549 = n3085 ^ n3064 ^ n1045 ;
  assign n4550 = n3832 & n4549 ;
  assign n4551 = n964 | n4550 ;
  assign n4552 = ( n1664 & ~n4548 ) | ( n1664 & n4551 ) | ( ~n4548 & n4551 ) ;
  assign n4556 = n2689 ^ n2422 ^ n1894 ;
  assign n4553 = ( n1006 & ~n2224 ) | ( n1006 & n2760 ) | ( ~n2224 & n2760 ) ;
  assign n4554 = n2724 ^ n2373 ^ 1'b0 ;
  assign n4555 = ( ~n3536 & n4553 ) | ( ~n3536 & n4554 ) | ( n4553 & n4554 ) ;
  assign n4557 = n4556 ^ n4555 ^ n4141 ;
  assign n4558 = ( ~n164 & n1159 ) | ( ~n164 & n2753 ) | ( n1159 & n2753 ) ;
  assign n4559 = n2025 ^ n1482 ^ n1428 ;
  assign n4560 = n4559 ^ n3751 ^ n1113 ;
  assign n4561 = ( x38 & n1663 ) | ( x38 & n2547 ) | ( n1663 & n2547 ) ;
  assign n4562 = ( n196 & n4560 ) | ( n196 & n4561 ) | ( n4560 & n4561 ) ;
  assign n4563 = ( ~n2783 & n4558 ) | ( ~n2783 & n4562 ) | ( n4558 & n4562 ) ;
  assign n4564 = n1560 ^ n1107 ^ 1'b0 ;
  assign n4569 = ( ~n381 & n1944 ) | ( ~n381 & n3518 ) | ( n1944 & n3518 ) ;
  assign n4570 = x84 & n4569 ;
  assign n4571 = n387 & n4570 ;
  assign n4572 = n3609 & ~n4571 ;
  assign n4573 = n2806 & n4572 ;
  assign n4565 = ~n613 & n3341 ;
  assign n4566 = n4174 | n4565 ;
  assign n4567 = n1577 & n4566 ;
  assign n4568 = n4567 ^ n3654 ^ 1'b0 ;
  assign n4574 = n4573 ^ n4568 ^ n2898 ;
  assign n4575 = ( ~n993 & n4564 ) | ( ~n993 & n4574 ) | ( n4564 & n4574 ) ;
  assign n4576 = n2354 & ~n3136 ;
  assign n4577 = n4576 ^ x116 ^ 1'b0 ;
  assign n4578 = n4577 ^ n4564 ^ n642 ;
  assign n4579 = n4578 ^ n3642 ^ n3090 ;
  assign n4586 = x7 & n1402 ;
  assign n4587 = n4586 ^ n782 ^ n572 ;
  assign n4588 = n771 ^ x106 ^ 1'b0 ;
  assign n4589 = n1288 & ~n4588 ;
  assign n4590 = n4587 & n4589 ;
  assign n4580 = n1534 ^ n287 ^ 1'b0 ;
  assign n4581 = ( n177 & ~n1503 ) | ( n177 & n1906 ) | ( ~n1503 & n1906 ) ;
  assign n4582 = n806 & ~n4581 ;
  assign n4583 = ~n3654 & n4582 ;
  assign n4584 = ( n1158 & n2256 ) | ( n1158 & ~n4583 ) | ( n2256 & ~n4583 ) ;
  assign n4585 = ( n1971 & n4580 ) | ( n1971 & ~n4584 ) | ( n4580 & ~n4584 ) ;
  assign n4591 = n4590 ^ n4585 ^ n1035 ;
  assign n4592 = x98 ^ x26 ^ 1'b0 ;
  assign n4593 = ~n676 & n4592 ;
  assign n4594 = n1929 ^ n1790 ^ 1'b0 ;
  assign n4595 = ~n985 & n4594 ;
  assign n4596 = ~n2036 & n4595 ;
  assign n4597 = ~n3616 & n4596 ;
  assign n4598 = n4597 ^ n2995 ^ n135 ;
  assign n4599 = ( n1284 & n2122 ) | ( n1284 & n4598 ) | ( n2122 & n4598 ) ;
  assign n4600 = n4599 ^ n2341 ^ n1300 ;
  assign n4601 = ( n3912 & ~n4593 ) | ( n3912 & n4600 ) | ( ~n4593 & n4600 ) ;
  assign n4604 = ( x56 & n138 ) | ( x56 & ~n1828 ) | ( n138 & ~n1828 ) ;
  assign n4605 = n4604 ^ n926 ^ 1'b0 ;
  assign n4602 = ~n191 & n3264 ;
  assign n4603 = n2355 & n4602 ;
  assign n4606 = n4605 ^ n4603 ^ n2517 ;
  assign n4607 = n3198 & n4606 ;
  assign n4608 = n4607 ^ n2789 ^ 1'b0 ;
  assign n4609 = n3673 ^ n3069 ^ n2330 ;
  assign n4610 = n3362 ^ n3226 ^ n2788 ;
  assign n4611 = n4609 & n4610 ;
  assign n4612 = ( n224 & n2633 ) | ( n224 & n3377 ) | ( n2633 & n3377 ) ;
  assign n4613 = ~n1264 & n2797 ;
  assign n4614 = n4613 ^ n4249 ^ 1'b0 ;
  assign n4615 = n1350 | n3518 ;
  assign n4616 = n2047 & ~n4615 ;
  assign n4617 = n2729 ^ n1034 ^ 1'b0 ;
  assign n4618 = n1084 & n4617 ;
  assign n4619 = ~x124 & n4618 ;
  assign n4620 = ( n654 & ~n4616 ) | ( n654 & n4619 ) | ( ~n4616 & n4619 ) ;
  assign n4621 = n3025 & n4620 ;
  assign n4622 = ~n4614 & n4621 ;
  assign n4623 = ( n947 & n4612 ) | ( n947 & ~n4622 ) | ( n4612 & ~n4622 ) ;
  assign n4624 = n3496 ^ n2096 ^ n1880 ;
  assign n4625 = n3188 | n4624 ;
  assign n4631 = n1926 ^ n1322 ^ n983 ;
  assign n4626 = ( n569 & n944 ) | ( n569 & ~n1371 ) | ( n944 & ~n1371 ) ;
  assign n4627 = n4626 ^ n1661 ^ n1171 ;
  assign n4628 = ( n360 & n3344 ) | ( n360 & ~n4627 ) | ( n3344 & ~n4627 ) ;
  assign n4629 = ( n1014 & n1271 ) | ( n1014 & n4628 ) | ( n1271 & n4628 ) ;
  assign n4630 = ( x47 & ~n2487 ) | ( x47 & n4629 ) | ( ~n2487 & n4629 ) ;
  assign n4632 = n4631 ^ n4630 ^ n1064 ;
  assign n4638 = n880 & n1367 ;
  assign n4639 = ~n2653 & n4638 ;
  assign n4637 = ( ~n448 & n2994 ) | ( ~n448 & n4421 ) | ( n2994 & n4421 ) ;
  assign n4635 = n142 & ~n2615 ;
  assign n4636 = ~n2880 & n4635 ;
  assign n4640 = n4639 ^ n4637 ^ n4636 ;
  assign n4641 = n4640 ^ n1567 ^ n878 ;
  assign n4642 = n4641 ^ n4340 ^ 1'b0 ;
  assign n4633 = ( n1123 & n2843 ) | ( n1123 & n2851 ) | ( n2843 & n2851 ) ;
  assign n4634 = n4200 & ~n4633 ;
  assign n4643 = n4642 ^ n4634 ^ 1'b0 ;
  assign n4644 = n206 ^ n149 ^ 1'b0 ;
  assign n4645 = n407 & n4644 ;
  assign n4646 = ( n1485 & n1767 ) | ( n1485 & ~n4645 ) | ( n1767 & ~n4645 ) ;
  assign n4647 = ( ~n178 & n465 ) | ( ~n178 & n3896 ) | ( n465 & n3896 ) ;
  assign n4648 = n2438 ^ n1280 ^ n510 ;
  assign n4649 = n3876 & ~n4648 ;
  assign n4650 = n4649 ^ n1485 ^ 1'b0 ;
  assign n4651 = ( n1215 & n3603 ) | ( n1215 & ~n4650 ) | ( n3603 & ~n4650 ) ;
  assign n4652 = ( n3921 & n4647 ) | ( n3921 & n4651 ) | ( n4647 & n4651 ) ;
  assign n4653 = ( n4444 & ~n4646 ) | ( n4444 & n4652 ) | ( ~n4646 & n4652 ) ;
  assign n4654 = ( x119 & ~n1702 ) | ( x119 & n2154 ) | ( ~n1702 & n2154 ) ;
  assign n4655 = n2677 ^ n142 ^ 1'b0 ;
  assign n4656 = n4655 ^ n1852 ^ 1'b0 ;
  assign n4657 = n4654 & n4656 ;
  assign n4658 = ( n4339 & ~n4653 ) | ( n4339 & n4657 ) | ( ~n4653 & n4657 ) ;
  assign n4659 = n3306 ^ n2761 ^ n198 ;
  assign n4673 = n1865 ^ n1233 ^ 1'b0 ;
  assign n4674 = n4673 ^ n1175 ^ n1120 ;
  assign n4675 = n4674 ^ n2985 ^ 1'b0 ;
  assign n4676 = ~n1136 & n4675 ;
  assign n4677 = n4676 ^ n2954 ^ n1413 ;
  assign n4668 = n2256 ^ n1639 ^ x47 ;
  assign n4669 = n4668 ^ n2313 ^ n1005 ;
  assign n4670 = n4669 ^ n292 ^ 1'b0 ;
  assign n4671 = n1383 & n4670 ;
  assign n4672 = n4671 ^ n4473 ^ n4207 ;
  assign n4660 = n1436 ^ n1035 ^ n554 ;
  assign n4661 = n1969 & ~n4660 ;
  assign n4662 = n2940 ^ n854 ^ n439 ;
  assign n4663 = n3664 ^ x81 ^ x32 ;
  assign n4664 = ( ~n922 & n3944 ) | ( ~n922 & n4663 ) | ( n3944 & n4663 ) ;
  assign n4665 = ( n229 & ~n2453 ) | ( n229 & n4664 ) | ( ~n2453 & n4664 ) ;
  assign n4666 = n4662 & ~n4665 ;
  assign n4667 = ( n2049 & n4661 ) | ( n2049 & ~n4666 ) | ( n4661 & ~n4666 ) ;
  assign n4678 = n4677 ^ n4672 ^ n4667 ;
  assign n4679 = n1855 ^ n545 ^ 1'b0 ;
  assign n4680 = n2821 & n4679 ;
  assign n4681 = n4680 ^ n4452 ^ n2343 ;
  assign n4682 = ( x29 & ~n1531 ) | ( x29 & n4681 ) | ( ~n1531 & n4681 ) ;
  assign n4683 = n2457 ^ n588 ^ 1'b0 ;
  assign n4707 = n3097 & ~n3270 ;
  assign n4708 = ( n191 & n3367 ) | ( n191 & n4707 ) | ( n3367 & n4707 ) ;
  assign n4693 = n2466 ^ n2361 ^ n255 ;
  assign n4694 = n2775 ^ n583 ^ 1'b0 ;
  assign n4695 = n4693 & ~n4694 ;
  assign n4691 = ( x22 & n184 ) | ( x22 & ~n1350 ) | ( n184 & ~n1350 ) ;
  assign n4688 = n4496 ^ n4222 ^ n986 ;
  assign n4687 = ~n188 & n1144 ;
  assign n4689 = n4688 ^ n4687 ^ 1'b0 ;
  assign n4684 = n1750 ^ n614 ^ x23 ;
  assign n4685 = ( n2912 & n4208 ) | ( n2912 & ~n4684 ) | ( n4208 & ~n4684 ) ;
  assign n4686 = n4292 | n4685 ;
  assign n4690 = n4689 ^ n4686 ^ 1'b0 ;
  assign n4692 = n4691 ^ n4690 ^ n4315 ;
  assign n4696 = n4695 ^ n4692 ^ n4651 ;
  assign n4697 = n4085 ^ n3882 ^ n2751 ;
  assign n4698 = ( n1048 & n1909 ) | ( n1048 & n4697 ) | ( n1909 & n4697 ) ;
  assign n4702 = n2689 ^ n2481 ^ x96 ;
  assign n4703 = ( ~n381 & n3526 ) | ( ~n381 & n4702 ) | ( n3526 & n4702 ) ;
  assign n4699 = n2461 ^ x75 ^ 1'b0 ;
  assign n4700 = n1028 | n4699 ;
  assign n4701 = n4700 ^ n469 ^ 1'b0 ;
  assign n4704 = n4703 ^ n4701 ^ n1313 ;
  assign n4705 = ( n4148 & n4698 ) | ( n4148 & n4704 ) | ( n4698 & n4704 ) ;
  assign n4706 = ~n4696 & n4705 ;
  assign n4709 = n4708 ^ n4706 ^ 1'b0 ;
  assign n4710 = n4709 ^ n3336 ^ n507 ;
  assign n4719 = n3584 ^ n2971 ^ 1'b0 ;
  assign n4713 = ~n251 & n2699 ;
  assign n4714 = n2890 & n4713 ;
  assign n4715 = n2173 ^ n1950 ^ n1908 ;
  assign n4716 = n406 & n4715 ;
  assign n4717 = n4714 & n4716 ;
  assign n4718 = ( n4036 & n4389 ) | ( n4036 & ~n4717 ) | ( n4389 & ~n4717 ) ;
  assign n4711 = ( n333 & n645 ) | ( n333 & ~n1313 ) | ( n645 & ~n1313 ) ;
  assign n4712 = n4711 ^ n3815 ^ n3621 ;
  assign n4720 = n4719 ^ n4718 ^ n4712 ;
  assign n4723 = n3121 ^ n1493 ^ 1'b0 ;
  assign n4724 = n4723 ^ n1046 ^ n512 ;
  assign n4725 = n3227 & ~n4724 ;
  assign n4721 = ( n255 & ~n1790 ) | ( n255 & n4605 ) | ( ~n1790 & n4605 ) ;
  assign n4722 = n4721 ^ n2236 ^ n1675 ;
  assign n4726 = n4725 ^ n4722 ^ n4721 ;
  assign n4727 = ~n223 & n2127 ;
  assign n4728 = n474 & n4727 ;
  assign n4729 = n4728 ^ n3210 ^ n958 ;
  assign n4730 = n4729 ^ n4587 ^ n2496 ;
  assign n4731 = ( ~n736 & n1245 ) | ( ~n736 & n4730 ) | ( n1245 & n4730 ) ;
  assign n4732 = n2739 ^ n1097 ^ n689 ;
  assign n4733 = ( ~n1582 & n4731 ) | ( ~n1582 & n4732 ) | ( n4731 & n4732 ) ;
  assign n4740 = n1806 ^ n1698 ^ 1'b0 ;
  assign n4738 = n1796 ^ n158 ^ 1'b0 ;
  assign n4739 = n1089 & ~n4738 ;
  assign n4741 = n4740 ^ n4739 ^ n339 ;
  assign n4734 = ( n906 & ~n1626 ) | ( n906 & n2729 ) | ( ~n1626 & n2729 ) ;
  assign n4735 = ( n131 & n2167 ) | ( n131 & ~n4734 ) | ( n2167 & ~n4734 ) ;
  assign n4736 = n4735 ^ n1119 ^ 1'b0 ;
  assign n4737 = n4172 & ~n4736 ;
  assign n4742 = n4741 ^ n4737 ^ n3078 ;
  assign n4743 = ( ~n2897 & n4733 ) | ( ~n2897 & n4742 ) | ( n4733 & n4742 ) ;
  assign n4744 = ( n1265 & n3769 ) | ( n1265 & ~n3993 ) | ( n3769 & ~n3993 ) ;
  assign n4745 = n2609 ^ n734 ^ x53 ;
  assign n4746 = ( n404 & ~n4744 ) | ( n404 & n4745 ) | ( ~n4744 & n4745 ) ;
  assign n4747 = n3341 ^ n2081 ^ 1'b0 ;
  assign n4748 = n508 ^ x33 ^ x21 ;
  assign n4749 = n4748 ^ n1659 ^ 1'b0 ;
  assign n4750 = ~n3246 & n4328 ;
  assign n4751 = n4750 ^ n2465 ^ 1'b0 ;
  assign n4757 = n2411 ^ n885 ^ n299 ;
  assign n4758 = n1410 & n4757 ;
  assign n4759 = n4758 ^ n3593 ^ 1'b0 ;
  assign n4752 = ( ~n411 & n681 ) | ( ~n411 & n1166 ) | ( n681 & n1166 ) ;
  assign n4753 = n3406 ^ n2885 ^ 1'b0 ;
  assign n4754 = n3766 & n4753 ;
  assign n4755 = ( n3854 & n4752 ) | ( n3854 & n4754 ) | ( n4752 & n4754 ) ;
  assign n4756 = n4755 ^ n2981 ^ n2019 ;
  assign n4760 = n4759 ^ n4756 ^ n1262 ;
  assign n4761 = n4760 ^ n4201 ^ 1'b0 ;
  assign n4764 = ( n292 & n811 ) | ( n292 & n1013 ) | ( n811 & n1013 ) ;
  assign n4763 = n3070 ^ n502 ^ 1'b0 ;
  assign n4765 = n4764 ^ n4763 ^ n173 ;
  assign n4762 = n692 ^ n580 ^ 1'b0 ;
  assign n4766 = n4765 ^ n4762 ^ 1'b0 ;
  assign n4769 = n3784 ^ n3128 ^ 1'b0 ;
  assign n4770 = n4769 ^ n1847 ^ n1105 ;
  assign n4767 = ( n859 & n887 ) | ( n859 & n922 ) | ( n887 & n922 ) ;
  assign n4768 = ( ~n588 & n2201 ) | ( ~n588 & n4767 ) | ( n2201 & n4767 ) ;
  assign n4771 = n4770 ^ n4768 ^ n502 ;
  assign n4772 = n4559 ^ n1822 ^ n1332 ;
  assign n4773 = n4772 ^ n3875 ^ n2730 ;
  assign n4774 = n4773 ^ n4023 ^ n2958 ;
  assign n4775 = n4774 ^ n2559 ^ 1'b0 ;
  assign n4776 = n2890 ^ n1138 ^ 1'b0 ;
  assign n4777 = n3882 ^ n886 ^ 1'b0 ;
  assign n4778 = n4777 ^ n3230 ^ n367 ;
  assign n4779 = n3020 & n4778 ;
  assign n4780 = n4779 ^ n3450 ^ 1'b0 ;
  assign n4781 = ( n833 & n1939 ) | ( n833 & ~n4780 ) | ( n1939 & ~n4780 ) ;
  assign n4782 = n4417 ^ n607 ^ n153 ;
  assign n4783 = ( n2458 & n3449 ) | ( n2458 & n4782 ) | ( n3449 & n4782 ) ;
  assign n4784 = n4783 ^ n2844 ^ x36 ;
  assign n4785 = n4784 ^ n3262 ^ n2403 ;
  assign n4792 = ( n865 & ~n1257 ) | ( n865 & n4444 ) | ( ~n1257 & n4444 ) ;
  assign n4793 = n611 ^ x0 ^ 1'b0 ;
  assign n4794 = n4792 & ~n4793 ;
  assign n4795 = n2277 & n4794 ;
  assign n4790 = n1867 & ~n3045 ;
  assign n4791 = n3111 & n4790 ;
  assign n4796 = n4795 ^ n4791 ^ n2338 ;
  assign n4797 = n2419 & n4796 ;
  assign n4798 = n4797 ^ n456 ^ 1'b0 ;
  assign n4786 = ( n2976 & n3012 ) | ( n2976 & ~n3860 ) | ( n3012 & ~n3860 ) ;
  assign n4787 = n2206 ^ n750 ^ 1'b0 ;
  assign n4788 = n4786 | n4787 ;
  assign n4789 = n4569 & ~n4788 ;
  assign n4799 = n4798 ^ n4789 ^ 1'b0 ;
  assign n4800 = n2222 ^ n425 ^ 1'b0 ;
  assign n4801 = x114 & ~n4800 ;
  assign n4802 = n4207 ^ n1563 ^ 1'b0 ;
  assign n4803 = n4802 ^ n4425 ^ n2183 ;
  assign n4804 = n4803 ^ n763 ^ n189 ;
  assign n4805 = n2235 & n3816 ;
  assign n4806 = n4804 & n4805 ;
  assign n4807 = ~n4370 & n4584 ;
  assign n4808 = n4806 & n4807 ;
  assign n4809 = n640 ^ n529 ^ n447 ;
  assign n4810 = n4809 ^ n4422 ^ n2038 ;
  assign n4811 = n2938 ^ n1073 ^ n432 ;
  assign n4812 = n4811 ^ n1971 ^ n1848 ;
  assign n4813 = ( n181 & ~n2609 ) | ( n181 & n4812 ) | ( ~n2609 & n4812 ) ;
  assign n4814 = n2425 & ~n4813 ;
  assign n4815 = n947 & n4814 ;
  assign n4816 = n436 ^ n232 ^ 1'b0 ;
  assign n4817 = ( ~n326 & n1174 ) | ( ~n326 & n4816 ) | ( n1174 & n4816 ) ;
  assign n4818 = n4817 ^ n697 ^ n394 ;
  assign n4819 = ( ~n180 & n3064 ) | ( ~n180 & n4818 ) | ( n3064 & n4818 ) ;
  assign n4820 = ~n1291 & n1438 ;
  assign n4821 = n2034 & n4820 ;
  assign n4822 = ( n4376 & n4819 ) | ( n4376 & ~n4821 ) | ( n4819 & ~n4821 ) ;
  assign n4823 = n3643 ^ n3024 ^ n268 ;
  assign n4824 = ( n714 & n1318 ) | ( n714 & ~n4823 ) | ( n1318 & ~n4823 ) ;
  assign n4825 = ~n676 & n1452 ;
  assign n4826 = ~n748 & n4825 ;
  assign n4827 = ~n2953 & n4647 ;
  assign n4828 = n4826 & n4827 ;
  assign n4829 = ( n1139 & ~n3499 ) | ( n1139 & n4828 ) | ( ~n3499 & n4828 ) ;
  assign n4830 = ( n157 & n2367 ) | ( n157 & n3621 ) | ( n2367 & n3621 ) ;
  assign n4831 = n4830 ^ n3070 ^ n1476 ;
  assign n4832 = ( ~n1217 & n3035 ) | ( ~n1217 & n4831 ) | ( n3035 & n4831 ) ;
  assign n4833 = n4829 | n4832 ;
  assign n4834 = n4824 & ~n4833 ;
  assign n4840 = n2973 ^ n409 ^ n291 ;
  assign n4841 = ( n3391 & ~n4779 ) | ( n3391 & n4840 ) | ( ~n4779 & n4840 ) ;
  assign n4836 = n2609 ^ n1657 ^ n1503 ;
  assign n4835 = n1322 ^ n1125 ^ n924 ;
  assign n4837 = n4836 ^ n4835 ^ n751 ;
  assign n4838 = ( n514 & ~n1262 ) | ( n514 & n1662 ) | ( ~n1262 & n1662 ) ;
  assign n4839 = ( ~n1406 & n4837 ) | ( ~n1406 & n4838 ) | ( n4837 & n4838 ) ;
  assign n4842 = n4841 ^ n4839 ^ n2830 ;
  assign n4843 = n841 ^ n769 ^ n655 ;
  assign n4844 = n4843 ^ n3158 ^ x27 ;
  assign n4857 = n4160 ^ n1789 ^ x56 ;
  assign n4852 = n2235 ^ n1866 ^ 1'b0 ;
  assign n4853 = ( n2165 & n2665 ) | ( n2165 & ~n4852 ) | ( n2665 & ~n4852 ) ;
  assign n4854 = n3330 ^ n3066 ^ 1'b0 ;
  assign n4855 = ~n4853 & n4854 ;
  assign n4849 = n4260 ^ n2255 ^ 1'b0 ;
  assign n4850 = n2901 | n4849 ;
  assign n4851 = ( n2481 & n2511 ) | ( n2481 & ~n4850 ) | ( n2511 & ~n4850 ) ;
  assign n4856 = n4855 ^ n4851 ^ x57 ;
  assign n4858 = n4857 ^ n4856 ^ n2735 ;
  assign n4845 = x77 & ~n3096 ;
  assign n4846 = ( n2924 & n3547 ) | ( n2924 & ~n4845 ) | ( n3547 & ~n4845 ) ;
  assign n4847 = n4846 ^ n4603 ^ n595 ;
  assign n4848 = n532 | n4847 ;
  assign n4859 = n4858 ^ n4848 ^ 1'b0 ;
  assign n4868 = ( ~n291 & n355 ) | ( ~n291 & n3721 ) | ( n355 & n3721 ) ;
  assign n4861 = n1022 ^ n500 ^ 1'b0 ;
  assign n4862 = ( ~n1391 & n1416 ) | ( ~n1391 & n4861 ) | ( n1416 & n4861 ) ;
  assign n4860 = n1379 ^ n958 ^ n644 ;
  assign n4863 = n4862 ^ n4860 ^ n2312 ;
  assign n4864 = ~x123 & n1084 ;
  assign n4865 = n4864 ^ n4863 ^ 1'b0 ;
  assign n4866 = n4863 | n4865 ;
  assign n4867 = n881 & n4866 ;
  assign n4869 = n4868 ^ n4867 ^ 1'b0 ;
  assign n4870 = ( x123 & n2275 ) | ( x123 & ~n2778 ) | ( n2275 & ~n2778 ) ;
  assign n4871 = n4870 ^ n4093 ^ n539 ;
  assign n4872 = n4871 ^ n4064 ^ 1'b0 ;
  assign n4873 = n4816 ^ n2644 ^ n1335 ;
  assign n4874 = n3176 & ~n4873 ;
  assign n4879 = n4165 ^ n3095 ^ n974 ;
  assign n4880 = ( x126 & n2021 ) | ( x126 & ~n4879 ) | ( n2021 & ~n4879 ) ;
  assign n4877 = n3135 ^ n549 ^ n131 ;
  assign n4878 = n4877 ^ n3106 ^ n1711 ;
  assign n4875 = n2464 & n4202 ;
  assign n4876 = n1607 & n4875 ;
  assign n4881 = n4880 ^ n4878 ^ n4876 ;
  assign n4887 = n2792 ^ n920 ^ 1'b0 ;
  assign n4888 = n1717 & n4887 ;
  assign n4884 = n1618 ^ n1508 ^ 1'b0 ;
  assign n4885 = ( n1352 & n1452 ) | ( n1352 & n4884 ) | ( n1452 & n4884 ) ;
  assign n4882 = ( n298 & n2037 ) | ( n298 & ~n3009 ) | ( n2037 & ~n3009 ) ;
  assign n4883 = n4882 ^ n1263 ^ x78 ;
  assign n4886 = n4885 ^ n4883 ^ n1635 ;
  assign n4889 = n4888 ^ n4886 ^ n2015 ;
  assign n4899 = n3102 ^ n1530 ^ x12 ;
  assign n4900 = n4899 ^ n1876 ^ x96 ;
  assign n4895 = n2237 ^ n1574 ^ 1'b0 ;
  assign n4896 = n4895 ^ n3162 ^ n2562 ;
  assign n4897 = n1259 & n4896 ;
  assign n4898 = n4897 ^ n2713 ^ 1'b0 ;
  assign n4901 = n4900 ^ n4898 ^ n4870 ;
  assign n4894 = ( x63 & n997 ) | ( x63 & n1265 ) | ( n997 & n1265 ) ;
  assign n4902 = n4901 ^ n4894 ^ n680 ;
  assign n4890 = n1198 & ~n2030 ;
  assign n4891 = ( ~n872 & n4078 ) | ( ~n872 & n4890 ) | ( n4078 & n4890 ) ;
  assign n4892 = ( n931 & ~n1064 ) | ( n931 & n1445 ) | ( ~n1064 & n1445 ) ;
  assign n4893 = ~n4891 & n4892 ;
  assign n4903 = n4902 ^ n4893 ^ 1'b0 ;
  assign n4905 = ( ~n1490 & n2878 ) | ( ~n1490 & n2897 ) | ( n2878 & n2897 ) ;
  assign n4906 = n3287 ^ n2388 ^ 1'b0 ;
  assign n4907 = n4905 | n4906 ;
  assign n4904 = n2305 | n4734 ;
  assign n4908 = n4907 ^ n4904 ^ 1'b0 ;
  assign n4909 = n3543 ^ n1582 ^ n1039 ;
  assign n4910 = ( n743 & ~n1873 ) | ( n743 & n4909 ) | ( ~n1873 & n4909 ) ;
  assign n4911 = ( n2271 & n4908 ) | ( n2271 & ~n4910 ) | ( n4908 & ~n4910 ) ;
  assign n4912 = ~n1927 & n2821 ;
  assign n4913 = ~n2609 & n4912 ;
  assign n4915 = ( n697 & n1584 ) | ( n697 & n2378 ) | ( n1584 & n2378 ) ;
  assign n4914 = ( n358 & ~n603 ) | ( n358 & n3480 ) | ( ~n603 & n3480 ) ;
  assign n4916 = n4915 ^ n4914 ^ 1'b0 ;
  assign n4917 = n4913 | n4916 ;
  assign n4918 = n1270 & n3573 ;
  assign n4919 = n575 & ~n3233 ;
  assign n4920 = n4919 ^ n2393 ^ 1'b0 ;
  assign n4921 = n4920 ^ n2157 ^ n677 ;
  assign n4922 = n2098 | n4921 ;
  assign n4923 = n4918 | n4922 ;
  assign n4924 = ( n1788 & n4644 ) | ( n1788 & n4923 ) | ( n4644 & n4923 ) ;
  assign n4925 = ( n2309 & n3519 ) | ( n2309 & n4924 ) | ( n3519 & n4924 ) ;
  assign n4926 = n4233 ^ n1847 ^ n1045 ;
  assign n4927 = n4926 ^ n4861 ^ n4451 ;
  assign n4933 = n3024 ^ n1292 ^ 1'b0 ;
  assign n4934 = n4898 | n4933 ;
  assign n4928 = n4068 ^ n3281 ^ n1704 ;
  assign n4929 = n978 | n3288 ;
  assign n4930 = n4929 ^ n3537 ^ 1'b0 ;
  assign n4931 = ( n828 & n3507 ) | ( n828 & n4930 ) | ( n3507 & n4930 ) ;
  assign n4932 = ~n4928 & n4931 ;
  assign n4935 = n4934 ^ n4932 ^ 1'b0 ;
  assign n4936 = n3451 ^ n3336 ^ n2257 ;
  assign n4937 = n1923 & ~n4936 ;
  assign n4944 = n583 & n3940 ;
  assign n4945 = n4944 ^ n1716 ^ 1'b0 ;
  assign n4946 = n4945 ^ n2294 ^ n1213 ;
  assign n4947 = ( x48 & n2525 ) | ( x48 & ~n4946 ) | ( n2525 & ~n4946 ) ;
  assign n4939 = n694 ^ n658 ^ n429 ;
  assign n4938 = x28 & n1679 ;
  assign n4940 = n4939 ^ n4938 ^ 1'b0 ;
  assign n4941 = n1392 & n4940 ;
  assign n4942 = ( n1510 & ~n3256 ) | ( n1510 & n4900 ) | ( ~n3256 & n4900 ) ;
  assign n4943 = n4941 & ~n4942 ;
  assign n4948 = n4947 ^ n4943 ^ 1'b0 ;
  assign n4949 = n4948 ^ n4263 ^ n1474 ;
  assign n4950 = n2789 ^ n800 ^ n456 ;
  assign n4951 = ( x22 & ~n2898 ) | ( x22 & n4950 ) | ( ~n2898 & n4950 ) ;
  assign n4952 = ( n187 & ~n951 ) | ( n187 & n1481 ) | ( ~n951 & n1481 ) ;
  assign n4953 = n4952 ^ n3219 ^ n2198 ;
  assign n4954 = ( n1984 & ~n4951 ) | ( n1984 & n4953 ) | ( ~n4951 & n4953 ) ;
  assign n4955 = ( n3209 & n3340 ) | ( n3209 & n4796 ) | ( n3340 & n4796 ) ;
  assign n4961 = ( ~n327 & n1307 ) | ( ~n327 & n4583 ) | ( n1307 & n4583 ) ;
  assign n4959 = n2784 ^ n1717 ^ n1474 ;
  assign n4957 = ~n451 & n3287 ;
  assign n4958 = n4957 ^ n1038 ^ 1'b0 ;
  assign n4960 = n4959 ^ n4958 ^ n2840 ;
  assign n4956 = n584 ^ n428 ^ 1'b0 ;
  assign n4962 = n4961 ^ n4960 ^ n4956 ;
  assign n4964 = ( x36 & n662 ) | ( x36 & n1808 ) | ( n662 & n1808 ) ;
  assign n4965 = ~x28 & n4964 ;
  assign n4963 = n2726 ^ n1695 ^ n1499 ;
  assign n4966 = n4965 ^ n4963 ^ n1232 ;
  assign n4967 = n4966 ^ n3901 ^ n838 ;
  assign n4968 = ( n1940 & ~n3845 ) | ( n1940 & n4967 ) | ( ~n3845 & n4967 ) ;
  assign n4969 = ( n813 & n4439 ) | ( n813 & ~n4721 ) | ( n4439 & ~n4721 ) ;
  assign n4970 = n4129 & ~n4969 ;
  assign n4971 = n1655 & n4970 ;
  assign n4972 = n4495 ^ n2188 ^ 1'b0 ;
  assign n4973 = n4972 ^ n4895 ^ n2373 ;
  assign n4974 = n4952 ^ n3952 ^ n2161 ;
  assign n4975 = ( n2124 & ~n3242 ) | ( n2124 & n4974 ) | ( ~n3242 & n4974 ) ;
  assign n4976 = n1326 ^ x29 ^ 1'b0 ;
  assign n4977 = n530 & n1392 ;
  assign n4978 = n4976 & n4977 ;
  assign n4979 = n4978 ^ n4017 ^ n3875 ;
  assign n4980 = n4975 | n4979 ;
  assign n4981 = n4973 & ~n4980 ;
  assign n4982 = n4586 & ~n4623 ;
  assign n4983 = ( ~n526 & n1438 ) | ( ~n526 & n3213 ) | ( n1438 & n3213 ) ;
  assign n4984 = n4983 ^ n1738 ^ 1'b0 ;
  assign n4985 = ( n1141 & n4398 ) | ( n1141 & n4640 ) | ( n4398 & n4640 ) ;
  assign n4986 = ( n1186 & n2982 ) | ( n1186 & ~n4985 ) | ( n2982 & ~n4985 ) ;
  assign n4987 = n1906 ^ n372 ^ n174 ;
  assign n4988 = n4987 ^ n211 ^ 1'b0 ;
  assign n4989 = n561 & ~n4988 ;
  assign n4990 = n1176 & n4989 ;
  assign n4991 = n3893 ^ n3866 ^ n186 ;
  assign n4992 = n2501 ^ n1115 ^ n438 ;
  assign n4993 = n2489 | n2494 ;
  assign n4994 = ( ~x91 & n959 ) | ( ~x91 & n2291 ) | ( n959 & n2291 ) ;
  assign n4995 = ( ~n770 & n1495 ) | ( ~n770 & n4994 ) | ( n1495 & n4994 ) ;
  assign n4996 = ( n2531 & n3553 ) | ( n2531 & n4995 ) | ( n3553 & n4995 ) ;
  assign n4997 = ( n4992 & n4993 ) | ( n4992 & ~n4996 ) | ( n4993 & ~n4996 ) ;
  assign n4998 = ( n4990 & n4991 ) | ( n4990 & n4997 ) | ( n4991 & n4997 ) ;
  assign n4999 = ( ~n1367 & n4453 ) | ( ~n1367 & n4798 ) | ( n4453 & n4798 ) ;
  assign n5000 = ( n718 & n2283 ) | ( n718 & ~n4999 ) | ( n2283 & ~n4999 ) ;
  assign n5001 = ( ~n2128 & n2565 ) | ( ~n2128 & n2769 ) | ( n2565 & n2769 ) ;
  assign n5002 = ( n304 & n2011 ) | ( n304 & n2443 ) | ( n2011 & n2443 ) ;
  assign n5003 = ( ~n3149 & n5001 ) | ( ~n3149 & n5002 ) | ( n5001 & n5002 ) ;
  assign n5007 = ( n223 & ~n386 ) | ( n223 & n3105 ) | ( ~n386 & n3105 ) ;
  assign n5004 = n2968 ^ n1717 ^ n731 ;
  assign n5005 = ( n3064 & n4302 ) | ( n3064 & n5004 ) | ( n4302 & n5004 ) ;
  assign n5006 = n5005 ^ n1546 ^ n214 ;
  assign n5008 = n5007 ^ n5006 ^ n4853 ;
  assign n5009 = n5008 ^ n1016 ^ 1'b0 ;
  assign n5010 = n1550 & ~n5009 ;
  assign n5011 = ( ~n5000 & n5003 ) | ( ~n5000 & n5010 ) | ( n5003 & n5010 ) ;
  assign n5039 = n4963 ^ n1528 ^ 1'b0 ;
  assign n5012 = n2551 | n4000 ;
  assign n5013 = ( n417 & n1576 ) | ( n417 & n5012 ) | ( n1576 & n5012 ) ;
  assign n5014 = n5013 ^ n736 ^ n502 ;
  assign n5035 = ~n2186 & n3009 ;
  assign n5015 = n3691 ^ n1752 ^ n598 ;
  assign n5019 = n1808 ^ n492 ^ n389 ;
  assign n5016 = n511 & ~n2130 ;
  assign n5017 = ~n502 & n5016 ;
  assign n5018 = ( n250 & n1802 ) | ( n250 & n5017 ) | ( n1802 & n5017 ) ;
  assign n5020 = n5019 ^ n5018 ^ n2851 ;
  assign n5021 = n4882 | n5020 ;
  assign n5022 = n5021 ^ n2384 ^ 1'b0 ;
  assign n5023 = ( ~n3609 & n5015 ) | ( ~n3609 & n5022 ) | ( n5015 & n5022 ) ;
  assign n5024 = ( x95 & n1889 ) | ( x95 & n2128 ) | ( n1889 & n2128 ) ;
  assign n5025 = n505 | n1738 ;
  assign n5026 = n607 & ~n5025 ;
  assign n5027 = ( x2 & n936 ) | ( x2 & ~n4407 ) | ( n936 & ~n4407 ) ;
  assign n5028 = ( n3806 & n5026 ) | ( n3806 & n5027 ) | ( n5026 & n5027 ) ;
  assign n5029 = ( n4424 & n5024 ) | ( n4424 & n5028 ) | ( n5024 & n5028 ) ;
  assign n5030 = n3045 ^ n2171 ^ n150 ;
  assign n5031 = ( n742 & n2671 ) | ( n742 & ~n5030 ) | ( n2671 & ~n5030 ) ;
  assign n5032 = n5029 | n5031 ;
  assign n5033 = n5032 ^ n4001 ^ 1'b0 ;
  assign n5034 = ( n2395 & n5023 ) | ( n2395 & ~n5033 ) | ( n5023 & ~n5033 ) ;
  assign n5036 = n5035 ^ n5034 ^ 1'b0 ;
  assign n5037 = n5014 & n5036 ;
  assign n5038 = n5037 ^ n2090 ^ 1'b0 ;
  assign n5040 = n5039 ^ n5038 ^ n4482 ;
  assign n5041 = ( n3216 & n4757 ) | ( n3216 & n4967 ) | ( n4757 & n4967 ) ;
  assign n5042 = n1124 ^ n814 ^ 1'b0 ;
  assign n5046 = x46 & x102 ;
  assign n5047 = n5046 ^ n1702 ^ 1'b0 ;
  assign n5048 = ( n559 & n3420 ) | ( n559 & n5047 ) | ( n3420 & n5047 ) ;
  assign n5045 = n4403 ^ n1759 ^ n990 ;
  assign n5049 = n5048 ^ n5045 ^ n1549 ;
  assign n5043 = n4546 ^ n1782 ^ n1703 ;
  assign n5044 = n5043 ^ n4058 ^ n2118 ;
  assign n5050 = n5049 ^ n5044 ^ n4056 ;
  assign n5051 = n5042 & n5050 ;
  assign n5053 = ( ~n487 & n3424 ) | ( ~n487 & n3943 ) | ( n3424 & n3943 ) ;
  assign n5052 = n4204 ^ n610 ^ 1'b0 ;
  assign n5054 = n5053 ^ n5052 ^ 1'b0 ;
  assign n5055 = n1039 | n5054 ;
  assign n5060 = ( x30 & ~n3185 ) | ( x30 & n3572 ) | ( ~n3185 & n3572 ) ;
  assign n5061 = n2818 | n5060 ;
  assign n5062 = ( n1534 & ~n2158 ) | ( n1534 & n5061 ) | ( ~n2158 & n5061 ) ;
  assign n5063 = ( n131 & n4840 ) | ( n131 & ~n5062 ) | ( n4840 & ~n5062 ) ;
  assign n5064 = n5063 ^ n2910 ^ n869 ;
  assign n5056 = n1433 ^ n672 ^ 1'b0 ;
  assign n5057 = n1740 & ~n5056 ;
  assign n5058 = n4952 & n5057 ;
  assign n5059 = n1179 | n5058 ;
  assign n5065 = n5064 ^ n5059 ^ 1'b0 ;
  assign n5066 = ( n1072 & ~n1451 ) | ( n1072 & n2222 ) | ( ~n1451 & n2222 ) ;
  assign n5067 = n3789 ^ n2391 ^ 1'b0 ;
  assign n5068 = ( x93 & n1151 ) | ( x93 & ~n2119 ) | ( n1151 & ~n2119 ) ;
  assign n5069 = ( n956 & n1170 ) | ( n956 & n2902 ) | ( n1170 & n2902 ) ;
  assign n5070 = ( x85 & n5068 ) | ( x85 & n5069 ) | ( n5068 & n5069 ) ;
  assign n5071 = n5070 ^ n4516 ^ n3628 ;
  assign n5076 = n4793 ^ n2976 ^ 1'b0 ;
  assign n5077 = ( n498 & ~n2082 ) | ( n498 & n5076 ) | ( ~n2082 & n5076 ) ;
  assign n5072 = n3222 ^ n2581 ^ n1690 ;
  assign n5073 = ~n320 & n5072 ;
  assign n5074 = ( n862 & n3182 ) | ( n862 & n5073 ) | ( n3182 & n5073 ) ;
  assign n5075 = ( n856 & n3294 ) | ( n856 & n5074 ) | ( n3294 & n5074 ) ;
  assign n5078 = n5077 ^ n5075 ^ 1'b0 ;
  assign n5079 = n1978 ^ n1101 ^ 1'b0 ;
  assign n5080 = n3355 & ~n5079 ;
  assign n5081 = ( n2438 & ~n4070 ) | ( n2438 & n5080 ) | ( ~n4070 & n5080 ) ;
  assign n5082 = n3023 ^ n2830 ^ n1259 ;
  assign n5083 = ( n4174 & n4502 ) | ( n4174 & ~n5082 ) | ( n4502 & ~n5082 ) ;
  assign n5084 = ~n1784 & n5083 ;
  assign n5085 = ~n2940 & n5084 ;
  assign n5088 = ( ~x22 & n778 ) | ( ~x22 & n3198 ) | ( n778 & n3198 ) ;
  assign n5089 = n1440 | n4861 ;
  assign n5090 = n5088 & ~n5089 ;
  assign n5091 = n5090 ^ n3624 ^ n1680 ;
  assign n5086 = n890 ^ x58 ^ 1'b0 ;
  assign n5087 = n1705 | n5086 ;
  assign n5092 = n5091 ^ n5087 ^ n2780 ;
  assign n5093 = n5092 ^ n4705 ^ n2455 ;
  assign n5094 = n2752 & ~n3600 ;
  assign n5095 = n5094 ^ n612 ^ 1'b0 ;
  assign n5096 = ( n268 & n670 ) | ( n268 & n955 ) | ( n670 & n955 ) ;
  assign n5097 = n3081 | n5096 ;
  assign n5098 = n5097 ^ n3053 ^ n1252 ;
  assign n5099 = ~n290 & n1493 ;
  assign n5100 = ~n5098 & n5099 ;
  assign n5101 = n5100 ^ n1747 ^ n1295 ;
  assign n5110 = n1187 & ~n3217 ;
  assign n5111 = n5110 ^ n1403 ^ 1'b0 ;
  assign n5109 = n2198 ^ n1561 ^ 1'b0 ;
  assign n5112 = n5111 ^ n5109 ^ n133 ;
  assign n5102 = n4277 ^ n197 ^ 1'b0 ;
  assign n5103 = n4816 & n5102 ;
  assign n5104 = ( ~n644 & n760 ) | ( ~n644 & n5103 ) | ( n760 & n5103 ) ;
  assign n5105 = n5104 ^ n539 ^ 1'b0 ;
  assign n5106 = ~n3882 & n5105 ;
  assign n5107 = ( n912 & ~n1779 ) | ( n912 & n5106 ) | ( ~n1779 & n5106 ) ;
  assign n5108 = n5107 ^ n841 ^ x46 ;
  assign n5113 = n5112 ^ n5108 ^ n1457 ;
  assign n5115 = n2704 ^ n2174 ^ x30 ;
  assign n5114 = n1102 ^ n201 ^ 1'b0 ;
  assign n5116 = n5115 ^ n5114 ^ 1'b0 ;
  assign n5117 = n5113 & n5116 ;
  assign n5118 = n1098 ^ n569 ^ n165 ;
  assign n5119 = n5118 ^ n1498 ^ 1'b0 ;
  assign n5120 = n2568 & ~n5119 ;
  assign n5121 = n3220 ^ n418 ^ 1'b0 ;
  assign n5122 = n5121 ^ n1923 ^ n624 ;
  assign n5123 = n2575 ^ n2051 ^ n1879 ;
  assign n5124 = n4606 & ~n5123 ;
  assign n5125 = n5124 ^ n3785 ^ 1'b0 ;
  assign n5126 = n1336 & n3762 ;
  assign n5127 = ( n3880 & ~n5125 ) | ( n3880 & n5126 ) | ( ~n5125 & n5126 ) ;
  assign n5128 = n3203 ^ n1287 ^ 1'b0 ;
  assign n5129 = n2415 & ~n5128 ;
  assign n5130 = ( n1995 & ~n3878 ) | ( n1995 & n5129 ) | ( ~n3878 & n5129 ) ;
  assign n5131 = ( n2157 & n2636 ) | ( n2157 & n4803 ) | ( n2636 & n4803 ) ;
  assign n5132 = ( n846 & n1909 ) | ( n846 & ~n5131 ) | ( n1909 & ~n5131 ) ;
  assign n5133 = n2389 | n5132 ;
  assign n5134 = n5133 ^ n495 ^ 1'b0 ;
  assign n5135 = n5134 ^ n890 ^ 1'b0 ;
  assign n5144 = n321 & ~n964 ;
  assign n5145 = n5144 ^ n4684 ^ 1'b0 ;
  assign n5136 = n3133 ^ n2982 ^ 1'b0 ;
  assign n5137 = n1150 | n5136 ;
  assign n5138 = ( n251 & n2465 ) | ( n251 & ~n3746 ) | ( n2465 & ~n3746 ) ;
  assign n5139 = n5138 ^ n3572 ^ 1'b0 ;
  assign n5140 = n5137 | n5139 ;
  assign n5141 = n1702 ^ n1354 ^ n997 ;
  assign n5142 = ( n4179 & ~n5140 ) | ( n4179 & n5141 ) | ( ~n5140 & n5141 ) ;
  assign n5143 = ~n2371 & n5142 ;
  assign n5146 = n5145 ^ n5143 ^ 1'b0 ;
  assign n5147 = n5146 ^ n4439 ^ 1'b0 ;
  assign n5148 = ( ~n1105 & n1491 ) | ( ~n1105 & n2529 ) | ( n1491 & n2529 ) ;
  assign n5149 = n5148 ^ n2164 ^ 1'b0 ;
  assign n5150 = n4463 | n5149 ;
  assign n5151 = ( ~n2241 & n3502 ) | ( ~n2241 & n5150 ) | ( n3502 & n5150 ) ;
  assign n5152 = ~n519 & n1249 ;
  assign n5153 = n2367 | n3106 ;
  assign n5154 = ( n4748 & n4951 ) | ( n4748 & ~n5153 ) | ( n4951 & ~n5153 ) ;
  assign n5155 = n5154 ^ n4860 ^ n4070 ;
  assign n5156 = n722 | n1071 ;
  assign n5157 = n5156 ^ x86 ^ 1'b0 ;
  assign n5158 = ( ~n976 & n3610 ) | ( ~n976 & n5157 ) | ( n3610 & n5157 ) ;
  assign n5159 = n2317 ^ n1306 ^ n670 ;
  assign n5160 = n5159 ^ n193 ^ 1'b0 ;
  assign n5162 = n3108 & n3251 ;
  assign n5161 = ( x53 & ~n961 ) | ( x53 & n2724 ) | ( ~n961 & n2724 ) ;
  assign n5163 = n5162 ^ n5161 ^ n569 ;
  assign n5164 = ( ~n1101 & n5160 ) | ( ~n1101 & n5163 ) | ( n5160 & n5163 ) ;
  assign n5166 = x70 & n2775 ;
  assign n5165 = n2445 ^ n1463 ^ 1'b0 ;
  assign n5167 = n5166 ^ n5165 ^ n4731 ;
  assign n5168 = n2573 | n5167 ;
  assign n5170 = ( n2455 & n3350 ) | ( n2455 & ~n3886 ) | ( n3350 & ~n3886 ) ;
  assign n5171 = ( n5030 & n5056 ) | ( n5030 & n5170 ) | ( n5056 & n5170 ) ;
  assign n5169 = n1375 & n1850 ;
  assign n5172 = n5171 ^ n5169 ^ 1'b0 ;
  assign n5173 = ( ~n140 & n1101 ) | ( ~n140 & n2186 ) | ( n1101 & n2186 ) ;
  assign n5174 = n2579 ^ n1251 ^ x87 ;
  assign n5175 = ( ~n456 & n639 ) | ( ~n456 & n716 ) | ( n639 & n716 ) ;
  assign n5176 = ( n3831 & n5174 ) | ( n3831 & ~n5175 ) | ( n5174 & ~n5175 ) ;
  assign n5177 = n3317 | n4346 ;
  assign n5178 = n841 & ~n5177 ;
  assign n5179 = ( ~n5173 & n5176 ) | ( ~n5173 & n5178 ) | ( n5176 & n5178 ) ;
  assign n5183 = ( n1028 & n1172 ) | ( n1028 & n2480 ) | ( n1172 & n2480 ) ;
  assign n5184 = n5183 ^ n2374 ^ n1456 ;
  assign n5180 = n1152 & ~n3622 ;
  assign n5181 = ~n1008 & n5180 ;
  assign n5182 = n5181 ^ n3374 ^ n1940 ;
  assign n5185 = n5184 ^ n5182 ^ 1'b0 ;
  assign n5186 = ( ~n647 & n2941 ) | ( ~n647 & n5185 ) | ( n2941 & n5185 ) ;
  assign n5187 = ( ~x61 & n1734 ) | ( ~x61 & n5186 ) | ( n1734 & n5186 ) ;
  assign n5190 = ( n268 & n486 ) | ( n268 & n2910 ) | ( n486 & n2910 ) ;
  assign n5188 = ~n1691 & n3774 ;
  assign n5189 = n5188 ^ n595 ^ 1'b0 ;
  assign n5191 = n5190 ^ n5189 ^ n526 ;
  assign n5192 = ( n852 & n1165 ) | ( n852 & n1792 ) | ( n1165 & n1792 ) ;
  assign n5193 = x61 & n5192 ;
  assign n5194 = n2701 ^ n2507 ^ n2281 ;
  assign n5195 = n953 & ~n5194 ;
  assign n5196 = n5195 ^ n162 ^ 1'b0 ;
  assign n5197 = n5196 ^ n3948 ^ 1'b0 ;
  assign n5199 = n3451 ^ n1069 ^ x30 ;
  assign n5198 = n717 & n2676 ;
  assign n5200 = n5199 ^ n5198 ^ 1'b0 ;
  assign n5201 = n5200 ^ n3262 ^ 1'b0 ;
  assign n5218 = n193 & n1807 ;
  assign n5216 = n4168 ^ n2010 ^ 1'b0 ;
  assign n5215 = n4495 ^ n1990 ^ 1'b0 ;
  assign n5217 = n5216 ^ n5215 ^ 1'b0 ;
  assign n5204 = n647 ^ n343 ^ 1'b0 ;
  assign n5205 = n1225 & ~n5204 ;
  assign n5206 = ~n2262 & n5205 ;
  assign n5207 = n3579 ^ n1923 ^ n1607 ;
  assign n5208 = ( ~x0 & n1987 ) | ( ~x0 & n4108 ) | ( n1987 & n4108 ) ;
  assign n5209 = n516 ^ n472 ^ n285 ;
  assign n5210 = n5209 ^ n3896 ^ n1149 ;
  assign n5211 = n5210 ^ n4763 ^ n2885 ;
  assign n5212 = ( n181 & n5208 ) | ( n181 & n5211 ) | ( n5208 & n5211 ) ;
  assign n5213 = ( n5206 & n5207 ) | ( n5206 & n5212 ) | ( n5207 & n5212 ) ;
  assign n5214 = n5213 ^ n3843 ^ n381 ;
  assign n5219 = n5218 ^ n5217 ^ n5214 ;
  assign n5202 = ~n1457 & n3096 ;
  assign n5203 = n426 & n5202 ;
  assign n5220 = n5219 ^ n5203 ^ 1'b0 ;
  assign n5224 = ( n425 & ~n1939 ) | ( n425 & n4294 ) | ( ~n1939 & n4294 ) ;
  assign n5221 = ( n840 & ~n1985 ) | ( n840 & n2421 ) | ( ~n1985 & n2421 ) ;
  assign n5222 = n863 & n5221 ;
  assign n5223 = ~n3692 & n5222 ;
  assign n5225 = n5224 ^ n5223 ^ n1101 ;
  assign n5226 = ( n738 & n860 ) | ( n738 & n4240 ) | ( n860 & n4240 ) ;
  assign n5227 = n3684 | n5226 ;
  assign n5229 = n3964 ^ n2601 ^ n949 ;
  assign n5230 = ( ~n1420 & n2235 ) | ( ~n1420 & n5229 ) | ( n2235 & n5229 ) ;
  assign n5231 = n5230 ^ n4728 ^ n2995 ;
  assign n5228 = n2075 & ~n2729 ;
  assign n5232 = n5231 ^ n5228 ^ 1'b0 ;
  assign n5233 = n411 | n3984 ;
  assign n5234 = n1708 | n5233 ;
  assign n5235 = n5234 ^ n3337 ^ n392 ;
  assign n5236 = n4148 & ~n5235 ;
  assign n5237 = n5232 & n5236 ;
  assign n5238 = n5237 ^ n2504 ^ 1'b0 ;
  assign n5239 = n5227 & ~n5238 ;
  assign n5240 = n2352 ^ n636 ^ 1'b0 ;
  assign n5241 = n4201 & n5240 ;
  assign n5242 = ( n1072 & n1268 ) | ( n1072 & ~n5241 ) | ( n1268 & ~n5241 ) ;
  assign n5243 = ( ~n1612 & n2663 ) | ( ~n1612 & n5242 ) | ( n2663 & n5242 ) ;
  assign n5244 = ( ~n940 & n1493 ) | ( ~n940 & n2764 ) | ( n1493 & n2764 ) ;
  assign n5245 = n1296 ^ n811 ^ 1'b0 ;
  assign n5246 = n2079 & ~n5245 ;
  assign n5247 = ( ~n1006 & n2960 ) | ( ~n1006 & n5246 ) | ( n2960 & n5246 ) ;
  assign n5248 = n5247 ^ n1214 ^ n247 ;
  assign n5249 = n3934 | n5248 ;
  assign n5250 = n5244 | n5249 ;
  assign n5254 = n3308 ^ n960 ^ 1'b0 ;
  assign n5255 = x92 & ~n5254 ;
  assign n5256 = ~n1209 & n5255 ;
  assign n5251 = ( n319 & n1585 ) | ( n319 & ~n3327 ) | ( n1585 & ~n3327 ) ;
  assign n5252 = x105 & ~n5251 ;
  assign n5253 = n5252 ^ n2722 ^ 1'b0 ;
  assign n5257 = n5256 ^ n5253 ^ n2979 ;
  assign n5259 = n1597 ^ n908 ^ 1'b0 ;
  assign n5258 = x86 & ~n1440 ;
  assign n5260 = n5259 ^ n5258 ^ 1'b0 ;
  assign n5261 = ~n5031 & n5260 ;
  assign n5262 = ( ~n5250 & n5257 ) | ( ~n5250 & n5261 ) | ( n5257 & n5261 ) ;
  assign n5263 = n3757 ^ n2216 ^ n258 ;
  assign n5264 = n3883 ^ n1677 ^ n216 ;
  assign n5265 = ( n4514 & n5141 ) | ( n4514 & ~n5264 ) | ( n5141 & ~n5264 ) ;
  assign n5266 = n3532 ^ n2182 ^ 1'b0 ;
  assign n5267 = n5266 ^ n3666 ^ 1'b0 ;
  assign n5268 = n5265 & ~n5267 ;
  assign n5269 = ( n305 & n1037 ) | ( n305 & ~n1747 ) | ( n1037 & ~n1747 ) ;
  assign n5270 = n2440 & ~n2606 ;
  assign n5271 = ( n4174 & ~n5269 ) | ( n4174 & n5270 ) | ( ~n5269 & n5270 ) ;
  assign n5272 = ( x102 & n159 ) | ( x102 & n1265 ) | ( n159 & n1265 ) ;
  assign n5273 = n5272 ^ n1822 ^ n1496 ;
  assign n5274 = ( n3403 & ~n3409 ) | ( n3403 & n5273 ) | ( ~n3409 & n5273 ) ;
  assign n5275 = n988 | n5274 ;
  assign n5276 = n5275 ^ n5231 ^ 1'b0 ;
  assign n5277 = n215 & ~n5276 ;
  assign n5278 = ( n794 & n3798 ) | ( n794 & n5277 ) | ( n3798 & n5277 ) ;
  assign n5279 = ( n299 & ~n1196 ) | ( n299 & n1907 ) | ( ~n1196 & n1907 ) ;
  assign n5280 = n5279 ^ n576 ^ n501 ;
  assign n5281 = ( ~n136 & n505 ) | ( ~n136 & n1004 ) | ( n505 & n1004 ) ;
  assign n5282 = ( ~x127 & n145 ) | ( ~x127 & n231 ) | ( n145 & n231 ) ;
  assign n5283 = n5282 ^ n1870 ^ x100 ;
  assign n5284 = ( n3676 & n5281 ) | ( n3676 & ~n5283 ) | ( n5281 & ~n5283 ) ;
  assign n5285 = ( n139 & n977 ) | ( n139 & n2201 ) | ( n977 & n2201 ) ;
  assign n5286 = ( n5280 & ~n5284 ) | ( n5280 & n5285 ) | ( ~n5284 & n5285 ) ;
  assign n5287 = n2323 ^ n470 ^ 1'b0 ;
  assign n5288 = ( n523 & n2825 ) | ( n523 & n5287 ) | ( n2825 & n5287 ) ;
  assign n5289 = n5288 ^ n2551 ^ n2344 ;
  assign n5290 = n5286 | n5289 ;
  assign n5292 = x39 & ~n294 ;
  assign n5293 = ( x88 & ~n469 ) | ( x88 & n5292 ) | ( ~n469 & n5292 ) ;
  assign n5291 = n2418 ^ n2224 ^ n1821 ;
  assign n5294 = n5293 ^ n5291 ^ n1110 ;
  assign n5295 = ( n1305 & n1727 ) | ( n1305 & n2032 ) | ( n1727 & n2032 ) ;
  assign n5296 = n2396 ^ n1712 ^ 1'b0 ;
  assign n5297 = ~n3797 & n5296 ;
  assign n5298 = n5295 & n5297 ;
  assign n5301 = n4809 ^ n873 ^ 1'b0 ;
  assign n5299 = ( n1231 & ~n2016 ) | ( n1231 & n2395 ) | ( ~n2016 & n2395 ) ;
  assign n5300 = n5299 ^ n3785 ^ n374 ;
  assign n5302 = n5301 ^ n5300 ^ n493 ;
  assign n5303 = n5302 ^ n4729 ^ n3459 ;
  assign n5304 = ( n601 & ~n5298 ) | ( n601 & n5303 ) | ( ~n5298 & n5303 ) ;
  assign n5319 = ( n736 & n1668 ) | ( n736 & n3200 ) | ( n1668 & n3200 ) ;
  assign n5320 = ( n1907 & n3590 ) | ( n1907 & ~n5319 ) | ( n3590 & ~n5319 ) ;
  assign n5316 = ( n129 & ~n621 ) | ( n129 & n4181 ) | ( ~n621 & n4181 ) ;
  assign n5317 = n5316 ^ n3276 ^ n2013 ;
  assign n5318 = n5317 ^ n3304 ^ n2469 ;
  assign n5306 = ( n765 & n1643 ) | ( n765 & n3069 ) | ( n1643 & n3069 ) ;
  assign n5305 = n2021 ^ n710 ^ x78 ;
  assign n5307 = n5306 ^ n5305 ^ n3230 ;
  assign n5308 = n5307 ^ n3344 ^ n2251 ;
  assign n5309 = ( n174 & ~n273 ) | ( n174 & n1691 ) | ( ~n273 & n1691 ) ;
  assign n5310 = n5309 ^ n2521 ^ n1084 ;
  assign n5311 = ( ~n2033 & n2186 ) | ( ~n2033 & n5310 ) | ( n2186 & n5310 ) ;
  assign n5312 = n2994 ^ n2143 ^ n669 ;
  assign n5313 = ( ~n1693 & n5311 ) | ( ~n1693 & n5312 ) | ( n5311 & n5312 ) ;
  assign n5314 = ( n3082 & n5308 ) | ( n3082 & n5313 ) | ( n5308 & n5313 ) ;
  assign n5315 = ( n820 & n4285 ) | ( n820 & n5314 ) | ( n4285 & n5314 ) ;
  assign n5321 = n5320 ^ n5318 ^ n5315 ;
  assign n5322 = ( n830 & n2816 ) | ( n830 & n3900 ) | ( n2816 & n3900 ) ;
  assign n5332 = n3579 ^ n730 ^ n360 ;
  assign n5333 = ( n2247 & ~n2821 ) | ( n2247 & n5332 ) | ( ~n2821 & n5332 ) ;
  assign n5328 = n273 | n1168 ;
  assign n5323 = n4850 ^ n2082 ^ n889 ;
  assign n5324 = ~n130 & n1643 ;
  assign n5325 = ~n1717 & n5324 ;
  assign n5326 = ( n860 & n5323 ) | ( n860 & ~n5325 ) | ( n5323 & ~n5325 ) ;
  assign n5327 = ~n3200 & n5326 ;
  assign n5329 = n5328 ^ n5327 ^ 1'b0 ;
  assign n5330 = ~n1787 & n5329 ;
  assign n5331 = n5330 ^ n5206 ^ 1'b0 ;
  assign n5334 = n5333 ^ n5331 ^ n2806 ;
  assign n5335 = n2046 ^ n912 ^ n529 ;
  assign n5336 = n3756 ^ n3297 ^ n985 ;
  assign n5337 = ( n1618 & ~n5335 ) | ( n1618 & n5336 ) | ( ~n5335 & n5336 ) ;
  assign n5338 = n5337 ^ n4610 ^ n1416 ;
  assign n5339 = n5015 ^ n2341 ^ 1'b0 ;
  assign n5340 = n2533 ^ n1697 ^ n1390 ;
  assign n5341 = n5340 ^ n990 ^ 1'b0 ;
  assign n5342 = n5341 ^ n4495 ^ 1'b0 ;
  assign n5343 = n3056 ^ n2770 ^ n1369 ;
  assign n5344 = ( n315 & n4231 ) | ( n315 & ~n4740 ) | ( n4231 & ~n4740 ) ;
  assign n5345 = n5344 ^ n5109 ^ n4737 ;
  assign n5346 = n828 ^ n577 ^ n287 ;
  assign n5347 = ( ~n3589 & n4519 ) | ( ~n3589 & n5346 ) | ( n4519 & n5346 ) ;
  assign n5348 = ( x73 & n699 ) | ( x73 & n2397 ) | ( n699 & n2397 ) ;
  assign n5349 = ( n2303 & ~n2973 ) | ( n2303 & n5348 ) | ( ~n2973 & n5348 ) ;
  assign n5350 = n1679 & n3425 ;
  assign n5351 = n5350 ^ n3539 ^ n1268 ;
  assign n5355 = n1612 ^ n1550 ^ n1080 ;
  assign n5352 = n3703 ^ n2589 ^ n2480 ;
  assign n5353 = n5352 ^ n4748 ^ 1'b0 ;
  assign n5354 = n566 | n5353 ;
  assign n5356 = n5355 ^ n5354 ^ x70 ;
  assign n5357 = ( n2233 & n5351 ) | ( n2233 & n5356 ) | ( n5351 & n5356 ) ;
  assign n5373 = n5252 ^ n1196 ^ n388 ;
  assign n5371 = ~n287 & n1632 ;
  assign n5372 = n2414 & n5371 ;
  assign n5374 = n5373 ^ n5372 ^ 1'b0 ;
  assign n5375 = n5162 | n5374 ;
  assign n5370 = n3607 ^ n3340 ^ n2320 ;
  assign n5376 = n5375 ^ n5370 ^ 1'b0 ;
  assign n5358 = ( n1717 & ~n4092 ) | ( n1717 & n4870 ) | ( ~n4092 & n4870 ) ;
  assign n5365 = ( ~n213 & n2752 ) | ( ~n213 & n3311 ) | ( n2752 & n3311 ) ;
  assign n5366 = ( n2989 & ~n3428 ) | ( n2989 & n5365 ) | ( ~n3428 & n5365 ) ;
  assign n5363 = n3536 ^ n226 ^ 1'b0 ;
  assign n5364 = n1526 | n5363 ;
  assign n5367 = n5366 ^ n5364 ^ n4959 ;
  assign n5360 = n1920 ^ n1143 ^ n1054 ;
  assign n5361 = n5360 ^ n2436 ^ n2373 ;
  assign n5359 = ( n568 & n1466 ) | ( n568 & ~n2549 ) | ( n1466 & ~n2549 ) ;
  assign n5362 = n5361 ^ n5359 ^ n1403 ;
  assign n5368 = n5367 ^ n5362 ^ n4041 ;
  assign n5369 = n5358 & ~n5368 ;
  assign n5377 = n5376 ^ n5369 ^ 1'b0 ;
  assign n5392 = n5306 ^ n3877 ^ 1'b0 ;
  assign n5386 = ( n1569 & ~n2849 ) | ( n1569 & n3377 ) | ( ~n2849 & n3377 ) ;
  assign n5387 = n247 & ~n1083 ;
  assign n5388 = n3984 & n5387 ;
  assign n5389 = ( ~n1249 & n5386 ) | ( ~n1249 & n5388 ) | ( n5386 & n5388 ) ;
  assign n5385 = n862 & ~n4232 ;
  assign n5390 = n5389 ^ n5385 ^ 1'b0 ;
  assign n5391 = ( n1822 & n2730 ) | ( n1822 & ~n5390 ) | ( n2730 & ~n5390 ) ;
  assign n5378 = n327 | n357 ;
  assign n5379 = n5378 ^ n1334 ^ 1'b0 ;
  assign n5380 = ( n2799 & n3690 ) | ( n2799 & n5379 ) | ( n3690 & n5379 ) ;
  assign n5381 = n5380 ^ n4645 ^ n916 ;
  assign n5382 = ( n238 & ~n1362 ) | ( n238 & n4235 ) | ( ~n1362 & n4235 ) ;
  assign n5383 = n5382 ^ n1025 ^ 1'b0 ;
  assign n5384 = ( n2379 & ~n5381 ) | ( n2379 & n5383 ) | ( ~n5381 & n5383 ) ;
  assign n5393 = n5392 ^ n5391 ^ n5384 ;
  assign n5394 = ( ~n350 & n477 ) | ( ~n350 & n3865 ) | ( n477 & n3865 ) ;
  assign n5395 = n5093 & ~n5394 ;
  assign n5396 = n2886 & n5395 ;
  assign n5397 = n2780 ^ n2655 ^ n374 ;
  assign n5398 = n2989 | n5397 ;
  assign n5400 = n4417 ^ n2375 ^ n1573 ;
  assign n5399 = n2615 ^ n1848 ^ 1'b0 ;
  assign n5401 = n5400 ^ n5399 ^ x124 ;
  assign n5402 = n4858 ^ n4781 ^ n159 ;
  assign n5403 = n1407 & ~n1946 ;
  assign n5404 = n430 & n5403 ;
  assign n5405 = ~n5402 & n5404 ;
  assign n5407 = ( n917 & n1110 ) | ( n917 & ~n1401 ) | ( n1110 & ~n1401 ) ;
  assign n5408 = n5407 ^ n163 ^ 1'b0 ;
  assign n5406 = n4676 ^ n2217 ^ 1'b0 ;
  assign n5409 = n5408 ^ n5406 ^ n5220 ;
  assign n5410 = n4303 ^ n235 ^ 1'b0 ;
  assign n5411 = n5410 ^ n2292 ^ n2145 ;
  assign n5413 = n246 | n426 ;
  assign n5414 = ~n1075 & n2542 ;
  assign n5415 = ~n5413 & n5414 ;
  assign n5412 = ( n334 & ~n1020 ) | ( n334 & n1874 ) | ( ~n1020 & n1874 ) ;
  assign n5416 = n5415 ^ n5412 ^ n2510 ;
  assign n5417 = ~n213 & n2829 ;
  assign n5418 = n5416 & ~n5417 ;
  assign n5419 = n5418 ^ n2277 ^ 1'b0 ;
  assign n5420 = n670 & n5419 ;
  assign n5421 = n5420 ^ n423 ^ 1'b0 ;
  assign n5422 = ( n914 & n5127 ) | ( n914 & n5421 ) | ( n5127 & n5421 ) ;
  assign n5423 = n4850 ^ n2674 ^ n640 ;
  assign n5424 = ( n521 & n674 ) | ( n521 & n5423 ) | ( n674 & n5423 ) ;
  assign n5425 = n3502 | n5424 ;
  assign n5426 = ( n231 & n2039 ) | ( n231 & ~n3603 ) | ( n2039 & ~n3603 ) ;
  assign n5427 = n5426 ^ n985 ^ x90 ;
  assign n5431 = n1744 ^ n1205 ^ n354 ;
  assign n5432 = ( n2994 & n3458 ) | ( n2994 & ~n5431 ) | ( n3458 & ~n5431 ) ;
  assign n5429 = ~n2364 & n3040 ;
  assign n5428 = n4619 ^ n4455 ^ 1'b0 ;
  assign n5430 = n5429 ^ n5428 ^ n1335 ;
  assign n5433 = n5432 ^ n5430 ^ 1'b0 ;
  assign n5434 = n5427 & ~n5433 ;
  assign n5438 = ~n486 & n4513 ;
  assign n5439 = n5438 ^ n5299 ^ 1'b0 ;
  assign n5440 = n5439 ^ n2127 ^ 1'b0 ;
  assign n5435 = n3616 ^ n3287 ^ n2587 ;
  assign n5436 = n5435 ^ n2872 ^ 1'b0 ;
  assign n5437 = ( ~n1369 & n2619 ) | ( ~n1369 & n5436 ) | ( n2619 & n5436 ) ;
  assign n5441 = n5440 ^ n5437 ^ 1'b0 ;
  assign n5445 = n3212 ^ n1864 ^ n1594 ;
  assign n5446 = n5445 ^ n1009 ^ n995 ;
  assign n5443 = n1005 ^ n750 ^ x5 ;
  assign n5444 = n5443 ^ n2924 ^ n2351 ;
  assign n5447 = n5446 ^ n5444 ^ x47 ;
  assign n5442 = n1713 | n1939 ;
  assign n5448 = n5447 ^ n5442 ^ n2754 ;
  assign n5449 = n5448 ^ n3624 ^ n1392 ;
  assign n5450 = n2186 ^ n889 ^ x99 ;
  assign n5451 = n4879 ^ n3988 ^ n3155 ;
  assign n5452 = n4253 ^ n2525 ^ n2112 ;
  assign n5453 = ( n1365 & n3423 ) | ( n1365 & ~n5452 ) | ( n3423 & ~n5452 ) ;
  assign n5454 = n5453 ^ n3334 ^ n981 ;
  assign n5455 = n5454 ^ n3418 ^ n2058 ;
  assign n5456 = ( n5450 & ~n5451 ) | ( n5450 & n5455 ) | ( ~n5451 & n5455 ) ;
  assign n5457 = ( n334 & n2784 ) | ( n334 & ~n3712 ) | ( n2784 & ~n3712 ) ;
  assign n5458 = ( ~n327 & n347 ) | ( ~n327 & n2022 ) | ( n347 & n2022 ) ;
  assign n5459 = n5458 ^ n3404 ^ n918 ;
  assign n5460 = n2705 ^ n1924 ^ n1680 ;
  assign n5461 = ( n391 & n3428 ) | ( n391 & n5460 ) | ( n3428 & n5460 ) ;
  assign n5462 = ( n1704 & n2360 ) | ( n1704 & ~n4880 ) | ( n2360 & ~n4880 ) ;
  assign n5463 = n5462 ^ n3258 ^ 1'b0 ;
  assign n5464 = n2061 | n5463 ;
  assign n5465 = n4641 ^ n1281 ^ 1'b0 ;
  assign n5466 = ( ~n1395 & n4844 ) | ( ~n1395 & n5465 ) | ( n4844 & n5465 ) ;
  assign n5467 = ( ~n1412 & n2661 ) | ( ~n1412 & n4627 ) | ( n2661 & n4627 ) ;
  assign n5468 = n3897 ^ n1715 ^ n439 ;
  assign n5469 = ( ~n257 & n4260 ) | ( ~n257 & n5468 ) | ( n4260 & n5468 ) ;
  assign n5470 = n5467 & ~n5469 ;
  assign n5471 = n2530 ^ n1781 ^ n521 ;
  assign n5472 = n2762 ^ n2151 ^ n1432 ;
  assign n5473 = n4473 ^ n1104 ^ 1'b0 ;
  assign n5474 = n2360 & n4818 ;
  assign n5475 = n1966 ^ n1395 ^ x28 ;
  assign n5476 = ( n3096 & n5474 ) | ( n3096 & ~n5475 ) | ( n5474 & ~n5475 ) ;
  assign n5477 = n5280 ^ n3868 ^ n2891 ;
  assign n5478 = ( n369 & n1481 ) | ( n369 & n5477 ) | ( n1481 & n5477 ) ;
  assign n5479 = ( n5295 & ~n5476 ) | ( n5295 & n5478 ) | ( ~n5476 & n5478 ) ;
  assign n5480 = n5473 | n5479 ;
  assign n5501 = x43 & n338 ;
  assign n5502 = ~n783 & n5501 ;
  assign n5503 = n852 | n5502 ;
  assign n5504 = n5503 ^ x116 ^ 1'b0 ;
  assign n5505 = n1142 & n5504 ;
  assign n5506 = n5505 ^ n1487 ^ 1'b0 ;
  assign n5507 = n5506 ^ n2311 ^ 1'b0 ;
  assign n5497 = n479 & ~n609 ;
  assign n5498 = n5497 ^ n2325 ^ 1'b0 ;
  assign n5499 = n5498 ^ n2546 ^ n974 ;
  assign n5481 = ( n877 & n1108 ) | ( n877 & n1380 ) | ( n1108 & n1380 ) ;
  assign n5482 = ( n1513 & n2070 ) | ( n1513 & ~n5481 ) | ( n2070 & ~n5481 ) ;
  assign n5494 = ( n1172 & n3668 ) | ( n1172 & n4157 ) | ( n3668 & n4157 ) ;
  assign n5486 = n3731 ^ n686 ^ x114 ;
  assign n5485 = n4793 ^ n3721 ^ n2134 ;
  assign n5487 = n5486 ^ n5485 ^ n3604 ;
  assign n5488 = n5487 ^ n4105 ^ x47 ;
  assign n5489 = ( n599 & n1011 ) | ( n599 & n2091 ) | ( n1011 & n2091 ) ;
  assign n5490 = ( x99 & n2575 ) | ( x99 & ~n5489 ) | ( n2575 & ~n5489 ) ;
  assign n5491 = ( n5092 & n5488 ) | ( n5092 & n5490 ) | ( n5488 & n5490 ) ;
  assign n5483 = n264 | n1189 ;
  assign n5484 = n5007 & ~n5483 ;
  assign n5492 = n5491 ^ n5484 ^ 1'b0 ;
  assign n5493 = ~n1674 & n5492 ;
  assign n5495 = n5494 ^ n5493 ^ n1103 ;
  assign n5496 = n5482 & n5495 ;
  assign n5500 = n5499 ^ n5496 ^ 1'b0 ;
  assign n5508 = n5507 ^ n5500 ^ 1'b0 ;
  assign n5509 = n4508 ^ n1586 ^ 1'b0 ;
  assign n5510 = n4383 & n5509 ;
  assign n5511 = n5510 ^ n4019 ^ n3967 ;
  assign n5512 = n5511 ^ n4232 ^ n1372 ;
  assign n5520 = ( n465 & n1191 ) | ( n465 & n3838 ) | ( n1191 & n3838 ) ;
  assign n5521 = n3138 & ~n3621 ;
  assign n5522 = ~n5520 & n5521 ;
  assign n5517 = n2843 ^ n2268 ^ n1983 ;
  assign n5518 = n5517 ^ n3970 ^ n893 ;
  assign n5513 = n3621 ^ n2855 ^ n2576 ;
  assign n5514 = n5513 ^ n2424 ^ n1644 ;
  assign n5515 = ~n1685 & n5514 ;
  assign n5516 = n2617 & n5515 ;
  assign n5519 = n5518 ^ n5516 ^ n2391 ;
  assign n5523 = n5522 ^ n5519 ^ n3521 ;
  assign n5524 = n4935 ^ n4432 ^ n3063 ;
  assign n5525 = n5524 ^ n4723 ^ n3557 ;
  assign n5526 = ( n524 & n1292 ) | ( n524 & ~n4094 ) | ( n1292 & ~n4094 ) ;
  assign n5527 = n5526 ^ n3215 ^ n2945 ;
  assign n5528 = n3540 ^ n1114 ^ x40 ;
  assign n5529 = ( n254 & n3305 ) | ( n254 & ~n4267 ) | ( n3305 & ~n4267 ) ;
  assign n5530 = n5528 & ~n5529 ;
  assign n5531 = ~n2430 & n5530 ;
  assign n5532 = n5531 ^ n4485 ^ n2189 ;
  assign n5535 = x3 & n3700 ;
  assign n5536 = ~n1084 & n5535 ;
  assign n5533 = ( ~n841 & n2729 ) | ( ~n841 & n3089 ) | ( n2729 & n3089 ) ;
  assign n5534 = n2098 | n5533 ;
  assign n5537 = n5536 ^ n5534 ^ 1'b0 ;
  assign n5538 = n385 | n3374 ;
  assign n5539 = n5538 ^ n3640 ^ 1'b0 ;
  assign n5540 = ( n449 & n921 ) | ( n449 & ~n1132 ) | ( n921 & ~n1132 ) ;
  assign n5541 = ( ~n815 & n1780 ) | ( ~n815 & n5540 ) | ( n1780 & n5540 ) ;
  assign n5542 = ( n1810 & n2220 ) | ( n1810 & ~n3371 ) | ( n2220 & ~n3371 ) ;
  assign n5543 = n5542 ^ n2558 ^ n1713 ;
  assign n5544 = ( n1961 & ~n3707 ) | ( n1961 & n5543 ) | ( ~n3707 & n5543 ) ;
  assign n5545 = ( n1799 & n3237 ) | ( n1799 & ~n5544 ) | ( n3237 & ~n5544 ) ;
  assign n5546 = n3367 ^ n1991 ^ n1792 ;
  assign n5547 = n5546 ^ n1818 ^ 1'b0 ;
  assign n5548 = n564 & n997 ;
  assign n5549 = n5548 ^ n2579 ^ n2065 ;
  assign n5550 = ( n4578 & ~n5547 ) | ( n4578 & n5549 ) | ( ~n5547 & n5549 ) ;
  assign n5551 = ( n1521 & n4616 ) | ( n1521 & ~n5488 ) | ( n4616 & ~n5488 ) ;
  assign n5552 = n5551 ^ n4320 ^ n505 ;
  assign n5553 = n5552 ^ n1645 ^ 1'b0 ;
  assign n5554 = x80 & ~n5553 ;
  assign n5555 = ( ~n246 & n452 ) | ( ~n246 & n2367 ) | ( n452 & n2367 ) ;
  assign n5556 = n5555 ^ n3932 ^ 1'b0 ;
  assign n5557 = n5554 & n5556 ;
  assign n5558 = n155 & ~n2599 ;
  assign n5559 = n5558 ^ n368 ^ 1'b0 ;
  assign n5560 = n1740 ^ n699 ^ n489 ;
  assign n5561 = ( n1517 & ~n2965 ) | ( n1517 & n5560 ) | ( ~n2965 & n5560 ) ;
  assign n5562 = n4784 ^ n3801 ^ n2117 ;
  assign n5563 = n234 | n5562 ;
  assign n5564 = ( n5559 & n5561 ) | ( n5559 & ~n5563 ) | ( n5561 & ~n5563 ) ;
  assign n5565 = n4587 ^ n2809 ^ n2780 ;
  assign n5566 = n2434 & ~n3989 ;
  assign n5567 = ( n2046 & ~n5565 ) | ( n2046 & n5566 ) | ( ~n5565 & n5566 ) ;
  assign n5568 = n5567 ^ n4989 ^ n4157 ;
  assign n5569 = ( n469 & n1336 ) | ( n469 & n3759 ) | ( n1336 & n3759 ) ;
  assign n5570 = n2743 | n4219 ;
  assign n5571 = n5570 ^ n4468 ^ 1'b0 ;
  assign n5572 = ( n1176 & n3432 ) | ( n1176 & n4830 ) | ( n3432 & n4830 ) ;
  assign n5573 = n5572 ^ n3396 ^ n1412 ;
  assign n5574 = ( n2508 & n2990 ) | ( n2508 & n5573 ) | ( n2990 & n5573 ) ;
  assign n5575 = ( n2447 & ~n5571 ) | ( n2447 & n5574 ) | ( ~n5571 & n5574 ) ;
  assign n5576 = n2869 ^ n1648 ^ n1247 ;
  assign n5577 = n5576 ^ n1212 ^ 1'b0 ;
  assign n5590 = ( n1433 & n1491 ) | ( n1433 & ~n3777 ) | ( n1491 & ~n3777 ) ;
  assign n5589 = ~n278 & n3701 ;
  assign n5578 = n3539 ^ n1285 ^ 1'b0 ;
  assign n5579 = ( n3039 & n3127 ) | ( n3039 & n5578 ) | ( n3127 & n5578 ) ;
  assign n5580 = n5579 ^ n1572 ^ 1'b0 ;
  assign n5581 = n3916 & ~n5580 ;
  assign n5582 = n1829 ^ n1165 ^ n359 ;
  assign n5583 = ( n637 & n863 ) | ( n637 & ~n1351 ) | ( n863 & ~n1351 ) ;
  assign n5584 = n5583 ^ n4326 ^ n3030 ;
  assign n5585 = ( n302 & n5582 ) | ( n302 & ~n5584 ) | ( n5582 & ~n5584 ) ;
  assign n5586 = ( n3614 & n5581 ) | ( n3614 & n5585 ) | ( n5581 & n5585 ) ;
  assign n5587 = n5586 ^ n3712 ^ n1354 ;
  assign n5588 = n5587 ^ n4339 ^ n558 ;
  assign n5591 = n5590 ^ n5589 ^ n5588 ;
  assign n5594 = n341 | n1860 ;
  assign n5595 = n5594 ^ n1299 ^ 1'b0 ;
  assign n5592 = ( ~n1214 & n1467 ) | ( ~n1214 & n1667 ) | ( n1467 & n1667 ) ;
  assign n5593 = ( n1021 & n4714 ) | ( n1021 & ~n5592 ) | ( n4714 & ~n5592 ) ;
  assign n5596 = n5595 ^ n5593 ^ n1667 ;
  assign n5597 = n3998 ^ n3539 ^ n2117 ;
  assign n5598 = n1010 & ~n5597 ;
  assign n5599 = ( x82 & ~n1357 ) | ( x82 & n1615 ) | ( ~n1357 & n1615 ) ;
  assign n5600 = ( n209 & ~n2861 ) | ( n209 & n5599 ) | ( ~n2861 & n5599 ) ;
  assign n5601 = ( n4664 & n5114 ) | ( n4664 & ~n5600 ) | ( n5114 & ~n5600 ) ;
  assign n5602 = n5601 ^ n1615 ^ 1'b0 ;
  assign n5603 = n1693 & ~n5602 ;
  assign n5604 = ( n3516 & n3882 ) | ( n3516 & n5603 ) | ( n3882 & n5603 ) ;
  assign n5605 = ( n1698 & n5598 ) | ( n1698 & ~n5604 ) | ( n5598 & ~n5604 ) ;
  assign n5606 = ( n183 & n2280 ) | ( n183 & n4510 ) | ( n2280 & n4510 ) ;
  assign n5607 = ( ~n2123 & n5514 ) | ( ~n2123 & n5606 ) | ( n5514 & n5606 ) ;
  assign n5609 = ( n974 & n3650 ) | ( n974 & n4243 ) | ( n3650 & n4243 ) ;
  assign n5608 = n3346 & ~n3669 ;
  assign n5610 = n5609 ^ n5608 ^ n3665 ;
  assign n5611 = ( ~n263 & n2183 ) | ( ~n263 & n5610 ) | ( n2183 & n5610 ) ;
  assign n5612 = n5223 | n5611 ;
  assign n5613 = n572 & ~n5612 ;
  assign n5614 = n1034 & ~n1044 ;
  assign n5615 = n5614 ^ n1359 ^ 1'b0 ;
  assign n5616 = ~n5613 & n5615 ;
  assign n5617 = n1786 | n4485 ;
  assign n5618 = n1020 | n5617 ;
  assign n5619 = ( n167 & n909 ) | ( n167 & n2538 ) | ( n909 & n2538 ) ;
  assign n5620 = n5618 & ~n5619 ;
  assign n5621 = n5620 ^ n3310 ^ 1'b0 ;
  assign n5622 = ( n886 & n1006 ) | ( n886 & n2879 ) | ( n1006 & n2879 ) ;
  assign n5624 = n1314 ^ n903 ^ x50 ;
  assign n5625 = ( n903 & ~n3236 ) | ( n903 & n5624 ) | ( ~n3236 & n5624 ) ;
  assign n5623 = n4946 ^ n4934 ^ n2902 ;
  assign n5626 = n5625 ^ n5623 ^ 1'b0 ;
  assign n5627 = n5622 & ~n5626 ;
  assign n5628 = ( ~n3217 & n3277 ) | ( ~n3217 & n3800 ) | ( n3277 & n3800 ) ;
  assign n5629 = ( n1569 & n3717 ) | ( n1569 & ~n4878 ) | ( n3717 & ~n4878 ) ;
  assign n5633 = n3896 ^ n2721 ^ 1'b0 ;
  assign n5634 = n5476 & n5633 ;
  assign n5630 = n2523 ^ n2256 ^ n244 ;
  assign n5631 = n5630 ^ n4377 ^ n2461 ;
  assign n5632 = ( n582 & n3403 ) | ( n582 & ~n5631 ) | ( n3403 & ~n5631 ) ;
  assign n5635 = n5634 ^ n5632 ^ n4966 ;
  assign n5636 = n3818 ^ n3450 ^ n3011 ;
  assign n5637 = n5636 ^ n2797 ^ n315 ;
  assign n5638 = n3753 ^ n3025 ^ n709 ;
  assign n5639 = ( n2402 & n5056 ) | ( n2402 & ~n5638 ) | ( n5056 & ~n5638 ) ;
  assign n5645 = n2291 ^ n1037 ^ n564 ;
  assign n5640 = ( n872 & n966 ) | ( n872 & ~n2047 ) | ( n966 & ~n2047 ) ;
  assign n5641 = ( n3880 & n5185 ) | ( n3880 & ~n5640 ) | ( n5185 & ~n5640 ) ;
  assign n5642 = n5641 ^ n1121 ^ x33 ;
  assign n5643 = n3203 | n5642 ;
  assign n5644 = ( ~n1179 & n2629 ) | ( ~n1179 & n5643 ) | ( n2629 & n5643 ) ;
  assign n5646 = n5645 ^ n5644 ^ 1'b0 ;
  assign n5647 = n5639 | n5646 ;
  assign n5648 = ( ~n800 & n1335 ) | ( ~n800 & n5336 ) | ( n1335 & n5336 ) ;
  assign n5649 = n3192 ^ n2712 ^ n393 ;
  assign n5650 = ( n3792 & n4791 ) | ( n3792 & n5649 ) | ( n4791 & n5649 ) ;
  assign n5651 = ~n5648 & n5650 ;
  assign n5652 = n5320 & n5651 ;
  assign n5653 = ~n3881 & n5652 ;
  assign n5654 = ( ~n662 & n3710 ) | ( ~n662 & n5653 ) | ( n3710 & n5653 ) ;
  assign n5655 = n1252 & n5200 ;
  assign n5656 = ~n4160 & n5655 ;
  assign n5658 = ( n394 & n2163 ) | ( n394 & n4850 ) | ( n2163 & n4850 ) ;
  assign n5657 = n5431 ^ n2658 ^ n790 ;
  assign n5659 = n5658 ^ n5657 ^ n1329 ;
  assign n5660 = n2829 ^ n1687 ^ 1'b0 ;
  assign n5661 = n5660 ^ n2260 ^ n1079 ;
  assign n5662 = ( n1469 & n3338 ) | ( n1469 & n5661 ) | ( n3338 & n5661 ) ;
  assign n5663 = n5662 ^ n493 ^ 1'b0 ;
  assign n5664 = n5659 & ~n5663 ;
  assign n5665 = n2177 ^ n1782 ^ 1'b0 ;
  assign n5666 = n4538 | n5665 ;
  assign n5671 = ( n1423 & ~n1467 ) | ( n1423 & n4549 ) | ( ~n1467 & n4549 ) ;
  assign n5672 = n5671 ^ n4085 ^ n1675 ;
  assign n5673 = n1478 ^ n819 ^ 1'b0 ;
  assign n5674 = n5672 & ~n5673 ;
  assign n5667 = ( ~x100 & n140 ) | ( ~x100 & n3105 ) | ( n140 & n3105 ) ;
  assign n5668 = n5667 ^ n3391 ^ n3179 ;
  assign n5669 = n1455 ^ n207 ^ 1'b0 ;
  assign n5670 = n5668 & ~n5669 ;
  assign n5675 = n5674 ^ n5670 ^ x53 ;
  assign n5676 = n5675 ^ n748 ^ n421 ;
  assign n5677 = n5676 ^ n1285 ^ n902 ;
  assign n5678 = n5489 ^ n3068 ^ n352 ;
  assign n5680 = ~n1206 & n1455 ;
  assign n5681 = n5015 ^ n2121 ^ n2089 ;
  assign n5682 = n5681 ^ n2507 ^ x43 ;
  assign n5683 = ( ~n3500 & n5680 ) | ( ~n3500 & n5682 ) | ( n5680 & n5682 ) ;
  assign n5679 = n1281 & ~n3222 ;
  assign n5684 = n5683 ^ n5679 ^ 1'b0 ;
  assign n5685 = n3160 ^ n149 ^ 1'b0 ;
  assign n5686 = n3888 | n5685 ;
  assign n5687 = ( n201 & ~n1899 ) | ( n201 & n5310 ) | ( ~n1899 & n5310 ) ;
  assign n5688 = n5687 ^ n3641 ^ n2174 ;
  assign n5689 = ( n5684 & ~n5686 ) | ( n5684 & n5688 ) | ( ~n5686 & n5688 ) ;
  assign n5690 = x123 & n2384 ;
  assign n5691 = n5690 ^ n317 ^ 1'b0 ;
  assign n5692 = ( n159 & ~n3610 ) | ( n159 & n5691 ) | ( ~n3610 & n5691 ) ;
  assign n5693 = n2396 & n4748 ;
  assign n5694 = n5693 ^ n2864 ^ n680 ;
  assign n5695 = n5694 ^ n1040 ^ n342 ;
  assign n5696 = ( n501 & ~n5692 ) | ( n501 & n5695 ) | ( ~n5692 & n5695 ) ;
  assign n5697 = n5696 ^ n1490 ^ n356 ;
  assign n5698 = ( n5678 & ~n5689 ) | ( n5678 & n5697 ) | ( ~n5689 & n5697 ) ;
  assign n5702 = ( ~n1045 & n1169 ) | ( ~n1045 & n4964 ) | ( n1169 & n4964 ) ;
  assign n5699 = n2529 ^ n1095 ^ 1'b0 ;
  assign n5700 = n929 & n5699 ;
  assign n5701 = n5700 ^ n561 ^ n319 ;
  assign n5703 = n5702 ^ n5701 ^ n5670 ;
  assign n5704 = n5703 ^ n1014 ^ x55 ;
  assign n5705 = n4217 ^ n329 ^ n179 ;
  assign n5707 = n5017 ^ n3023 ^ n582 ;
  assign n5706 = ( n1302 & ~n2663 ) | ( n1302 & n3136 ) | ( ~n2663 & n3136 ) ;
  assign n5708 = n5707 ^ n5706 ^ n772 ;
  assign n5710 = n1872 & ~n3111 ;
  assign n5709 = ( n1254 & n2175 ) | ( n1254 & n4217 ) | ( n2175 & n4217 ) ;
  assign n5711 = n5710 ^ n5709 ^ 1'b0 ;
  assign n5712 = n5708 & ~n5711 ;
  assign n5713 = ( n3171 & ~n5705 ) | ( n3171 & n5712 ) | ( ~n5705 & n5712 ) ;
  assign n5715 = n4375 ^ n1837 ^ n1614 ;
  assign n5714 = ( ~n742 & n1745 ) | ( ~n742 & n2363 ) | ( n1745 & n2363 ) ;
  assign n5716 = n5715 ^ n5714 ^ n2637 ;
  assign n5717 = n5713 & n5716 ;
  assign n5718 = n5704 & n5717 ;
  assign n5719 = n1643 & ~n2121 ;
  assign n5720 = ( n2077 & n4100 ) | ( n2077 & n5719 ) | ( n4100 & n5719 ) ;
  assign n5721 = n2030 ^ n130 ^ x11 ;
  assign n5722 = n5721 ^ n2762 ^ n749 ;
  assign n5723 = n5720 | n5722 ;
  assign n5724 = n2443 | n3105 ;
  assign n5726 = n2619 ^ n1397 ^ x2 ;
  assign n5727 = n3088 | n5726 ;
  assign n5728 = n1549 & n5727 ;
  assign n5729 = n5728 ^ x14 ^ 1'b0 ;
  assign n5730 = ( n3460 & n4583 ) | ( n3460 & n5729 ) | ( n4583 & n5729 ) ;
  assign n5731 = n2175 ^ n1960 ^ 1'b0 ;
  assign n5732 = n5731 ^ n2900 ^ n1254 ;
  assign n5733 = n5732 ^ n5390 ^ n2659 ;
  assign n5734 = ( n4031 & ~n5730 ) | ( n4031 & n5733 ) | ( ~n5730 & n5733 ) ;
  assign n5725 = n4645 ^ n4260 ^ 1'b0 ;
  assign n5735 = n5734 ^ n5725 ^ n4339 ;
  assign n5736 = ( n1421 & n1971 ) | ( n1421 & ~n4934 ) | ( n1971 & ~n4934 ) ;
  assign n5738 = ( n613 & n3791 ) | ( n613 & n4588 ) | ( n3791 & n4588 ) ;
  assign n5739 = n5738 ^ n4277 ^ 1'b0 ;
  assign n5740 = n2855 & n5739 ;
  assign n5741 = n4657 ^ n1444 ^ 1'b0 ;
  assign n5742 = ~n3754 & n5741 ;
  assign n5743 = ( n2754 & n5740 ) | ( n2754 & ~n5742 ) | ( n5740 & ~n5742 ) ;
  assign n5737 = n4550 & ~n5100 ;
  assign n5744 = n5743 ^ n5737 ^ 1'b0 ;
  assign n5745 = ( n199 & n5736 ) | ( n199 & ~n5744 ) | ( n5736 & ~n5744 ) ;
  assign n5749 = ( ~n2130 & n2730 ) | ( ~n2130 & n5610 ) | ( n2730 & n5610 ) ;
  assign n5746 = ~n2350 & n4782 ;
  assign n5747 = n922 & n5746 ;
  assign n5748 = ( n369 & ~n2019 ) | ( n369 & n5747 ) | ( ~n2019 & n5747 ) ;
  assign n5750 = n5749 ^ n5748 ^ n3262 ;
  assign n5751 = ( ~n1206 & n4885 ) | ( ~n1206 & n5593 ) | ( n4885 & n5593 ) ;
  assign n5760 = ( ~n996 & n1834 ) | ( ~n996 & n4375 ) | ( n1834 & n4375 ) ;
  assign n5761 = n5760 ^ n2291 ^ x27 ;
  assign n5752 = ( n1998 & n2157 ) | ( n1998 & n4144 ) | ( n2157 & n4144 ) ;
  assign n5753 = ( ~n1904 & n2268 ) | ( ~n1904 & n2406 ) | ( n2268 & n2406 ) ;
  assign n5754 = n5753 ^ n667 ^ n263 ;
  assign n5755 = n963 ^ n893 ^ 1'b0 ;
  assign n5756 = n5754 | n5755 ;
  assign n5757 = ~n5752 & n5756 ;
  assign n5758 = n5757 ^ n3120 ^ 1'b0 ;
  assign n5759 = n2139 | n5758 ;
  assign n5762 = n5761 ^ n5759 ^ n4769 ;
  assign n5763 = n3020 ^ n1150 ^ n578 ;
  assign n5764 = n2702 | n5763 ;
  assign n5765 = n5764 ^ n753 ^ 1'b0 ;
  assign n5766 = n3576 ^ n387 ^ 1'b0 ;
  assign n5767 = ~n769 & n3684 ;
  assign n5768 = ~n2436 & n5767 ;
  assign n5769 = n2562 ^ n2073 ^ n1431 ;
  assign n5770 = n4657 ^ n987 ^ n273 ;
  assign n5771 = n5769 & n5770 ;
  assign n5772 = ~x104 & n5771 ;
  assign n5773 = ( n249 & n735 ) | ( n249 & ~n3441 ) | ( n735 & ~n3441 ) ;
  assign n5774 = ( n2843 & n2918 ) | ( n2843 & n5307 ) | ( n2918 & n5307 ) ;
  assign n5775 = ( ~n1636 & n5773 ) | ( ~n1636 & n5774 ) | ( n5773 & n5774 ) ;
  assign n5776 = ~n1544 & n3892 ;
  assign n5777 = n5776 ^ n3225 ^ 1'b0 ;
  assign n5778 = ~n972 & n2936 ;
  assign n5779 = n5778 ^ n3480 ^ 1'b0 ;
  assign n5780 = n5779 ^ n4968 ^ n4891 ;
  assign n5781 = ~n2262 & n2466 ;
  assign n5784 = n2721 ^ n2049 ^ n1176 ;
  assign n5782 = n3652 ^ n1610 ^ n944 ;
  assign n5783 = n5782 ^ n3111 ^ n2050 ;
  assign n5785 = n5784 ^ n5783 ^ 1'b0 ;
  assign n5786 = n3547 ^ n896 ^ 1'b0 ;
  assign n5787 = ( n1756 & n5785 ) | ( n1756 & n5786 ) | ( n5785 & n5786 ) ;
  assign n5788 = n1251 & ~n5295 ;
  assign n5789 = n5566 & n5788 ;
  assign n5791 = n5226 ^ n2450 ^ 1'b0 ;
  assign n5790 = n2680 ^ n1709 ^ n994 ;
  assign n5792 = n5791 ^ n5790 ^ 1'b0 ;
  assign n5796 = ( n1115 & n1580 ) | ( n1115 & ~n3131 ) | ( n1580 & ~n3131 ) ;
  assign n5795 = n3561 ^ n2157 ^ n1420 ;
  assign n5794 = n3972 ^ n3606 ^ n2930 ;
  assign n5797 = n5796 ^ n5795 ^ n5794 ;
  assign n5793 = ( n2745 & ~n2754 ) | ( n2745 & n5276 ) | ( ~n2754 & n5276 ) ;
  assign n5798 = n5797 ^ n5793 ^ n1709 ;
  assign n5799 = ( x121 & n1091 ) | ( x121 & n2311 ) | ( n1091 & n2311 ) ;
  assign n5800 = ( n966 & ~n1351 ) | ( n966 & n1464 ) | ( ~n1351 & n1464 ) ;
  assign n5801 = ( n160 & n247 ) | ( n160 & n5800 ) | ( n247 & n5800 ) ;
  assign n5802 = ( n1778 & ~n5799 ) | ( n1778 & n5801 ) | ( ~n5799 & n5801 ) ;
  assign n5803 = ( ~n1502 & n3272 ) | ( ~n1502 & n3624 ) | ( n3272 & n3624 ) ;
  assign n5804 = ( n1154 & n3742 ) | ( n1154 & ~n5803 ) | ( n3742 & ~n5803 ) ;
  assign n5805 = ( n306 & n5802 ) | ( n306 & ~n5804 ) | ( n5802 & ~n5804 ) ;
  assign n5806 = n5411 | n5805 ;
  assign n5807 = n2872 | n5806 ;
  assign n5808 = n2540 ^ n2225 ^ n2132 ;
  assign n5809 = ( n1101 & n3219 ) | ( n1101 & n5808 ) | ( n3219 & n5808 ) ;
  assign n5810 = ( n5214 & n5391 ) | ( n5214 & ~n5809 ) | ( n5391 & ~n5809 ) ;
  assign n5811 = ( n1046 & n3331 ) | ( n1046 & ~n4061 ) | ( n3331 & ~n4061 ) ;
  assign n5812 = n5254 ^ n3646 ^ 1'b0 ;
  assign n5814 = ( ~n1731 & n1912 ) | ( ~n1731 & n3164 ) | ( n1912 & n3164 ) ;
  assign n5813 = n830 & ~n1064 ;
  assign n5815 = n5814 ^ n5813 ^ n4947 ;
  assign n5818 = ( n470 & ~n1395 ) | ( n470 & n1451 ) | ( ~n1395 & n1451 ) ;
  assign n5816 = ( n2488 & n3507 ) | ( n2488 & n5097 ) | ( n3507 & n5097 ) ;
  assign n5817 = n1948 | n5816 ;
  assign n5819 = n5818 ^ n5817 ^ 1'b0 ;
  assign n5820 = n3731 & n4439 ;
  assign n5821 = n1417 & n3425 ;
  assign n5825 = ( x122 & ~n2249 ) | ( x122 & n4791 ) | ( ~n2249 & n4791 ) ;
  assign n5822 = ( ~n1767 & n3026 ) | ( ~n1767 & n5088 ) | ( n3026 & n5088 ) ;
  assign n5823 = n3278 & ~n5822 ;
  assign n5824 = n5823 ^ n2124 ^ 1'b0 ;
  assign n5826 = n5825 ^ n5824 ^ n688 ;
  assign n5827 = ( n596 & n3389 ) | ( n596 & ~n4641 ) | ( n3389 & ~n4641 ) ;
  assign n5828 = n2579 ^ n2409 ^ n951 ;
  assign n5829 = ~n1674 & n3792 ;
  assign n5830 = n5829 ^ n1337 ^ 1'b0 ;
  assign n5831 = ( n3345 & n5828 ) | ( n3345 & ~n5830 ) | ( n5828 & ~n5830 ) ;
  assign n5832 = n5831 ^ n5727 ^ 1'b0 ;
  assign n5833 = ~n471 & n5832 ;
  assign n5834 = ~n291 & n2877 ;
  assign n5835 = n5834 ^ n5598 ^ n337 ;
  assign n5836 = n549 & n885 ;
  assign n5837 = n4296 ^ n3805 ^ n3755 ;
  assign n5838 = ( n3405 & n5836 ) | ( n3405 & n5837 ) | ( n5836 & n5837 ) ;
  assign n5839 = ( n3977 & n5567 ) | ( n3977 & ~n5838 ) | ( n5567 & ~n5838 ) ;
  assign n5840 = ( n2754 & n5835 ) | ( n2754 & ~n5839 ) | ( n5835 & ~n5839 ) ;
  assign n5844 = n1895 ^ n1374 ^ n1146 ;
  assign n5841 = n1865 ^ n805 ^ n500 ;
  assign n5842 = n4813 ^ n4360 ^ 1'b0 ;
  assign n5843 = ~n5841 & n5842 ;
  assign n5845 = n5844 ^ n5843 ^ 1'b0 ;
  assign n5846 = n3403 & ~n5845 ;
  assign n5847 = ( n536 & n1799 ) | ( n536 & ~n5018 ) | ( n1799 & ~n5018 ) ;
  assign n5848 = n1617 ^ n564 ^ 1'b0 ;
  assign n5849 = n3093 | n5848 ;
  assign n5853 = ~n782 & n4417 ;
  assign n5854 = n5853 ^ n5340 ^ 1'b0 ;
  assign n5852 = n4231 ^ n2088 ^ n1216 ;
  assign n5851 = n1990 ^ n1425 ^ n250 ;
  assign n5855 = n5854 ^ n5852 ^ n5851 ;
  assign n5850 = ( n2483 & n3048 ) | ( n2483 & ~n3484 ) | ( n3048 & ~n3484 ) ;
  assign n5856 = n5855 ^ n5850 ^ 1'b0 ;
  assign n5857 = n3941 ^ n3361 ^ 1'b0 ;
  assign n5858 = n2834 & ~n5857 ;
  assign n5859 = ( ~x17 & n1675 ) | ( ~x17 & n1745 ) | ( n1675 & n1745 ) ;
  assign n5860 = ( ~n372 & n5858 ) | ( ~n372 & n5859 ) | ( n5858 & n5859 ) ;
  assign n5870 = n2510 ^ n1941 ^ x28 ;
  assign n5871 = ( ~n4400 & n5259 ) | ( ~n4400 & n5870 ) | ( n5259 & n5870 ) ;
  assign n5872 = n4357 ^ n3782 ^ n478 ;
  assign n5873 = ( n3192 & ~n5871 ) | ( n3192 & n5872 ) | ( ~n5871 & n5872 ) ;
  assign n5861 = n806 ^ n665 ^ 1'b0 ;
  assign n5862 = n382 | n5861 ;
  assign n5863 = n2609 & n3137 ;
  assign n5864 = ~n1637 & n5863 ;
  assign n5865 = ( ~n351 & n1549 ) | ( ~n351 & n5864 ) | ( n1549 & n5864 ) ;
  assign n5866 = n5865 ^ n3115 ^ n2333 ;
  assign n5867 = x30 & n5866 ;
  assign n5868 = n5862 & n5867 ;
  assign n5869 = ( n1657 & n5273 ) | ( n1657 & ~n5868 ) | ( n5273 & ~n5868 ) ;
  assign n5874 = n5873 ^ n5869 ^ 1'b0 ;
  assign n5875 = n1112 ^ n369 ^ n202 ;
  assign n5876 = ( n1589 & n4546 ) | ( n1589 & ~n5875 ) | ( n4546 & ~n5875 ) ;
  assign n5877 = n5876 ^ n4891 ^ 1'b0 ;
  assign n5878 = n3112 ^ n2368 ^ 1'b0 ;
  assign n5879 = ( n1765 & n3471 ) | ( n1765 & n5878 ) | ( n3471 & n5878 ) ;
  assign n5880 = ( n2231 & ~n4213 ) | ( n2231 & n4260 ) | ( ~n4213 & n4260 ) ;
  assign n5881 = ( ~n1365 & n5879 ) | ( ~n1365 & n5880 ) | ( n5879 & n5880 ) ;
  assign n5882 = n5881 ^ n2663 ^ 1'b0 ;
  assign n5883 = n2130 ^ n1557 ^ 1'b0 ;
  assign n5884 = n448 & ~n5883 ;
  assign n5885 = n5884 ^ n2384 ^ n1584 ;
  assign n5886 = ( n1502 & n4613 ) | ( n1502 & ~n5885 ) | ( n4613 & ~n5885 ) ;
  assign n5887 = ( n2307 & n5882 ) | ( n2307 & ~n5886 ) | ( n5882 & ~n5886 ) ;
  assign n5888 = n1503 & n1627 ;
  assign n5889 = n5888 ^ n3452 ^ n3392 ;
  assign n5891 = n777 & ~n4950 ;
  assign n5892 = n5891 ^ n2436 ^ 1'b0 ;
  assign n5893 = n5892 ^ n3693 ^ n3046 ;
  assign n5890 = n1288 & n5708 ;
  assign n5894 = n5893 ^ n5890 ^ 1'b0 ;
  assign n5895 = ( ~n1589 & n4194 ) | ( ~n1589 & n5601 ) | ( n4194 & n5601 ) ;
  assign n5912 = n4976 ^ n3773 ^ n466 ;
  assign n5908 = ( n472 & n737 ) | ( n472 & n2859 ) | ( n737 & n2859 ) ;
  assign n5905 = ( n502 & n1504 ) | ( n502 & ~n2086 ) | ( n1504 & ~n2086 ) ;
  assign n5906 = n5905 ^ n1460 ^ n1265 ;
  assign n5907 = ~n769 & n5906 ;
  assign n5909 = n5908 ^ n5907 ^ 1'b0 ;
  assign n5903 = ( n1065 & n2165 ) | ( n1065 & ~n3997 ) | ( n2165 & ~n3997 ) ;
  assign n5904 = n5903 ^ n3229 ^ n675 ;
  assign n5910 = n5909 ^ n5904 ^ n3594 ;
  assign n5911 = n5910 ^ n2594 ^ n2499 ;
  assign n5899 = n4260 ^ n2885 ^ n852 ;
  assign n5900 = n5899 ^ n2832 ^ 1'b0 ;
  assign n5901 = n4689 | n5900 ;
  assign n5896 = n3292 ^ n3155 ^ n1124 ;
  assign n5897 = n4987 ^ n2105 ^ 1'b0 ;
  assign n5898 = ~n5896 & n5897 ;
  assign n5902 = n5901 ^ n5898 ^ n1290 ;
  assign n5913 = n5912 ^ n5911 ^ n5902 ;
  assign n5914 = n1502 ^ n1411 ^ 1'b0 ;
  assign n5915 = ( ~n1533 & n1724 ) | ( ~n1533 & n3361 ) | ( n1724 & n3361 ) ;
  assign n5916 = ( ~n3690 & n5914 ) | ( ~n3690 & n5915 ) | ( n5914 & n5915 ) ;
  assign n5917 = ( n3193 & n4267 ) | ( n3193 & ~n5916 ) | ( n4267 & ~n5916 ) ;
  assign n5920 = n3573 ^ n2809 ^ n2022 ;
  assign n5918 = n153 & ~n1663 ;
  assign n5919 = n5918 ^ n4502 ^ 1'b0 ;
  assign n5921 = n5920 ^ n5919 ^ n4880 ;
  assign n5922 = n5917 & n5921 ;
  assign n5923 = n5922 ^ n4286 ^ n453 ;
  assign n5933 = n4586 ^ n878 ^ n509 ;
  assign n5930 = n5295 ^ n5061 ^ n4877 ;
  assign n5931 = ( n1405 & n2726 ) | ( n1405 & n5930 ) | ( n2726 & n5930 ) ;
  assign n5932 = ( n1879 & ~n1896 ) | ( n1879 & n5931 ) | ( ~n1896 & n5931 ) ;
  assign n5924 = n2397 ^ n1464 ^ n905 ;
  assign n5925 = n1022 | n5924 ;
  assign n5926 = n1542 ^ n935 ^ n192 ;
  assign n5927 = n4511 & n5926 ;
  assign n5928 = ~n5925 & n5927 ;
  assign n5929 = n5928 ^ n2664 ^ 1'b0 ;
  assign n5934 = n5933 ^ n5932 ^ n5929 ;
  assign n5936 = n3111 ^ n1444 ^ 1'b0 ;
  assign n5937 = n1057 & ~n5936 ;
  assign n5935 = ~n2701 & n5705 ;
  assign n5938 = n5937 ^ n5935 ^ n3800 ;
  assign n5939 = n4093 ^ n3247 ^ n2696 ;
  assign n5940 = ( ~x83 & n1870 ) | ( ~x83 & n5939 ) | ( n1870 & n5939 ) ;
  assign n5941 = x89 & n780 ;
  assign n5942 = n5941 ^ n4294 ^ 1'b0 ;
  assign n5943 = ( n719 & n3487 ) | ( n719 & ~n5942 ) | ( n3487 & ~n5942 ) ;
  assign n5944 = n2751 & n3360 ;
  assign n5945 = n5943 & n5944 ;
  assign n5946 = ( n2521 & ~n4804 ) | ( n2521 & n5945 ) | ( ~n4804 & n5945 ) ;
  assign n5947 = x121 & ~n5946 ;
  assign n5948 = ~n2525 & n5947 ;
  assign n5949 = ( ~n665 & n1274 ) | ( ~n665 & n3341 ) | ( n1274 & n3341 ) ;
  assign n5950 = ( n2554 & ~n4500 ) | ( n2554 & n5949 ) | ( ~n4500 & n5949 ) ;
  assign n5951 = ( n4177 & ~n4186 ) | ( n4177 & n5950 ) | ( ~n4186 & n5950 ) ;
  assign n5952 = n216 | n3452 ;
  assign n5953 = n772 & ~n5952 ;
  assign n5962 = ( ~n163 & n1225 ) | ( ~n163 & n3287 ) | ( n1225 & n3287 ) ;
  assign n5960 = ( ~n793 & n1860 ) | ( ~n793 & n3146 ) | ( n1860 & n3146 ) ;
  assign n5961 = n5960 ^ n3984 ^ n1676 ;
  assign n5958 = n3669 ^ n2838 ^ n1187 ;
  assign n5954 = ( ~n1700 & n2690 ) | ( ~n1700 & n4662 ) | ( n2690 & n4662 ) ;
  assign n5955 = ( n508 & n4158 ) | ( n508 & n5954 ) | ( n4158 & n5954 ) ;
  assign n5956 = n1928 ^ n1893 ^ n1438 ;
  assign n5957 = n5955 & ~n5956 ;
  assign n5959 = n5958 ^ n5957 ^ 1'b0 ;
  assign n5963 = n5962 ^ n5961 ^ n5959 ;
  assign n5964 = n3241 ^ n2327 ^ x3 ;
  assign n5965 = n4097 ^ n3477 ^ n1539 ;
  assign n5966 = ( n441 & n5964 ) | ( n441 & ~n5965 ) | ( n5964 & ~n5965 ) ;
  assign n5967 = n2724 ^ n1168 ^ n232 ;
  assign n5968 = ( ~n619 & n1446 ) | ( ~n619 & n5967 ) | ( n1446 & n5967 ) ;
  assign n5969 = ( n3481 & n5966 ) | ( n3481 & ~n5968 ) | ( n5966 & ~n5968 ) ;
  assign n5970 = ( n5953 & ~n5963 ) | ( n5953 & n5969 ) | ( ~n5963 & n5969 ) ;
  assign n5971 = ( n1068 & n3012 ) | ( n1068 & n4764 ) | ( n3012 & n4764 ) ;
  assign n5989 = ( n709 & n945 ) | ( n709 & n3761 ) | ( n945 & n3761 ) ;
  assign n5990 = n5989 ^ n943 ^ n919 ;
  assign n5986 = n426 & ~n2285 ;
  assign n5987 = n5072 & n5986 ;
  assign n5982 = ( x123 & n1784 ) | ( x123 & n2869 ) | ( n1784 & n2869 ) ;
  assign n5983 = n5982 ^ n1121 ^ 1'b0 ;
  assign n5984 = n5983 ^ n2089 ^ n1022 ;
  assign n5985 = n4557 | n5984 ;
  assign n5988 = n5987 ^ n5985 ^ 1'b0 ;
  assign n5979 = n1680 ^ n379 ^ 1'b0 ;
  assign n5977 = ( n778 & n1030 ) | ( n778 & n2539 ) | ( n1030 & n2539 ) ;
  assign n5975 = ( n255 & ~n2509 ) | ( n255 & n3622 ) | ( ~n2509 & n3622 ) ;
  assign n5976 = n3062 & ~n5975 ;
  assign n5978 = n5977 ^ n5976 ^ 1'b0 ;
  assign n5980 = n5979 ^ n5978 ^ 1'b0 ;
  assign n5972 = n3126 ^ n3040 ^ n235 ;
  assign n5973 = n5972 ^ n2773 ^ n987 ;
  assign n5974 = ( n4538 & ~n4793 ) | ( n4538 & n5973 ) | ( ~n4793 & n5973 ) ;
  assign n5981 = n5980 ^ n5974 ^ n4852 ;
  assign n5991 = n5990 ^ n5988 ^ n5981 ;
  assign n5992 = ( n5804 & ~n5971 ) | ( n5804 & n5991 ) | ( ~n5971 & n5991 ) ;
  assign n5993 = n5006 ^ n3953 ^ n347 ;
  assign n5994 = n2959 | n5993 ;
  assign n5995 = n5994 ^ n918 ^ 1'b0 ;
  assign n5996 = ~n373 & n2094 ;
  assign n5997 = n5996 ^ x58 ^ 1'b0 ;
  assign n5998 = n1284 | n5997 ;
  assign n5999 = n1180 | n2132 ;
  assign n6000 = n4934 & ~n5999 ;
  assign n6001 = n6000 ^ n5413 ^ 1'b0 ;
  assign n6002 = n736 & ~n1405 ;
  assign n6003 = n517 | n2405 ;
  assign n6004 = n6003 ^ n3170 ^ 1'b0 ;
  assign n6008 = ( n1983 & n4580 ) | ( n1983 & n5783 ) | ( n4580 & n5783 ) ;
  assign n6009 = ( n694 & n5560 ) | ( n694 & ~n6008 ) | ( n5560 & ~n6008 ) ;
  assign n6005 = n2940 ^ n1857 ^ 1'b0 ;
  assign n6006 = ( n1203 & n2479 ) | ( n1203 & ~n6005 ) | ( n2479 & ~n6005 ) ;
  assign n6007 = ( ~n3093 & n4907 ) | ( ~n3093 & n6006 ) | ( n4907 & n6006 ) ;
  assign n6010 = n6009 ^ n6007 ^ 1'b0 ;
  assign n6011 = n6004 & n6010 ;
  assign n6012 = n2737 ^ n545 ^ 1'b0 ;
  assign n6013 = n2596 & n6012 ;
  assign n6014 = n6013 ^ n1213 ^ 1'b0 ;
  assign n6015 = ~n4075 & n6014 ;
  assign n6016 = n864 & n6015 ;
  assign n6017 = n6007 | n6016 ;
  assign n6018 = n882 & ~n6017 ;
  assign n6019 = ( n180 & n2088 ) | ( n180 & ~n3967 ) | ( n2088 & ~n3967 ) ;
  assign n6020 = ( n261 & ~n808 ) | ( n261 & n3143 ) | ( ~n808 & n3143 ) ;
  assign n6021 = n6020 ^ n1513 ^ n245 ;
  assign n6022 = ( ~n3733 & n5834 ) | ( ~n3733 & n6021 ) | ( n5834 & n6021 ) ;
  assign n6023 = n250 & n582 ;
  assign n6024 = ~n2358 & n6023 ;
  assign n6025 = n2957 | n6024 ;
  assign n6026 = n6025 ^ n1329 ^ 1'b0 ;
  assign n6027 = n6026 ^ n5341 ^ n2396 ;
  assign n6028 = n1166 & n3526 ;
  assign n6029 = ~n404 & n6028 ;
  assign n6030 = n4294 ^ n3593 ^ n724 ;
  assign n6031 = n384 & ~n3402 ;
  assign n6032 = n6031 ^ n1791 ^ 1'b0 ;
  assign n6033 = ( n6029 & n6030 ) | ( n6029 & ~n6032 ) | ( n6030 & ~n6032 ) ;
  assign n6034 = ( n2209 & n2563 ) | ( n2209 & n6033 ) | ( n2563 & n6033 ) ;
  assign n6035 = ( n822 & n6027 ) | ( n822 & ~n6034 ) | ( n6027 & ~n6034 ) ;
  assign n6036 = n2900 ^ n1997 ^ n539 ;
  assign n6037 = n1621 ^ n829 ^ 1'b0 ;
  assign n6038 = n4853 | n6037 ;
  assign n6039 = ( n2953 & n3885 ) | ( n2953 & ~n6038 ) | ( n3885 & ~n6038 ) ;
  assign n6040 = n4495 ^ x124 ^ 1'b0 ;
  assign n6041 = ( n5346 & n5925 ) | ( n5346 & n6040 ) | ( n5925 & n6040 ) ;
  assign n6042 = ( n442 & n4936 ) | ( n442 & ~n5250 ) | ( n4936 & ~n5250 ) ;
  assign n6048 = n1777 & ~n2603 ;
  assign n6049 = n918 & ~n6048 ;
  assign n6050 = ~n4190 & n6049 ;
  assign n6043 = n1923 ^ n1603 ^ n930 ;
  assign n6044 = n3666 ^ n2900 ^ n1103 ;
  assign n6045 = ( ~x119 & n6043 ) | ( ~x119 & n6044 ) | ( n6043 & n6044 ) ;
  assign n6046 = ( n2626 & n5854 ) | ( n2626 & n6045 ) | ( n5854 & n6045 ) ;
  assign n6047 = n6046 ^ n5943 ^ n1419 ;
  assign n6051 = n6050 ^ n6047 ^ n5352 ;
  assign n6052 = n5813 ^ n4640 ^ n231 ;
  assign n6053 = n3988 & n6052 ;
  assign n6054 = n6053 ^ x81 ^ 1'b0 ;
  assign n6055 = n5002 ^ n2378 ^ n1369 ;
  assign n6056 = n6055 ^ n5520 ^ n1636 ;
  assign n6057 = ( n397 & ~n416 ) | ( n397 & n3827 ) | ( ~n416 & n3827 ) ;
  assign n6060 = n5005 ^ n3003 ^ x118 ;
  assign n6058 = n5710 ^ n3536 ^ n2552 ;
  assign n6059 = ( ~n1134 & n3087 ) | ( ~n1134 & n6058 ) | ( n3087 & n6058 ) ;
  assign n6061 = n6060 ^ n6059 ^ 1'b0 ;
  assign n6062 = ~n3106 & n6061 ;
  assign n6063 = ( n1228 & n6057 ) | ( n1228 & n6062 ) | ( n6057 & n6062 ) ;
  assign n6084 = ( n1792 & n2697 ) | ( n1792 & n3777 ) | ( n2697 & n3777 ) ;
  assign n6067 = ( n772 & n926 ) | ( n772 & ~n3720 ) | ( n926 & ~n3720 ) ;
  assign n6068 = n1956 & ~n6067 ;
  assign n6069 = n6068 ^ n5333 ^ 1'b0 ;
  assign n6064 = n5458 ^ n2087 ^ 1'b0 ;
  assign n6065 = n1777 | n6064 ;
  assign n6066 = n5107 & ~n6065 ;
  assign n6070 = n6069 ^ n6066 ^ 1'b0 ;
  assign n6072 = n3854 ^ n3372 ^ 1'b0 ;
  assign n6071 = ~n421 & n2809 ;
  assign n6073 = n6072 ^ n6071 ^ n5478 ;
  assign n6076 = n3119 ^ n2373 ^ n1419 ;
  assign n6074 = n458 & n5209 ;
  assign n6075 = n6074 ^ n2274 ^ 1'b0 ;
  assign n6077 = n6076 ^ n6075 ^ n209 ;
  assign n6078 = n6077 ^ n4369 ^ n3841 ;
  assign n6079 = ( n1409 & n4995 ) | ( n1409 & n6078 ) | ( n4995 & n6078 ) ;
  assign n6080 = ( ~n2146 & n5386 ) | ( ~n2146 & n6079 ) | ( n5386 & n6079 ) ;
  assign n6081 = n4013 | n6080 ;
  assign n6082 = n6081 ^ n3734 ^ 1'b0 ;
  assign n6083 = ( n6070 & n6073 ) | ( n6070 & n6082 ) | ( n6073 & n6082 ) ;
  assign n6085 = n6084 ^ n6083 ^ n536 ;
  assign n6086 = n4910 ^ n2178 ^ n1059 ;
  assign n6087 = n2170 ^ n1093 ^ 1'b0 ;
  assign n6088 = n4821 & ~n5173 ;
  assign n6089 = ( n3371 & n4158 ) | ( n3371 & n6088 ) | ( n4158 & n6088 ) ;
  assign n6091 = n1332 ^ n489 ^ 1'b0 ;
  assign n6092 = n6091 ^ n3345 ^ n3154 ;
  assign n6093 = n2650 & n4612 ;
  assign n6094 = n6092 & n6093 ;
  assign n6090 = n4190 ^ n515 ^ x67 ;
  assign n6095 = n6094 ^ n6090 ^ n3487 ;
  assign n6096 = ( n6087 & n6089 ) | ( n6087 & ~n6095 ) | ( n6089 & ~n6095 ) ;
  assign n6097 = n6096 ^ n4136 ^ 1'b0 ;
  assign n6098 = ( n1446 & ~n1469 ) | ( n1446 & n3562 ) | ( ~n1469 & n3562 ) ;
  assign n6099 = n6098 ^ n3594 ^ n1143 ;
  assign n6100 = n6099 ^ n4588 ^ n4371 ;
  assign n6101 = ( n3230 & n5606 ) | ( n3230 & ~n6100 ) | ( n5606 & ~n6100 ) ;
  assign n6102 = n355 & n4598 ;
  assign n6103 = n5474 ^ n1725 ^ n1342 ;
  assign n6104 = ( n139 & n2804 ) | ( n139 & ~n6103 ) | ( n2804 & ~n6103 ) ;
  assign n6105 = n830 | n4458 ;
  assign n6106 = n4413 | n6105 ;
  assign n6107 = ( n6102 & n6104 ) | ( n6102 & n6106 ) | ( n6104 & n6106 ) ;
  assign n6108 = ( n1976 & n6101 ) | ( n1976 & ~n6107 ) | ( n6101 & ~n6107 ) ;
  assign n6109 = ( n1985 & n3251 ) | ( n1985 & ~n6108 ) | ( n3251 & ~n6108 ) ;
  assign n6112 = n1290 | n4711 ;
  assign n6113 = n6112 ^ n3639 ^ 1'b0 ;
  assign n6114 = ~n3522 & n6113 ;
  assign n6110 = n3322 ^ n3198 ^ n1375 ;
  assign n6111 = n6110 ^ n1476 ^ n280 ;
  assign n6115 = n6114 ^ n6111 ^ 1'b0 ;
  assign n6129 = n319 | n932 ;
  assign n6130 = n6129 ^ n233 ^ 1'b0 ;
  assign n6131 = n2821 ^ n1200 ^ 1'b0 ;
  assign n6132 = ( ~n646 & n6130 ) | ( ~n646 & n6131 ) | ( n6130 & n6131 ) ;
  assign n6133 = ( n1516 & ~n3121 ) | ( n1516 & n6132 ) | ( ~n3121 & n6132 ) ;
  assign n6127 = ( n1913 & ~n3641 ) | ( n1913 & n5260 ) | ( ~n3641 & n5260 ) ;
  assign n6128 = ( ~n4115 & n4203 ) | ( ~n4115 & n6127 ) | ( n4203 & n6127 ) ;
  assign n6134 = n6133 ^ n6128 ^ n1069 ;
  assign n6138 = ( ~n3171 & n4406 ) | ( ~n3171 & n5730 ) | ( n4406 & n5730 ) ;
  assign n6137 = n4644 ^ n4262 ^ 1'b0 ;
  assign n6139 = n6138 ^ n6137 ^ x108 ;
  assign n6135 = n2449 ^ x76 ^ 1'b0 ;
  assign n6136 = n4409 & n6135 ;
  assign n6140 = n6139 ^ n6136 ^ 1'b0 ;
  assign n6141 = n6140 ^ n3654 ^ n2385 ;
  assign n6142 = ~n6134 & n6141 ;
  assign n6143 = ~n4688 & n6142 ;
  assign n6118 = x16 & n1084 ;
  assign n6119 = n6118 ^ n2737 ^ 1'b0 ;
  assign n6120 = n6119 ^ n4278 ^ n1582 ;
  assign n6121 = ( n1921 & n2427 ) | ( n1921 & ~n4845 ) | ( n2427 & ~n4845 ) ;
  assign n6122 = n1224 & ~n6121 ;
  assign n6123 = ~n6120 & n6122 ;
  assign n6116 = n1777 ^ n1195 ^ n254 ;
  assign n6117 = n6116 ^ n3588 ^ n3429 ;
  assign n6124 = n6123 ^ n6117 ^ n3477 ;
  assign n6125 = n2073 & n6124 ;
  assign n6126 = n6125 ^ n2495 ^ 1'b0 ;
  assign n6144 = n6143 ^ n6126 ^ n408 ;
  assign n6149 = ( ~n238 & n1044 ) | ( ~n238 & n1051 ) | ( n1044 & n1051 ) ;
  assign n6150 = ( n1298 & n4919 ) | ( n1298 & n6149 ) | ( n4919 & n6149 ) ;
  assign n6145 = n1113 | n5920 ;
  assign n6146 = n6145 ^ n713 ^ 1'b0 ;
  assign n6147 = n6146 ^ n648 ^ 1'b0 ;
  assign n6148 = ( n208 & ~n3205 ) | ( n208 & n6147 ) | ( ~n3205 & n6147 ) ;
  assign n6151 = n6150 ^ n6148 ^ n2950 ;
  assign n6152 = ( n1220 & ~n3171 ) | ( n1220 & n5430 ) | ( ~n3171 & n5430 ) ;
  assign n6153 = n6152 ^ n1912 ^ n1759 ;
  assign n6154 = n3878 ^ n1056 ^ n194 ;
  assign n6155 = ( n2210 & n4473 ) | ( n2210 & ~n6154 ) | ( n4473 & ~n6154 ) ;
  assign n6180 = ~n2749 & n3110 ;
  assign n6166 = ~n1091 & n3573 ;
  assign n6167 = n6166 ^ n1390 ^ 1'b0 ;
  assign n6168 = n6167 ^ n2615 ^ 1'b0 ;
  assign n6169 = n2088 & ~n6168 ;
  assign n6170 = n6169 ^ n2439 ^ n558 ;
  assign n6171 = ( ~n4527 & n4532 ) | ( ~n4527 & n6170 ) | ( n4532 & n6170 ) ;
  assign n6172 = ( ~n2949 & n5424 ) | ( ~n2949 & n6171 ) | ( n5424 & n6171 ) ;
  assign n6173 = ( x39 & n1066 ) | ( x39 & n2242 ) | ( n1066 & n2242 ) ;
  assign n6174 = x116 & n6173 ;
  assign n6175 = n6174 ^ n5468 ^ 1'b0 ;
  assign n6176 = n3796 & ~n4423 ;
  assign n6177 = ~n6175 & n6176 ;
  assign n6178 = n3748 & ~n6177 ;
  assign n6179 = ~n6172 & n6178 ;
  assign n6157 = n5450 ^ n1661 ^ 1'b0 ;
  assign n6158 = ( n1388 & n3568 ) | ( n1388 & ~n6157 ) | ( n3568 & ~n6157 ) ;
  assign n6156 = n3639 ^ n3622 ^ n551 ;
  assign n6159 = n6158 ^ n6156 ^ 1'b0 ;
  assign n6160 = n5969 & ~n6159 ;
  assign n6161 = n6160 ^ n1691 ^ 1'b0 ;
  assign n6162 = ( ~n557 & n776 ) | ( ~n557 & n1978 ) | ( n776 & n1978 ) ;
  assign n6163 = n4081 ^ n3336 ^ 1'b0 ;
  assign n6164 = n6162 | n6163 ;
  assign n6165 = n6161 | n6164 ;
  assign n6181 = n6180 ^ n6179 ^ n6165 ;
  assign n6182 = n5063 ^ n3541 ^ 1'b0 ;
  assign n6183 = n2305 & n2539 ;
  assign n6184 = ( n820 & n1107 ) | ( n820 & n6183 ) | ( n1107 & n6183 ) ;
  assign n6190 = n2720 & n3327 ;
  assign n6186 = n3910 ^ n1675 ^ n270 ;
  assign n6185 = n5419 ^ n1040 ^ n975 ;
  assign n6187 = n6186 ^ n6185 ^ 1'b0 ;
  assign n6188 = ( n2015 & n5919 ) | ( n2015 & n6187 ) | ( n5919 & n6187 ) ;
  assign n6189 = ( x70 & n4388 ) | ( x70 & ~n6188 ) | ( n4388 & ~n6188 ) ;
  assign n6191 = n6190 ^ n6189 ^ n4719 ;
  assign n6192 = ~n6184 & n6191 ;
  assign n6194 = ( n408 & n1479 ) | ( n408 & n1803 ) | ( n1479 & n1803 ) ;
  assign n6193 = ~n488 & n1981 ;
  assign n6195 = n6194 ^ n6193 ^ 1'b0 ;
  assign n6196 = ~n232 & n1161 ;
  assign n6197 = n925 & n6196 ;
  assign n6198 = n4199 ^ n1398 ^ n408 ;
  assign n6199 = ( n449 & n2093 ) | ( n449 & ~n6198 ) | ( n2093 & ~n6198 ) ;
  assign n6200 = ( n5192 & n6197 ) | ( n5192 & n6199 ) | ( n6197 & n6199 ) ;
  assign n6201 = n1055 & ~n2997 ;
  assign n6202 = ~n3240 & n6201 ;
  assign n6203 = n352 & n1465 ;
  assign n6204 = ( n1749 & ~n6202 ) | ( n1749 & n6203 ) | ( ~n6202 & n6203 ) ;
  assign n6205 = n6204 ^ n2191 ^ n1069 ;
  assign n6206 = n2610 ^ n1569 ^ 1'b0 ;
  assign n6207 = n5289 | n6206 ;
  assign n6208 = n572 ^ x72 ^ 1'b0 ;
  assign n6209 = ( n2662 & n3480 ) | ( n2662 & ~n6208 ) | ( n3480 & ~n6208 ) ;
  assign n6211 = ( ~n197 & n1412 ) | ( ~n197 & n1932 ) | ( n1412 & n1932 ) ;
  assign n6210 = ( n233 & ~n611 ) | ( n233 & n2480 ) | ( ~n611 & n2480 ) ;
  assign n6212 = n6211 ^ n6210 ^ n1103 ;
  assign n6213 = n6209 & n6212 ;
  assign n6221 = ( n773 & n943 ) | ( n773 & ~n1894 ) | ( n943 & ~n1894 ) ;
  assign n6220 = n3025 ^ n2058 ^ n1940 ;
  assign n6216 = n3053 ^ n1813 ^ n319 ;
  assign n6217 = n1209 & ~n6216 ;
  assign n6218 = n6217 ^ n4684 ^ 1'b0 ;
  assign n6214 = n3574 ^ n1058 ^ n919 ;
  assign n6215 = ( n3639 & ~n4121 ) | ( n3639 & n6214 ) | ( ~n4121 & n6214 ) ;
  assign n6219 = n6218 ^ n6215 ^ n5392 ;
  assign n6222 = n6221 ^ n6220 ^ n6219 ;
  assign n6223 = n818 & n3626 ;
  assign n6224 = n6223 ^ n3593 ^ 1'b0 ;
  assign n6225 = n1473 | n6224 ;
  assign n6226 = n1294 & n1419 ;
  assign n6227 = ( n2868 & n4764 ) | ( n2868 & ~n5307 ) | ( n4764 & ~n5307 ) ;
  assign n6228 = n6227 ^ n4400 ^ n460 ;
  assign n6229 = ( n416 & n1045 ) | ( n416 & n1617 ) | ( n1045 & n1617 ) ;
  assign n6230 = n6229 ^ n6029 ^ n577 ;
  assign n6231 = n5234 ^ n2268 ^ n733 ;
  assign n6232 = ( n3617 & ~n3660 ) | ( n3617 & n6231 ) | ( ~n3660 & n6231 ) ;
  assign n6233 = ( n6228 & ~n6230 ) | ( n6228 & n6232 ) | ( ~n6230 & n6232 ) ;
  assign n6234 = ( x96 & n1065 ) | ( x96 & ~n6233 ) | ( n1065 & ~n6233 ) ;
  assign n6235 = n6226 & ~n6234 ;
  assign n6236 = n6225 & n6235 ;
  assign n6237 = n2971 & ~n6236 ;
  assign n6238 = n6237 ^ n1810 ^ 1'b0 ;
  assign n6239 = ( n530 & n5288 ) | ( n530 & ~n5956 ) | ( n5288 & ~n5956 ) ;
  assign n6240 = ( ~x49 & n857 ) | ( ~x49 & n6239 ) | ( n857 & n6239 ) ;
  assign n6241 = ( n1076 & n1508 ) | ( n1076 & ~n2819 ) | ( n1508 & ~n2819 ) ;
  assign n6242 = ( ~n187 & n4636 ) | ( ~n187 & n6241 ) | ( n4636 & n6241 ) ;
  assign n6243 = n2281 & ~n3389 ;
  assign n6244 = ~n5244 & n6243 ;
  assign n6245 = n6244 ^ n4285 ^ 1'b0 ;
  assign n6246 = ~n3655 & n6245 ;
  assign n6247 = n6246 ^ n993 ^ 1'b0 ;
  assign n6248 = ( n336 & n3478 ) | ( n336 & ~n6247 ) | ( n3478 & ~n6247 ) ;
  assign n6249 = ~n1053 & n1437 ;
  assign n6250 = ( ~n5045 & n5459 ) | ( ~n5045 & n6249 ) | ( n5459 & n6249 ) ;
  assign n6251 = n2519 ^ n408 ^ 1'b0 ;
  assign n6252 = ( n582 & ~n1095 ) | ( n582 & n1505 ) | ( ~n1095 & n1505 ) ;
  assign n6253 = n6252 ^ n4541 ^ 1'b0 ;
  assign n6254 = n2345 & n3845 ;
  assign n6255 = n6254 ^ n2050 ^ 1'b0 ;
  assign n6256 = ( n6251 & ~n6253 ) | ( n6251 & n6255 ) | ( ~n6253 & n6255 ) ;
  assign n6257 = n6256 ^ n2901 ^ 1'b0 ;
  assign n6258 = ( n1735 & n5031 ) | ( n1735 & ~n6230 ) | ( n5031 & ~n6230 ) ;
  assign n6259 = n5311 ^ n3744 ^ 1'b0 ;
  assign n6260 = ~n1584 & n6259 ;
  assign n6261 = n5026 ^ n2328 ^ n1923 ;
  assign n6262 = ( n1122 & ~n1186 ) | ( n1122 & n6261 ) | ( ~n1186 & n6261 ) ;
  assign n6263 = n6262 ^ n4695 ^ 1'b0 ;
  assign n6264 = n3118 | n6263 ;
  assign n6265 = ( ~n4196 & n6260 ) | ( ~n4196 & n6264 ) | ( n6260 & n6264 ) ;
  assign n6266 = x119 & ~n353 ;
  assign n6267 = n6266 ^ n334 ^ 1'b0 ;
  assign n6268 = ( n188 & n1708 ) | ( n188 & n6267 ) | ( n1708 & n6267 ) ;
  assign n6269 = n6268 ^ n326 ^ 1'b0 ;
  assign n6270 = n2378 & n6269 ;
  assign n6271 = n6270 ^ n3295 ^ n2456 ;
  assign n6272 = ( x57 & n6265 ) | ( x57 & n6271 ) | ( n6265 & n6271 ) ;
  assign n6273 = ( n285 & n2659 ) | ( n285 & n3943 ) | ( n2659 & n3943 ) ;
  assign n6274 = n6273 ^ n5578 ^ n358 ;
  assign n6284 = ~n1299 & n1367 ;
  assign n6285 = n6284 ^ n1585 ^ 1'b0 ;
  assign n6283 = ( n688 & ~n2397 ) | ( n688 & n2636 ) | ( ~n2397 & n2636 ) ;
  assign n6286 = n6285 ^ n6283 ^ 1'b0 ;
  assign n6287 = ~n2272 & n6286 ;
  assign n6280 = ( n3427 & ~n3495 ) | ( n3427 & n3882 ) | ( ~n3495 & n3882 ) ;
  assign n6281 = n6280 ^ n2927 ^ 1'b0 ;
  assign n6282 = ~n2901 & n6281 ;
  assign n6275 = n5668 ^ n2066 ^ 1'b0 ;
  assign n6276 = n4653 & n6275 ;
  assign n6277 = ~n289 & n6276 ;
  assign n6278 = n6277 ^ n146 ^ 1'b0 ;
  assign n6279 = ~n3449 & n6278 ;
  assign n6288 = n6287 ^ n6282 ^ n6279 ;
  assign n6289 = n1164 ^ n320 ^ 1'b0 ;
  assign n6290 = n2049 & ~n6289 ;
  assign n6291 = ( n2193 & n4006 ) | ( n2193 & ~n6290 ) | ( n4006 & ~n6290 ) ;
  assign n6292 = n6291 ^ n2448 ^ n2089 ;
  assign n6293 = x93 & n3400 ;
  assign n6294 = n6292 & n6293 ;
  assign n6295 = n2989 ^ n423 ^ 1'b0 ;
  assign n6296 = n2902 ^ n1069 ^ 1'b0 ;
  assign n6297 = n2698 | n6296 ;
  assign n6298 = n6297 ^ n5730 ^ n4623 ;
  assign n6299 = ( ~x13 & n2715 ) | ( ~x13 & n4513 ) | ( n2715 & n4513 ) ;
  assign n6307 = n2606 & ~n2716 ;
  assign n6308 = n6307 ^ n597 ^ 1'b0 ;
  assign n6309 = ( n808 & ~n1796 ) | ( n808 & n2142 ) | ( ~n1796 & n2142 ) ;
  assign n6310 = ( n1189 & n6308 ) | ( n1189 & n6309 ) | ( n6308 & n6309 ) ;
  assign n6311 = n2980 | n6310 ;
  assign n6312 = n6311 ^ n5510 ^ 1'b0 ;
  assign n6313 = n6312 ^ n3522 ^ n3091 ;
  assign n6305 = n5803 & ~n6277 ;
  assign n6306 = n6305 ^ n3733 ^ 1'b0 ;
  assign n6314 = n6313 ^ n6306 ^ n2386 ;
  assign n6300 = n6251 ^ n1863 ^ 1'b0 ;
  assign n6301 = n3086 & ~n6300 ;
  assign n6302 = n6156 ^ n5183 ^ n3164 ;
  assign n6303 = ( n3156 & n6301 ) | ( n3156 & n6302 ) | ( n6301 & n6302 ) ;
  assign n6304 = n168 & n6303 ;
  assign n6315 = n6314 ^ n6304 ^ 1'b0 ;
  assign n6316 = ( n3269 & n6299 ) | ( n3269 & ~n6315 ) | ( n6299 & ~n6315 ) ;
  assign n6317 = n6315 ^ n5207 ^ n5160 ;
  assign n6318 = ( x123 & n2376 ) | ( x123 & n3884 ) | ( n2376 & n3884 ) ;
  assign n6319 = n4214 ^ n2412 ^ 1'b0 ;
  assign n6320 = n2137 & n6319 ;
  assign n6321 = ~n4456 & n6320 ;
  assign n6322 = n3193 ^ n1017 ^ n130 ;
  assign n6323 = ( n956 & n1026 ) | ( n956 & ~n5419 ) | ( n1026 & ~n5419 ) ;
  assign n6324 = n6322 | n6323 ;
  assign n6325 = n144 | n6324 ;
  assign n6326 = n5908 ^ n2806 ^ n528 ;
  assign n6327 = n829 & n6326 ;
  assign n6328 = n186 & ~n4296 ;
  assign n6329 = n6327 & n6328 ;
  assign n6330 = n2728 ^ n309 ^ 1'b0 ;
  assign n6331 = ( ~n3920 & n4468 ) | ( ~n3920 & n6330 ) | ( n4468 & n6330 ) ;
  assign n6332 = ( n6325 & n6329 ) | ( n6325 & n6331 ) | ( n6329 & n6331 ) ;
  assign n6335 = ~x43 & n323 ;
  assign n6336 = ( x99 & ~n1216 ) | ( x99 & n2719 ) | ( ~n1216 & n2719 ) ;
  assign n6337 = ( ~n2770 & n2955 ) | ( ~n2770 & n6336 ) | ( n2955 & n6336 ) ;
  assign n6338 = ( n496 & n6335 ) | ( n496 & n6337 ) | ( n6335 & n6337 ) ;
  assign n6333 = n2985 ^ n1693 ^ 1'b0 ;
  assign n6334 = n4185 & n6333 ;
  assign n6339 = n6338 ^ n6334 ^ 1'b0 ;
  assign n6340 = n549 & ~n1119 ;
  assign n6341 = ( n412 & n1214 ) | ( n412 & ~n6340 ) | ( n1214 & ~n6340 ) ;
  assign n6342 = n6341 ^ n2445 ^ 1'b0 ;
  assign n6343 = n2855 & ~n6342 ;
  assign n6344 = n1873 & ~n3400 ;
  assign n6345 = ( ~n1641 & n2757 ) | ( ~n1641 & n6344 ) | ( n2757 & n6344 ) ;
  assign n6346 = ( n4211 & n6343 ) | ( n4211 & ~n6345 ) | ( n6343 & ~n6345 ) ;
  assign n6347 = n214 | n4660 ;
  assign n6348 = n6347 ^ n5791 ^ 1'b0 ;
  assign n6349 = n4323 ^ n4004 ^ n2392 ;
  assign n6350 = n2856 & n4655 ;
  assign n6351 = n6350 ^ n5507 ^ n909 ;
  assign n6352 = ( n4390 & ~n6349 ) | ( n4390 & n6351 ) | ( ~n6349 & n6351 ) ;
  assign n6362 = x52 & ~n309 ;
  assign n6363 = n6362 ^ n3297 ^ 1'b0 ;
  assign n6357 = n2183 ^ n1334 ^ n1258 ;
  assign n6358 = ( ~n585 & n5204 ) | ( ~n585 & n6357 ) | ( n5204 & n6357 ) ;
  assign n6359 = n6358 ^ n959 ^ 1'b0 ;
  assign n6360 = n5012 | n6359 ;
  assign n6361 = n6360 ^ n3631 ^ n1265 ;
  assign n6353 = n1548 | n4087 ;
  assign n6354 = n6353 ^ n3878 ^ 1'b0 ;
  assign n6355 = ~n6293 & n6354 ;
  assign n6356 = ~n2160 & n6355 ;
  assign n6364 = n6363 ^ n6361 ^ n6356 ;
  assign n6365 = n2769 ^ n2544 ^ n1211 ;
  assign n6366 = n6365 ^ n1774 ^ x11 ;
  assign n6367 = n6366 ^ n4695 ^ n2691 ;
  assign n6368 = n4705 ^ n258 ^ 1'b0 ;
  assign n6373 = n654 & ~n1041 ;
  assign n6370 = n3873 ^ n3082 ^ n1120 ;
  assign n6369 = n6340 ^ n4731 ^ n730 ;
  assign n6371 = n6370 ^ n6369 ^ n3178 ;
  assign n6372 = ( n1649 & n2033 ) | ( n1649 & ~n6371 ) | ( n2033 & ~n6371 ) ;
  assign n6374 = n6373 ^ n6372 ^ n2412 ;
  assign n6375 = ( n6367 & n6368 ) | ( n6367 & n6374 ) | ( n6368 & n6374 ) ;
  assign n6376 = ~n4029 & n6120 ;
  assign n6377 = n6376 ^ n786 ^ 1'b0 ;
  assign n6378 = n292 | n2601 ;
  assign n6379 = ( n3130 & ~n4461 ) | ( n3130 & n6378 ) | ( ~n4461 & n6378 ) ;
  assign n6380 = ~n3222 & n6379 ;
  assign n6386 = ( ~n4144 & n5657 ) | ( ~n4144 & n5681 ) | ( n5657 & n5681 ) ;
  assign n6382 = ( n1467 & ~n2619 ) | ( n1467 & n2697 ) | ( ~n2619 & n2697 ) ;
  assign n6383 = n3979 ^ n908 ^ 1'b0 ;
  assign n6384 = ( n5828 & n6382 ) | ( n5828 & ~n6383 ) | ( n6382 & ~n6383 ) ;
  assign n6381 = n2178 & ~n2521 ;
  assign n6385 = n6384 ^ n6381 ^ 1'b0 ;
  assign n6387 = n6386 ^ n6385 ^ n375 ;
  assign n6390 = n5247 ^ n3025 ^ n1682 ;
  assign n6391 = ( ~n2285 & n5613 ) | ( ~n2285 & n6390 ) | ( n5613 & n6390 ) ;
  assign n6388 = n5073 ^ n2663 ^ 1'b0 ;
  assign n6389 = x81 & n6388 ;
  assign n6392 = n6391 ^ n6389 ^ 1'b0 ;
  assign n6393 = n4419 ^ n1462 ^ n702 ;
  assign n6394 = n913 & n6393 ;
  assign n6395 = n6394 ^ n345 ^ 1'b0 ;
  assign n6396 = n3243 ^ n2910 ^ n1064 ;
  assign n6397 = ( n1492 & n2356 ) | ( n1492 & n2965 ) | ( n2356 & n2965 ) ;
  assign n6398 = ( n520 & n6396 ) | ( n520 & n6397 ) | ( n6396 & n6397 ) ;
  assign n6401 = n1178 | n5358 ;
  assign n6402 = ( n532 & n4410 ) | ( n532 & n6401 ) | ( n4410 & n6401 ) ;
  assign n6399 = n2496 & ~n2806 ;
  assign n6400 = n6399 ^ n2123 ^ 1'b0 ;
  assign n6403 = n6402 ^ n6400 ^ n2083 ;
  assign n6404 = n6182 ^ n2701 ^ n1704 ;
  assign n6406 = ( n1026 & n1076 ) | ( n1026 & ~n1431 ) | ( n1076 & ~n1431 ) ;
  assign n6405 = ( n1079 & n1243 ) | ( n1079 & ~n2314 ) | ( n1243 & ~n2314 ) ;
  assign n6407 = n6406 ^ n6405 ^ n2206 ;
  assign n6408 = ( n1064 & ~n4695 ) | ( n1064 & n6407 ) | ( ~n4695 & n6407 ) ;
  assign n6409 = n4154 ^ n1179 ^ 1'b0 ;
  assign n6410 = n5682 | n6409 ;
  assign n6419 = ( ~n2425 & n2437 ) | ( ~n2425 & n3642 ) | ( n2437 & n3642 ) ;
  assign n6418 = n5529 ^ n3104 ^ n464 ;
  assign n6414 = n1030 ^ n1028 ^ n603 ;
  assign n6415 = ( n3868 & n4812 ) | ( n3868 & n6414 ) | ( n4812 & n6414 ) ;
  assign n6416 = ( n3008 & n3714 ) | ( n3008 & n6415 ) | ( n3714 & n6415 ) ;
  assign n6411 = n1479 ^ x75 ^ 1'b0 ;
  assign n6412 = ( x127 & n1180 ) | ( x127 & n6411 ) | ( n1180 & n6411 ) ;
  assign n6413 = n6412 ^ n2563 ^ 1'b0 ;
  assign n6417 = n6416 ^ n6413 ^ n2771 ;
  assign n6420 = n6419 ^ n6418 ^ n6417 ;
  assign n6421 = n6310 ^ n3168 ^ n521 ;
  assign n6422 = ( x49 & n3160 ) | ( x49 & ~n4918 ) | ( n3160 & ~n4918 ) ;
  assign n6423 = n1614 & ~n6422 ;
  assign n6424 = ( ~n1932 & n6421 ) | ( ~n1932 & n6423 ) | ( n6421 & n6423 ) ;
  assign n6429 = n3126 ^ n2659 ^ n148 ;
  assign n6430 = ( n2953 & ~n3423 ) | ( n2953 & n6429 ) | ( ~n3423 & n6429 ) ;
  assign n6425 = n4908 ^ n3890 ^ n1079 ;
  assign n6426 = n2485 ^ n2058 ^ n999 ;
  assign n6427 = n6426 ^ n2190 ^ n917 ;
  assign n6428 = n6425 & ~n6427 ;
  assign n6431 = n6430 ^ n6428 ^ 1'b0 ;
  assign n6432 = ( ~n2705 & n3803 ) | ( ~n2705 & n5803 ) | ( n3803 & n5803 ) ;
  assign n6440 = n2499 ^ n1076 ^ n983 ;
  assign n6438 = ( n188 & n1280 ) | ( n188 & ~n4861 ) | ( n1280 & ~n4861 ) ;
  assign n6434 = n4626 ^ n3451 ^ 1'b0 ;
  assign n6435 = n1322 | n6434 ;
  assign n6436 = n2981 ^ n529 ^ 1'b0 ;
  assign n6437 = n6435 | n6436 ;
  assign n6439 = n6438 ^ n6437 ^ n3613 ;
  assign n6441 = n6440 ^ n6439 ^ n1422 ;
  assign n6433 = ( n3782 & n5624 ) | ( n3782 & ~n6127 ) | ( n5624 & ~n6127 ) ;
  assign n6442 = n6441 ^ n6433 ^ n5939 ;
  assign n6443 = n6244 ^ n3997 ^ 1'b0 ;
  assign n6444 = n6443 ^ n6372 ^ n1621 ;
  assign n6453 = x80 & ~n1182 ;
  assign n6454 = ~n829 & n6453 ;
  assign n6448 = n1895 ^ n649 ^ 1'b0 ;
  assign n6449 = n1750 | n6448 ;
  assign n6450 = n6449 ^ n4817 ^ n2061 ;
  assign n6451 = n6450 ^ n6405 ^ x0 ;
  assign n6452 = n908 & ~n6451 ;
  assign n6455 = n6454 ^ n6452 ^ 1'b0 ;
  assign n6447 = n4303 ^ n1488 ^ n1138 ;
  assign n6456 = n6455 ^ n6447 ^ n3992 ;
  assign n6445 = ~n4261 & n4856 ;
  assign n6446 = n6445 ^ n4494 ^ 1'b0 ;
  assign n6457 = n6456 ^ n6446 ^ n5557 ;
  assign n6458 = n391 & n3635 ;
  assign n6459 = ~x61 & n6458 ;
  assign n6460 = n6459 ^ n511 ^ 1'b0 ;
  assign n6461 = n5930 ^ n1469 ^ 1'b0 ;
  assign n6462 = n6460 | n6461 ;
  assign n6463 = n5531 ^ n1597 ^ 1'b0 ;
  assign n6464 = n1430 & ~n3777 ;
  assign n6465 = n6464 ^ n3694 ^ n1068 ;
  assign n6466 = ( n940 & n2629 ) | ( n940 & ~n6465 ) | ( n2629 & ~n6465 ) ;
  assign n6467 = ( n2676 & n4707 ) | ( n2676 & n6466 ) | ( n4707 & n6466 ) ;
  assign n6468 = ( ~n4659 & n6029 ) | ( ~n4659 & n6467 ) | ( n6029 & n6467 ) ;
  assign n6470 = ( n3304 & ~n4325 ) | ( n3304 & n5088 ) | ( ~n4325 & n5088 ) ;
  assign n6471 = n3015 ^ n628 ^ n472 ;
  assign n6472 = n6471 ^ n2046 ^ 1'b0 ;
  assign n6473 = n6470 & n6472 ;
  assign n6469 = n4770 ^ n2537 ^ n1141 ;
  assign n6474 = n6473 ^ n6469 ^ n2262 ;
  assign n6475 = n3896 ^ n1848 ^ n712 ;
  assign n6476 = ( n855 & n4210 ) | ( n855 & n6475 ) | ( n4210 & n6475 ) ;
  assign n6477 = n6358 ^ n2956 ^ 1'b0 ;
  assign n6478 = ( x52 & n1056 ) | ( x52 & n2047 ) | ( n1056 & n2047 ) ;
  assign n6479 = n3325 ^ n2552 ^ n862 ;
  assign n6480 = n3243 ^ n970 ^ 1'b0 ;
  assign n6481 = ( n1153 & n6479 ) | ( n1153 & ~n6480 ) | ( n6479 & ~n6480 ) ;
  assign n6482 = ( n2110 & n4960 ) | ( n2110 & n6481 ) | ( n4960 & n6481 ) ;
  assign n6483 = ( n2609 & ~n6478 ) | ( n2609 & n6482 ) | ( ~n6478 & n6482 ) ;
  assign n6484 = n5917 ^ n5244 ^ n1586 ;
  assign n6485 = n448 & n3430 ;
  assign n6486 = n6485 ^ n2979 ^ 1'b0 ;
  assign n6487 = x24 & n6486 ;
  assign n6488 = n6487 ^ n2801 ^ 1'b0 ;
  assign n6489 = n4433 ^ n4132 ^ n2189 ;
  assign n6490 = n6489 ^ n3852 ^ n2061 ;
  assign n6491 = n2084 | n4260 ;
  assign n6492 = n3035 & ~n6491 ;
  assign n6493 = n6492 ^ n5744 ^ n4037 ;
  assign n6494 = ( ~n5155 & n6490 ) | ( ~n5155 & n6493 ) | ( n6490 & n6493 ) ;
  assign n6495 = n5017 ^ n529 ^ n255 ;
  assign n6496 = ~n2573 & n2604 ;
  assign n6497 = n6495 & n6496 ;
  assign n6504 = n168 & n6268 ;
  assign n6505 = n6504 ^ n981 ^ 1'b0 ;
  assign n6500 = n4116 ^ n3707 ^ n264 ;
  assign n6501 = n6473 ^ n3449 ^ n437 ;
  assign n6502 = ( n1242 & n6500 ) | ( n1242 & n6501 ) | ( n6500 & n6501 ) ;
  assign n6498 = n5332 ^ n4950 ^ n2626 ;
  assign n6499 = n6498 ^ n2082 ^ n516 ;
  assign n6503 = n6502 ^ n6499 ^ n3880 ;
  assign n6506 = n6505 ^ n6503 ^ n2393 ;
  assign n6508 = n5859 ^ n3635 ^ n1168 ;
  assign n6507 = ( n559 & ~n2502 ) | ( n559 & n3025 ) | ( ~n2502 & n3025 ) ;
  assign n6509 = n6508 ^ n6507 ^ n4791 ;
  assign n6510 = n1346 & n6267 ;
  assign n6511 = n6510 ^ n5096 ^ n130 ;
  assign n6512 = n6511 ^ n5317 ^ n3084 ;
  assign n6514 = n2724 ^ n928 ^ 1'b0 ;
  assign n6515 = n6190 ^ n2849 ^ n478 ;
  assign n6516 = ( n668 & n1598 ) | ( n668 & ~n2858 ) | ( n1598 & ~n2858 ) ;
  assign n6517 = ( n1834 & ~n4732 ) | ( n1834 & n6516 ) | ( ~n4732 & n6516 ) ;
  assign n6518 = ( ~n948 & n6515 ) | ( ~n948 & n6517 ) | ( n6515 & n6517 ) ;
  assign n6519 = ( n5799 & n6514 ) | ( n5799 & n6518 ) | ( n6514 & n6518 ) ;
  assign n6513 = n314 & n4210 ;
  assign n6520 = n6519 ^ n6513 ^ 1'b0 ;
  assign n6521 = ~n731 & n1196 ;
  assign n6522 = n4341 & n6030 ;
  assign n6523 = n6521 & n6522 ;
  assign n6524 = ( n1232 & ~n4510 ) | ( n1232 & n6523 ) | ( ~n4510 & n6523 ) ;
  assign n6532 = n3704 | n6100 ;
  assign n6529 = ( n377 & n1191 ) | ( n377 & ~n1214 ) | ( n1191 & ~n1214 ) ;
  assign n6530 = n6529 ^ n2556 ^ n1065 ;
  assign n6525 = ~n397 & n5210 ;
  assign n6526 = ( n1510 & n2812 ) | ( n1510 & n6525 ) | ( n2812 & n6525 ) ;
  assign n6527 = n6526 ^ n2276 ^ n834 ;
  assign n6528 = n6527 ^ n2955 ^ x69 ;
  assign n6531 = n6530 ^ n6528 ^ n5974 ;
  assign n6533 = n6532 ^ n6531 ^ n4107 ;
  assign n6534 = n670 & n2390 ;
  assign n6535 = n1093 & n1867 ;
  assign n6536 = ( n4655 & n5668 ) | ( n4655 & n6535 ) | ( n5668 & n6535 ) ;
  assign n6537 = ~n340 & n3576 ;
  assign n6538 = ~n6536 & n6537 ;
  assign n6539 = ( ~n713 & n6534 ) | ( ~n713 & n6538 ) | ( n6534 & n6538 ) ;
  assign n6540 = n2618 ^ n2593 ^ 1'b0 ;
  assign n6541 = ( n1191 & n3873 ) | ( n1191 & ~n6540 ) | ( n3873 & ~n6540 ) ;
  assign n6542 = n5581 ^ n3449 ^ n3221 ;
  assign n6543 = ( ~x71 & n6541 ) | ( ~x71 & n6542 ) | ( n6541 & n6542 ) ;
  assign n6544 = ( x64 & n4101 ) | ( x64 & n5334 ) | ( n4101 & n5334 ) ;
  assign n6545 = ( ~n1400 & n2064 ) | ( ~n1400 & n5709 ) | ( n2064 & n5709 ) ;
  assign n6546 = n6545 ^ n3583 ^ n1499 ;
  assign n6547 = ( n3020 & n4574 ) | ( n3020 & n6546 ) | ( n4574 & n6546 ) ;
  assign n6548 = ( n247 & ~n605 ) | ( n247 & n998 ) | ( ~n605 & n998 ) ;
  assign n6553 = ( ~n1830 & n2607 ) | ( ~n1830 & n3189 ) | ( n2607 & n3189 ) ;
  assign n6549 = n2022 & n2577 ;
  assign n6550 = n1852 & n6549 ;
  assign n6551 = n6550 ^ n5162 ^ n3998 ;
  assign n6552 = n6551 ^ n4039 ^ n2483 ;
  assign n6554 = n6553 ^ n6552 ^ 1'b0 ;
  assign n6555 = ( ~n1206 & n6548 ) | ( ~n1206 & n6554 ) | ( n6548 & n6554 ) ;
  assign n6559 = n6407 ^ n2386 ^ n1005 ;
  assign n6560 = ( n167 & n4898 ) | ( n167 & n6559 ) | ( n4898 & n6559 ) ;
  assign n6556 = ( ~n1308 & n3603 ) | ( ~n1308 & n4934 ) | ( n3603 & n4934 ) ;
  assign n6557 = ( n1521 & n5392 ) | ( n1521 & n6556 ) | ( n5392 & n6556 ) ;
  assign n6558 = n6557 ^ n2821 ^ n661 ;
  assign n6561 = n6560 ^ n6558 ^ n4597 ;
  assign n6562 = n3005 ^ n2692 ^ n1908 ;
  assign n6563 = ( n1652 & n4473 ) | ( n1652 & ~n6562 ) | ( n4473 & ~n6562 ) ;
  assign n6564 = n5439 ^ n4710 ^ n3593 ;
  assign n6565 = ( n4755 & n4882 ) | ( n4755 & ~n5271 ) | ( n4882 & ~n5271 ) ;
  assign n6566 = n3375 ^ n2878 ^ n1791 ;
  assign n6567 = ( n5311 & ~n6553 ) | ( n5311 & n6566 ) | ( ~n6553 & n6566 ) ;
  assign n6568 = n4855 ^ n762 ^ 1'b0 ;
  assign n6569 = n6568 ^ n2138 ^ n1719 ;
  assign n6572 = ( n1282 & n1698 ) | ( n1282 & ~n1972 ) | ( n1698 & ~n1972 ) ;
  assign n6573 = n6572 ^ n4254 ^ n691 ;
  assign n6574 = n3980 ^ n754 ^ 1'b0 ;
  assign n6575 = ~n1072 & n6574 ;
  assign n6576 = ( n3832 & n6573 ) | ( n3832 & n6575 ) | ( n6573 & n6575 ) ;
  assign n6570 = ( n646 & ~n5285 ) | ( n646 & n5814 ) | ( ~n5285 & n5814 ) ;
  assign n6571 = ( n2616 & ~n3319 ) | ( n2616 & n6570 ) | ( ~n3319 & n6570 ) ;
  assign n6577 = n6576 ^ n6571 ^ 1'b0 ;
  assign n6578 = ( n6567 & n6569 ) | ( n6567 & ~n6577 ) | ( n6569 & ~n6577 ) ;
  assign n6591 = n3665 ^ n2485 ^ n844 ;
  assign n6589 = n3423 & ~n5993 ;
  assign n6590 = n6589 ^ n2809 ^ 1'b0 ;
  assign n6586 = ( n591 & n1419 ) | ( n591 & n4134 ) | ( n1419 & n4134 ) ;
  assign n6587 = n6586 ^ n5163 ^ n3522 ;
  assign n6585 = x67 & ~n3308 ;
  assign n6588 = n6587 ^ n6585 ^ 1'b0 ;
  assign n6592 = n6591 ^ n6590 ^ n6588 ;
  assign n6579 = n6231 ^ n4096 ^ n2777 ;
  assign n6580 = n1813 | n6579 ;
  assign n6581 = ~n351 & n1433 ;
  assign n6582 = n6581 ^ n2723 ^ n2701 ;
  assign n6583 = n6582 ^ n6270 ^ n5049 ;
  assign n6584 = n6580 & ~n6583 ;
  assign n6593 = n6592 ^ n6584 ^ 1'b0 ;
  assign n6596 = n2562 & n4914 ;
  assign n6597 = n6596 ^ n152 ^ 1'b0 ;
  assign n6594 = n2096 ^ n749 ^ n353 ;
  assign n6595 = ( n196 & ~n5283 ) | ( n196 & n6594 ) | ( ~n5283 & n6594 ) ;
  assign n6598 = n6597 ^ n6595 ^ 1'b0 ;
  assign n6600 = n4389 ^ n1453 ^ x15 ;
  assign n6599 = ~n2190 & n3536 ;
  assign n6601 = n6600 ^ n6599 ^ 1'b0 ;
  assign n6602 = n2354 ^ n605 ^ 1'b0 ;
  assign n6603 = n6601 | n6602 ;
  assign n6604 = ( ~n3483 & n5377 ) | ( ~n3483 & n6603 ) | ( n5377 & n6603 ) ;
  assign n6605 = n1344 & n4723 ;
  assign n6606 = n5871 & n6605 ;
  assign n6607 = x29 & x85 ;
  assign n6608 = ~n936 & n6607 ;
  assign n6609 = n5310 & ~n6608 ;
  assign n6610 = n6609 ^ n5392 ^ n4166 ;
  assign n6611 = n5319 ^ n2853 ^ n2289 ;
  assign n6612 = n6611 ^ n2390 ^ n1194 ;
  assign n6613 = n4246 ^ n222 ^ 1'b0 ;
  assign n6614 = n6613 ^ n2452 ^ n2426 ;
  assign n6615 = n3728 & ~n3954 ;
  assign n6616 = ( n1609 & n4488 ) | ( n1609 & ~n6615 ) | ( n4488 & ~n6615 ) ;
  assign n6617 = ( x64 & n2420 ) | ( x64 & ~n6616 ) | ( n2420 & ~n6616 ) ;
  assign n6618 = n6617 ^ n937 ^ 1'b0 ;
  assign n6619 = n589 & n6618 ;
  assign n6620 = n6614 & n6619 ;
  assign n6621 = n4919 ^ n1721 ^ n1296 ;
  assign n6622 = n6621 ^ n2305 ^ 1'b0 ;
  assign n6625 = x81 & x111 ;
  assign n6626 = n6625 ^ n1957 ^ 1'b0 ;
  assign n6627 = n3337 & ~n6626 ;
  assign n6623 = n2686 ^ n2650 ^ n803 ;
  assign n6624 = ( n3682 & ~n4443 ) | ( n3682 & n6623 ) | ( ~n4443 & n6623 ) ;
  assign n6628 = n6627 ^ n6624 ^ n931 ;
  assign n6629 = n4108 ^ n3564 ^ 1'b0 ;
  assign n6630 = n1402 & ~n6629 ;
  assign n6631 = n6630 ^ x107 ^ 1'b0 ;
  assign n6632 = n1922 & n6631 ;
  assign n6633 = n6579 ^ n5961 ^ n2813 ;
  assign n6634 = n3895 ^ n2725 ^ n239 ;
  assign n6635 = n4535 ^ n4474 ^ 1'b0 ;
  assign n6636 = n1320 ^ n858 ^ n243 ;
  assign n6637 = n6636 ^ n3137 ^ n2051 ;
  assign n6638 = ~n2112 & n2493 ;
  assign n6639 = n6638 ^ n1834 ^ 1'b0 ;
  assign n6640 = n6639 ^ n2985 ^ n242 ;
  assign n6641 = ( n6175 & ~n6637 ) | ( n6175 & n6640 ) | ( ~n6637 & n6640 ) ;
  assign n6642 = ( n659 & ~n2338 ) | ( n659 & n4038 ) | ( ~n2338 & n4038 ) ;
  assign n6643 = ( ~n6635 & n6641 ) | ( ~n6635 & n6642 ) | ( n6641 & n6642 ) ;
  assign n6644 = n2973 ^ n2636 ^ 1'b0 ;
  assign n6645 = ~n1661 & n6644 ;
  assign n6646 = n3610 | n6645 ;
  assign n6647 = n6646 ^ n4202 ^ n2157 ;
  assign n6648 = n2546 ^ n1363 ^ 1'b0 ;
  assign n6649 = n1721 & ~n6648 ;
  assign n6650 = n3346 & ~n6218 ;
  assign n6651 = ( ~n373 & n6649 ) | ( ~n373 & n6650 ) | ( n6649 & n6650 ) ;
  assign n6652 = ( n2489 & ~n3993 ) | ( n2489 & n6651 ) | ( ~n3993 & n6651 ) ;
  assign n6655 = n1431 ^ n900 ^ n702 ;
  assign n6653 = n1972 ^ n1854 ^ x5 ;
  assign n6654 = n6653 ^ n1574 ^ 1'b0 ;
  assign n6656 = n6655 ^ n6654 ^ 1'b0 ;
  assign n6657 = n1351 & n2079 ;
  assign n6658 = ( n413 & ~n1507 ) | ( n413 & n4178 ) | ( ~n1507 & n4178 ) ;
  assign n6659 = n1377 & n5346 ;
  assign n6660 = n6659 ^ n1747 ^ n182 ;
  assign n6661 = ( ~n6657 & n6658 ) | ( ~n6657 & n6660 ) | ( n6658 & n6660 ) ;
  assign n6662 = n5109 & ~n6661 ;
  assign n6663 = n6662 ^ n6261 ^ n4057 ;
  assign n6664 = n202 & ~n2131 ;
  assign n6668 = ( ~n306 & n1924 ) | ( ~n306 & n2189 ) | ( n1924 & n2189 ) ;
  assign n6666 = n363 | n2054 ;
  assign n6667 = n4604 | n6666 ;
  assign n6665 = n4489 ^ n2686 ^ n1987 ;
  assign n6669 = n6668 ^ n6667 ^ n6665 ;
  assign n6670 = n4976 ^ n1413 ^ n605 ;
  assign n6671 = n4600 & ~n6670 ;
  assign n6672 = n6671 ^ n3907 ^ n3847 ;
  assign n6673 = ( n917 & ~n4327 ) | ( n917 & n6672 ) | ( ~n4327 & n6672 ) ;
  assign n6674 = ( n1970 & n4124 ) | ( n1970 & n6595 ) | ( n4124 & n6595 ) ;
  assign n6675 = n1473 | n1716 ;
  assign n6676 = n6675 ^ n1294 ^ 1'b0 ;
  assign n6677 = ( n4144 & n6030 ) | ( n4144 & ~n6676 ) | ( n6030 & ~n6676 ) ;
  assign n6678 = n6677 ^ n2431 ^ 1'b0 ;
  assign n6679 = n2104 & n6678 ;
  assign n6680 = ~n1781 & n2562 ;
  assign n6681 = ~n6679 & n6680 ;
  assign n6682 = n4913 | n6681 ;
  assign n6683 = n5498 & ~n6682 ;
  assign n6684 = n6115 ^ n1114 ^ n338 ;
  assign n6688 = n4900 ^ n2853 ^ n447 ;
  assign n6689 = ( ~n890 & n1882 ) | ( ~n890 & n6688 ) | ( n1882 & n6688 ) ;
  assign n6690 = ~n2389 & n6689 ;
  assign n6691 = n6690 ^ n644 ^ 1'b0 ;
  assign n6692 = n6302 ^ n1788 ^ 1'b0 ;
  assign n6693 = ~n5802 & n6692 ;
  assign n6694 = ( n4371 & n6691 ) | ( n4371 & n6693 ) | ( n6691 & n6693 ) ;
  assign n6686 = ( n1095 & ~n2487 ) | ( n1095 & n2775 ) | ( ~n2487 & n2775 ) ;
  assign n6685 = n3873 ^ n1597 ^ n180 ;
  assign n6687 = n6686 ^ n6685 ^ n1377 ;
  assign n6695 = n6694 ^ n6687 ^ n6660 ;
  assign n6696 = ( n3430 & ~n6133 ) | ( n3430 & n6695 ) | ( ~n6133 & n6695 ) ;
  assign n6699 = x100 & n3142 ;
  assign n6700 = n6699 ^ n4571 ^ 1'b0 ;
  assign n6701 = ( ~n1295 & n1703 ) | ( ~n1295 & n6700 ) | ( n1703 & n6700 ) ;
  assign n6697 = ( n648 & n1131 ) | ( n648 & ~n1565 ) | ( n1131 & ~n1565 ) ;
  assign n6698 = n6697 ^ n1080 ^ n476 ;
  assign n6702 = n6701 ^ n6698 ^ n1545 ;
  assign n6707 = ( n409 & n1368 ) | ( n409 & ~n2092 ) | ( n1368 & ~n2092 ) ;
  assign n6705 = ( n1954 & n2525 ) | ( n1954 & n5559 ) | ( n2525 & n5559 ) ;
  assign n6703 = ( n1195 & n1367 ) | ( n1195 & ~n1940 ) | ( n1367 & ~n1940 ) ;
  assign n6704 = n4723 & n6703 ;
  assign n6706 = n6705 ^ n6704 ^ 1'b0 ;
  assign n6708 = n6707 ^ n6706 ^ n2412 ;
  assign n6711 = x107 & n4792 ;
  assign n6712 = ~n141 & n6711 ;
  assign n6713 = ( n3987 & n5103 ) | ( n3987 & n6685 ) | ( n5103 & n6685 ) ;
  assign n6714 = n6713 ^ n5803 ^ 1'b0 ;
  assign n6715 = n3407 & n6714 ;
  assign n6716 = ~n913 & n6715 ;
  assign n6717 = ( n1961 & n6712 ) | ( n1961 & n6716 ) | ( n6712 & n6716 ) ;
  assign n6709 = n5223 ^ n731 ^ 1'b0 ;
  assign n6710 = n5453 & n6709 ;
  assign n6718 = n6717 ^ n6710 ^ 1'b0 ;
  assign n6724 = ( n554 & ~n2941 ) | ( n554 & n4882 ) | ( ~n2941 & n4882 ) ;
  assign n6720 = n3585 ^ n2830 ^ n2191 ;
  assign n6721 = n6720 ^ n4928 ^ n4782 ;
  assign n6722 = ( n465 & ~n3219 ) | ( n465 & n6721 ) | ( ~n3219 & n6721 ) ;
  assign n6719 = n4505 ^ n3419 ^ n3147 ;
  assign n6723 = n6722 ^ n6719 ^ n1032 ;
  assign n6725 = n6724 ^ n6723 ^ n5431 ;
  assign n6726 = n1181 ^ n598 ^ 1'b0 ;
  assign n6727 = ~n2835 & n6726 ;
  assign n6728 = ( n3928 & n6529 ) | ( n3928 & ~n6727 ) | ( n6529 & ~n6727 ) ;
  assign n6729 = n2910 ^ n2224 ^ n1154 ;
  assign n6730 = ( n1269 & n6728 ) | ( n1269 & ~n6729 ) | ( n6728 & ~n6729 ) ;
  assign n6731 = n6730 ^ n5650 ^ n1058 ;
  assign n6732 = n5920 ^ n3805 ^ n547 ;
  assign n6733 = ( n2316 & ~n3640 ) | ( n2316 & n6732 ) | ( ~n3640 & n6732 ) ;
  assign n6734 = n6733 ^ n6469 ^ n5134 ;
  assign n6735 = n387 & n3346 ;
  assign n6742 = n4321 ^ n733 ^ n333 ;
  assign n6739 = n2910 ^ n2422 ^ n810 ;
  assign n6740 = n6739 ^ n1168 ^ n144 ;
  assign n6741 = n6740 ^ n5971 ^ n256 ;
  assign n6743 = n6742 ^ n6741 ^ n3121 ;
  assign n6736 = ( n808 & ~n1017 ) | ( n808 & n3115 ) | ( ~n1017 & n3115 ) ;
  assign n6737 = n6736 ^ n367 ^ 1'b0 ;
  assign n6738 = ( x119 & n2179 ) | ( x119 & n6737 ) | ( n2179 & n6737 ) ;
  assign n6744 = n6743 ^ n6738 ^ n4865 ;
  assign n6745 = n1052 | n2425 ;
  assign n6746 = n6639 ^ n3471 ^ 1'b0 ;
  assign n6747 = n6745 | n6746 ;
  assign n6748 = ~n640 & n4211 ;
  assign n6749 = n981 & n6748 ;
  assign n6750 = ( n3127 & ~n3545 ) | ( n3127 & n6749 ) | ( ~n3545 & n6749 ) ;
  assign n6751 = ( n3119 & n6747 ) | ( n3119 & ~n6750 ) | ( n6747 & ~n6750 ) ;
  assign n6752 = n748 & ~n2758 ;
  assign n6753 = n6752 ^ n2436 ^ 1'b0 ;
  assign n6754 = n6753 ^ n3350 ^ n3088 ;
  assign n6755 = n6754 ^ n3756 ^ n3488 ;
  assign n6756 = n3849 & ~n6755 ;
  assign n6757 = n6751 & n6756 ;
  assign n6758 = n422 & n1057 ;
  assign n6759 = n6758 ^ n6521 ^ 1'b0 ;
  assign n6760 = n2447 & n2916 ;
  assign n6761 = n3590 & n6760 ;
  assign n6762 = n6761 ^ n3210 ^ 1'b0 ;
  assign n6763 = ( ~n539 & n3542 ) | ( ~n539 & n4178 ) | ( n3542 & n4178 ) ;
  assign n6764 = ( n828 & n6762 ) | ( n828 & n6763 ) | ( n6762 & n6763 ) ;
  assign n6765 = n6764 ^ n5546 ^ n2216 ;
  assign n6766 = ( ~n150 & n953 ) | ( ~n150 & n6765 ) | ( n953 & n6765 ) ;
  assign n6773 = n5287 ^ n1435 ^ n439 ;
  assign n6774 = n6773 ^ n2872 ^ 1'b0 ;
  assign n6775 = ~n1896 & n6774 ;
  assign n6767 = ( n374 & ~n1504 ) | ( n374 & n4243 ) | ( ~n1504 & n4243 ) ;
  assign n6768 = n143 | n1559 ;
  assign n6769 = n6767 | n6768 ;
  assign n6770 = n457 & ~n826 ;
  assign n6771 = n6770 ^ n3931 ^ 1'b0 ;
  assign n6772 = ( n5157 & ~n6769 ) | ( n5157 & n6771 ) | ( ~n6769 & n6771 ) ;
  assign n6776 = n6775 ^ n6772 ^ n6441 ;
  assign n6777 = ( n5159 & n6024 ) | ( n5159 & n6776 ) | ( n6024 & n6776 ) ;
  assign n6783 = n5083 ^ n1535 ^ x98 ;
  assign n6778 = ~n642 & n3212 ;
  assign n6779 = ( ~n215 & n4899 ) | ( ~n215 & n6778 ) | ( n4899 & n6778 ) ;
  assign n6780 = n5924 ^ n1394 ^ 1'b0 ;
  assign n6781 = n1271 & ~n6780 ;
  assign n6782 = ( ~n6419 & n6779 ) | ( ~n6419 & n6781 ) | ( n6779 & n6781 ) ;
  assign n6784 = n6783 ^ n6782 ^ n5763 ;
  assign n6785 = n3176 ^ n2104 ^ n629 ;
  assign n6786 = ( n946 & n3270 ) | ( n946 & ~n6098 ) | ( n3270 & ~n6098 ) ;
  assign n6787 = ( n370 & n2302 ) | ( n370 & n6572 ) | ( n2302 & n6572 ) ;
  assign n6788 = n5424 & ~n6787 ;
  assign n6789 = n6788 ^ n3928 ^ 1'b0 ;
  assign n6790 = ( n1081 & ~n2799 ) | ( n1081 & n6789 ) | ( ~n2799 & n6789 ) ;
  assign n6793 = ( ~n1012 & n1278 ) | ( ~n1012 & n4900 ) | ( n1278 & n4900 ) ;
  assign n6794 = n6793 ^ n5458 ^ 1'b0 ;
  assign n6791 = n931 ^ x122 ^ 1'b0 ;
  assign n6792 = n5582 | n6791 ;
  assign n6795 = n6794 ^ n6792 ^ n995 ;
  assign n6796 = n4650 ^ x62 ^ 1'b0 ;
  assign n6811 = n2272 | n6742 ;
  assign n6812 = n6811 ^ n5151 ^ 1'b0 ;
  assign n6805 = n1790 & n5622 ;
  assign n6806 = n6805 ^ n5310 ^ 1'b0 ;
  assign n6807 = n6806 ^ n6131 ^ n675 ;
  assign n6802 = ( ~n348 & n863 ) | ( ~n348 & n2670 ) | ( n863 & n2670 ) ;
  assign n6803 = x126 & n6802 ;
  assign n6804 = n6803 ^ n1577 ^ 1'b0 ;
  assign n6800 = n5060 ^ n4728 ^ n1350 ;
  assign n6801 = ( n1320 & n3759 ) | ( n1320 & ~n6800 ) | ( n3759 & ~n6800 ) ;
  assign n6808 = n6807 ^ n6804 ^ n6801 ;
  assign n6797 = n6479 ^ n3514 ^ n599 ;
  assign n6798 = ( n2325 & n3130 ) | ( n2325 & ~n6797 ) | ( n3130 & ~n6797 ) ;
  assign n6799 = n2449 & ~n6798 ;
  assign n6809 = n6808 ^ n6799 ^ 1'b0 ;
  assign n6810 = n5443 | n6809 ;
  assign n6813 = n6812 ^ n6810 ^ 1'b0 ;
  assign n6814 = ( n926 & n2775 ) | ( n926 & n3281 ) | ( n2775 & n3281 ) ;
  assign n6815 = n6542 | n6814 ;
  assign n6816 = x1 | n6815 ;
  assign n6817 = ( n438 & n735 ) | ( n438 & ~n1958 ) | ( n735 & ~n1958 ) ;
  assign n6823 = ( n573 & n678 ) | ( n573 & ~n5668 ) | ( n678 & ~n5668 ) ;
  assign n6820 = ~n161 & n872 ;
  assign n6821 = n1200 & ~n6820 ;
  assign n6822 = n6821 ^ n2477 ^ 1'b0 ;
  assign n6818 = x115 & ~n4864 ;
  assign n6819 = ( n1233 & n1995 ) | ( n1233 & ~n6818 ) | ( n1995 & ~n6818 ) ;
  assign n6824 = n6823 ^ n6822 ^ n6819 ;
  assign n6825 = n6824 ^ n4770 ^ 1'b0 ;
  assign n6826 = ~n6817 & n6825 ;
  assign n6827 = ( n816 & n2663 ) | ( n816 & ~n4544 ) | ( n2663 & ~n4544 ) ;
  assign n6828 = n4486 | n6827 ;
  assign n6829 = n1572 | n6828 ;
  assign n6830 = n5406 ^ n3542 ^ n3179 ;
  assign n6831 = n6830 ^ n3134 ^ 1'b0 ;
  assign n6832 = ~n4482 & n6831 ;
  assign n6833 = n6832 ^ n3101 ^ 1'b0 ;
  assign n6834 = n6829 & n6833 ;
  assign n6837 = ( n827 & n1392 ) | ( n827 & n1680 ) | ( n1392 & n1680 ) ;
  assign n6836 = n2388 ^ n1579 ^ 1'b0 ;
  assign n6835 = n167 & n5209 ;
  assign n6838 = n6837 ^ n6836 ^ n6835 ;
  assign n6839 = n5637 ^ n5458 ^ n2869 ;
  assign n6840 = ( n1165 & n5303 ) | ( n1165 & n6839 ) | ( n5303 & n6839 ) ;
  assign n6843 = n6402 ^ n4390 ^ n254 ;
  assign n6844 = n6247 ^ n3773 ^ n3340 ;
  assign n6845 = ( ~n3886 & n6843 ) | ( ~n3886 & n6844 ) | ( n6843 & n6844 ) ;
  assign n6841 = n2854 ^ n896 ^ 1'b0 ;
  assign n6842 = n2170 & ~n6841 ;
  assign n6846 = n6845 ^ n6842 ^ 1'b0 ;
  assign n6847 = n2546 & n4911 ;
  assign n6848 = n5227 ^ n1494 ^ x2 ;
  assign n6849 = ( n1574 & n3247 ) | ( n1574 & ~n4091 ) | ( n3247 & ~n4091 ) ;
  assign n6850 = n6849 ^ n6640 ^ 1'b0 ;
  assign n6851 = n3189 | n6850 ;
  assign n6852 = n6851 ^ n1721 ^ n1119 ;
  assign n6853 = ( ~n6327 & n6848 ) | ( ~n6327 & n6852 ) | ( n6848 & n6852 ) ;
  assign n6854 = ~n4060 & n5733 ;
  assign n6855 = ( n1549 & ~n5252 ) | ( n1549 & n6613 ) | ( ~n5252 & n6613 ) ;
  assign n6856 = n6855 ^ n3218 ^ 1'b0 ;
  assign n6858 = n4318 ^ n1705 ^ 1'b0 ;
  assign n6857 = ( n1144 & n1502 ) | ( n1144 & n5129 ) | ( n1502 & n5129 ) ;
  assign n6859 = n6858 ^ n6857 ^ n4408 ;
  assign n6863 = n2493 ^ n2229 ^ 1'b0 ;
  assign n6864 = n3102 & n6863 ;
  assign n6865 = n2652 & n6864 ;
  assign n6860 = n6400 ^ n4472 ^ n1747 ;
  assign n6861 = n6860 ^ n320 ^ 1'b0 ;
  assign n6862 = ( n865 & ~n3486 ) | ( n865 & n6861 ) | ( ~n3486 & n6861 ) ;
  assign n6866 = n6865 ^ n6862 ^ n6520 ;
  assign n6867 = n3825 ^ n1920 ^ n1056 ;
  assign n6868 = n5630 ^ n4591 ^ n3919 ;
  assign n6869 = ( n175 & n6867 ) | ( n175 & n6868 ) | ( n6867 & n6868 ) ;
  assign n6879 = n372 ^ x124 ^ 1'b0 ;
  assign n6880 = n1786 | n6879 ;
  assign n6881 = n2376 | n6880 ;
  assign n6870 = ( n1132 & n1434 ) | ( n1132 & ~n2106 ) | ( n1434 & ~n2106 ) ;
  assign n6871 = n4028 & ~n6870 ;
  assign n6872 = n2783 & n6871 ;
  assign n6873 = n1066 ^ n665 ^ n653 ;
  assign n6874 = ( n1820 & n2302 ) | ( n1820 & ~n6873 ) | ( n2302 & ~n6873 ) ;
  assign n6875 = n2713 & n4059 ;
  assign n6876 = n3755 & n6875 ;
  assign n6877 = n6874 & n6876 ;
  assign n6878 = n6872 | n6877 ;
  assign n6882 = n6881 ^ n6878 ^ 1'b0 ;
  assign n6883 = n5042 ^ n3805 ^ n1971 ;
  assign n6884 = ( n155 & n3317 ) | ( n155 & ~n6883 ) | ( n3317 & ~n6883 ) ;
  assign n6886 = ~n2147 & n4044 ;
  assign n6885 = n5595 ^ n2629 ^ n1971 ;
  assign n6887 = n6886 ^ n6885 ^ n1063 ;
  assign n6888 = ( n6282 & ~n6884 ) | ( n6282 & n6887 ) | ( ~n6884 & n6887 ) ;
  assign n6889 = n2762 ^ n2163 ^ n1676 ;
  assign n6890 = n6889 ^ n5808 ^ n1022 ;
  assign n6891 = ( n1727 & n5814 ) | ( n1727 & n6890 ) | ( n5814 & n6890 ) ;
  assign n6892 = ( n931 & ~n2196 ) | ( n931 & n6891 ) | ( ~n2196 & n6891 ) ;
  assign n6893 = ( x66 & n2208 ) | ( x66 & n2987 ) | ( n2208 & n2987 ) ;
  assign n6894 = n4918 ^ n2513 ^ n774 ;
  assign n6895 = n6894 ^ n1841 ^ x48 ;
  assign n6896 = n6895 ^ n3697 ^ n1474 ;
  assign n6897 = ~n2748 & n3863 ;
  assign n6898 = n2262 ^ n1584 ^ 1'b0 ;
  assign n6899 = n6897 | n6898 ;
  assign n6900 = ( n1395 & n6896 ) | ( n1395 & ~n6899 ) | ( n6896 & ~n6899 ) ;
  assign n6901 = n2617 & ~n6900 ;
  assign n6902 = n1400 | n1854 ;
  assign n6903 = n3396 & ~n6902 ;
  assign n6904 = n1647 & ~n6903 ;
  assign n6905 = ( n903 & n2922 ) | ( n903 & ~n6904 ) | ( n2922 & ~n6904 ) ;
  assign n6906 = n6905 ^ n2640 ^ 1'b0 ;
  assign n6907 = ~n4590 & n6906 ;
  assign n6908 = n6247 ^ n4116 ^ n3450 ;
  assign n6909 = n6908 ^ n3634 ^ 1'b0 ;
  assign n6910 = n6907 & ~n6909 ;
  assign n6911 = ~n5303 & n6910 ;
  assign n6912 = ~n6697 & n6911 ;
  assign n6913 = n2163 & n6559 ;
  assign n6919 = n3929 ^ n677 ^ 1'b0 ;
  assign n6920 = ~n3882 & n6919 ;
  assign n6921 = n6920 ^ n5181 ^ n1399 ;
  assign n6918 = n661 | n4150 ;
  assign n6917 = n6541 ^ n1163 ^ n143 ;
  assign n6922 = n6921 ^ n6918 ^ n6917 ;
  assign n6914 = n3231 ^ n2279 ^ n1423 ;
  assign n6915 = ( n1649 & n3555 ) | ( n1649 & ~n6914 ) | ( n3555 & ~n6914 ) ;
  assign n6916 = n5879 & ~n6915 ;
  assign n6923 = n6922 ^ n6916 ^ 1'b0 ;
  assign n6937 = ~n444 & n1259 ;
  assign n6938 = n6937 ^ x122 ^ 1'b0 ;
  assign n6939 = ( ~n564 & n4603 ) | ( ~n564 & n6938 ) | ( n4603 & n6938 ) ;
  assign n6933 = n2733 ^ n1356 ^ 1'b0 ;
  assign n6934 = n6933 ^ n1480 ^ n1050 ;
  assign n6931 = n984 | n1778 ;
  assign n6932 = n6931 ^ n456 ^ 1'b0 ;
  assign n6930 = ( n3534 & n3551 ) | ( n3534 & ~n4437 ) | ( n3551 & ~n4437 ) ;
  assign n6935 = n6934 ^ n6932 ^ n6930 ;
  assign n6936 = n3133 | n6935 ;
  assign n6940 = n6939 ^ n6936 ^ 1'b0 ;
  assign n6941 = n4216 | n6940 ;
  assign n6924 = n1821 ^ n762 ^ n619 ;
  assign n6925 = n6924 ^ n1848 ^ 1'b0 ;
  assign n6926 = ( n306 & ~n794 ) | ( n306 & n3491 ) | ( ~n794 & n3491 ) ;
  assign n6927 = ~n3655 & n6926 ;
  assign n6928 = n6927 ^ n1451 ^ 1'b0 ;
  assign n6929 = n6925 & n6928 ;
  assign n6942 = n6941 ^ n6929 ^ n2487 ;
  assign n6943 = ( n320 & n2570 ) | ( n320 & ~n3210 ) | ( n2570 & ~n3210 ) ;
  assign n6944 = ( ~n4619 & n6550 ) | ( ~n4619 & n6943 ) | ( n6550 & n6943 ) ;
  assign n6945 = n2709 ^ n346 ^ 1'b0 ;
  assign n6946 = n6944 & n6945 ;
  assign n6947 = n6946 ^ n692 ^ 1'b0 ;
  assign n6951 = ( ~n1093 & n1962 ) | ( ~n1093 & n2000 ) | ( n1962 & n2000 ) ;
  assign n6948 = ( ~n1725 & n3124 ) | ( ~n1725 & n6030 ) | ( n3124 & n6030 ) ;
  assign n6949 = n6281 ^ n5014 ^ n1083 ;
  assign n6950 = ( n6340 & n6948 ) | ( n6340 & n6949 ) | ( n6948 & n6949 ) ;
  assign n6952 = n6951 ^ n6950 ^ n4834 ;
  assign n6953 = n4667 ^ n4617 ^ n529 ;
  assign n6954 = n6953 ^ n2196 ^ 1'b0 ;
  assign n6955 = n1281 & ~n2719 ;
  assign n6956 = ~n279 & n6955 ;
  assign n6957 = n4184 & n4721 ;
  assign n6958 = ~n1812 & n4326 ;
  assign n6959 = n6958 ^ n404 ^ 1'b0 ;
  assign n6960 = n6959 ^ n3684 ^ n1012 ;
  assign n6961 = n1073 & ~n3740 ;
  assign n6962 = ( n5710 & n6960 ) | ( n5710 & n6961 ) | ( n6960 & n6961 ) ;
  assign n6963 = ( n4987 & n6957 ) | ( n4987 & ~n6962 ) | ( n6957 & ~n6962 ) ;
  assign n6964 = ( n2297 & n6956 ) | ( n2297 & n6963 ) | ( n6956 & n6963 ) ;
  assign n6965 = n3480 ^ n511 ^ 1'b0 ;
  assign n6966 = ( n2017 & n6216 ) | ( n2017 & n6965 ) | ( n6216 & n6965 ) ;
  assign n6967 = ~n3178 & n6966 ;
  assign n6968 = n6967 ^ n1538 ^ 1'b0 ;
  assign n6969 = ( n3614 & ~n4251 ) | ( n3614 & n6968 ) | ( ~n4251 & n6968 ) ;
  assign n6970 = n3594 ^ n2532 ^ n2164 ;
  assign n6971 = ~x55 & n3012 ;
  assign n6972 = n4009 ^ n3684 ^ n589 ;
  assign n6973 = ( n1842 & n6971 ) | ( n1842 & ~n6972 ) | ( n6971 & ~n6972 ) ;
  assign n6974 = ( ~n3227 & n4257 ) | ( ~n3227 & n6973 ) | ( n4257 & n6973 ) ;
  assign n6975 = n6974 ^ n5990 ^ n2788 ;
  assign n6976 = ( n509 & n1432 ) | ( n509 & n4899 ) | ( n1432 & n4899 ) ;
  assign n6977 = n4802 ^ n4495 ^ n1910 ;
  assign n6978 = n6977 ^ n4321 ^ n943 ;
  assign n6979 = ( n6204 & ~n6976 ) | ( n6204 & n6978 ) | ( ~n6976 & n6978 ) ;
  assign n6980 = ( ~n1830 & n3263 ) | ( ~n1830 & n5111 ) | ( n3263 & n5111 ) ;
  assign n6981 = ( n2603 & ~n4195 ) | ( n2603 & n6980 ) | ( ~n4195 & n6980 ) ;
  assign n6982 = ( n2733 & n6979 ) | ( n2733 & n6981 ) | ( n6979 & n6981 ) ;
  assign n6983 = n4806 ^ n4450 ^ 1'b0 ;
  assign n6984 = n6983 ^ n2489 ^ 1'b0 ;
  assign n6985 = n5358 ^ n4487 ^ n2255 ;
  assign n6986 = n6985 ^ n3609 ^ 1'b0 ;
  assign n6987 = n3255 ^ n2926 ^ n2527 ;
  assign n6988 = ( n2236 & n4120 ) | ( n2236 & ~n6987 ) | ( n4120 & ~n6987 ) ;
  assign n6989 = n6988 ^ n5018 ^ x25 ;
  assign n6990 = ( n4222 & ~n6986 ) | ( n4222 & n6989 ) | ( ~n6986 & n6989 ) ;
  assign n6991 = n6695 ^ n3112 ^ 1'b0 ;
  assign n6992 = n3021 & n6991 ;
  assign n6993 = ( n3923 & n4862 ) | ( n3923 & ~n6992 ) | ( n4862 & ~n6992 ) ;
  assign n6994 = ( ~n201 & n2517 ) | ( ~n201 & n3079 ) | ( n2517 & n3079 ) ;
  assign n6996 = ~n778 & n1310 ;
  assign n6997 = n6996 ^ n3131 ^ n2269 ;
  assign n6995 = ( ~n1970 & n3214 ) | ( ~n1970 & n4504 ) | ( n3214 & n4504 ) ;
  assign n6998 = n6997 ^ n6995 ^ n5759 ;
  assign n6999 = n5296 ^ n2293 ^ n1912 ;
  assign n7002 = n500 & n3684 ;
  assign n7003 = n5828 | n7002 ;
  assign n7000 = n4071 & n4792 ;
  assign n7001 = n7000 ^ x68 ^ 1'b0 ;
  assign n7004 = n7003 ^ n7001 ^ n2849 ;
  assign n7005 = ( n6020 & n6999 ) | ( n6020 & n7004 ) | ( n6999 & n7004 ) ;
  assign n7006 = n4421 ^ n2871 ^ n1350 ;
  assign n7007 = n7006 ^ n3088 ^ n1806 ;
  assign n7008 = ( n2694 & ~n6302 ) | ( n2694 & n7007 ) | ( ~n6302 & n7007 ) ;
  assign n7009 = n2913 ^ n1120 ^ n730 ;
  assign n7010 = n3047 | n7009 ;
  assign n7011 = n1672 & ~n7010 ;
  assign n7012 = n3199 | n7011 ;
  assign n7013 = n3264 | n7012 ;
  assign n7014 = ( n4172 & n7008 ) | ( n4172 & n7013 ) | ( n7008 & n7013 ) ;
  assign n7016 = ( n1168 & n3773 ) | ( n1168 & ~n5061 ) | ( n3773 & ~n5061 ) ;
  assign n7015 = n3477 ^ n2380 ^ n1731 ;
  assign n7017 = n7016 ^ n7015 ^ n2661 ;
  assign n7018 = n2091 & n4143 ;
  assign n7019 = n7018 ^ n6949 ^ 1'b0 ;
  assign n7020 = n2305 ^ x70 ^ 1'b0 ;
  assign n7021 = ( n5091 & n6366 ) | ( n5091 & ~n7020 ) | ( n6366 & ~n7020 ) ;
  assign n7022 = n1310 & ~n7021 ;
  assign n7023 = ( x2 & n2034 ) | ( x2 & ~n3581 ) | ( n2034 & ~n3581 ) ;
  assign n7024 = ( ~n2026 & n6971 ) | ( ~n2026 & n7023 ) | ( n6971 & n7023 ) ;
  assign n7025 = n7024 ^ n6984 ^ 1'b0 ;
  assign n7026 = ~n7022 & n7025 ;
  assign n7031 = n6657 ^ n6572 ^ n4817 ;
  assign n7032 = ( ~n218 & n5803 ) | ( ~n218 & n7031 ) | ( n5803 & n7031 ) ;
  assign n7027 = n688 | n4156 ;
  assign n7028 = n2471 | n7027 ;
  assign n7029 = ( n3362 & ~n3967 ) | ( n3362 & n4587 ) | ( ~n3967 & n4587 ) ;
  assign n7030 = n7028 | n7029 ;
  assign n7033 = n7032 ^ n7030 ^ n873 ;
  assign n7034 = ( n425 & n2925 ) | ( n425 & n3033 ) | ( n2925 & n3033 ) ;
  assign n7035 = n7034 ^ n6383 ^ n5649 ;
  assign n7036 = n209 | n7035 ;
  assign n7037 = n707 & ~n7011 ;
  assign n7038 = n7037 ^ n1544 ^ 1'b0 ;
  assign n7041 = ( n704 & ~n1606 ) | ( n704 & n1733 ) | ( ~n1606 & n1733 ) ;
  assign n7039 = n1265 ^ n735 ^ 1'b0 ;
  assign n7040 = ( n1675 & ~n4690 ) | ( n1675 & n7039 ) | ( ~n4690 & n7039 ) ;
  assign n7042 = n7041 ^ n7040 ^ n2623 ;
  assign n7043 = n7042 ^ n4096 ^ n2037 ;
  assign n7044 = n913 | n4207 ;
  assign n7045 = ~n734 & n7044 ;
  assign n7046 = n7045 ^ n2924 ^ 1'b0 ;
  assign n7048 = ~n1448 & n4183 ;
  assign n7049 = n3220 & n7048 ;
  assign n7047 = n784 & ~n5488 ;
  assign n7050 = n7049 ^ n7047 ^ 1'b0 ;
  assign n7051 = n141 & n7050 ;
  assign n7052 = n7051 ^ n1644 ^ n711 ;
  assign n7053 = n7052 ^ n3303 ^ 1'b0 ;
  assign n7054 = ( ~n3559 & n4196 ) | ( ~n3559 & n4519 ) | ( n4196 & n4519 ) ;
  assign n7055 = n7054 ^ n2040 ^ 1'b0 ;
  assign n7056 = n402 & n1874 ;
  assign n7057 = n6110 & n7056 ;
  assign n7058 = ( n4281 & n5702 ) | ( n4281 & ~n7057 ) | ( n5702 & ~n7057 ) ;
  assign n7059 = n1550 & n4707 ;
  assign n7060 = n3791 ^ n130 ^ x11 ;
  assign n7061 = n7060 ^ n6459 ^ 1'b0 ;
  assign n7062 = n7059 & ~n7061 ;
  assign n7063 = n7062 ^ n5183 ^ n1268 ;
  assign n7064 = n1466 | n2626 ;
  assign n7065 = n1143 & ~n7064 ;
  assign n7072 = n3566 ^ n2107 ^ 1'b0 ;
  assign n7073 = n4346 ^ n2098 ^ n1942 ;
  assign n7074 = ( n3707 & n7072 ) | ( n3707 & ~n7073 ) | ( n7072 & ~n7073 ) ;
  assign n7069 = n930 & n2778 ;
  assign n7070 = n566 & n7069 ;
  assign n7071 = n7070 ^ n2621 ^ n1201 ;
  assign n7075 = n7074 ^ n7071 ^ n3757 ;
  assign n7066 = ( n1216 & ~n2337 ) | ( n1216 & n2402 ) | ( ~n2337 & n2402 ) ;
  assign n7067 = n3317 ^ n878 ^ n799 ;
  assign n7068 = n7066 | n7067 ;
  assign n7076 = n7075 ^ n7068 ^ n4176 ;
  assign n7077 = ( ~n4059 & n7065 ) | ( ~n4059 & n7076 ) | ( n7065 & n7076 ) ;
  assign n7078 = n4774 & ~n7077 ;
  assign n7079 = n5965 ^ n2697 ^ n1335 ;
  assign n7080 = ~n2127 & n7079 ;
  assign n7081 = n7080 ^ n2032 ^ n1072 ;
  assign n7082 = n7081 ^ n3475 ^ 1'b0 ;
  assign n7083 = n1837 ^ n385 ^ n149 ;
  assign n7084 = n1929 & n7083 ;
  assign n7085 = n7084 ^ n5348 ^ 1'b0 ;
  assign n7086 = n6175 ^ n5165 ^ n4302 ;
  assign n7087 = ~n583 & n7086 ;
  assign n7088 = ( ~x65 & n1656 ) | ( ~x65 & n3266 ) | ( n1656 & n3266 ) ;
  assign n7090 = n2862 ^ n727 ^ 1'b0 ;
  assign n7091 = x70 & n7090 ;
  assign n7089 = n6951 ^ n6863 ^ n597 ;
  assign n7092 = n7091 ^ n7089 ^ n543 ;
  assign n7093 = n4855 ^ n4691 ^ n3890 ;
  assign n7094 = n7093 ^ n2855 ^ 1'b0 ;
  assign n7098 = ( n1164 & ~n3904 ) | ( n1164 & n5154 ) | ( ~n3904 & n5154 ) ;
  assign n7095 = n5712 ^ x115 ^ 1'b0 ;
  assign n7096 = n326 & n7095 ;
  assign n7097 = n7096 ^ n6277 ^ 1'b0 ;
  assign n7099 = n7098 ^ n7097 ^ n618 ;
  assign n7100 = n6260 ^ n2203 ^ 1'b0 ;
  assign n7101 = n5899 ^ n3651 ^ n3121 ;
  assign n7102 = n7101 ^ n6651 ^ x65 ;
  assign n7103 = n5251 ^ n2858 ^ n1153 ;
  assign n7104 = n761 & n1124 ;
  assign n7105 = n7104 ^ n3286 ^ 1'b0 ;
  assign n7106 = ~n6903 & n7105 ;
  assign n7107 = n3107 ^ n2561 ^ 1'b0 ;
  assign n7108 = n7106 & n7107 ;
  assign n7109 = ~n7103 & n7108 ;
  assign n7110 = ~n3097 & n7109 ;
  assign n7115 = n2659 ^ n2397 ^ 1'b0 ;
  assign n7116 = n344 & ~n7115 ;
  assign n7111 = n2150 ^ n1675 ^ n1652 ;
  assign n7112 = n4437 & ~n7111 ;
  assign n7113 = n7112 ^ n4798 ^ n4015 ;
  assign n7114 = ~n4063 & n7113 ;
  assign n7117 = n7116 ^ n7114 ^ 1'b0 ;
  assign n7119 = ( n399 & n1663 ) | ( n399 & ~n3276 ) | ( n1663 & ~n3276 ) ;
  assign n7120 = ( n4668 & n4958 ) | ( n4668 & ~n7119 ) | ( n4958 & ~n7119 ) ;
  assign n7118 = ~n964 & n2925 ;
  assign n7121 = n7120 ^ n7118 ^ 1'b0 ;
  assign n7122 = n7117 | n7121 ;
  assign n7125 = n6987 ^ n3562 ^ n1476 ;
  assign n7123 = ( ~n3844 & n4689 ) | ( ~n3844 & n5015 ) | ( n4689 & n5015 ) ;
  assign n7124 = ( n3424 & n5173 ) | ( n3424 & ~n7123 ) | ( n5173 & ~n7123 ) ;
  assign n7126 = n7125 ^ n7124 ^ 1'b0 ;
  assign n7127 = n3053 & ~n7126 ;
  assign n7138 = ~n1274 & n1377 ;
  assign n7129 = n2837 ^ n2234 ^ 1'b0 ;
  assign n7128 = n4711 ^ n2161 ^ n935 ;
  assign n7130 = n7129 ^ n7128 ^ n2993 ;
  assign n7132 = ( n1544 & n4296 ) | ( n1544 & n4914 ) | ( n4296 & n4914 ) ;
  assign n7133 = n7132 ^ n6088 ^ n5162 ;
  assign n7134 = ( ~n6265 & n6556 ) | ( ~n6265 & n7133 ) | ( n6556 & n7133 ) ;
  assign n7131 = ~n4157 & n5731 ;
  assign n7135 = n7134 ^ n7131 ^ 1'b0 ;
  assign n7136 = n6872 | n7135 ;
  assign n7137 = n7130 | n7136 ;
  assign n7139 = n7138 ^ n7137 ^ n350 ;
  assign n7140 = ( n822 & n2291 ) | ( n822 & n6979 ) | ( n2291 & n6979 ) ;
  assign n7141 = ( n1458 & ~n2718 ) | ( n1458 & n7140 ) | ( ~n2718 & n7140 ) ;
  assign n7150 = n1071 | n3805 ;
  assign n7151 = n556 & ~n7150 ;
  assign n7147 = n3560 ^ n1263 ^ n987 ;
  assign n7146 = ( n2979 & n3180 ) | ( n2979 & ~n4533 ) | ( n3180 & ~n4533 ) ;
  assign n7148 = n7147 ^ n7146 ^ n5973 ;
  assign n7149 = n7148 ^ n374 ^ 1'b0 ;
  assign n7142 = n5042 ^ n3483 ^ n3320 ;
  assign n7143 = n7142 ^ n3750 ^ n1531 ;
  assign n7144 = n4270 | n7143 ;
  assign n7145 = n7144 ^ n2744 ^ 1'b0 ;
  assign n7152 = n7151 ^ n7149 ^ n7145 ;
  assign n7153 = ( n1116 & n1263 ) | ( n1116 & ~n1271 ) | ( n1263 & ~n1271 ) ;
  assign n7154 = n7153 ^ n4928 ^ n2413 ;
  assign n7155 = ( n144 & n4004 ) | ( n144 & n7154 ) | ( n4004 & n7154 ) ;
  assign n7156 = ( n149 & n3121 ) | ( n149 & ~n7155 ) | ( n3121 & ~n7155 ) ;
  assign n7157 = ( n2539 & n2716 ) | ( n2539 & n2851 ) | ( n2716 & n2851 ) ;
  assign n7158 = n5315 & ~n6281 ;
  assign n7159 = ~n7157 & n7158 ;
  assign n7160 = ( n1894 & n7156 ) | ( n1894 & n7159 ) | ( n7156 & n7159 ) ;
  assign n7161 = n5068 ^ n4929 ^ 1'b0 ;
  assign n7162 = n560 & ~n7161 ;
  assign n7163 = n7162 ^ n4018 ^ 1'b0 ;
  assign n7164 = n3717 ^ n1563 ^ 1'b0 ;
  assign n7165 = n7164 ^ n4837 ^ n4714 ;
  assign n7166 = ( n332 & n1163 ) | ( n332 & n1530 ) | ( n1163 & n1530 ) ;
  assign n7167 = ( n2236 & ~n4428 ) | ( n2236 & n7166 ) | ( ~n4428 & n7166 ) ;
  assign n7168 = n889 | n2267 ;
  assign n7169 = n7168 ^ n1226 ^ 1'b0 ;
  assign n7170 = n648 & ~n3361 ;
  assign n7171 = n5361 & n7170 ;
  assign n7172 = n7171 ^ n1028 ^ 1'b0 ;
  assign n7186 = ( ~n951 & n1395 ) | ( ~n951 & n3589 ) | ( n1395 & n3589 ) ;
  assign n7184 = ( n1471 & n2562 ) | ( n1471 & ~n4945 ) | ( n2562 & ~n4945 ) ;
  assign n7185 = ( ~n3417 & n4368 ) | ( ~n3417 & n7184 ) | ( n4368 & n7184 ) ;
  assign n7173 = n3670 ^ n3084 ^ n1607 ;
  assign n7174 = n7173 ^ n1248 ^ n1009 ;
  assign n7175 = n1541 & n2442 ;
  assign n7181 = n2091 ^ n1585 ^ n1020 ;
  assign n7176 = n6197 ^ n3784 ^ n736 ;
  assign n7177 = ( n249 & n4868 ) | ( n249 & ~n7176 ) | ( n4868 & ~n7176 ) ;
  assign n7178 = ( n2949 & ~n4097 ) | ( n2949 & n7112 ) | ( ~n4097 & n7112 ) ;
  assign n7179 = n4590 | n7178 ;
  assign n7180 = n7177 | n7179 ;
  assign n7182 = n7181 ^ n7180 ^ 1'b0 ;
  assign n7183 = ( n7174 & n7175 ) | ( n7174 & ~n7182 ) | ( n7175 & ~n7182 ) ;
  assign n7187 = n7186 ^ n7185 ^ n7183 ;
  assign n7188 = n7187 ^ n6454 ^ 1'b0 ;
  assign n7189 = ~n5585 & n7188 ;
  assign n7190 = x40 & n2660 ;
  assign n7191 = ( n3435 & ~n4802 ) | ( n3435 & n7190 ) | ( ~n4802 & n7190 ) ;
  assign n7192 = n7191 ^ n4474 ^ n2083 ;
  assign n7193 = n4340 | n7192 ;
  assign n7194 = n7193 ^ n1576 ^ 1'b0 ;
  assign n7201 = n3481 ^ n1516 ^ n385 ;
  assign n7195 = n1109 ^ n926 ^ 1'b0 ;
  assign n7197 = n1306 ^ n692 ^ 1'b0 ;
  assign n7198 = n3467 & n7197 ;
  assign n7196 = ( n2389 & n3178 ) | ( n2389 & ~n5091 ) | ( n3178 & ~n5091 ) ;
  assign n7199 = n7198 ^ n7196 ^ n4213 ;
  assign n7200 = ( x41 & n7195 ) | ( x41 & ~n7199 ) | ( n7195 & ~n7199 ) ;
  assign n7202 = n7201 ^ n7200 ^ n423 ;
  assign n7203 = n451 & n2690 ;
  assign n7204 = n4277 & ~n7203 ;
  assign n7205 = n7204 ^ n4620 ^ n2888 ;
  assign n7206 = n7205 ^ n1373 ^ n186 ;
  assign n7207 = n2022 ^ n893 ^ n434 ;
  assign n7208 = n7207 ^ n2105 ^ n2006 ;
  assign n7209 = ( ~n3857 & n5526 ) | ( ~n3857 & n7208 ) | ( n5526 & n7208 ) ;
  assign n7210 = n1572 & n5624 ;
  assign n7211 = n7210 ^ n5763 ^ 1'b0 ;
  assign n7212 = n2976 ^ n1876 ^ 1'b0 ;
  assign n7213 = n4102 & n7212 ;
  assign n7214 = n4087 ^ n1565 ^ n1348 ;
  assign n7215 = n7214 ^ n5352 ^ n3285 ;
  assign n7216 = n5574 & ~n7215 ;
  assign n7217 = n4009 & n7216 ;
  assign n7229 = n3201 ^ n3074 ^ n772 ;
  assign n7230 = n3294 ^ n3068 ^ n775 ;
  assign n7231 = n7230 ^ n551 ^ 1'b0 ;
  assign n7232 = n7229 & n7231 ;
  assign n7233 = n3734 & n7232 ;
  assign n7226 = ( n846 & n1904 ) | ( n846 & n5161 ) | ( n1904 & n5161 ) ;
  assign n7227 = ( ~n1959 & n2022 ) | ( ~n1959 & n7226 ) | ( n2022 & n7226 ) ;
  assign n7223 = n1228 & n4520 ;
  assign n7224 = n5933 & n7223 ;
  assign n7225 = n7224 ^ n3640 ^ n1737 ;
  assign n7218 = ( ~n716 & n952 ) | ( ~n716 & n2873 ) | ( n952 & n2873 ) ;
  assign n7219 = n3664 ^ n2055 ^ n815 ;
  assign n7220 = ~n7218 & n7219 ;
  assign n7221 = x22 & ~n3375 ;
  assign n7222 = n7220 & n7221 ;
  assign n7228 = n7227 ^ n7225 ^ n7222 ;
  assign n7234 = n7233 ^ n7228 ^ 1'b0 ;
  assign n7235 = n7217 | n7234 ;
  assign n7236 = n3079 ^ n1656 ^ n1200 ;
  assign n7237 = n3496 & n7236 ;
  assign n7238 = n7237 ^ n2016 ^ 1'b0 ;
  assign n7239 = n7238 ^ n3342 ^ 1'b0 ;
  assign n7240 = n5624 | n7239 ;
  assign n7241 = n2018 & n2043 ;
  assign n7242 = n2094 ^ n1338 ^ 1'b0 ;
  assign n7243 = ~n7241 & n7242 ;
  assign n7244 = n7243 ^ n4895 ^ 1'b0 ;
  assign n7246 = n2191 ^ n635 ^ 1'b0 ;
  assign n7247 = n7246 ^ n5090 ^ 1'b0 ;
  assign n7248 = n4663 | n7247 ;
  assign n7245 = ~n1630 & n2826 ;
  assign n7249 = n7248 ^ n7245 ^ n497 ;
  assign n7250 = ~n1575 & n7249 ;
  assign n7251 = n3045 ^ n1038 ^ n941 ;
  assign n7256 = n3023 ^ n1281 ^ 1'b0 ;
  assign n7257 = n1205 & ~n7256 ;
  assign n7252 = n3623 ^ n3182 ^ 1'b0 ;
  assign n7253 = n678 & ~n7252 ;
  assign n7254 = ( ~n539 & n6976 ) | ( ~n539 & n7253 ) | ( n6976 & n7253 ) ;
  assign n7255 = n7254 ^ n3983 ^ n837 ;
  assign n7258 = n7257 ^ n7255 ^ n1272 ;
  assign n7259 = n7251 & ~n7258 ;
  assign n7260 = n4705 ^ n139 ^ 1'b0 ;
  assign n7261 = n5279 ^ n795 ^ 1'b0 ;
  assign n7262 = ~n7022 & n7261 ;
  assign n7263 = n7260 & n7262 ;
  assign n7277 = n5049 & ~n7024 ;
  assign n7278 = n3659 & n7277 ;
  assign n7270 = ( n2782 & ~n2923 ) | ( n2782 & n3232 ) | ( ~n2923 & n3232 ) ;
  assign n7266 = n6789 ^ n4900 ^ n2648 ;
  assign n7265 = n2239 & n6401 ;
  assign n7267 = n7266 ^ n7265 ^ 1'b0 ;
  assign n7264 = n1346 ^ n280 ^ 1'b0 ;
  assign n7268 = n7267 ^ n7264 ^ n2385 ;
  assign n7269 = n7268 ^ n3920 ^ n3854 ;
  assign n7271 = n7270 ^ n7269 ^ n2481 ;
  assign n7272 = n4783 ^ n4549 ^ n2712 ;
  assign n7273 = ( n4959 & n5700 ) | ( n4959 & ~n7272 ) | ( n5700 & ~n7272 ) ;
  assign n7274 = ( n2018 & n7271 ) | ( n2018 & ~n7273 ) | ( n7271 & ~n7273 ) ;
  assign n7275 = n1988 | n7274 ;
  assign n7276 = n7275 ^ n2912 ^ 1'b0 ;
  assign n7279 = n7278 ^ n7276 ^ n4810 ;
  assign n7280 = ( n997 & n5318 ) | ( n997 & ~n5624 ) | ( n5318 & ~n5624 ) ;
  assign n7281 = ~n592 & n4484 ;
  assign n7282 = ( n1198 & n2621 ) | ( n1198 & n7281 ) | ( n2621 & n7281 ) ;
  assign n7283 = ( n2527 & n4233 ) | ( n2527 & n7282 ) | ( n4233 & n7282 ) ;
  assign n7286 = n2615 | n2735 ;
  assign n7287 = n3523 | n7286 ;
  assign n7284 = ( n476 & n2135 ) | ( n476 & n3107 ) | ( n2135 & n3107 ) ;
  assign n7285 = ~n3566 & n7284 ;
  assign n7288 = n7287 ^ n7285 ^ 1'b0 ;
  assign n7289 = n7288 ^ n4834 ^ n2337 ;
  assign n7290 = n3096 ^ n2479 ^ n1929 ;
  assign n7291 = n6976 & n7290 ;
  assign n7292 = n7291 ^ n1601 ^ 1'b0 ;
  assign n7294 = n3990 ^ n1635 ^ x67 ;
  assign n7295 = ( ~n1019 & n5260 ) | ( ~n1019 & n7151 ) | ( n5260 & n7151 ) ;
  assign n7296 = ( ~n3073 & n7294 ) | ( ~n3073 & n7295 ) | ( n7294 & n7295 ) ;
  assign n7293 = n2664 & n3976 ;
  assign n7297 = n7296 ^ n7293 ^ 1'b0 ;
  assign n7298 = n4685 ^ n2320 ^ 1'b0 ;
  assign n7299 = n174 & n7298 ;
  assign n7300 = n7299 ^ n6924 ^ n2365 ;
  assign n7301 = n2009 | n6302 ;
  assign n7302 = n7300 & ~n7301 ;
  assign n7303 = ( n1414 & n5839 ) | ( n1414 & ~n7302 ) | ( n5839 & ~n7302 ) ;
  assign n7304 = ( ~n6856 & n7297 ) | ( ~n6856 & n7303 ) | ( n7297 & n7303 ) ;
  assign n7305 = ( n2535 & ~n3064 ) | ( n2535 & n4389 ) | ( ~n3064 & n4389 ) ;
  assign n7306 = n1591 & ~n4535 ;
  assign n7307 = ~n1184 & n7306 ;
  assign n7308 = n7307 ^ n2037 ^ n1108 ;
  assign n7309 = n4793 | n7308 ;
  assign n7310 = ( n282 & n704 ) | ( n282 & n3068 ) | ( n704 & n3068 ) ;
  assign n7311 = n6945 & n7310 ;
  assign n7312 = n7311 ^ n2501 ^ 1'b0 ;
  assign n7313 = ( n7305 & ~n7309 ) | ( n7305 & n7312 ) | ( ~n7309 & n7312 ) ;
  assign n7314 = n3008 ^ n551 ^ 1'b0 ;
  assign n7315 = n7314 ^ n7079 ^ n3651 ;
  assign n7316 = n1116 & n7315 ;
  assign n7317 = n7316 ^ n6464 ^ 1'b0 ;
  assign n7318 = ~n1423 & n7317 ;
  assign n7319 = n7318 ^ n6476 ^ 1'b0 ;
  assign n7320 = n3156 ^ n200 ^ 1'b0 ;
  assign n7321 = n7320 ^ n2982 ^ 1'b0 ;
  assign n7332 = n3040 ^ n2096 ^ 1'b0 ;
  assign n7333 = ~n5012 & n7332 ;
  assign n7334 = n3392 ^ n1340 ^ 1'b0 ;
  assign n7335 = n7333 & n7334 ;
  assign n7336 = n7284 ^ n4796 ^ n4450 ;
  assign n7337 = n7335 & n7336 ;
  assign n7338 = n2875 & n7337 ;
  assign n7328 = ( n1045 & n1835 ) | ( n1045 & ~n3384 ) | ( n1835 & ~n3384 ) ;
  assign n7329 = n7328 ^ n1679 ^ n474 ;
  assign n7330 = n7329 ^ n3721 ^ 1'b0 ;
  assign n7331 = n1230 | n7330 ;
  assign n7325 = n4762 ^ n2305 ^ n2289 ;
  assign n7326 = n7325 ^ n6275 ^ 1'b0 ;
  assign n7322 = n2463 ^ n1059 ^ n664 ;
  assign n7323 = ( n873 & n5090 ) | ( n873 & n5547 ) | ( n5090 & n5547 ) ;
  assign n7324 = ( n846 & ~n7322 ) | ( n846 & n7323 ) | ( ~n7322 & n7323 ) ;
  assign n7327 = n7326 ^ n7324 ^ n4208 ;
  assign n7339 = n7338 ^ n7331 ^ n7327 ;
  assign n7345 = n3631 ^ n2458 ^ n1601 ;
  assign n7340 = n6976 ^ n2558 ^ n749 ;
  assign n7341 = n7340 ^ n3761 ^ 1'b0 ;
  assign n7342 = n991 & ~n7341 ;
  assign n7343 = n1674 & ~n4828 ;
  assign n7344 = ( n3944 & ~n7342 ) | ( n3944 & n7343 ) | ( ~n7342 & n7343 ) ;
  assign n7346 = n7345 ^ n7344 ^ n3815 ;
  assign n7347 = n2516 ^ n809 ^ 1'b0 ;
  assign n7348 = ~n2639 & n7347 ;
  assign n7349 = ( n3797 & n4601 ) | ( n3797 & n7348 ) | ( n4601 & n7348 ) ;
  assign n7350 = ( ~n828 & n1009 ) | ( ~n828 & n7349 ) | ( n1009 & n7349 ) ;
  assign n7351 = n3221 ^ n1418 ^ n974 ;
  assign n7352 = n7351 ^ n5056 ^ n2547 ;
  assign n7353 = n1759 | n7352 ;
  assign n7354 = n4642 ^ n714 ^ n425 ;
  assign n7355 = n3919 & ~n7354 ;
  assign n7356 = ~n7353 & n7355 ;
  assign n7357 = n4899 ^ n3909 ^ n2934 ;
  assign n7358 = ~n623 & n6822 ;
  assign n7359 = ( n1211 & n1246 ) | ( n1211 & n1805 ) | ( n1246 & n1805 ) ;
  assign n7360 = n7359 ^ n2028 ^ n611 ;
  assign n7361 = n1269 ^ n861 ^ 1'b0 ;
  assign n7362 = ( n6192 & ~n6951 ) | ( n6192 & n7361 ) | ( ~n6951 & n7361 ) ;
  assign n7363 = ( n5060 & ~n5092 ) | ( n5060 & n5332 ) | ( ~n5092 & n5332 ) ;
  assign n7364 = n761 & n2152 ;
  assign n7365 = ( n2241 & n3499 ) | ( n2241 & ~n5142 ) | ( n3499 & ~n5142 ) ;
  assign n7366 = ( ~n396 & n3015 ) | ( ~n396 & n7365 ) | ( n3015 & n7365 ) ;
  assign n7367 = n5361 ^ n2252 ^ n1083 ;
  assign n7368 = ( ~n7364 & n7366 ) | ( ~n7364 & n7367 ) | ( n7366 & n7367 ) ;
  assign n7369 = n7214 ^ n4399 ^ n665 ;
  assign n7370 = ( n1258 & n1782 ) | ( n1258 & ~n4324 ) | ( n1782 & ~n4324 ) ;
  assign n7371 = n7370 ^ n3756 ^ 1'b0 ;
  assign n7372 = ( n4191 & n7369 ) | ( n4191 & n7371 ) | ( n7369 & n7371 ) ;
  assign n7373 = ( n2571 & n6753 ) | ( n2571 & n7372 ) | ( n6753 & n7372 ) ;
  assign n7374 = n1255 & ~n7373 ;
  assign n7375 = n7374 ^ n3523 ^ 1'b0 ;
  assign n7376 = x68 & ~n676 ;
  assign n7377 = n7376 ^ n765 ^ 1'b0 ;
  assign n7378 = n3195 ^ n2792 ^ n1519 ;
  assign n7379 = n2891 & n7378 ;
  assign n7380 = ( n2509 & ~n4655 ) | ( n2509 & n5039 ) | ( ~n4655 & n5039 ) ;
  assign n7381 = n7380 ^ n5763 ^ n2732 ;
  assign n7382 = n1431 ^ n1083 ^ 1'b0 ;
  assign n7383 = n7382 ^ n2396 ^ n1339 ;
  assign n7384 = n3430 & ~n5417 ;
  assign n7385 = ~n2577 & n7384 ;
  assign n7386 = n2173 ^ n2123 ^ n1296 ;
  assign n7387 = ~n1248 & n7386 ;
  assign n7388 = n763 & n7387 ;
  assign n7389 = n7385 & n7388 ;
  assign n7390 = n2076 | n7389 ;
  assign n7391 = ( n7381 & n7383 ) | ( n7381 & n7390 ) | ( n7383 & n7390 ) ;
  assign n7392 = ( n835 & n3452 ) | ( n835 & n6978 ) | ( n3452 & n6978 ) ;
  assign n7399 = n5386 ^ n465 ^ 1'b0 ;
  assign n7393 = n6130 ^ n3206 ^ n1290 ;
  assign n7394 = ( n2609 & ~n2834 ) | ( n2609 & n3660 ) | ( ~n2834 & n3660 ) ;
  assign n7395 = n7393 & n7394 ;
  assign n7396 = n4983 ^ n1402 ^ 1'b0 ;
  assign n7397 = ~x110 & n7396 ;
  assign n7398 = ~n7395 & n7397 ;
  assign n7400 = n7399 ^ n7398 ^ 1'b0 ;
  assign n7401 = ~n915 & n4421 ;
  assign n7402 = n5058 & n7401 ;
  assign n7403 = n4079 ^ n791 ^ n252 ;
  assign n7404 = ( n564 & ~n676 ) | ( n564 & n7403 ) | ( ~n676 & n7403 ) ;
  assign n7405 = n7404 ^ n5283 ^ n3150 ;
  assign n7406 = n1944 & n4804 ;
  assign n7407 = n7406 ^ n4154 ^ n671 ;
  assign n7408 = n3525 ^ n1728 ^ n1158 ;
  assign n7409 = ~n149 & n2036 ;
  assign n7410 = ( n3046 & n7408 ) | ( n3046 & ~n7409 ) | ( n7408 & ~n7409 ) ;
  assign n7411 = ( ~n5171 & n7300 ) | ( ~n5171 & n7410 ) | ( n7300 & n7410 ) ;
  assign n7412 = ( ~n7405 & n7407 ) | ( ~n7405 & n7411 ) | ( n7407 & n7411 ) ;
  assign n7422 = ~n1265 & n3643 ;
  assign n7421 = n3702 ^ n3457 ^ n2842 ;
  assign n7413 = n278 & ~n1705 ;
  assign n7414 = n2953 & n7413 ;
  assign n7415 = n1946 ^ n1340 ^ n208 ;
  assign n7416 = n7415 ^ n581 ^ 1'b0 ;
  assign n7417 = ~n2717 & n7416 ;
  assign n7418 = n7417 ^ n3307 ^ n2191 ;
  assign n7419 = ( n3286 & n7414 ) | ( n3286 & ~n7418 ) | ( n7414 & ~n7418 ) ;
  assign n7420 = ~n2167 & n7419 ;
  assign n7423 = n7422 ^ n7421 ^ n7420 ;
  assign n7424 = ~n1006 & n1882 ;
  assign n7425 = ( ~n3429 & n5977 ) | ( ~n3429 & n7424 ) | ( n5977 & n7424 ) ;
  assign n7426 = n7284 ^ n906 ^ n421 ;
  assign n7427 = n7426 ^ n2297 ^ n461 ;
  assign n7428 = n7427 ^ n2480 ^ 1'b0 ;
  assign n7433 = ( ~n2198 & n5282 ) | ( ~n2198 & n6285 ) | ( n5282 & n6285 ) ;
  assign n7429 = n2353 ^ n216 ^ 1'b0 ;
  assign n7430 = ~n3279 & n7429 ;
  assign n7431 = n7430 ^ n2496 ^ 1'b0 ;
  assign n7432 = n7431 ^ n1591 ^ n1415 ;
  assign n7434 = n7433 ^ n7432 ^ n1305 ;
  assign n7435 = ( n7425 & n7428 ) | ( n7425 & n7434 ) | ( n7428 & n7434 ) ;
  assign n7436 = ( n1723 & n2734 ) | ( n1723 & n3844 ) | ( n2734 & n3844 ) ;
  assign n7437 = n7436 ^ n3491 ^ n3117 ;
  assign n7438 = ~n5641 & n7437 ;
  assign n7439 = ~n4190 & n7438 ;
  assign n7440 = n7439 ^ n3145 ^ n2272 ;
  assign n7441 = n1842 ^ n1235 ^ 1'b0 ;
  assign n7447 = x78 & n2602 ;
  assign n7442 = ~n588 & n5336 ;
  assign n7443 = n7074 ^ n2756 ^ 1'b0 ;
  assign n7444 = n5150 ^ n3908 ^ n1765 ;
  assign n7445 = ( n5167 & n7443 ) | ( n5167 & ~n7444 ) | ( n7443 & ~n7444 ) ;
  assign n7446 = ( ~n778 & n7442 ) | ( ~n778 & n7445 ) | ( n7442 & n7445 ) ;
  assign n7448 = n7447 ^ n7446 ^ n2977 ;
  assign n7449 = ( ~n351 & n1743 ) | ( ~n351 & n2226 ) | ( n1743 & n2226 ) ;
  assign n7450 = n7449 ^ n7166 ^ n2181 ;
  assign n7451 = ( n381 & ~n829 ) | ( n381 & n7450 ) | ( ~n829 & n7450 ) ;
  assign n7452 = ( ~n2302 & n3878 ) | ( ~n2302 & n5060 ) | ( n3878 & n5060 ) ;
  assign n7453 = ( n6778 & n7451 ) | ( n6778 & n7452 ) | ( n7451 & n7452 ) ;
  assign n7454 = ( n1205 & n1335 ) | ( n1205 & ~n7453 ) | ( n1335 & ~n7453 ) ;
  assign n7455 = ( n558 & ~n3430 ) | ( n558 & n5524 ) | ( ~n3430 & n5524 ) ;
  assign n7471 = n1652 ^ n382 ^ x20 ;
  assign n7472 = ( n5026 & ~n6253 ) | ( n5026 & n7471 ) | ( ~n6253 & n7471 ) ;
  assign n7469 = ~n290 & n6299 ;
  assign n7470 = n7469 ^ n3863 ^ n423 ;
  assign n7456 = n3886 ^ n2259 ^ 1'b0 ;
  assign n7457 = n7456 ^ n2170 ^ n1936 ;
  assign n7458 = ( ~n248 & n2506 ) | ( ~n248 & n5379 ) | ( n2506 & n5379 ) ;
  assign n7459 = n295 & ~n7458 ;
  assign n7460 = ~x4 & n7459 ;
  assign n7461 = n1579 ^ n1530 ^ n486 ;
  assign n7462 = n7460 & ~n7461 ;
  assign n7465 = ( n422 & ~n1496 ) | ( n422 & n5708 ) | ( ~n1496 & n5708 ) ;
  assign n7463 = n4741 | n5802 ;
  assign n7464 = n681 & ~n7463 ;
  assign n7466 = n7465 ^ n7464 ^ n2269 ;
  assign n7467 = n3997 | n7466 ;
  assign n7468 = ( ~n7457 & n7462 ) | ( ~n7457 & n7467 ) | ( n7462 & n7467 ) ;
  assign n7473 = n7472 ^ n7470 ^ n7468 ;
  assign n7482 = n5513 ^ n3483 ^ n2028 ;
  assign n7483 = ~n1985 & n7482 ;
  assign n7477 = n2551 ^ n450 ^ 1'b0 ;
  assign n7478 = n4064 ^ n3933 ^ n780 ;
  assign n7479 = ( n1295 & ~n7477 ) | ( n1295 & n7478 ) | ( ~n7477 & n7478 ) ;
  assign n7480 = n7479 ^ n4008 ^ 1'b0 ;
  assign n7475 = ( ~n2624 & n4923 ) | ( ~n2624 & n5641 ) | ( n4923 & n5641 ) ;
  assign n7474 = n2403 ^ n2279 ^ 1'b0 ;
  assign n7476 = n7475 ^ n7474 ^ n5926 ;
  assign n7481 = n7480 ^ n7476 ^ n5389 ;
  assign n7484 = n7483 ^ n7481 ^ n6048 ;
  assign n7485 = n6905 ^ n5476 ^ n2089 ;
  assign n7486 = ( ~n3012 & n6443 ) | ( ~n3012 & n7485 ) | ( n6443 & n7485 ) ;
  assign n7487 = ( x31 & ~n2307 ) | ( x31 & n3989 ) | ( ~n2307 & n3989 ) ;
  assign n7488 = n1874 & n4235 ;
  assign n7489 = n2900 & n7488 ;
  assign n7490 = n7009 ^ n3035 ^ n145 ;
  assign n7491 = n7489 | n7490 ;
  assign n7492 = n7487 & ~n7491 ;
  assign n7494 = n6503 ^ n2346 ^ n1009 ;
  assign n7493 = n6738 ^ n5963 ^ n1244 ;
  assign n7495 = n7494 ^ n7493 ^ n4389 ;
  assign n7496 = ( ~n219 & n1688 ) | ( ~n219 & n1767 ) | ( n1688 & n1767 ) ;
  assign n7497 = n7496 ^ n3603 ^ 1'b0 ;
  assign n7498 = n1092 & ~n7497 ;
  assign n7499 = ( n2466 & n3709 ) | ( n2466 & n5311 ) | ( n3709 & n5311 ) ;
  assign n7500 = n7499 ^ n6696 ^ 1'b0 ;
  assign n7501 = n7498 & n7500 ;
  assign n7502 = n6378 & n6553 ;
  assign n7503 = ~n177 & n5549 ;
  assign n7504 = n7503 ^ n3896 ^ 1'b0 ;
  assign n7505 = n1304 & n1324 ;
  assign n7511 = ( ~n3488 & n4830 ) | ( ~n3488 & n7264 ) | ( n4830 & n7264 ) ;
  assign n7512 = n1572 & n1874 ;
  assign n7513 = n5423 & n7512 ;
  assign n7514 = ~n425 & n6098 ;
  assign n7515 = ( n4588 & n7513 ) | ( n4588 & n7514 ) | ( n7513 & n7514 ) ;
  assign n7516 = ( ~n3939 & n7511 ) | ( ~n3939 & n7515 ) | ( n7511 & n7515 ) ;
  assign n7506 = n2838 & n4046 ;
  assign n7507 = n4978 ^ n4476 ^ 1'b0 ;
  assign n7508 = n1304 & ~n7507 ;
  assign n7509 = ~n4000 & n7508 ;
  assign n7510 = n7506 | n7509 ;
  assign n7517 = n7516 ^ n7510 ^ 1'b0 ;
  assign n7518 = ( n1606 & n2019 ) | ( n1606 & ~n2598 ) | ( n2019 & ~n2598 ) ;
  assign n7519 = n7518 ^ n4930 ^ n2397 ;
  assign n7520 = ( n3617 & n6642 ) | ( n3617 & n7519 ) | ( n6642 & n7519 ) ;
  assign n7521 = n5410 ^ n5404 ^ n541 ;
  assign n7522 = n7521 ^ n5568 ^ n5518 ;
  assign n7523 = n3933 | n5564 ;
  assign n7524 = n7523 ^ n3423 ^ 1'b0 ;
  assign n7525 = n3117 ^ n2667 ^ n1541 ;
  assign n7526 = n7525 ^ n1863 ^ n1077 ;
  assign n7527 = n3259 & n4877 ;
  assign n7528 = n3953 & n7527 ;
  assign n7529 = n7528 ^ n3020 ^ n301 ;
  assign n7530 = ( n3677 & n7526 ) | ( n3677 & ~n7529 ) | ( n7526 & ~n7529 ) ;
  assign n7533 = ~n505 & n3876 ;
  assign n7534 = n7533 ^ n547 ^ 1'b0 ;
  assign n7531 = ( n699 & ~n3264 ) | ( n699 & n5424 ) | ( ~n3264 & n5424 ) ;
  assign n7532 = ( n1251 & n1925 ) | ( n1251 & ~n7531 ) | ( n1925 & ~n7531 ) ;
  assign n7535 = n7534 ^ n7532 ^ n2663 ;
  assign n7538 = n680 ^ n138 ^ x72 ;
  assign n7536 = n5047 ^ n4702 ^ n4383 ;
  assign n7537 = n1536 & ~n7536 ;
  assign n7539 = n7538 ^ n7537 ^ n2157 ;
  assign n7540 = n913 | n7147 ;
  assign n7541 = ( n1996 & ~n4213 ) | ( n1996 & n7540 ) | ( ~n4213 & n7540 ) ;
  assign n7542 = n161 | n3560 ;
  assign n7543 = n7542 ^ n649 ^ 1'b0 ;
  assign n7544 = n331 & n7543 ;
  assign n7545 = n4685 ^ x58 ^ 1'b0 ;
  assign n7546 = n988 | n7545 ;
  assign n7547 = n7544 & ~n7546 ;
  assign n7548 = n252 & n7547 ;
  assign n7549 = n7548 ^ n1563 ^ n1451 ;
  assign n7550 = ( ~n448 & n7541 ) | ( ~n448 & n7549 ) | ( n7541 & n7549 ) ;
  assign n7551 = n2154 ^ n1369 ^ 1'b0 ;
  assign n7552 = n733 | n7551 ;
  assign n7553 = n3801 & ~n7552 ;
  assign n7554 = n2866 ^ n2265 ^ n1364 ;
  assign n7555 = ( n1465 & n1921 ) | ( n1465 & n2007 ) | ( n1921 & n2007 ) ;
  assign n7556 = ( n3646 & n7554 ) | ( n3646 & ~n7555 ) | ( n7554 & ~n7555 ) ;
  assign n7557 = ( n3285 & n3621 ) | ( n3285 & ~n5083 ) | ( n3621 & ~n5083 ) ;
  assign n7558 = n6024 ^ n1271 ^ 1'b0 ;
  assign n7559 = n7149 ^ n5668 ^ n5519 ;
  assign n7560 = ( ~n7557 & n7558 ) | ( ~n7557 & n7559 ) | ( n7558 & n7559 ) ;
  assign n7565 = ( n195 & n1141 ) | ( n195 & ~n2132 ) | ( n1141 & ~n2132 ) ;
  assign n7562 = n2879 ^ n1752 ^ 1'b0 ;
  assign n7563 = n1550 & n7562 ;
  assign n7564 = n7563 ^ n3545 ^ n1932 ;
  assign n7566 = n7565 ^ n7564 ^ n4701 ;
  assign n7561 = n7146 ^ n4973 ^ n3283 ;
  assign n7567 = n7566 ^ n7561 ^ n5308 ;
  assign n7568 = ( ~n7556 & n7560 ) | ( ~n7556 & n7567 ) | ( n7560 & n7567 ) ;
  assign n7569 = n2733 ^ n1804 ^ x21 ;
  assign n7570 = n7569 ^ n5930 ^ n5226 ;
  assign n7578 = n7328 ^ n4043 ^ n3805 ;
  assign n7579 = ( ~n1095 & n1290 ) | ( ~n1095 & n7578 ) | ( n1290 & n7578 ) ;
  assign n7580 = ~n1317 & n1383 ;
  assign n7581 = ~n7579 & n7580 ;
  assign n7582 = n5961 ^ n1798 ^ 1'b0 ;
  assign n7583 = n7581 | n7582 ;
  assign n7571 = ( n760 & n2711 ) | ( n760 & n5800 ) | ( n2711 & n5800 ) ;
  assign n7572 = n7571 ^ n5073 ^ n3062 ;
  assign n7573 = n7204 | n7572 ;
  assign n7574 = n6313 & ~n7573 ;
  assign n7575 = n7574 ^ n5552 ^ n154 ;
  assign n7576 = n7575 ^ n4578 ^ 1'b0 ;
  assign n7577 = ~n2864 & n7576 ;
  assign n7584 = n7583 ^ n7577 ^ n2053 ;
  assign n7588 = ( x113 & ~n3396 ) | ( x113 & n4590 ) | ( ~n3396 & n4590 ) ;
  assign n7589 = n7588 ^ n4028 ^ n1726 ;
  assign n7590 = n7589 ^ n2333 ^ n1939 ;
  assign n7585 = n4321 ^ n562 ^ n497 ;
  assign n7586 = n7585 ^ n7049 ^ n2397 ;
  assign n7587 = n5657 & ~n7586 ;
  assign n7591 = n7590 ^ n7587 ^ 1'b0 ;
  assign n7592 = n5407 ^ n3981 ^ n639 ;
  assign n7593 = ( ~n165 & n1276 ) | ( ~n165 & n7592 ) | ( n1276 & n7592 ) ;
  assign n7594 = ~n348 & n5979 ;
  assign n7595 = ~n1146 & n7594 ;
  assign n7596 = n3179 ^ n1873 ^ 1'b0 ;
  assign n7597 = n6076 & n7596 ;
  assign n7598 = n7597 ^ n7450 ^ 1'b0 ;
  assign n7599 = ( ~n1685 & n2621 ) | ( ~n1685 & n3296 ) | ( n2621 & n3296 ) ;
  assign n7600 = n7599 ^ n1757 ^ n908 ;
  assign n7601 = ( n2084 & n7598 ) | ( n2084 & n7600 ) | ( n7598 & n7600 ) ;
  assign n7602 = ( x27 & n1324 ) | ( x27 & n7601 ) | ( n1324 & n7601 ) ;
  assign n7604 = n7212 ^ n2473 ^ 1'b0 ;
  assign n7605 = n4748 & ~n7604 ;
  assign n7603 = n5308 ^ n4160 ^ n404 ;
  assign n7606 = n7605 ^ n7603 ^ n3626 ;
  assign n7609 = n7290 ^ n3794 ^ 1'b0 ;
  assign n7607 = ( n1494 & n1799 ) | ( n1494 & ~n1981 ) | ( n1799 & ~n1981 ) ;
  assign n7608 = n3117 & n7607 ;
  assign n7610 = n7609 ^ n7608 ^ n435 ;
  assign n7611 = ( ~n1904 & n4975 ) | ( ~n1904 & n7610 ) | ( n4975 & n7610 ) ;
  assign n7612 = ( ~n153 & n2041 ) | ( ~n153 & n2387 ) | ( n2041 & n2387 ) ;
  assign n7613 = n4155 ^ n4079 ^ 1'b0 ;
  assign n7614 = ( n3254 & ~n7612 ) | ( n3254 & n7613 ) | ( ~n7612 & n7613 ) ;
  assign n7615 = n2331 ^ n1294 ^ n388 ;
  assign n7616 = n4263 ^ n2171 ^ 1'b0 ;
  assign n7618 = n5528 ^ n3070 ^ 1'b0 ;
  assign n7617 = n4992 ^ n1161 ^ x109 ;
  assign n7619 = n7618 ^ n7617 ^ n2132 ;
  assign n7620 = ( ~n510 & n7616 ) | ( ~n510 & n7619 ) | ( n7616 & n7619 ) ;
  assign n7621 = ~n2268 & n4374 ;
  assign n7622 = ~n5235 & n7621 ;
  assign n7623 = n7622 ^ n1296 ^ 1'b0 ;
  assign n7624 = n7620 & ~n7623 ;
  assign n7625 = ( n2976 & n7615 ) | ( n2976 & n7624 ) | ( n7615 & n7624 ) ;
  assign n7626 = n4266 ^ n3313 ^ n1914 ;
  assign n7627 = ~n6225 & n7626 ;
  assign n7628 = n7627 ^ n5547 ^ n2661 ;
  assign n7629 = ( n1708 & n5647 ) | ( n1708 & n7057 ) | ( n5647 & n7057 ) ;
  assign n7630 = n6103 ^ n354 ^ 1'b0 ;
  assign n7631 = n3302 & ~n7630 ;
  assign n7632 = n7631 ^ n6340 ^ n872 ;
  assign n7633 = ( n1567 & n2055 ) | ( n1567 & n7632 ) | ( n2055 & n7632 ) ;
  assign n7634 = ( ~n437 & n2424 ) | ( ~n437 & n2470 ) | ( n2424 & n2470 ) ;
  assign n7635 = ( n3066 & n3690 ) | ( n3066 & n3987 ) | ( n3690 & n3987 ) ;
  assign n7636 = ( n3149 & n7634 ) | ( n3149 & ~n7635 ) | ( n7634 & ~n7635 ) ;
  assign n7643 = n2997 ^ n1688 ^ n346 ;
  assign n7642 = n944 | n1612 ;
  assign n7644 = n7643 ^ n7642 ^ 1'b0 ;
  assign n7645 = n7644 ^ n3075 ^ 1'b0 ;
  assign n7646 = ( n495 & n3928 ) | ( n495 & ~n7645 ) | ( n3928 & ~n7645 ) ;
  assign n7637 = n5450 ^ n674 ^ 1'b0 ;
  assign n7638 = n760 & ~n7637 ;
  assign n7639 = ( n3545 & ~n3753 ) | ( n3545 & n7638 ) | ( ~n3753 & n7638 ) ;
  assign n7640 = n7639 ^ n3395 ^ 1'b0 ;
  assign n7641 = ~n6740 & n7640 ;
  assign n7647 = n7646 ^ n7641 ^ n959 ;
  assign n7648 = ( n5990 & n7636 ) | ( n5990 & ~n7647 ) | ( n7636 & ~n7647 ) ;
  assign n7649 = n392 & n760 ;
  assign n7650 = ~n4551 & n7649 ;
  assign n7651 = n3970 ^ n2274 ^ 1'b0 ;
  assign n7652 = ( ~n4976 & n7650 ) | ( ~n4976 & n7651 ) | ( n7650 & n7651 ) ;
  assign n7653 = n497 | n871 ;
  assign n7654 = n1264 | n2551 ;
  assign n7655 = n4829 ^ n4187 ^ n3185 ;
  assign n7656 = ~n7654 & n7655 ;
  assign n7657 = n7656 ^ n4866 ^ 1'b0 ;
  assign n7658 = ( n3072 & n7653 ) | ( n3072 & ~n7657 ) | ( n7653 & ~n7657 ) ;
  assign n7659 = n3525 ^ n3521 ^ 1'b0 ;
  assign n7660 = n5555 & n7659 ;
  assign n7661 = n7660 ^ n6645 ^ n2425 ;
  assign n7662 = n1452 & ~n7661 ;
  assign n7663 = n7662 ^ n2079 ^ 1'b0 ;
  assign n7664 = n7443 ^ n5779 ^ n5404 ;
  assign n7665 = n5460 ^ n597 ^ 1'b0 ;
  assign n7666 = ~n4014 & n7665 ;
  assign n7667 = n7666 ^ n4522 ^ 1'b0 ;
  assign n7668 = n1674 | n1977 ;
  assign n7669 = n5802 | n7668 ;
  assign n7670 = n7669 ^ n4303 ^ 1'b0 ;
  assign n7671 = n6229 ^ n917 ^ 1'b0 ;
  assign n7672 = n7671 ^ n4058 ^ n340 ;
  assign n7673 = n5263 ^ n3983 ^ 1'b0 ;
  assign n7674 = ( ~x93 & n2424 ) | ( ~x93 & n2760 ) | ( n2424 & n2760 ) ;
  assign n7675 = ~n275 & n3470 ;
  assign n7676 = n4439 | n7675 ;
  assign n7677 = n7676 ^ n4728 ^ 1'b0 ;
  assign n7678 = n5386 ^ n4725 ^ n4702 ;
  assign n7679 = ~n3515 & n7678 ;
  assign n7680 = ~n7677 & n7679 ;
  assign n7681 = n7674 & n7680 ;
  assign n7683 = n4189 ^ n680 ^ 1'b0 ;
  assign n7682 = n3528 ^ n390 ^ 1'b0 ;
  assign n7684 = n7683 ^ n7682 ^ n3200 ;
  assign n7694 = n2488 ^ n1886 ^ n1342 ;
  assign n7695 = n1786 & n7694 ;
  assign n7691 = n5624 ^ n5394 ^ n4034 ;
  assign n7692 = n7691 ^ n2815 ^ n1691 ;
  assign n7685 = n3642 ^ n345 ^ x17 ;
  assign n7686 = n4929 & ~n7685 ;
  assign n7687 = n4286 ^ n3845 ^ n1464 ;
  assign n7688 = ( n627 & n7686 ) | ( n627 & ~n7687 ) | ( n7686 & ~n7687 ) ;
  assign n7689 = n4022 ^ n2289 ^ 1'b0 ;
  assign n7690 = n7688 & ~n7689 ;
  assign n7693 = n7692 ^ n7690 ^ n1742 ;
  assign n7696 = n7695 ^ n7693 ^ n209 ;
  assign n7697 = n6521 ^ n2754 ^ 1'b0 ;
  assign n7698 = n4326 & ~n7697 ;
  assign n7699 = ~n5777 & n7698 ;
  assign n7700 = ( n3088 & ~n5769 ) | ( n3088 & n7699 ) | ( ~n5769 & n7699 ) ;
  assign n7701 = n4608 | n7632 ;
  assign n7702 = n2487 & ~n7701 ;
  assign n7703 = n3700 ^ n1623 ^ n698 ;
  assign n7704 = n6591 ^ n6437 ^ n4486 ;
  assign n7705 = ( n4251 & ~n4950 ) | ( n4251 & n5024 ) | ( ~n4950 & n5024 ) ;
  assign n7706 = ( n4218 & ~n7704 ) | ( n4218 & n7705 ) | ( ~n7704 & n7705 ) ;
  assign n7707 = ( n1612 & ~n4905 ) | ( n1612 & n7706 ) | ( ~n4905 & n7706 ) ;
  assign n7708 = n4155 & ~n4400 ;
  assign n7709 = n7708 ^ n6858 ^ 1'b0 ;
  assign n7710 = n7709 ^ n3634 ^ n3402 ;
  assign n7711 = n1969 & n7710 ;
  assign n7712 = n4949 & n7711 ;
  assign n7713 = n2358 ^ n801 ^ n595 ;
  assign n7714 = n7713 ^ n2465 ^ 1'b0 ;
  assign n7715 = n4453 ^ n4444 ^ n2482 ;
  assign n7716 = n3316 & ~n7715 ;
  assign n7717 = n5494 ^ n4506 ^ 1'b0 ;
  assign n7718 = n7716 | n7717 ;
  assign n7719 = ( n1362 & ~n7714 ) | ( n1362 & n7718 ) | ( ~n7714 & n7718 ) ;
  assign n7721 = ~n3483 & n4579 ;
  assign n7720 = n205 | n5176 ;
  assign n7722 = n7721 ^ n7720 ^ 1'b0 ;
  assign n7723 = ~n2021 & n3516 ;
  assign n7724 = n7723 ^ n3335 ^ 1'b0 ;
  assign n7725 = ( ~n4828 & n5417 ) | ( ~n4828 & n7724 ) | ( n5417 & n7724 ) ;
  assign n7726 = n1890 ^ x91 ^ 1'b0 ;
  assign n7727 = ~n1041 & n5622 ;
  assign n7728 = n7727 ^ n5705 ^ n4167 ;
  assign n7730 = n1723 ^ n1251 ^ n1249 ;
  assign n7729 = ~n2891 & n7257 ;
  assign n7731 = n7730 ^ n7729 ^ 1'b0 ;
  assign n7732 = ( n7726 & n7728 ) | ( n7726 & ~n7731 ) | ( n7728 & ~n7731 ) ;
  assign n7738 = n7218 ^ n4525 ^ n1883 ;
  assign n7733 = n4520 ^ n2697 ^ 1'b0 ;
  assign n7734 = n5335 ^ n4364 ^ 1'b0 ;
  assign n7735 = n829 & n7734 ;
  assign n7736 = ( ~n4286 & n6459 ) | ( ~n4286 & n7735 ) | ( n6459 & n7735 ) ;
  assign n7737 = n7733 | n7736 ;
  assign n7739 = n7738 ^ n7737 ^ n1799 ;
  assign n7740 = ( n3217 & n4990 ) | ( n3217 & n7739 ) | ( n4990 & n7739 ) ;
  assign n7741 = n903 | n4418 ;
  assign n7742 = n7741 ^ n5838 ^ n5636 ;
  assign n7743 = n7742 ^ n5700 ^ 1'b0 ;
  assign n7744 = ( n1065 & ~n1704 ) | ( n1065 & n2088 ) | ( ~n1704 & n2088 ) ;
  assign n7745 = n2210 & ~n2286 ;
  assign n7746 = n2891 & n7745 ;
  assign n7747 = n2751 & ~n7746 ;
  assign n7748 = ~n3049 & n7747 ;
  assign n7749 = ~n7744 & n7748 ;
  assign n7750 = n7373 ^ n5270 ^ n4577 ;
  assign n7751 = n1928 & ~n4116 ;
  assign n7759 = n254 & n3435 ;
  assign n7760 = n7759 ^ n868 ^ 1'b0 ;
  assign n7761 = ( n1471 & n5488 ) | ( n1471 & ~n7760 ) | ( n5488 & ~n7760 ) ;
  assign n7762 = n7761 ^ n5526 ^ n3218 ;
  assign n7763 = n7762 ^ n1484 ^ n458 ;
  assign n7752 = n3677 ^ n3224 ^ n1419 ;
  assign n7753 = n7752 ^ n4243 ^ n964 ;
  assign n7754 = n5281 ^ n3514 ^ n3345 ;
  assign n7755 = n2245 & ~n5645 ;
  assign n7756 = ~n3352 & n7755 ;
  assign n7757 = n3833 | n7756 ;
  assign n7758 = ( n7753 & ~n7754 ) | ( n7753 & n7757 ) | ( ~n7754 & n7757 ) ;
  assign n7764 = n7763 ^ n7758 ^ n4847 ;
  assign n7765 = n7521 ^ n1126 ^ x99 ;
  assign n7766 = ( n294 & n1252 ) | ( n294 & n1469 ) | ( n1252 & n1469 ) ;
  assign n7767 = n7766 ^ n6967 ^ n4243 ;
  assign n7768 = n5697 ^ n4202 ^ 1'b0 ;
  assign n7773 = ( n1360 & n2812 ) | ( n1360 & ~n4240 ) | ( n2812 & ~n4240 ) ;
  assign n7770 = n3257 ^ n788 ^ 1'b0 ;
  assign n7771 = ~n860 & n7770 ;
  assign n7769 = ( n3860 & ~n6156 ) | ( n3860 & n7744 ) | ( ~n6156 & n7744 ) ;
  assign n7772 = n7771 ^ n7769 ^ n2211 ;
  assign n7774 = n7773 ^ n7772 ^ n7324 ;
  assign n7775 = ( n1677 & ~n2024 ) | ( n1677 & n4961 ) | ( ~n2024 & n4961 ) ;
  assign n7776 = ( n5955 & ~n7198 ) | ( n5955 & n7775 ) | ( ~n7198 & n7775 ) ;
  assign n7777 = n7776 ^ n4259 ^ n4255 ;
  assign n7780 = n6308 ^ n4587 ^ n414 ;
  assign n7778 = n3927 ^ n3794 ^ 1'b0 ;
  assign n7779 = n5458 & ~n7778 ;
  assign n7781 = n7780 ^ n7779 ^ n3079 ;
  assign n7782 = n1798 & ~n7781 ;
  assign n7783 = n7782 ^ n5412 ^ 1'b0 ;
  assign n7792 = n4398 ^ n873 ^ n396 ;
  assign n7787 = n2746 ^ n581 ^ 1'b0 ;
  assign n7788 = n4668 & ~n7787 ;
  assign n7789 = n4752 ^ n4093 ^ 1'b0 ;
  assign n7790 = n7788 & ~n7789 ;
  assign n7791 = n7790 ^ n4311 ^ 1'b0 ;
  assign n7784 = ( x61 & ~n462 ) | ( x61 & n1944 ) | ( ~n462 & n1944 ) ;
  assign n7785 = n7784 ^ n4566 ^ 1'b0 ;
  assign n7786 = n5681 & n7785 ;
  assign n7793 = n7792 ^ n7791 ^ n7786 ;
  assign n7798 = ( n161 & ~n3379 ) | ( n161 & n3882 ) | ( ~n3379 & n3882 ) ;
  assign n7797 = n2754 | n5693 ;
  assign n7799 = n7798 ^ n7797 ^ 1'b0 ;
  assign n7795 = ( n168 & n2783 ) | ( n168 & ~n3061 ) | ( n2783 & ~n3061 ) ;
  assign n7794 = n5964 ^ n3610 ^ 1'b0 ;
  assign n7796 = n7795 ^ n7794 ^ n1848 ;
  assign n7800 = n7799 ^ n7796 ^ n817 ;
  assign n7801 = n2689 ^ n768 ^ 1'b0 ;
  assign n7802 = n994 | n7801 ;
  assign n7803 = n7802 ^ n6931 ^ n2819 ;
  assign n7804 = n2960 ^ n2931 ^ 1'b0 ;
  assign n7805 = ( n2766 & n6413 ) | ( n2766 & n7804 ) | ( n6413 & n7804 ) ;
  assign n7806 = n4636 ^ n4036 ^ n3912 ;
  assign n7807 = n7806 ^ n7741 ^ 1'b0 ;
  assign n7808 = n6192 | n7807 ;
  assign n7809 = n270 & ~n634 ;
  assign n7810 = n5256 & n7809 ;
  assign n7811 = n7810 ^ n5394 ^ x107 ;
  assign n7812 = n4125 ^ n2640 ^ 1'b0 ;
  assign n7813 = n7812 ^ n4042 ^ n1768 ;
  assign n7814 = n4224 | n7813 ;
  assign n7815 = ( n5200 & n7811 ) | ( n5200 & ~n7814 ) | ( n7811 & ~n7814 ) ;
  assign n7816 = n5841 ^ n1377 ^ n1271 ;
  assign n7817 = ( n1205 & n7057 ) | ( n1205 & ~n7816 ) | ( n7057 & ~n7816 ) ;
  assign n7818 = n7817 ^ n6547 ^ n2254 ;
  assign n7819 = n5662 ^ n2982 ^ n889 ;
  assign n7820 = n7819 ^ n6953 ^ n3133 ;
  assign n7821 = ( n2781 & ~n3816 ) | ( n2781 & n5261 ) | ( ~n3816 & n5261 ) ;
  assign n7822 = ( n3515 & n5142 ) | ( n3515 & ~n7821 ) | ( n5142 & ~n7821 ) ;
  assign n7823 = ( n6822 & n7820 ) | ( n6822 & ~n7822 ) | ( n7820 & ~n7822 ) ;
  assign n7824 = n6241 ^ n2279 ^ n589 ;
  assign n7825 = ( n188 & ~n4870 ) | ( n188 & n7824 ) | ( ~n4870 & n7824 ) ;
  assign n7826 = n953 ^ n862 ^ 1'b0 ;
  assign n7827 = n7826 ^ n724 ^ n722 ;
  assign n7828 = x104 & n7827 ;
  assign n7829 = n7828 ^ n3876 ^ 1'b0 ;
  assign n7830 = n2777 ^ n2704 ^ 1'b0 ;
  assign n7831 = n7830 ^ n4196 ^ n4166 ;
  assign n7832 = ( ~n6601 & n6793 ) | ( ~n6601 & n7831 ) | ( n6793 & n7831 ) ;
  assign n7833 = ( ~n252 & n1361 ) | ( ~n252 & n7832 ) | ( n1361 & n7832 ) ;
  assign n7834 = ( n1674 & ~n7829 ) | ( n1674 & n7833 ) | ( ~n7829 & n7833 ) ;
  assign n7835 = n3331 ^ n1476 ^ 1'b0 ;
  assign n7836 = n7428 ^ n6295 ^ n3685 ;
  assign n7837 = n3182 ^ n636 ^ x48 ;
  assign n7838 = ( n1470 & ~n3319 ) | ( n1470 & n7837 ) | ( ~n3319 & n7837 ) ;
  assign n7839 = ( n336 & ~n7716 ) | ( n336 & n7838 ) | ( ~n7716 & n7838 ) ;
  assign n7840 = n7839 ^ n6285 ^ n2158 ;
  assign n7841 = ( n1245 & ~n2493 ) | ( n1245 & n7840 ) | ( ~n2493 & n7840 ) ;
  assign n7842 = ( n306 & n2783 ) | ( n306 & n3213 ) | ( n2783 & n3213 ) ;
  assign n7843 = n5239 & ~n7842 ;
  assign n7844 = n1574 & n7843 ;
  assign n7852 = ( x88 & ~n2074 ) | ( x88 & n5783 ) | ( ~n2074 & n5783 ) ;
  assign n7846 = ( ~n2995 & n5264 ) | ( ~n2995 & n6940 ) | ( n5264 & n6940 ) ;
  assign n7847 = ( n1783 & n3210 ) | ( n1783 & ~n3525 ) | ( n3210 & ~n3525 ) ;
  assign n7848 = ( n681 & n4109 ) | ( n681 & ~n5232 ) | ( n4109 & ~n5232 ) ;
  assign n7849 = ( n1008 & n7847 ) | ( n1008 & ~n7848 ) | ( n7847 & ~n7848 ) ;
  assign n7850 = ( n1864 & n6712 ) | ( n1864 & n7849 ) | ( n6712 & n7849 ) ;
  assign n7851 = n7846 & n7850 ;
  assign n7853 = n7852 ^ n7851 ^ n7569 ;
  assign n7845 = n6875 & ~n7308 ;
  assign n7854 = n7853 ^ n7845 ^ 1'b0 ;
  assign n7858 = n140 & ~n556 ;
  assign n7859 = n7858 ^ n491 ^ 1'b0 ;
  assign n7860 = n7859 ^ n6691 ^ 1'b0 ;
  assign n7855 = ( n1682 & n2506 ) | ( n1682 & ~n3017 ) | ( n2506 & ~n3017 ) ;
  assign n7856 = ( n5235 & n7336 ) | ( n5235 & n7855 ) | ( n7336 & n7855 ) ;
  assign n7857 = n5434 & ~n7856 ;
  assign n7861 = n7860 ^ n7857 ^ 1'b0 ;
  assign n7866 = n4945 ^ n943 ^ 1'b0 ;
  assign n7867 = n7310 & ~n7866 ;
  assign n7862 = ( n731 & ~n1268 ) | ( n731 & n1421 ) | ( ~n1268 & n1421 ) ;
  assign n7863 = ( ~n249 & n2076 ) | ( ~n249 & n7862 ) | ( n2076 & n7862 ) ;
  assign n7864 = n7863 ^ n5145 ^ 1'b0 ;
  assign n7865 = n277 & n7864 ;
  assign n7868 = n7867 ^ n7865 ^ n7763 ;
  assign n7869 = n1617 & n7868 ;
  assign n7870 = ( ~n3669 & n5357 ) | ( ~n3669 & n7869 ) | ( n5357 & n7869 ) ;
  assign n7871 = n7870 ^ n908 ^ 1'b0 ;
  assign n7872 = n935 & ~n7871 ;
  assign n7878 = n4038 & ~n7852 ;
  assign n7873 = ( n1380 & n3706 ) | ( n1380 & n4597 ) | ( n3706 & n4597 ) ;
  assign n7874 = ( n5279 & n7451 ) | ( n5279 & ~n7873 ) | ( n7451 & ~n7873 ) ;
  assign n7875 = n7762 & n7874 ;
  assign n7876 = n7875 ^ n4480 ^ 1'b0 ;
  assign n7877 = n1237 | n7876 ;
  assign n7879 = n7878 ^ n7877 ^ 1'b0 ;
  assign n7880 = n952 & n1798 ;
  assign n7881 = n7880 ^ n3450 ^ 1'b0 ;
  assign n7882 = ( n168 & n5994 ) | ( n168 & ~n7881 ) | ( n5994 & ~n7881 ) ;
  assign n7887 = n6886 ^ n5280 ^ n964 ;
  assign n7888 = n7887 ^ n3258 ^ n471 ;
  assign n7889 = n3983 & n7888 ;
  assign n7885 = n2615 ^ n2106 ^ n383 ;
  assign n7886 = n7885 ^ n978 ^ 1'b0 ;
  assign n7890 = n7889 ^ n7886 ^ n6275 ;
  assign n7891 = ( n4812 & ~n7496 ) | ( n4812 & n7890 ) | ( ~n7496 & n7890 ) ;
  assign n7883 = n3361 ^ n3094 ^ n2480 ;
  assign n7884 = ( n2793 & ~n5814 ) | ( n2793 & n7883 ) | ( ~n5814 & n7883 ) ;
  assign n7892 = n7891 ^ n7884 ^ n5382 ;
  assign n7895 = n2307 ^ n2123 ^ 1'b0 ;
  assign n7894 = n5364 ^ n901 ^ 1'b0 ;
  assign n7893 = ( ~n772 & n1088 ) | ( ~n772 & n5060 ) | ( n1088 & n5060 ) ;
  assign n7896 = n7895 ^ n7894 ^ n7893 ;
  assign n7898 = ( n352 & n3791 ) | ( n352 & n3972 ) | ( n3791 & n3972 ) ;
  assign n7897 = n4295 ^ n1610 ^ n1581 ;
  assign n7899 = n7898 ^ n7897 ^ n3646 ;
  assign n7900 = n2606 ^ n899 ^ 1'b0 ;
  assign n7901 = n7899 & ~n7900 ;
  assign n7902 = n7896 & n7901 ;
  assign n7903 = n3100 | n3124 ;
  assign n7904 = ( n768 & n4059 ) | ( n768 & n5702 ) | ( n4059 & n5702 ) ;
  assign n7905 = n4429 & ~n7613 ;
  assign n7906 = ( n7903 & n7904 ) | ( n7903 & n7905 ) | ( n7904 & n7905 ) ;
  assign n7907 = ( ~n3177 & n4782 ) | ( ~n3177 & n7906 ) | ( n4782 & n7906 ) ;
  assign n7908 = ( n896 & n3015 ) | ( n896 & n7020 ) | ( n3015 & n7020 ) ;
  assign n7909 = ( n414 & ~n2806 ) | ( n414 & n2830 ) | ( ~n2806 & n2830 ) ;
  assign n7910 = ( ~n357 & n7908 ) | ( ~n357 & n7909 ) | ( n7908 & n7909 ) ;
  assign n7911 = n7910 ^ n3642 ^ n2746 ;
  assign n7912 = n4321 & ~n7911 ;
  assign n7913 = n2787 & n7912 ;
  assign n7914 = ( n1144 & ~n1207 ) | ( n1144 & n3316 ) | ( ~n1207 & n3316 ) ;
  assign n7915 = n7914 ^ n1411 ^ 1'b0 ;
  assign n7916 = n4548 & ~n7915 ;
  assign n7917 = ( n3114 & n6419 ) | ( n3114 & n7916 ) | ( n6419 & n7916 ) ;
  assign n7918 = ( ~n852 & n1171 ) | ( ~n852 & n2556 ) | ( n1171 & n2556 ) ;
  assign n7919 = n7918 ^ n2932 ^ n2546 ;
  assign n7920 = n7919 ^ n1124 ^ 1'b0 ;
  assign n7921 = n7917 & n7920 ;
  assign n7922 = n6197 ^ n3704 ^ n548 ;
  assign n7923 = n7922 ^ n1675 ^ n1027 ;
  assign n7924 = n7923 ^ n5640 ^ n3919 ;
  assign n7926 = n6397 ^ n541 ^ 1'b0 ;
  assign n7927 = n685 | n7926 ;
  assign n7928 = n7927 ^ n2746 ^ 1'b0 ;
  assign n7925 = ( n3534 & n7147 ) | ( n3534 & n7353 ) | ( n7147 & n7353 ) ;
  assign n7929 = n7928 ^ n7925 ^ 1'b0 ;
  assign n7930 = ( ~n5186 & n7924 ) | ( ~n5186 & n7929 ) | ( n7924 & n7929 ) ;
  assign n7931 = n3623 ^ n1523 ^ n167 ;
  assign n7932 = ( n1052 & n2050 ) | ( n1052 & ~n4068 ) | ( n2050 & ~n4068 ) ;
  assign n7933 = n7932 ^ n2882 ^ n2654 ;
  assign n7934 = n1853 | n7933 ;
  assign n7935 = n7931 & ~n7934 ;
  assign n7939 = ~n5283 & n7201 ;
  assign n7936 = n7219 ^ n3382 ^ 1'b0 ;
  assign n7937 = n7936 ^ n5719 ^ n2658 ;
  assign n7938 = n2122 & n7937 ;
  assign n7940 = n7939 ^ n7938 ^ n1632 ;
  assign n7941 = n1549 & n5033 ;
  assign n7942 = n6686 & n7941 ;
  assign n7943 = n3087 ^ n1411 ^ 1'b0 ;
  assign n7944 = n7943 ^ n3172 ^ n1607 ;
  assign n7945 = ( n6352 & n7942 ) | ( n6352 & n7944 ) | ( n7942 & n7944 ) ;
  assign n7946 = ~n1012 & n6389 ;
  assign n7947 = n326 & n3486 ;
  assign n7948 = ~n7946 & n7947 ;
  assign n7952 = ( n752 & n2322 ) | ( n752 & ~n5252 ) | ( n2322 & ~n5252 ) ;
  assign n7949 = n3609 & n5926 ;
  assign n7950 = n7949 ^ x40 ^ 1'b0 ;
  assign n7951 = n1175 | n7950 ;
  assign n7953 = n7952 ^ n7951 ^ n5262 ;
  assign n7954 = n7953 ^ n7051 ^ n4728 ;
  assign n7955 = n2012 ^ n1892 ^ 1'b0 ;
  assign n7956 = n3119 & ~n7955 ;
  assign n7957 = n7956 ^ n4992 ^ n1550 ;
  assign n7958 = n7957 ^ n6306 ^ n3005 ;
  assign n7959 = ( n1805 & ~n1901 ) | ( n1805 & n2164 ) | ( ~n1901 & n2164 ) ;
  assign n7960 = ( n367 & n3983 ) | ( n367 & n7959 ) | ( n3983 & n7959 ) ;
  assign n7963 = ~n4728 & n5061 ;
  assign n7961 = n803 & ~n4287 ;
  assign n7962 = n5072 & n7961 ;
  assign n7964 = n7963 ^ n7962 ^ 1'b0 ;
  assign n7965 = ( ~n2839 & n7960 ) | ( ~n2839 & n7964 ) | ( n7960 & n7964 ) ;
  assign n7966 = n658 & ~n1552 ;
  assign n7967 = ( x13 & ~n1401 ) | ( x13 & n7966 ) | ( ~n1401 & n7966 ) ;
  assign n7968 = n7967 ^ n7959 ^ n440 ;
  assign n7969 = ( ~n2138 & n6627 ) | ( ~n2138 & n7968 ) | ( n6627 & n7968 ) ;
  assign n7970 = ( n7958 & n7965 ) | ( n7958 & n7969 ) | ( n7965 & n7969 ) ;
  assign n7971 = n2995 | n7675 ;
  assign n7972 = n742 & ~n7971 ;
  assign n7973 = n7972 ^ n4186 ^ x38 ;
  assign n7974 = ( ~n3297 & n4488 ) | ( ~n3297 & n7973 ) | ( n4488 & n7973 ) ;
  assign n7975 = n6043 ^ n2478 ^ n648 ;
  assign n7976 = n2144 & ~n4236 ;
  assign n7977 = n7975 & n7976 ;
  assign n7978 = n7974 & n7977 ;
  assign n7979 = n1411 ^ n806 ^ 1'b0 ;
  assign n7980 = n7979 ^ n5966 ^ n5282 ;
  assign n7981 = n4636 ^ n3734 ^ n3451 ;
  assign n7982 = n7980 | n7981 ;
  assign n7983 = n5111 & ~n7982 ;
  assign n7984 = n4326 ^ n2353 ^ x21 ;
  assign n7985 = ( n520 & n1600 ) | ( n520 & ~n2117 ) | ( n1600 & ~n2117 ) ;
  assign n7986 = ( n798 & n4097 ) | ( n798 & n7985 ) | ( n4097 & n7985 ) ;
  assign n7987 = n3452 | n4127 ;
  assign n7988 = ~n5850 & n7987 ;
  assign n7989 = ( n7984 & n7986 ) | ( n7984 & ~n7988 ) | ( n7986 & ~n7988 ) ;
  assign n7990 = ( n761 & n4166 ) | ( n761 & ~n5269 ) | ( n4166 & ~n5269 ) ;
  assign n7991 = ( n2220 & ~n3215 ) | ( n2220 & n5924 ) | ( ~n3215 & n5924 ) ;
  assign n7992 = ( n2342 & n7990 ) | ( n2342 & n7991 ) | ( n7990 & n7991 ) ;
  assign n7993 = n2378 ^ n528 ^ 1'b0 ;
  assign n7994 = n5814 ^ n5326 ^ n4318 ;
  assign n7995 = n2716 | n5908 ;
  assign n7996 = n634 & ~n7995 ;
  assign n7997 = ( n7993 & n7994 ) | ( n7993 & ~n7996 ) | ( n7994 & ~n7996 ) ;
  assign n8004 = n7176 ^ n2667 ^ n2512 ;
  assign n8000 = ( x117 & n852 ) | ( x117 & n1753 ) | ( n852 & n1753 ) ;
  assign n8001 = ~n6414 & n8000 ;
  assign n8002 = ~n1962 & n8001 ;
  assign n7998 = ( x49 & ~x91 ) | ( x49 & n990 ) | ( ~x91 & n990 ) ;
  assign n7999 = n7998 ^ n2676 ^ x73 ;
  assign n8003 = n8002 ^ n7999 ^ n1400 ;
  assign n8005 = n8004 ^ n8003 ^ n4073 ;
  assign n8006 = n2422 ^ n505 ^ 1'b0 ;
  assign n8007 = n8006 ^ n6942 ^ n954 ;
  assign n8008 = n2854 | n6776 ;
  assign n8009 = ~n2893 & n5017 ;
  assign n8010 = n8009 ^ n3047 ^ n1586 ;
  assign n8011 = ( n3704 & n8008 ) | ( n3704 & ~n8010 ) | ( n8008 & ~n8010 ) ;
  assign n8012 = ( ~n179 & n1470 ) | ( ~n179 & n5259 ) | ( n1470 & n5259 ) ;
  assign n8013 = ( n1983 & n2494 ) | ( n1983 & ~n8012 ) | ( n2494 & ~n8012 ) ;
  assign n8014 = n6280 ^ n4406 ^ n3331 ;
  assign n8015 = ~n4813 & n8014 ;
  assign n8016 = ~n2722 & n8015 ;
  assign n8017 = ( n458 & n636 ) | ( n458 & n8016 ) | ( n636 & n8016 ) ;
  assign n8018 = n8017 ^ n3986 ^ n1077 ;
  assign n8019 = ( ~n1652 & n3015 ) | ( ~n1652 & n8018 ) | ( n3015 & n8018 ) ;
  assign n8020 = n6454 & ~n8019 ;
  assign n8021 = n3337 ^ n2856 ^ 1'b0 ;
  assign n8022 = ~n3063 & n8021 ;
  assign n8023 = n3653 ^ n3646 ^ 1'b0 ;
  assign n8024 = n8023 ^ n4751 ^ n4025 ;
  assign n8025 = ( ~n129 & n8022 ) | ( ~n129 & n8024 ) | ( n8022 & n8024 ) ;
  assign n8026 = n6592 ^ n1262 ^ 1'b0 ;
  assign n8027 = n4258 ^ n641 ^ 1'b0 ;
  assign n8028 = ( n5966 & ~n8026 ) | ( n5966 & n8027 ) | ( ~n8026 & n8027 ) ;
  assign n8039 = ( ~n576 & n985 ) | ( ~n576 & n2579 ) | ( n985 & n2579 ) ;
  assign n8040 = n8039 ^ n5560 ^ 1'b0 ;
  assign n8041 = n1006 & n8040 ;
  assign n8042 = ( n1675 & n2116 ) | ( n1675 & n8041 ) | ( n2116 & n8041 ) ;
  assign n8043 = n8042 ^ n5077 ^ n980 ;
  assign n8044 = n8043 ^ n2954 ^ n1970 ;
  assign n8037 = ~n2623 & n3485 ;
  assign n8038 = n8037 ^ n6962 ^ 1'b0 ;
  assign n8035 = n3607 ^ n2577 ^ x36 ;
  assign n8032 = n1740 ^ n1452 ^ n905 ;
  assign n8029 = ( ~n1627 & n1991 ) | ( ~n1627 & n2061 ) | ( n1991 & n2061 ) ;
  assign n8030 = n3313 & ~n8029 ;
  assign n8031 = ~n3012 & n8030 ;
  assign n8033 = n8032 ^ n8031 ^ n3053 ;
  assign n8034 = ( n248 & ~n3214 ) | ( n248 & n8033 ) | ( ~n3214 & n8033 ) ;
  assign n8036 = n8035 ^ n8034 ^ 1'b0 ;
  assign n8045 = n8044 ^ n8038 ^ n8036 ;
  assign n8046 = n1853 ^ n248 ^ 1'b0 ;
  assign n8047 = n1857 & ~n8046 ;
  assign n8048 = ~n723 & n8047 ;
  assign n8049 = n5661 & n8048 ;
  assign n8051 = ( n1290 & ~n3420 ) | ( n1290 & n7842 ) | ( ~n3420 & n7842 ) ;
  assign n8050 = n7031 ^ n1838 ^ n1104 ;
  assign n8052 = n8051 ^ n8050 ^ 1'b0 ;
  assign n8053 = ( n3374 & n8049 ) | ( n3374 & ~n8052 ) | ( n8049 & ~n8052 ) ;
  assign n8054 = ( n735 & n2178 ) | ( n735 & n4092 ) | ( n2178 & n4092 ) ;
  assign n8055 = n8054 ^ n1916 ^ 1'b0 ;
  assign n8056 = ~n1212 & n8055 ;
  assign n8057 = n5687 & ~n8056 ;
  assign n8058 = ( n624 & n1021 ) | ( n624 & ~n3030 ) | ( n1021 & ~n3030 ) ;
  assign n8059 = n2437 & ~n8058 ;
  assign n8060 = n8057 & n8059 ;
  assign n8061 = n8060 ^ n4959 ^ n4597 ;
  assign n8062 = n2004 ^ n570 ^ 1'b0 ;
  assign n8063 = n2114 & n8062 ;
  assign n8064 = ( ~n4079 & n5815 ) | ( ~n4079 & n8063 ) | ( n5815 & n8063 ) ;
  assign n8065 = n4107 ^ n655 ^ 1'b0 ;
  assign n8066 = n6325 & ~n8065 ;
  assign n8067 = n8066 ^ n6685 ^ 1'b0 ;
  assign n8068 = n8067 ^ n4178 ^ n3353 ;
  assign n8074 = ( ~n581 & n3596 ) | ( ~n581 & n7190 ) | ( n3596 & n7190 ) ;
  assign n8071 = n4514 & n6024 ;
  assign n8069 = ( n326 & n4254 ) | ( n326 & ~n5919 ) | ( n4254 & ~n5919 ) ;
  assign n8070 = n3876 & ~n8069 ;
  assign n8072 = n8071 ^ n8070 ^ 1'b0 ;
  assign n8073 = n6108 & ~n8072 ;
  assign n8075 = n8074 ^ n8073 ^ n5142 ;
  assign n8076 = ( n1271 & n3626 ) | ( n1271 & n8075 ) | ( n3626 & n8075 ) ;
  assign n8077 = n1300 ^ n1250 ^ n717 ;
  assign n8078 = n4581 ^ n3146 ^ n1781 ;
  assign n8079 = n8077 & ~n8078 ;
  assign n8086 = n1248 ^ x38 ^ 1'b0 ;
  assign n8087 = n6229 & ~n8086 ;
  assign n8084 = ( n1888 & n7393 ) | ( n1888 & ~n7752 ) | ( n7393 & ~n7752 ) ;
  assign n8085 = n7445 & ~n8084 ;
  assign n8080 = ( n734 & ~n2649 ) | ( n734 & n2683 ) | ( ~n2649 & n2683 ) ;
  assign n8081 = n1908 & ~n8080 ;
  assign n8082 = n8081 ^ n4780 ^ 1'b0 ;
  assign n8083 = n3242 & n8082 ;
  assign n8088 = n8087 ^ n8085 ^ n8083 ;
  assign n8089 = n8088 ^ n1972 ^ n1516 ;
  assign n8090 = ( n2417 & n3003 ) | ( n2417 & ~n5454 ) | ( n3003 & ~n5454 ) ;
  assign n8100 = n4900 ^ n4663 ^ 1'b0 ;
  assign n8091 = n2978 & n4202 ;
  assign n8092 = n8091 ^ n3115 ^ 1'b0 ;
  assign n8093 = n6256 & n8092 ;
  assign n8094 = n8093 ^ n4125 ^ 1'b0 ;
  assign n8095 = n5163 ^ n1040 ^ 1'b0 ;
  assign n8096 = n7016 | n8095 ;
  assign n8097 = n6314 ^ n1504 ^ n146 ;
  assign n8098 = ( ~n1792 & n5742 ) | ( ~n1792 & n8097 ) | ( n5742 & n8097 ) ;
  assign n8099 = ( n8094 & n8096 ) | ( n8094 & ~n8098 ) | ( n8096 & ~n8098 ) ;
  assign n8101 = n8100 ^ n8099 ^ n4378 ;
  assign n8102 = n7078 ^ n5400 ^ n4640 ;
  assign n8103 = n395 | n7780 ;
  assign n8104 = n1844 & ~n8103 ;
  assign n8105 = n8104 ^ n5216 ^ n5096 ;
  assign n8106 = ( ~n3536 & n5030 ) | ( ~n3536 & n8105 ) | ( n5030 & n8105 ) ;
  assign n8107 = n8106 ^ n2463 ^ x85 ;
  assign n8108 = n8107 ^ n381 ^ 1'b0 ;
  assign n8109 = n6501 & n8108 ;
  assign n8110 = ( n798 & n6358 ) | ( n798 & n8109 ) | ( n6358 & n8109 ) ;
  assign n8111 = n2690 ^ n1982 ^ 1'b0 ;
  assign n8112 = ( ~n1477 & n1890 ) | ( ~n1477 & n7832 ) | ( n1890 & n7832 ) ;
  assign n8113 = n994 & ~n2912 ;
  assign n8114 = n6921 & ~n8113 ;
  assign n8115 = ~n7320 & n8114 ;
  assign n8116 = n5786 ^ n2472 ^ 1'b0 ;
  assign n8117 = n2430 & ~n8116 ;
  assign n8148 = n3648 ^ n508 ^ n256 ;
  assign n8149 = ( ~n2914 & n3445 ) | ( ~n2914 & n8148 ) | ( n3445 & n8148 ) ;
  assign n8147 = n4166 ^ n2009 ^ n1196 ;
  assign n8136 = ( n603 & ~n1308 ) | ( n603 & n1527 ) | ( ~n1308 & n1527 ) ;
  assign n8137 = ( n2719 & n7543 ) | ( n2719 & ~n8136 ) | ( n7543 & ~n8136 ) ;
  assign n8138 = ( n2860 & n3176 ) | ( n2860 & n6939 ) | ( n3176 & n6939 ) ;
  assign n8139 = ( n1841 & n2874 ) | ( n1841 & ~n8138 ) | ( n2874 & ~n8138 ) ;
  assign n8140 = ( n4883 & n8137 ) | ( n4883 & ~n8139 ) | ( n8137 & ~n8139 ) ;
  assign n8141 = ~n951 & n3195 ;
  assign n8142 = n8141 ^ n2827 ^ 1'b0 ;
  assign n8143 = ( ~n319 & n5494 ) | ( ~n319 & n8142 ) | ( n5494 & n8142 ) ;
  assign n8144 = ~n5254 & n8143 ;
  assign n8145 = n8140 | n8144 ;
  assign n8133 = n5243 | n5543 ;
  assign n8134 = n1287 | n8133 ;
  assign n8129 = ( ~n2272 & n2403 ) | ( ~n2272 & n6212 ) | ( n2403 & n6212 ) ;
  assign n8130 = n1913 & ~n8129 ;
  assign n8126 = n2653 & n5565 ;
  assign n8127 = ~n810 & n8126 ;
  assign n8128 = n570 & ~n8127 ;
  assign n8131 = n8130 ^ n8128 ^ n3667 ;
  assign n8124 = ( n1445 & ~n1592 ) | ( n1445 & n4603 ) | ( ~n1592 & n4603 ) ;
  assign n8125 = n8124 ^ n972 ^ 1'b0 ;
  assign n8132 = n8131 ^ n8125 ^ n2394 ;
  assign n8135 = n8134 ^ n8132 ^ n4657 ;
  assign n8118 = ( ~n358 & n2891 ) | ( ~n358 & n2958 ) | ( n2891 & n2958 ) ;
  assign n8119 = ( ~n1826 & n5131 ) | ( ~n1826 & n8118 ) | ( n5131 & n8118 ) ;
  assign n8120 = ( n2026 & n5281 ) | ( n2026 & n7704 ) | ( n5281 & n7704 ) ;
  assign n8121 = ( ~n2062 & n3766 ) | ( ~n2062 & n8120 ) | ( n3766 & n8120 ) ;
  assign n8122 = n8121 ^ n2437 ^ n284 ;
  assign n8123 = ( ~n2855 & n8119 ) | ( ~n2855 & n8122 ) | ( n8119 & n8122 ) ;
  assign n8146 = n8145 ^ n8135 ^ n8123 ;
  assign n8150 = n8149 ^ n8147 ^ n8146 ;
  assign n8151 = n6686 ^ n3070 ^ n2667 ;
  assign n8152 = n3518 | n3572 ;
  assign n8153 = ( n5688 & n8151 ) | ( n5688 & n8152 ) | ( n8151 & n8152 ) ;
  assign n8154 = n4598 ^ n4280 ^ 1'b0 ;
  assign n8155 = n657 ^ n275 ^ n139 ;
  assign n8156 = ( n8153 & n8154 ) | ( n8153 & ~n8155 ) | ( n8154 & ~n8155 ) ;
  assign n8158 = ( n2539 & ~n2570 ) | ( n2539 & n2826 ) | ( ~n2570 & n2826 ) ;
  assign n8157 = n1980 ^ n510 ^ 1'b0 ;
  assign n8159 = n8158 ^ n8157 ^ n1430 ;
  assign n8160 = n8156 & n8159 ;
  assign n8161 = ( n2445 & n3576 ) | ( n2445 & ~n7806 ) | ( n3576 & ~n7806 ) ;
  assign n8162 = n5634 & ~n8161 ;
  assign n8163 = ~n7698 & n8162 ;
  assign n8167 = n7671 ^ n3217 ^ n1239 ;
  assign n8168 = n8167 ^ n6301 ^ n4884 ;
  assign n8164 = n6535 ^ n6500 ^ n1719 ;
  assign n8165 = ( n5611 & ~n6639 ) | ( n5611 & n8164 ) | ( ~n6639 & n8164 ) ;
  assign n8166 = n8165 ^ n198 ^ 1'b0 ;
  assign n8169 = n8168 ^ n8166 ^ n2832 ;
  assign n8170 = n8169 ^ n140 ^ x60 ;
  assign n8171 = ( n294 & n2122 ) | ( n294 & n2642 ) | ( n2122 & n2642 ) ;
  assign n8172 = n6131 ^ n4160 ^ n2169 ;
  assign n8173 = n3637 & n8172 ;
  assign n8174 = n8173 ^ n1343 ^ 1'b0 ;
  assign n8175 = ( x42 & ~n867 ) | ( x42 & n2307 ) | ( ~n867 & n2307 ) ;
  assign n8176 = ( n680 & n1441 ) | ( n680 & n2002 ) | ( n1441 & n2002 ) ;
  assign n8177 = ~n2575 & n8176 ;
  assign n8178 = n8177 ^ n1451 ^ 1'b0 ;
  assign n8179 = n8175 & n8178 ;
  assign n8180 = ~n8174 & n8179 ;
  assign n8181 = ( n350 & n553 ) | ( n350 & n8100 ) | ( n553 & n8100 ) ;
  assign n8182 = ( n887 & n1902 ) | ( n887 & ~n3380 ) | ( n1902 & ~n3380 ) ;
  assign n8183 = n8182 ^ n4497 ^ n3938 ;
  assign n8189 = ( n5053 & ~n5662 ) | ( n5053 & n6411 ) | ( ~n5662 & n6411 ) ;
  assign n8184 = ( ~n3912 & n3918 ) | ( ~n3912 & n4496 ) | ( n3918 & n4496 ) ;
  assign n8185 = ~n2656 & n3717 ;
  assign n8186 = ( n5413 & ~n5828 ) | ( n5413 & n8185 ) | ( ~n5828 & n8185 ) ;
  assign n8187 = n8186 ^ n2941 ^ n2489 ;
  assign n8188 = ( ~n4734 & n8184 ) | ( ~n4734 & n8187 ) | ( n8184 & n8187 ) ;
  assign n8190 = n8189 ^ n8188 ^ n3051 ;
  assign n8191 = n8190 ^ n7731 ^ n5273 ;
  assign n8192 = ~n1254 & n3074 ;
  assign n8193 = n8192 ^ n2970 ^ n1490 ;
  assign n8194 = n3585 & n6783 ;
  assign n8195 = n1001 & ~n8194 ;
  assign n8196 = ( ~n1788 & n6097 ) | ( ~n1788 & n8195 ) | ( n6097 & n8195 ) ;
  assign n8198 = n191 | n5375 ;
  assign n8199 = n8198 ^ n691 ^ 1'b0 ;
  assign n8197 = n4707 ^ n3451 ^ n1491 ;
  assign n8200 = n8199 ^ n8197 ^ n2055 ;
  assign n8201 = n7302 ^ n3773 ^ x11 ;
  assign n8202 = ( ~n1469 & n7015 ) | ( ~n1469 & n8201 ) | ( n7015 & n8201 ) ;
  assign n8203 = ( ~n3096 & n3539 ) | ( ~n3096 & n8202 ) | ( n3539 & n8202 ) ;
  assign n8208 = ( n816 & n2313 ) | ( n816 & n6530 ) | ( n2313 & n6530 ) ;
  assign n8206 = ~n2702 & n2872 ;
  assign n8207 = ~n3677 & n8206 ;
  assign n8204 = ~n147 & n2516 ;
  assign n8205 = ~n3965 & n8204 ;
  assign n8209 = n8208 ^ n8207 ^ n8205 ;
  assign n8210 = ~n3582 & n6407 ;
  assign n8213 = ( n2989 & n3101 ) | ( n2989 & n5320 ) | ( n3101 & n5320 ) ;
  assign n8211 = ( n2276 & n6293 ) | ( n2276 & n7403 ) | ( n6293 & n7403 ) ;
  assign n8212 = n8211 ^ n1351 ^ x123 ;
  assign n8214 = n8213 ^ n8212 ^ n6773 ;
  assign n8215 = ~n8210 & n8214 ;
  assign n8216 = ~n5241 & n8215 ;
  assign n8217 = ( n219 & n3573 ) | ( n219 & n4277 ) | ( n3573 & n4277 ) ;
  assign n8218 = n8217 ^ n7113 ^ n2479 ;
  assign n8219 = n6681 ^ n6401 ^ n2896 ;
  assign n8220 = n8219 ^ n3973 ^ n1828 ;
  assign n8221 = ~n8218 & n8220 ;
  assign n8222 = n852 | n4295 ;
  assign n8223 = n8222 ^ n396 ^ 1'b0 ;
  assign n8224 = n4344 | n8223 ;
  assign n8225 = n385 & ~n8224 ;
  assign n8226 = ( ~n734 & n7287 ) | ( ~n734 & n8225 ) | ( n7287 & n8225 ) ;
  assign n8227 = ( n188 & ~n1762 ) | ( n188 & n5672 ) | ( ~n1762 & n5672 ) ;
  assign n8228 = n6274 | n8227 ;
  assign n8229 = n1332 & ~n8228 ;
  assign n8230 = n8137 ^ n2762 ^ n964 ;
  assign n8231 = n8230 ^ n7737 ^ n1296 ;
  assign n8238 = ( n1277 & ~n1281 ) | ( n1277 & n1645 ) | ( ~n1281 & n1645 ) ;
  assign n8239 = n8238 ^ n3277 ^ 1'b0 ;
  assign n8237 = ( n850 & n1462 ) | ( n850 & ~n2968 ) | ( n1462 & ~n2968 ) ;
  assign n8232 = n5721 | n5753 ;
  assign n8233 = n8232 ^ n1007 ^ 1'b0 ;
  assign n8234 = ( ~n1150 & n1504 ) | ( ~n1150 & n5419 ) | ( n1504 & n5419 ) ;
  assign n8235 = n3416 ^ n1883 ^ n746 ;
  assign n8236 = ( n8233 & ~n8234 ) | ( n8233 & n8235 ) | ( ~n8234 & n8235 ) ;
  assign n8240 = n8239 ^ n8237 ^ n8236 ;
  assign n8241 = ( n6301 & n8231 ) | ( n6301 & n8240 ) | ( n8231 & n8240 ) ;
  assign n8242 = n7310 ^ n6894 ^ 1'b0 ;
  assign n8243 = ~n2481 & n8242 ;
  assign n8244 = n8243 ^ n4851 ^ 1'b0 ;
  assign n8245 = ( n3012 & ~n4321 ) | ( n3012 & n6265 ) | ( ~n4321 & n6265 ) ;
  assign n8246 = n2095 & n3101 ;
  assign n8247 = n8246 ^ n4178 ^ 1'b0 ;
  assign n8248 = n3981 ^ n1920 ^ 1'b0 ;
  assign n8249 = ~n2313 & n8248 ;
  assign n8250 = n8249 ^ n6934 ^ n3845 ;
  assign n8251 = ( ~n3124 & n8247 ) | ( ~n3124 & n8250 ) | ( n8247 & n8250 ) ;
  assign n8252 = n2755 | n4473 ;
  assign n8253 = n2021 & ~n8252 ;
  assign n8255 = n4386 ^ n2131 ^ n159 ;
  assign n8254 = n2150 & n4802 ;
  assign n8256 = n8255 ^ n8254 ^ n1471 ;
  assign n8257 = ( ~n8251 & n8253 ) | ( ~n8251 & n8256 ) | ( n8253 & n8256 ) ;
  assign n8258 = ( n989 & ~n7424 ) | ( n989 & n7661 ) | ( ~n7424 & n7661 ) ;
  assign n8259 = n5279 ^ n2291 ^ n1420 ;
  assign n8260 = n3424 ^ n2556 ^ n2081 ;
  assign n8261 = n8260 ^ n7526 ^ n2572 ;
  assign n8262 = n8261 ^ n7214 ^ 1'b0 ;
  assign n8263 = ~n8259 & n8262 ;
  assign n8265 = ( n585 & n2174 ) | ( n585 & ~n3905 ) | ( n2174 & ~n3905 ) ;
  assign n8264 = n4872 ^ n2914 ^ 1'b0 ;
  assign n8266 = n8265 ^ n8264 ^ 1'b0 ;
  assign n8267 = n6721 ^ n2923 ^ n707 ;
  assign n8268 = n6992 ^ n2540 ^ n873 ;
  assign n8269 = ( x121 & ~n5540 ) | ( x121 & n6939 ) | ( ~n5540 & n6939 ) ;
  assign n8270 = ( n2537 & n8268 ) | ( n2537 & n8269 ) | ( n8268 & n8269 ) ;
  assign n8271 = n8270 ^ n5192 ^ n1291 ;
  assign n8272 = ( n2906 & n8267 ) | ( n2906 & n8271 ) | ( n8267 & n8271 ) ;
  assign n8273 = n4406 ^ n2581 ^ n512 ;
  assign n8274 = n657 | n8273 ;
  assign n8275 = ( n818 & n1488 ) | ( n818 & n4796 ) | ( n1488 & n4796 ) ;
  assign n8276 = ( n379 & ~n2481 ) | ( n379 & n8275 ) | ( ~n2481 & n8275 ) ;
  assign n8279 = ( n763 & n3325 ) | ( n763 & n3636 ) | ( n3325 & n3636 ) ;
  assign n8277 = n1008 | n4466 ;
  assign n8278 = ~n3663 & n8277 ;
  assign n8280 = n8279 ^ n8278 ^ 1'b0 ;
  assign n8281 = ( n2211 & n2363 ) | ( n2211 & ~n6643 ) | ( n2363 & ~n6643 ) ;
  assign n8282 = n3842 ^ n2235 ^ n1458 ;
  assign n8283 = ( ~n2753 & n2923 ) | ( ~n2753 & n8282 ) | ( n2923 & n8282 ) ;
  assign n8285 = n1113 ^ n1056 ^ x92 ;
  assign n8286 = n760 & ~n4890 ;
  assign n8287 = n2032 & n8286 ;
  assign n8288 = ( n1032 & n8285 ) | ( n1032 & ~n8287 ) | ( n8285 & ~n8287 ) ;
  assign n8284 = n1520 & n5557 ;
  assign n8289 = n8288 ^ n8284 ^ 1'b0 ;
  assign n8290 = n1511 | n7271 ;
  assign n8291 = ( ~n234 & n3948 ) | ( ~n234 & n7891 ) | ( n3948 & n7891 ) ;
  assign n8292 = n4121 ^ n2744 ^ n1145 ;
  assign n8295 = ( ~n397 & n556 ) | ( ~n397 & n3547 ) | ( n556 & n3547 ) ;
  assign n8296 = ( ~n826 & n1925 ) | ( ~n826 & n3507 ) | ( n1925 & n3507 ) ;
  assign n8297 = n8295 | n8296 ;
  assign n8293 = ( n171 & n1154 ) | ( n171 & n1580 ) | ( n1154 & n1580 ) ;
  assign n8294 = ( ~n1638 & n3420 ) | ( ~n1638 & n8293 ) | ( n3420 & n8293 ) ;
  assign n8298 = n8297 ^ n8294 ^ 1'b0 ;
  assign n8299 = n8292 & n8298 ;
  assign n8300 = n855 & ~n2618 ;
  assign n8301 = ( n498 & ~n1287 ) | ( n498 & n8300 ) | ( ~n1287 & n8300 ) ;
  assign n8302 = ( n1733 & ~n6077 ) | ( n1733 & n8301 ) | ( ~n6077 & n8301 ) ;
  assign n8303 = n8302 ^ n5579 ^ n4707 ;
  assign n8304 = n6380 ^ n4995 ^ n3782 ;
  assign n8305 = n7328 ^ n1927 ^ n1463 ;
  assign n8306 = ( n2156 & n4556 ) | ( n2156 & ~n8305 ) | ( n4556 & ~n8305 ) ;
  assign n8307 = ( x53 & n740 ) | ( x53 & ~n859 ) | ( n740 & ~n859 ) ;
  assign n8308 = ( n1820 & n1946 ) | ( n1820 & ~n8307 ) | ( n1946 & ~n8307 ) ;
  assign n8309 = n8308 ^ n4488 ^ n1565 ;
  assign n8310 = ~n7532 & n8309 ;
  assign n8311 = ( n2560 & n4384 ) | ( n2560 & ~n8310 ) | ( n4384 & ~n8310 ) ;
  assign n8312 = n7283 | n8311 ;
  assign n8313 = n2096 ^ n835 ^ n665 ;
  assign n8314 = n5885 ^ n2948 ^ 1'b0 ;
  assign n8315 = ~n8313 & n8314 ;
  assign n8316 = ( ~n1158 & n5244 ) | ( ~n1158 & n6357 ) | ( n5244 & n6357 ) ;
  assign n8317 = n8316 ^ n1979 ^ n662 ;
  assign n8318 = n778 | n5870 ;
  assign n8319 = n8318 ^ n3542 ^ 1'b0 ;
  assign n8323 = n4368 ^ n1727 ^ n1490 ;
  assign n8324 = n5348 | n7613 ;
  assign n8325 = n8323 & ~n8324 ;
  assign n8320 = n951 & ~n6309 ;
  assign n8321 = n8320 ^ n7462 ^ n507 ;
  assign n8322 = ( n2204 & n6354 ) | ( n2204 & ~n8321 ) | ( n6354 & ~n8321 ) ;
  assign n8326 = n8325 ^ n8322 ^ 1'b0 ;
  assign n8327 = ( n8317 & n8319 ) | ( n8317 & n8326 ) | ( n8319 & n8326 ) ;
  assign n8328 = n3101 ^ n2952 ^ n386 ;
  assign n8329 = ~n1674 & n3406 ;
  assign n8330 = ( n7309 & n8328 ) | ( n7309 & ~n8329 ) | ( n8328 & ~n8329 ) ;
  assign n8331 = ( n2893 & n6863 ) | ( n2893 & n8330 ) | ( n6863 & n8330 ) ;
  assign n8332 = n1664 & ~n6262 ;
  assign n8333 = n1318 & n8332 ;
  assign n8334 = n8333 ^ n6939 ^ n4196 ;
  assign n8337 = n5103 ^ n761 ^ 1'b0 ;
  assign n8335 = x97 & ~n3626 ;
  assign n8336 = n2988 & n8335 ;
  assign n8338 = n8337 ^ n8336 ^ n6214 ;
  assign n8339 = n3742 ^ n3435 ^ n195 ;
  assign n8340 = n8338 | n8339 ;
  assign n8341 = n8340 ^ n5908 ^ 1'b0 ;
  assign n8342 = ( n8178 & n8334 ) | ( n8178 & n8341 ) | ( n8334 & n8341 ) ;
  assign n8343 = n7802 ^ n2568 ^ n2358 ;
  assign n8344 = n2855 ^ n1960 ^ n562 ;
  assign n8345 = ( ~n4423 & n7297 ) | ( ~n4423 & n8344 ) | ( n7297 & n8344 ) ;
  assign n8346 = ( n4207 & n8343 ) | ( n4207 & n8345 ) | ( n8343 & n8345 ) ;
  assign n8347 = ( n7424 & ~n8342 ) | ( n7424 & n8346 ) | ( ~n8342 & n8346 ) ;
  assign n8349 = n2569 ^ n2186 ^ n2016 ;
  assign n8348 = n3375 ^ n809 ^ 1'b0 ;
  assign n8350 = n8349 ^ n8348 ^ n2977 ;
  assign n8351 = n6676 ^ n5381 ^ n1903 ;
  assign n8352 = ( n774 & n8348 ) | ( n774 & ~n8351 ) | ( n8348 & ~n8351 ) ;
  assign n8353 = ( ~n7294 & n8350 ) | ( ~n7294 & n8352 ) | ( n8350 & n8352 ) ;
  assign n8354 = ( n1317 & n2232 ) | ( n1317 & n5866 ) | ( n2232 & n5866 ) ;
  assign n8355 = ( n1541 & n7065 ) | ( n1541 & n8354 ) | ( n7065 & n8354 ) ;
  assign n8360 = n577 & n3189 ;
  assign n8356 = n6880 ^ n1064 ^ 1'b0 ;
  assign n8357 = ~n3733 & n8356 ;
  assign n8358 = n1334 & n5221 ;
  assign n8359 = n8357 & n8358 ;
  assign n8361 = n8360 ^ n8359 ^ 1'b0 ;
  assign n8362 = n6498 ^ n1777 ^ n1520 ;
  assign n8363 = n8362 ^ n3988 ^ 1'b0 ;
  assign n8364 = n8361 & n8363 ;
  assign n8365 = ( ~n2738 & n8355 ) | ( ~n2738 & n8364 ) | ( n8355 & n8364 ) ;
  assign n8366 = n8365 ^ n6730 ^ n171 ;
  assign n8367 = ( n572 & ~n2468 ) | ( n572 & n3222 ) | ( ~n2468 & n3222 ) ;
  assign n8368 = ( n4037 & n4559 ) | ( n4037 & n8367 ) | ( n4559 & n8367 ) ;
  assign n8369 = n8368 ^ n8089 ^ n5707 ;
  assign n8375 = n3717 ^ n3365 ^ 1'b0 ;
  assign n8376 = n8375 ^ n2047 ^ n1932 ;
  assign n8377 = ( n4357 & ~n6147 ) | ( n4357 & n8376 ) | ( ~n6147 & n8376 ) ;
  assign n8371 = x86 & ~n759 ;
  assign n8372 = ~n1294 & n8371 ;
  assign n8370 = ( n1675 & ~n2952 ) | ( n1675 & n7671 ) | ( ~n2952 & n7671 ) ;
  assign n8373 = n8372 ^ n8370 ^ n3201 ;
  assign n8374 = ( ~n3696 & n7556 ) | ( ~n3696 & n8373 ) | ( n7556 & n8373 ) ;
  assign n8378 = n8377 ^ n8374 ^ n1716 ;
  assign n8379 = n430 | n6713 ;
  assign n8380 = n487 & ~n8379 ;
  assign n8381 = n4196 ^ n373 ^ 1'b0 ;
  assign n8382 = n8012 | n8381 ;
  assign n8384 = ( n1167 & ~n1411 ) | ( n1167 & n2348 ) | ( ~n1411 & n2348 ) ;
  assign n8383 = ( x66 & n4783 ) | ( x66 & ~n8217 ) | ( n4783 & ~n8217 ) ;
  assign n8385 = n8384 ^ n8383 ^ n5140 ;
  assign n8386 = ( n8380 & ~n8382 ) | ( n8380 & n8385 ) | ( ~n8382 & n8385 ) ;
  assign n8387 = n8386 ^ n5019 ^ n3688 ;
  assign n8388 = ( ~n425 & n2119 ) | ( ~n425 & n3357 ) | ( n2119 & n3357 ) ;
  assign n8389 = n8388 ^ n773 ^ n222 ;
  assign n8390 = n8389 ^ n5684 ^ n5407 ;
  assign n8391 = n7963 & n8128 ;
  assign n8392 = ~n1152 & n8391 ;
  assign n8393 = n8392 ^ n3453 ^ n2943 ;
  assign n8394 = n1868 ^ n1648 ^ 1'b0 ;
  assign n8395 = x71 & ~n8394 ;
  assign n8396 = n8393 & ~n8395 ;
  assign n8404 = n3281 | n6268 ;
  assign n8405 = n4029 ^ n2464 ^ 1'b0 ;
  assign n8406 = n8404 & ~n8405 ;
  assign n8407 = n8406 ^ n5977 ^ n2338 ;
  assign n8401 = n2971 & n8307 ;
  assign n8402 = n8401 ^ n2042 ^ 1'b0 ;
  assign n8397 = n1668 & ~n3982 ;
  assign n8398 = n8397 ^ n1901 ^ 1'b0 ;
  assign n8399 = n8398 ^ n3193 ^ n1617 ;
  assign n8400 = n8399 ^ n4515 ^ n1565 ;
  assign n8403 = n8402 ^ n8400 ^ n175 ;
  assign n8408 = n8407 ^ n8403 ^ 1'b0 ;
  assign n8411 = ( n4071 & ~n4222 ) | ( n4071 & n5599 ) | ( ~n4222 & n5599 ) ;
  assign n8412 = n8411 ^ n5993 ^ n2186 ;
  assign n8409 = n402 & ~n3134 ;
  assign n8410 = n8409 ^ n5975 ^ 1'b0 ;
  assign n8413 = n8412 ^ n8410 ^ n4421 ;
  assign n8414 = n1906 ^ n1842 ^ n648 ;
  assign n8415 = n2475 & n6091 ;
  assign n8416 = n8415 ^ n1484 ^ 1'b0 ;
  assign n8417 = ( n1994 & n8414 ) | ( n1994 & ~n8416 ) | ( n8414 & ~n8416 ) ;
  assign n8418 = n421 & ~n8417 ;
  assign n8419 = n7229 | n8418 ;
  assign n8420 = ( n447 & n1038 ) | ( n447 & ~n2376 ) | ( n1038 & ~n2376 ) ;
  assign n8421 = ( n4172 & ~n8419 ) | ( n4172 & n8420 ) | ( ~n8419 & n8420 ) ;
  assign n8422 = ( n1612 & n1701 ) | ( n1612 & n1777 ) | ( n1701 & n1777 ) ;
  assign n8423 = ( n164 & ~n976 ) | ( n164 & n4101 ) | ( ~n976 & n4101 ) ;
  assign n8424 = ( n234 & n996 ) | ( n234 & n8423 ) | ( n996 & n8423 ) ;
  assign n8425 = n8422 | n8424 ;
  assign n8426 = n8270 ^ n6996 ^ x6 ;
  assign n8427 = n424 | n610 ;
  assign n8428 = n8427 ^ n277 ^ 1'b0 ;
  assign n8429 = ( n1919 & n2384 ) | ( n1919 & ~n8428 ) | ( n2384 & ~n8428 ) ;
  assign n8430 = n8429 ^ n3363 ^ n2444 ;
  assign n8431 = ( ~n3081 & n4571 ) | ( ~n3081 & n8430 ) | ( n4571 & n8430 ) ;
  assign n8432 = n7003 | n8431 ;
  assign n8433 = ( ~n529 & n4309 ) | ( ~n529 & n5901 ) | ( n4309 & n5901 ) ;
  assign n8434 = n8433 ^ n1464 ^ n461 ;
  assign n8435 = ( n1649 & n4472 ) | ( n1649 & ~n5607 ) | ( n4472 & ~n5607 ) ;
  assign n8436 = ( n740 & n8434 ) | ( n740 & ~n8435 ) | ( n8434 & ~n8435 ) ;
  assign n8437 = n3157 | n3515 ;
  assign n8438 = n8437 ^ x89 ^ 1'b0 ;
  assign n8439 = ( n7062 & n7919 ) | ( n7062 & n8438 ) | ( n7919 & n8438 ) ;
  assign n8440 = n8439 ^ n1627 ^ n675 ;
  assign n8441 = n8440 ^ n6891 ^ n338 ;
  assign n8442 = ( n765 & n3451 ) | ( n765 & ~n8441 ) | ( n3451 & ~n8441 ) ;
  assign n8443 = ( x37 & n2783 ) | ( x37 & ~n7710 ) | ( n2783 & ~n7710 ) ;
  assign n8444 = ( n1415 & n2869 ) | ( n1415 & n3307 ) | ( n2869 & n3307 ) ;
  assign n8445 = n8444 ^ n181 ^ 1'b0 ;
  assign n8448 = n4665 ^ n4495 ^ 1'b0 ;
  assign n8449 = n4022 & ~n8448 ;
  assign n8446 = n7837 ^ n2618 ^ n204 ;
  assign n8447 = n8446 ^ n1016 ^ 1'b0 ;
  assign n8450 = n8449 ^ n8447 ^ n7586 ;
  assign n8451 = n3911 ^ n2868 ^ n1398 ;
  assign n8452 = n3614 ^ n1397 ^ n1042 ;
  assign n8453 = n8452 ^ n3398 ^ n1818 ;
  assign n8454 = ~n3463 & n8453 ;
  assign n8455 = n3001 & n8454 ;
  assign n8456 = ( n898 & ~n8451 ) | ( n898 & n8455 ) | ( ~n8451 & n8455 ) ;
  assign n8457 = n1058 ^ n1020 ^ x110 ;
  assign n8458 = ( n817 & ~n3191 ) | ( n817 & n8457 ) | ( ~n3191 & n8457 ) ;
  assign n8459 = n7638 ^ n5582 ^ 1'b0 ;
  assign n8469 = ( n1016 & n4793 ) | ( n1016 & n8265 ) | ( n4793 & n8265 ) ;
  assign n8470 = n8469 ^ n3567 ^ n1848 ;
  assign n8471 = ( n1035 & ~n4828 ) | ( n1035 & n8470 ) | ( ~n4828 & n8470 ) ;
  assign n8468 = n1791 ^ n1356 ^ n1231 ;
  assign n8460 = ( n1058 & n2716 ) | ( n1058 & n2838 ) | ( n2716 & n2838 ) ;
  assign n8461 = n8338 ^ n3222 ^ 1'b0 ;
  assign n8462 = n4891 ^ n3070 ^ 1'b0 ;
  assign n8463 = n5919 & n8462 ;
  assign n8464 = n8461 & n8463 ;
  assign n8465 = n8460 & n8464 ;
  assign n8466 = n3182 & ~n8465 ;
  assign n8467 = n8466 ^ n6322 ^ 1'b0 ;
  assign n8472 = n8471 ^ n8468 ^ n8467 ;
  assign n8473 = n6883 ^ n6059 ^ n2727 ;
  assign n8474 = ( n2153 & ~n2224 ) | ( n2153 & n4194 ) | ( ~n2224 & n4194 ) ;
  assign n8475 = n8474 ^ n5415 ^ n1585 ;
  assign n8476 = n1028 & n8475 ;
  assign n8477 = n4018 ^ n3073 ^ 1'b0 ;
  assign n8482 = ~n1573 & n3402 ;
  assign n8483 = n2533 & ~n8482 ;
  assign n8484 = n8483 ^ n1735 ^ 1'b0 ;
  assign n8485 = n8484 ^ n6670 ^ n5536 ;
  assign n8478 = n7162 ^ n3582 ^ n1126 ;
  assign n8479 = n4731 ^ n255 ^ 1'b0 ;
  assign n8480 = ( ~n5323 & n5518 ) | ( ~n5323 & n8479 ) | ( n5518 & n8479 ) ;
  assign n8481 = ( n2656 & n8478 ) | ( n2656 & n8480 ) | ( n8478 & n8480 ) ;
  assign n8486 = n8485 ^ n8481 ^ 1'b0 ;
  assign n8487 = ( n2215 & n3106 ) | ( n2215 & n4202 ) | ( n3106 & n4202 ) ;
  assign n8488 = n1498 & ~n8451 ;
  assign n8489 = n8488 ^ n387 ^ 1'b0 ;
  assign n8490 = n8489 ^ n3642 ^ n409 ;
  assign n8491 = ( n384 & n2581 ) | ( n384 & ~n8295 ) | ( n2581 & ~n8295 ) ;
  assign n8492 = n8491 ^ n1456 ^ 1'b0 ;
  assign n8493 = ~n8032 & n8492 ;
  assign n8494 = ( n6538 & ~n7001 ) | ( n6538 & n7655 ) | ( ~n7001 & n7655 ) ;
  assign n8496 = ( n1437 & n2330 ) | ( n1437 & n4185 ) | ( n2330 & n4185 ) ;
  assign n8495 = n2502 & n2608 ;
  assign n8497 = n8496 ^ n8495 ^ n6703 ;
  assign n8498 = n8497 ^ n3702 ^ 1'b0 ;
  assign n8499 = n5068 & n6548 ;
  assign n8500 = n3666 & n8499 ;
  assign n8501 = n4252 & n8500 ;
  assign n8502 = ( ~n978 & n1166 ) | ( ~n978 & n5526 ) | ( n1166 & n5526 ) ;
  assign n8503 = n5293 ^ n3631 ^ n1652 ;
  assign n8504 = ( n751 & n7821 ) | ( n751 & n8503 ) | ( n7821 & n8503 ) ;
  assign n8505 = ( n1876 & n8502 ) | ( n1876 & ~n8504 ) | ( n8502 & ~n8504 ) ;
  assign n8513 = ( n2165 & n2302 ) | ( n2165 & ~n7487 ) | ( n2302 & ~n7487 ) ;
  assign n8514 = n3498 | n8513 ;
  assign n8508 = n8000 ^ n3880 ^ n476 ;
  assign n8506 = n1435 | n4015 ;
  assign n8507 = n8506 ^ n2202 ^ 1'b0 ;
  assign n8509 = n8508 ^ n8507 ^ 1'b0 ;
  assign n8510 = ~n7555 & n8509 ;
  assign n8511 = n6313 ^ n5893 ^ n3120 ;
  assign n8512 = ( n5799 & n8510 ) | ( n5799 & ~n8511 ) | ( n8510 & ~n8511 ) ;
  assign n8515 = n8514 ^ n8512 ^ n1143 ;
  assign n8516 = ( ~n1073 & n1642 ) | ( ~n1073 & n7950 ) | ( n1642 & n7950 ) ;
  assign n8517 = n4266 ^ n1156 ^ n1129 ;
  assign n8518 = n8517 ^ n7013 ^ n4793 ;
  assign n8519 = ( ~n4271 & n8516 ) | ( ~n4271 & n8518 ) | ( n8516 & n8518 ) ;
  assign n8520 = ( ~n1402 & n2989 ) | ( ~n1402 & n8519 ) | ( n2989 & n8519 ) ;
  assign n8521 = n6697 ^ n5178 ^ n2480 ;
  assign n8527 = ( ~n503 & n1406 ) | ( ~n503 & n2424 ) | ( n1406 & n2424 ) ;
  assign n8528 = ~n6422 & n8527 ;
  assign n8522 = n7781 ^ n1324 ^ n738 ;
  assign n8523 = ~n1507 & n8522 ;
  assign n8524 = n8523 ^ n4267 ^ 1'b0 ;
  assign n8525 = n8524 ^ n8104 ^ n1350 ;
  assign n8526 = n8525 ^ n739 ^ x6 ;
  assign n8529 = n8528 ^ n8526 ^ n133 ;
  assign n8530 = n2091 & n3325 ;
  assign n8531 = ~n3435 & n8530 ;
  assign n8532 = n8531 ^ n4648 ^ n1052 ;
  assign n8533 = n3532 ^ n784 ^ n655 ;
  assign n8534 = n8533 ^ n2982 ^ n1513 ;
  assign n8535 = n8532 & n8534 ;
  assign n8536 = n8535 ^ n674 ^ 1'b0 ;
  assign n8544 = n3432 ^ n2292 ^ n251 ;
  assign n8545 = n4413 ^ n576 ^ n305 ;
  assign n8546 = n8544 & n8545 ;
  assign n8547 = n8546 ^ n1068 ^ 1'b0 ;
  assign n8537 = n5366 ^ n4905 ^ n2826 ;
  assign n8538 = n8537 ^ n4534 ^ n1069 ;
  assign n8539 = ( ~n2432 & n4298 ) | ( ~n2432 & n8538 ) | ( n4298 & n8538 ) ;
  assign n8540 = n8539 ^ n5484 ^ 1'b0 ;
  assign n8541 = n2163 & n4060 ;
  assign n8542 = n4177 & ~n8541 ;
  assign n8543 = n8540 & n8542 ;
  assign n8548 = n8547 ^ n8543 ^ n4283 ;
  assign n8549 = n4700 ^ n3064 ^ 1'b0 ;
  assign n8550 = ( n1698 & ~n3876 ) | ( n1698 & n5452 ) | ( ~n3876 & n5452 ) ;
  assign n8551 = ~n2557 & n3822 ;
  assign n8552 = n8550 & n8551 ;
  assign n8557 = n1580 ^ n1525 ^ 1'b0 ;
  assign n8558 = ~n916 & n8557 ;
  assign n8553 = n5903 ^ n1365 ^ 1'b0 ;
  assign n8554 = n3237 & ~n8553 ;
  assign n8555 = n8554 ^ n4463 ^ 1'b0 ;
  assign n8556 = n2837 | n8555 ;
  assign n8559 = n8558 ^ n8556 ^ n8132 ;
  assign n8560 = ( n935 & ~n1059 ) | ( n935 & n8559 ) | ( ~n1059 & n8559 ) ;
  assign n8561 = n4012 & n8560 ;
  assign n8562 = ~n2201 & n3822 ;
  assign n8563 = n800 ^ n675 ^ 1'b0 ;
  assign n8564 = ~n8562 & n8563 ;
  assign n8565 = n6741 & ~n7799 ;
  assign n8566 = ~n2157 & n8565 ;
  assign n8567 = n578 & ~n3081 ;
  assign n8568 = n8567 ^ n888 ^ 1'b0 ;
  assign n8569 = n2875 ^ n2108 ^ x119 ;
  assign n8570 = ( n1328 & ~n5200 ) | ( n1328 & n8569 ) | ( ~n5200 & n8569 ) ;
  assign n8571 = n8570 ^ n4244 ^ 1'b0 ;
  assign n8572 = n8568 | n8571 ;
  assign n8573 = n3769 & ~n5583 ;
  assign n8574 = n6096 & ~n7812 ;
  assign n8575 = n8574 ^ n5469 ^ 1'b0 ;
  assign n8576 = n4995 ^ n4826 ^ n400 ;
  assign n8577 = ( n2488 & n5373 ) | ( n2488 & n6767 ) | ( n5373 & n6767 ) ;
  assign n8578 = n8577 ^ n7469 ^ n3818 ;
  assign n8579 = ( n1738 & n4888 ) | ( n1738 & n8578 ) | ( n4888 & n8578 ) ;
  assign n8580 = n4013 | n7312 ;
  assign n8581 = n3580 & ~n8580 ;
  assign n8582 = n3789 ^ n3445 ^ 1'b0 ;
  assign n8583 = ( n1870 & ~n2225 ) | ( n1870 & n8582 ) | ( ~n2225 & n8582 ) ;
  assign n8584 = n1195 & ~n5073 ;
  assign n8585 = n8584 ^ n8503 ^ 1'b0 ;
  assign n8586 = n7564 ^ n4054 ^ 1'b0 ;
  assign n8587 = n8440 ^ n5485 ^ 1'b0 ;
  assign n8588 = ( n676 & ~n2819 ) | ( n676 & n3967 ) | ( ~n2819 & n3967 ) ;
  assign n8589 = ( ~n3986 & n4828 ) | ( ~n3986 & n6501 ) | ( n4828 & n6501 ) ;
  assign n8590 = n3551 ^ n1220 ^ 1'b0 ;
  assign n8591 = n3177 | n8590 ;
  assign n8592 = ( ~n1126 & n4969 ) | ( ~n1126 & n8591 ) | ( n4969 & n8591 ) ;
  assign n8593 = ( n4419 & n5175 ) | ( n4419 & n8592 ) | ( n5175 & n8592 ) ;
  assign n8594 = ( n2581 & n8589 ) | ( n2581 & ~n8593 ) | ( n8589 & ~n8593 ) ;
  assign n8595 = ( ~n7718 & n8588 ) | ( ~n7718 & n8594 ) | ( n8588 & n8594 ) ;
  assign n8596 = n520 & n3525 ;
  assign n8597 = n8596 ^ n2240 ^ 1'b0 ;
  assign n8598 = n8597 ^ n856 ^ 1'b0 ;
  assign n8599 = n4643 & ~n8598 ;
  assign n8600 = n6220 & n8599 ;
  assign n8601 = n8600 ^ n3096 ^ 1'b0 ;
  assign n8602 = n7464 ^ n5370 ^ n2869 ;
  assign n8603 = n6149 ^ n5997 ^ n923 ;
  assign n8604 = n5131 ^ n441 ^ n317 ;
  assign n8605 = ( n357 & ~n2642 ) | ( n357 & n8604 ) | ( ~n2642 & n8604 ) ;
  assign n8606 = n8605 ^ n966 ^ 1'b0 ;
  assign n8607 = ( n7436 & n8603 ) | ( n7436 & ~n8606 ) | ( n8603 & ~n8606 ) ;
  assign n8608 = n8607 ^ n5993 ^ n381 ;
  assign n8613 = n7804 ^ n3117 ^ n516 ;
  assign n8609 = n4122 ^ n3248 ^ n1627 ;
  assign n8610 = n8609 ^ n6935 ^ n2185 ;
  assign n8611 = ( n5386 & n5988 ) | ( n5386 & n8610 ) | ( n5988 & n8610 ) ;
  assign n8612 = n3970 & ~n8611 ;
  assign n8614 = n8613 ^ n8612 ^ 1'b0 ;
  assign n8615 = ( n3221 & ~n3294 ) | ( n3221 & n3936 ) | ( ~n3294 & n3936 ) ;
  assign n8616 = n1814 & ~n8615 ;
  assign n8617 = ~n8149 & n8616 ;
  assign n8620 = n7162 ^ n3484 ^ n2055 ;
  assign n8621 = n8620 ^ n4037 ^ n2060 ;
  assign n8619 = ( n507 & n1388 ) | ( n507 & n4306 ) | ( n1388 & n4306 ) ;
  assign n8618 = n8275 ^ n635 ^ x72 ;
  assign n8622 = n8621 ^ n8619 ^ n8618 ;
  assign n8624 = ( n1388 & n3091 ) | ( n1388 & ~n6571 ) | ( n3091 & ~n6571 ) ;
  assign n8623 = ( ~n1016 & n1436 ) | ( ~n1016 & n5311 ) | ( n1436 & n5311 ) ;
  assign n8625 = n8624 ^ n8623 ^ 1'b0 ;
  assign n8626 = n4398 ^ n2038 ^ n1730 ;
  assign n8627 = n8626 ^ n8308 ^ n7324 ;
  assign n8628 = ( n1052 & n1799 ) | ( n1052 & n2812 ) | ( n1799 & n2812 ) ;
  assign n8629 = n664 | n1245 ;
  assign n8630 = ( n911 & ~n8628 ) | ( n911 & n8629 ) | ( ~n8628 & n8629 ) ;
  assign n8631 = n8627 & ~n8630 ;
  assign n8632 = n6009 & n7860 ;
  assign n8633 = n8632 ^ n2744 ^ 1'b0 ;
  assign n8634 = ( n3209 & n3682 ) | ( n3209 & ~n8251 ) | ( n3682 & ~n8251 ) ;
  assign n8635 = n8634 ^ n3193 ^ 1'b0 ;
  assign n8636 = n2262 & n8635 ;
  assign n8637 = n458 | n751 ;
  assign n8638 = n6817 ^ n2340 ^ n1568 ;
  assign n8639 = n6639 ^ n2594 ^ n564 ;
  assign n8640 = ( n6568 & n8638 ) | ( n6568 & ~n8639 ) | ( n8638 & ~n8639 ) ;
  assign n8641 = ( n506 & ~n8637 ) | ( n506 & n8640 ) | ( ~n8637 & n8640 ) ;
  assign n8642 = n7930 & ~n8641 ;
  assign n8643 = n3905 ^ n2782 ^ n2181 ;
  assign n8644 = n7747 & ~n7994 ;
  assign n8645 = ( n8556 & n8643 ) | ( n8556 & n8644 ) | ( n8643 & n8644 ) ;
  assign n8646 = n3363 ^ n2793 ^ 1'b0 ;
  assign n8650 = ~n327 & n1609 ;
  assign n8651 = n8650 ^ n1196 ^ 1'b0 ;
  assign n8649 = ( ~n3987 & n5473 ) | ( ~n3987 & n7128 ) | ( n5473 & n7128 ) ;
  assign n8652 = n8651 ^ n8649 ^ n5151 ;
  assign n8653 = n8652 ^ n5262 ^ n3838 ;
  assign n8647 = n4376 & n5020 ;
  assign n8648 = n252 | n8647 ;
  assign n8654 = n8653 ^ n8648 ^ n6198 ;
  assign n8655 = ( ~n1894 & n8646 ) | ( ~n1894 & n8654 ) | ( n8646 & n8654 ) ;
  assign n8656 = n7474 ^ n6047 ^ 1'b0 ;
  assign n8657 = n6119 ^ n3923 ^ 1'b0 ;
  assign n8658 = n2358 & n8657 ;
  assign n8659 = ~n4859 & n8658 ;
  assign n8660 = ~n4484 & n8659 ;
  assign n8661 = n8092 ^ n6724 ^ n1942 ;
  assign n8665 = ( ~n605 & n4740 ) | ( ~n605 & n6194 ) | ( n4740 & n6194 ) ;
  assign n8666 = ( n2821 & ~n7460 ) | ( n2821 & n8665 ) | ( ~n7460 & n8665 ) ;
  assign n8667 = n8666 ^ n2165 ^ 1'b0 ;
  assign n8668 = n3179 & n8667 ;
  assign n8662 = n4310 ^ n3584 ^ n2393 ;
  assign n8663 = n4645 ^ n3633 ^ 1'b0 ;
  assign n8664 = ~n8662 & n8663 ;
  assign n8669 = n8668 ^ n8664 ^ 1'b0 ;
  assign n8670 = n6976 ^ n6855 ^ n1113 ;
  assign n8671 = ( n355 & ~n8669 ) | ( n355 & n8670 ) | ( ~n8669 & n8670 ) ;
  assign n8672 = ( n314 & ~n2289 ) | ( n314 & n5526 ) | ( ~n2289 & n5526 ) ;
  assign n8673 = n1385 & n3897 ;
  assign n8678 = ( n209 & n1510 ) | ( n209 & ~n7788 ) | ( n1510 & ~n7788 ) ;
  assign n8674 = ( n1110 & n1690 ) | ( n1110 & n4793 ) | ( n1690 & n4793 ) ;
  assign n8675 = n8674 ^ n4303 ^ 1'b0 ;
  assign n8676 = n2395 & n8675 ;
  assign n8677 = n8676 ^ n4267 ^ n3970 ;
  assign n8679 = n8678 ^ n8677 ^ n4878 ;
  assign n8680 = ( n6495 & n8673 ) | ( n6495 & n8679 ) | ( n8673 & n8679 ) ;
  assign n8681 = ( n6282 & n8672 ) | ( n6282 & ~n8680 ) | ( n8672 & ~n8680 ) ;
  assign n8684 = n2426 ^ n1280 ^ x123 ;
  assign n8682 = n3337 ^ n327 ^ x3 ;
  assign n8683 = ( n3712 & n7918 ) | ( n3712 & n8682 ) | ( n7918 & n8682 ) ;
  assign n8685 = n8684 ^ n8683 ^ n628 ;
  assign n8686 = n1942 | n8685 ;
  assign n8687 = n2653 ^ n776 ^ n693 ;
  assign n8688 = ( n2563 & n6228 ) | ( n2563 & ~n8687 ) | ( n6228 & ~n8687 ) ;
  assign n8689 = n8688 ^ n7713 ^ n5974 ;
  assign n8691 = n3920 ^ n1614 ^ n1284 ;
  assign n8692 = n8691 ^ n1675 ^ n596 ;
  assign n8690 = ( ~n2365 & n4410 ) | ( ~n2365 & n4721 ) | ( n4410 & n4721 ) ;
  assign n8693 = n8692 ^ n8690 ^ n698 ;
  assign n8694 = n2562 ^ n1591 ^ n1392 ;
  assign n8695 = ( n528 & n1709 ) | ( n528 & n8694 ) | ( n1709 & n8694 ) ;
  assign n8696 = n2348 ^ n1327 ^ 1'b0 ;
  assign n8697 = n8696 ^ n1609 ^ 1'b0 ;
  assign n8698 = n6396 & ~n8697 ;
  assign n8701 = ( n499 & ~n1834 ) | ( n499 & n2822 ) | ( ~n1834 & n2822 ) ;
  assign n8702 = n1580 & ~n8701 ;
  assign n8703 = ~n2540 & n8702 ;
  assign n8699 = ( ~n1798 & n3597 ) | ( ~n1798 & n7299 ) | ( n3597 & n7299 ) ;
  assign n8700 = n1310 & n8699 ;
  assign n8704 = n8703 ^ n8700 ^ 1'b0 ;
  assign n8705 = ( n818 & n8698 ) | ( n818 & ~n8704 ) | ( n8698 & ~n8704 ) ;
  assign n8706 = ( n1012 & ~n8695 ) | ( n1012 & n8705 ) | ( ~n8695 & n8705 ) ;
  assign n8707 = ( n8689 & n8693 ) | ( n8689 & ~n8706 ) | ( n8693 & ~n8706 ) ;
  assign n8713 = n6454 ^ n3967 ^ n1037 ;
  assign n8708 = ( n4093 & n5131 ) | ( n4093 & ~n7378 ) | ( n5131 & ~n7378 ) ;
  assign n8710 = n3536 ^ n1315 ^ n995 ;
  assign n8709 = ( n944 & ~n1076 ) | ( n944 & n7333 ) | ( ~n1076 & n7333 ) ;
  assign n8711 = n8710 ^ n8709 ^ n841 ;
  assign n8712 = ~n8708 & n8711 ;
  assign n8714 = n8713 ^ n8712 ^ 1'b0 ;
  assign n8716 = n1991 ^ n1052 ^ n414 ;
  assign n8717 = ~n5067 & n8716 ;
  assign n8718 = ~n8109 & n8717 ;
  assign n8715 = n3295 & n5229 ;
  assign n8719 = n8718 ^ n8715 ^ n5407 ;
  assign n8722 = n1451 | n2107 ;
  assign n8723 = n1926 | n8722 ;
  assign n8724 = n8723 ^ n4044 ^ 1'b0 ;
  assign n8725 = ( n4168 & ~n4508 ) | ( n4168 & n8724 ) | ( ~n4508 & n8724 ) ;
  assign n8726 = n8725 ^ n7184 ^ n1625 ;
  assign n8720 = ~n136 & n8470 ;
  assign n8721 = ~n3532 & n8720 ;
  assign n8727 = n8726 ^ n8721 ^ n2846 ;
  assign n8729 = ( x3 & n4267 ) | ( x3 & n8428 ) | ( n4267 & n8428 ) ;
  assign n8728 = ~n1107 & n7335 ;
  assign n8730 = n8729 ^ n8728 ^ n4786 ;
  assign n8731 = n8730 ^ n2702 ^ n1246 ;
  assign n8732 = n8731 ^ n6460 ^ n2218 ;
  assign n8733 = n8732 ^ n1089 ^ 1'b0 ;
  assign n8734 = n662 & ~n8733 ;
  assign n8735 = n8734 ^ n6626 ^ n6364 ;
  assign n8736 = n6291 ^ n2119 ^ 1'b0 ;
  assign n8737 = n3724 | n8736 ;
  assign n8738 = ( x71 & n4995 ) | ( x71 & n8737 ) | ( n4995 & n8737 ) ;
  assign n8739 = n8738 ^ n7780 ^ n6763 ;
  assign n8740 = n1718 ^ n771 ^ x46 ;
  assign n8741 = n3498 & n5342 ;
  assign n8742 = n7081 ^ n4598 ^ n1113 ;
  assign n8743 = ( ~n5682 & n8741 ) | ( ~n5682 & n8742 ) | ( n8741 & n8742 ) ;
  assign n8744 = ( n3971 & n8740 ) | ( n3971 & n8743 ) | ( n8740 & n8743 ) ;
  assign n8745 = ~n3222 & n7172 ;
  assign n8746 = n278 ^ x115 ^ 1'b0 ;
  assign n8747 = n8745 & n8746 ;
  assign n8748 = n4037 ^ n1371 ^ 1'b0 ;
  assign n8749 = ( ~n3352 & n5390 ) | ( ~n3352 & n5721 ) | ( n5390 & n5721 ) ;
  assign n8751 = n5997 ^ n5504 ^ n3797 ;
  assign n8750 = n5674 ^ n5431 ^ 1'b0 ;
  assign n8752 = n8751 ^ n8750 ^ n5023 ;
  assign n8753 = ( n4154 & n4714 ) | ( n4154 & ~n8752 ) | ( n4714 & ~n8752 ) ;
  assign n8754 = n3573 ^ n2239 ^ 1'b0 ;
  assign n8755 = ( n1093 & n4030 ) | ( n1093 & n5458 ) | ( n4030 & n5458 ) ;
  assign n8756 = ( ~n4899 & n5915 ) | ( ~n4899 & n7059 ) | ( n5915 & n7059 ) ;
  assign n8757 = n7296 & n7830 ;
  assign n8758 = ~n8756 & n8757 ;
  assign n8759 = ~n8755 & n8758 ;
  assign n8760 = ( ~n8276 & n8476 ) | ( ~n8276 & n8759 ) | ( n8476 & n8759 ) ;
  assign n8761 = n1597 | n3481 ;
  assign n8762 = n1982 | n8761 ;
  assign n8763 = n8762 ^ n5269 ^ 1'b0 ;
  assign n8764 = n2346 ^ n475 ^ 1'b0 ;
  assign n8765 = n8764 ^ n6540 ^ 1'b0 ;
  assign n8766 = n8763 & n8765 ;
  assign n8767 = n8766 ^ n6945 ^ n6114 ;
  assign n8768 = n7646 ^ n1732 ^ n1331 ;
  assign n8769 = ( n642 & n1924 ) | ( n642 & ~n2081 ) | ( n1924 & ~n2081 ) ;
  assign n8770 = n1470 | n7718 ;
  assign n8771 = n8769 | n8770 ;
  assign n8774 = ( n2821 & n5106 ) | ( n2821 & n6479 ) | ( n5106 & n6479 ) ;
  assign n8772 = n1440 | n2900 ;
  assign n8773 = n8772 ^ n5915 ^ 1'b0 ;
  assign n8775 = n8774 ^ n8773 ^ n4890 ;
  assign n8776 = n4513 ^ n3357 ^ 1'b0 ;
  assign n8777 = n5436 | n8776 ;
  assign n8778 = n8777 ^ n4127 ^ 1'b0 ;
  assign n8779 = n8775 | n8778 ;
  assign n8780 = n2073 & ~n8779 ;
  assign n8781 = n893 & n8780 ;
  assign n8782 = n8781 ^ n2721 ^ n2471 ;
  assign n8783 = n8782 ^ n7924 ^ 1'b0 ;
  assign n8784 = ( ~n2793 & n3618 ) | ( ~n2793 & n4730 ) | ( n3618 & n4730 ) ;
  assign n8785 = n3236 ^ n1797 ^ n923 ;
  assign n8786 = n8785 ^ n6670 ^ n6500 ;
  assign n8787 = x65 & n796 ;
  assign n8788 = ( ~n3759 & n5042 ) | ( ~n3759 & n8787 ) | ( n5042 & n8787 ) ;
  assign n8789 = n8788 ^ n901 ^ n680 ;
  assign n8790 = ( n8784 & n8786 ) | ( n8784 & n8789 ) | ( n8786 & n8789 ) ;
  assign n8792 = n8604 ^ n7164 ^ n4336 ;
  assign n8793 = n8792 ^ n3277 ^ 1'b0 ;
  assign n8791 = ( ~n2766 & n3444 ) | ( ~n2766 & n7798 ) | ( n3444 & n7798 ) ;
  assign n8794 = n8793 ^ n8791 ^ 1'b0 ;
  assign n8795 = ( n2269 & ~n5051 ) | ( n2269 & n5074 ) | ( ~n5051 & n5074 ) ;
  assign n8796 = ~n1884 & n3040 ;
  assign n8797 = ~n3798 & n8796 ;
  assign n8798 = ( ~n2787 & n7372 ) | ( ~n2787 & n8797 ) | ( n7372 & n8797 ) ;
  assign n8799 = ( n3143 & n8795 ) | ( n3143 & n8798 ) | ( n8795 & n8798 ) ;
  assign n8800 = n8799 ^ n5422 ^ n3873 ;
  assign n8801 = ( n862 & ~n2471 ) | ( n862 & n3324 ) | ( ~n2471 & n3324 ) ;
  assign n8802 = n5217 & n7824 ;
  assign n8803 = n3483 & n8802 ;
  assign n8804 = n8803 ^ n8032 ^ n2206 ;
  assign n8805 = ( n235 & n8801 ) | ( n235 & n8804 ) | ( n8801 & n8804 ) ;
  assign n8806 = n3642 ^ n3105 ^ n2546 ;
  assign n8807 = ( n2549 & n5114 ) | ( n2549 & n8806 ) | ( n5114 & n8806 ) ;
  assign n8808 = n8186 ^ n7040 ^ n3983 ;
  assign n8809 = n7039 ^ n4076 ^ n2428 ;
  assign n8810 = n201 & n2891 ;
  assign n8811 = ( n2050 & ~n5069 ) | ( n2050 & n8810 ) | ( ~n5069 & n8810 ) ;
  assign n8812 = n8811 ^ n2962 ^ 1'b0 ;
  assign n8813 = n8809 & n8812 ;
  assign n8814 = ( ~n691 & n4156 ) | ( ~n691 & n8568 ) | ( n4156 & n8568 ) ;
  assign n8815 = ( n3422 & ~n6335 ) | ( n3422 & n7303 ) | ( ~n6335 & n7303 ) ;
  assign n8816 = n1079 ^ n793 ^ x85 ;
  assign n8817 = n8816 ^ n6727 ^ n1478 ;
  assign n8818 = n8817 ^ n3481 ^ n975 ;
  assign n8819 = ( n7201 & n7938 ) | ( n7201 & n8818 ) | ( n7938 & n8818 ) ;
  assign n8823 = ( ~n1077 & n4104 ) | ( ~n1077 & n5713 ) | ( n4104 & n5713 ) ;
  assign n8820 = ( n553 & n1150 ) | ( n553 & n4174 ) | ( n1150 & n4174 ) ;
  assign n8821 = ( ~n601 & n2023 ) | ( ~n601 & n8820 ) | ( n2023 & n8820 ) ;
  assign n8822 = n8821 ^ n8031 ^ n5312 ;
  assign n8824 = n8823 ^ n8822 ^ n8129 ;
  assign n8825 = ( n142 & n6004 ) | ( n142 & ~n7757 ) | ( n6004 & ~n7757 ) ;
  assign n8826 = n3205 ^ n2486 ^ 1'b0 ;
  assign n8827 = ( n351 & ~n2702 ) | ( n351 & n3276 ) | ( ~n2702 & n3276 ) ;
  assign n8828 = n7465 & n8827 ;
  assign n8829 = n3091 & n8828 ;
  assign n8830 = n5112 | n5223 ;
  assign n8831 = n1119 & ~n8830 ;
  assign n8832 = n5288 ^ n2485 ^ n1761 ;
  assign n8833 = n6707 & ~n8832 ;
  assign n8834 = n3924 & n8833 ;
  assign n8835 = n8834 ^ n4842 ^ 1'b0 ;
  assign n8836 = n4022 & n8835 ;
  assign n8837 = ( n837 & n1886 ) | ( n837 & n6435 ) | ( n1886 & n6435 ) ;
  assign n8839 = n4382 ^ n3927 ^ n1803 ;
  assign n8838 = ( ~n448 & n2457 ) | ( ~n448 & n3311 ) | ( n2457 & n3311 ) ;
  assign n8840 = n8839 ^ n8838 ^ n1562 ;
  assign n8841 = ( n4925 & n8837 ) | ( n4925 & ~n8840 ) | ( n8837 & ~n8840 ) ;
  assign n8842 = ( n6529 & n8836 ) | ( n6529 & n8841 ) | ( n8836 & n8841 ) ;
  assign n8843 = n8517 ^ n5581 ^ 1'b0 ;
  assign n8847 = ( n199 & n693 ) | ( n199 & n8412 ) | ( n693 & n8412 ) ;
  assign n8846 = n5224 ^ n4945 ^ n4783 ;
  assign n8844 = n5012 ^ n4381 ^ 1'b0 ;
  assign n8845 = n2502 | n8844 ;
  assign n8848 = n8847 ^ n8846 ^ n8845 ;
  assign n8849 = n8848 ^ n5291 ^ n1775 ;
  assign n8850 = ( ~n1187 & n8843 ) | ( ~n1187 & n8849 ) | ( n8843 & n8849 ) ;
  assign n8851 = n8850 ^ n6264 ^ 1'b0 ;
  assign n8853 = n695 & n5068 ;
  assign n8854 = n8853 ^ n1324 ^ 1'b0 ;
  assign n8852 = ( n667 & n4363 ) | ( n667 & ~n5769 ) | ( n4363 & ~n5769 ) ;
  assign n8855 = n8854 ^ n8852 ^ n5634 ;
  assign n8858 = ~n1227 & n4302 ;
  assign n8856 = n5682 ^ n4124 ^ 1'b0 ;
  assign n8857 = n808 & ~n8856 ;
  assign n8859 = n8858 ^ n8857 ^ 1'b0 ;
  assign n8862 = n7326 ^ n5671 ^ n2445 ;
  assign n8863 = n8862 ^ n3842 ^ n1198 ;
  assign n8860 = n8357 ^ n1254 ^ 1'b0 ;
  assign n8861 = n8860 ^ n6114 ^ n3253 ;
  assign n8864 = n8863 ^ n8861 ^ n8457 ;
  assign n8865 = n5533 & ~n8864 ;
  assign n8866 = n1446 ^ n639 ^ n208 ;
  assign n8867 = n8866 ^ n5425 ^ n1697 ;
  assign n8870 = n4248 ^ n996 ^ 1'b0 ;
  assign n8871 = n8870 ^ n1471 ^ n1172 ;
  assign n8868 = n3286 ^ n3228 ^ n1934 ;
  assign n8869 = n8868 ^ n7869 ^ n1569 ;
  assign n8872 = n8871 ^ n8869 ^ n7932 ;
  assign n8873 = n4057 ^ n759 ^ 1'b0 ;
  assign n8874 = n3206 ^ n458 ^ 1'b0 ;
  assign n8875 = n857 & n8874 ;
  assign n8876 = n8875 ^ n3114 ^ 1'b0 ;
  assign n8877 = ( n6809 & n7479 ) | ( n6809 & ~n8068 ) | ( n7479 & ~n8068 ) ;
  assign n8890 = n1892 ^ n719 ^ n418 ;
  assign n8889 = n6525 ^ n2139 ^ 1'b0 ;
  assign n8878 = ( ~n4240 & n7195 ) | ( ~n4240 & n7850 ) | ( n7195 & n7850 ) ;
  assign n8879 = ( ~n1716 & n5852 ) | ( ~n1716 & n8878 ) | ( n5852 & n8878 ) ;
  assign n8883 = n3812 ^ n2463 ^ n1267 ;
  assign n8884 = n8883 ^ n4976 ^ n1279 ;
  assign n8881 = n3817 ^ n3325 ^ n2201 ;
  assign n8880 = n7130 & n7149 ;
  assign n8882 = n8881 ^ n8880 ^ 1'b0 ;
  assign n8885 = n8884 ^ n8882 ^ n2680 ;
  assign n8886 = ~n8879 & n8885 ;
  assign n8887 = n8150 ^ n4555 ^ 1'b0 ;
  assign n8888 = ~n8886 & n8887 ;
  assign n8891 = n8890 ^ n8889 ^ n8888 ;
  assign n8899 = n2297 ^ n1836 ^ 1'b0 ;
  assign n8900 = n1228 & ~n8899 ;
  assign n8892 = ~n5548 & n6312 ;
  assign n8893 = n2363 & n8892 ;
  assign n8894 = n6495 ^ n3660 ^ n1806 ;
  assign n8895 = ~n8893 & n8894 ;
  assign n8896 = n8895 ^ n5365 ^ 1'b0 ;
  assign n8897 = n8896 ^ n4495 ^ 1'b0 ;
  assign n8898 = ( n2291 & ~n7929 ) | ( n2291 & n8897 ) | ( ~n7929 & n8897 ) ;
  assign n8901 = n8900 ^ n8898 ^ n2279 ;
  assign n8905 = x115 & ~n751 ;
  assign n8906 = n1044 & n8905 ;
  assign n8903 = ( n1733 & ~n1978 ) | ( n1733 & n3640 ) | ( ~n1978 & n3640 ) ;
  assign n8904 = n8903 ^ n2775 ^ n2028 ;
  assign n8907 = n8906 ^ n8904 ^ n3303 ;
  assign n8902 = n7698 ^ n7433 ^ n3923 ;
  assign n8908 = n8907 ^ n8902 ^ n4410 ;
  assign n8909 = ( n2608 & n2764 ) | ( n2608 & ~n5328 ) | ( n2764 & ~n5328 ) ;
  assign n8910 = n4195 ^ n3976 ^ n3855 ;
  assign n8911 = n4968 & ~n8910 ;
  assign n8912 = ~n8909 & n8911 ;
  assign n8913 = ( ~n1319 & n4304 ) | ( ~n1319 & n6008 ) | ( n4304 & n6008 ) ;
  assign n8914 = n8913 ^ n3094 ^ n216 ;
  assign n8915 = n6818 ^ n2708 ^ n2006 ;
  assign n8916 = n4987 ^ n2512 ^ n2177 ;
  assign n8917 = ~n6231 & n8916 ;
  assign n8918 = ~n5702 & n8917 ;
  assign n8919 = n7998 ^ n3980 ^ n2936 ;
  assign n8924 = ( n2342 & ~n3912 ) | ( n2342 & n7184 ) | ( ~n3912 & n7184 ) ;
  assign n8925 = n8924 ^ n4357 ^ n1669 ;
  assign n8920 = n6639 ^ n5332 ^ n4668 ;
  assign n8921 = ( n509 & n1472 ) | ( n509 & ~n2265 ) | ( n1472 & ~n2265 ) ;
  assign n8922 = n8921 ^ n3023 ^ 1'b0 ;
  assign n8923 = ( ~n658 & n8920 ) | ( ~n658 & n8922 ) | ( n8920 & n8922 ) ;
  assign n8926 = n8925 ^ n8923 ^ n4036 ;
  assign n8927 = n6078 ^ n5494 ^ n5045 ;
  assign n8928 = n822 | n8927 ;
  assign n8929 = n8926 | n8928 ;
  assign n8930 = n8300 ^ n2895 ^ n1229 ;
  assign n8931 = n2512 & ~n8930 ;
  assign n8932 = n8931 ^ n5202 ^ n209 ;
  assign n8933 = n8932 ^ n7476 ^ 1'b0 ;
  assign n8934 = n734 & n5955 ;
  assign n8935 = n2135 ^ n1511 ^ 1'b0 ;
  assign n8936 = n8935 ^ n5232 ^ 1'b0 ;
  assign n8937 = n4671 ^ n3599 ^ n2375 ;
  assign n8938 = n3294 ^ n1996 ^ n468 ;
  assign n8939 = ( n6413 & n7931 ) | ( n6413 & ~n8938 ) | ( n7931 & ~n8938 ) ;
  assign n8940 = ( n6621 & n8937 ) | ( n6621 & n8939 ) | ( n8937 & n8939 ) ;
  assign n8941 = n8764 ^ n5014 ^ n1346 ;
  assign n8942 = ( n3766 & n6482 ) | ( n3766 & ~n8941 ) | ( n6482 & ~n8941 ) ;
  assign n8943 = ( n7152 & n8940 ) | ( n7152 & n8942 ) | ( n8940 & n8942 ) ;
  assign n8944 = n5416 ^ n4148 ^ x41 ;
  assign n8945 = n8944 ^ n7312 ^ n3459 ;
  assign n8950 = n3010 & ~n5578 ;
  assign n8946 = n5514 ^ n344 ^ 1'b0 ;
  assign n8947 = ~n2624 & n8946 ;
  assign n8948 = ( n646 & n2377 ) | ( n646 & ~n8947 ) | ( n2377 & ~n8947 ) ;
  assign n8949 = n8948 ^ n7588 ^ x101 ;
  assign n8951 = n8950 ^ n8949 ^ n2441 ;
  assign n8952 = n1458 ^ n949 ^ 1'b0 ;
  assign n8953 = n3481 | n7101 ;
  assign n8954 = n8953 ^ n1657 ^ 1'b0 ;
  assign n8955 = n8954 ^ n7718 ^ n6660 ;
  assign n8956 = n2980 & n3860 ;
  assign n8965 = ( n565 & n2637 ) | ( n565 & n4695 ) | ( n2637 & n4695 ) ;
  assign n8966 = n8965 ^ n3825 ^ n237 ;
  assign n8960 = x47 & n1910 ;
  assign n8961 = n8960 ^ n8319 ^ 1'b0 ;
  assign n8962 = n8961 ^ n4691 ^ 1'b0 ;
  assign n8959 = n3154 & ~n8832 ;
  assign n8963 = n8962 ^ n8959 ^ 1'b0 ;
  assign n8957 = n6770 ^ n4243 ^ 1'b0 ;
  assign n8958 = ( ~n4555 & n7424 ) | ( ~n4555 & n8957 ) | ( n7424 & n8957 ) ;
  assign n8964 = n8963 ^ n8958 ^ n3384 ;
  assign n8967 = n8966 ^ n8964 ^ 1'b0 ;
  assign n8968 = ~n8956 & n8967 ;
  assign n8970 = n978 ^ n834 ^ 1'b0 ;
  assign n8969 = ( n4485 & ~n4585 ) | ( n4485 & n7665 ) | ( ~n4585 & n7665 ) ;
  assign n8971 = n8970 ^ n8969 ^ n7953 ;
  assign n8975 = n1959 ^ n865 ^ 1'b0 ;
  assign n8976 = n1186 & n8975 ;
  assign n8972 = n1277 | n6679 ;
  assign n8973 = ( n357 & ~n5338 ) | ( n357 & n8972 ) | ( ~n5338 & n8972 ) ;
  assign n8974 = ( ~n1977 & n6972 ) | ( ~n1977 & n8973 ) | ( n6972 & n8973 ) ;
  assign n8977 = n8976 ^ n8974 ^ n8732 ;
  assign n8978 = n8867 ^ n1697 ^ 1'b0 ;
  assign n8979 = n8977 & n8978 ;
  assign n8980 = n6824 ^ n1291 ^ n718 ;
  assign n8984 = n3361 ^ n2095 ^ n1655 ;
  assign n8985 = n8984 ^ n3397 ^ n3370 ;
  assign n8986 = n8985 ^ n7151 ^ n5752 ;
  assign n8987 = n8296 ^ n8014 ^ 1'b0 ;
  assign n8988 = n8986 | n8987 ;
  assign n8981 = n8264 ^ n5973 ^ 1'b0 ;
  assign n8982 = n2465 & n8981 ;
  assign n8983 = n2507 & n8982 ;
  assign n8989 = n8988 ^ n8983 ^ n180 ;
  assign n8990 = n7308 ^ n2716 ^ n753 ;
  assign n8991 = n3514 ^ n1412 ^ 1'b0 ;
  assign n8992 = n2492 | n8991 ;
  assign n8993 = n3299 & ~n8992 ;
  assign n8994 = n8993 ^ n4514 ^ n1560 ;
  assign n8995 = n5194 ^ n3993 ^ 1'b0 ;
  assign n8996 = n3004 & n8995 ;
  assign n8997 = ( n2360 & n5630 ) | ( n2360 & ~n6397 ) | ( n5630 & ~n6397 ) ;
  assign n8998 = n6951 & n8997 ;
  assign n8999 = ( ~x113 & n8996 ) | ( ~x113 & n8998 ) | ( n8996 & n8998 ) ;
  assign n9010 = n6338 ^ n4828 ^ n1497 ;
  assign n9011 = n9010 ^ n8199 ^ n6465 ;
  assign n9004 = n4784 ^ n2313 ^ 1'b0 ;
  assign n9005 = n7918 & n9004 ;
  assign n9006 = ( n2635 & n2987 ) | ( n2635 & n9005 ) | ( n2987 & n9005 ) ;
  assign n9007 = n4008 | n9006 ;
  assign n9000 = n4821 ^ n3338 ^ 1'b0 ;
  assign n9001 = n2066 & ~n9000 ;
  assign n9002 = ( ~n933 & n1243 ) | ( ~n933 & n9001 ) | ( n1243 & n9001 ) ;
  assign n9003 = n1219 & n9002 ;
  assign n9008 = n9007 ^ n9003 ^ 1'b0 ;
  assign n9009 = ( n1013 & n3808 ) | ( n1013 & ~n9008 ) | ( n3808 & ~n9008 ) ;
  assign n9012 = n9011 ^ n9009 ^ n4254 ;
  assign n9013 = n7112 | n9012 ;
  assign n9014 = n8801 ^ n8178 ^ 1'b0 ;
  assign n9015 = n2965 & ~n8955 ;
  assign n9016 = ~n9014 & n9015 ;
  assign n9018 = n5502 ^ n5072 ^ n2802 ;
  assign n9017 = n1016 ^ n177 ^ n142 ;
  assign n9019 = n9018 ^ n9017 ^ n5687 ;
  assign n9024 = n2643 & n2677 ;
  assign n9025 = ( n1228 & ~n4966 ) | ( n1228 & n9024 ) | ( ~n4966 & n9024 ) ;
  assign n9020 = n1868 ^ n147 ^ 1'b0 ;
  assign n9021 = n800 & n2089 ;
  assign n9022 = n187 & n9021 ;
  assign n9023 = ( n2651 & n9020 ) | ( n2651 & n9022 ) | ( n9020 & n9022 ) ;
  assign n9026 = n9025 ^ n9023 ^ n3706 ;
  assign n9027 = n9026 ^ n6120 ^ n1025 ;
  assign n9028 = ( n3606 & n7588 ) | ( n3606 & n7716 ) | ( n7588 & n7716 ) ;
  assign n9029 = ( n4721 & n8316 ) | ( n4721 & n9028 ) | ( n8316 & n9028 ) ;
  assign n9030 = ( n811 & n3928 ) | ( n811 & ~n5504 ) | ( n3928 & ~n5504 ) ;
  assign n9031 = n8227 ^ n6309 ^ n3800 ;
  assign n9032 = ( ~n558 & n1804 ) | ( ~n558 & n2960 ) | ( n1804 & n2960 ) ;
  assign n9033 = n9032 ^ n4913 ^ n986 ;
  assign n9034 = ( n9030 & ~n9031 ) | ( n9030 & n9033 ) | ( ~n9031 & n9033 ) ;
  assign n9035 = ( n389 & ~n4161 ) | ( n389 & n5115 ) | ( ~n4161 & n5115 ) ;
  assign n9036 = ( n877 & n4096 ) | ( n877 & n4203 ) | ( n4096 & n4203 ) ;
  assign n9037 = ( n191 & n9035 ) | ( n191 & ~n9036 ) | ( n9035 & ~n9036 ) ;
  assign n9038 = ( ~n3620 & n4168 ) | ( ~n3620 & n9037 ) | ( n4168 & n9037 ) ;
  assign n9039 = n9038 ^ n9018 ^ n5253 ;
  assign n9040 = n9039 ^ n5321 ^ n1740 ;
  assign n9041 = n7307 ^ n6830 ^ 1'b0 ;
  assign n9042 = n8444 ^ n2940 ^ n651 ;
  assign n9043 = n2920 & n4744 ;
  assign n9044 = n9043 ^ n2307 ^ n1049 ;
  assign n9045 = n9044 ^ n7898 ^ n876 ;
  assign n9046 = ( n844 & n1262 ) | ( n844 & ~n7310 ) | ( n1262 & ~n7310 ) ;
  assign n9047 = ( n1054 & n3802 ) | ( n1054 & n9046 ) | ( n3802 & n9046 ) ;
  assign n9048 = ( ~n238 & n1778 ) | ( ~n238 & n9047 ) | ( n1778 & n9047 ) ;
  assign n9049 = ( ~n9042 & n9045 ) | ( ~n9042 & n9048 ) | ( n9045 & n9048 ) ;
  assign n9057 = ~n2175 & n5658 ;
  assign n9058 = n9057 ^ n2764 ^ 1'b0 ;
  assign n9050 = n8414 ^ n285 ^ 1'b0 ;
  assign n9051 = n3899 ^ n2821 ^ 1'b0 ;
  assign n9052 = n9051 ^ n654 ^ 1'b0 ;
  assign n9053 = n9050 | n9052 ;
  assign n9054 = n280 | n3112 ;
  assign n9055 = n9054 ^ n2906 ^ 1'b0 ;
  assign n9056 = n9053 | n9055 ;
  assign n9059 = n9058 ^ n9056 ^ n8368 ;
  assign n9060 = n9059 ^ n5183 ^ n4373 ;
  assign n9063 = n8508 ^ n4995 ^ 1'b0 ;
  assign n9064 = n198 & ~n9063 ;
  assign n9061 = ( n453 & n1189 ) | ( n453 & n4819 ) | ( n1189 & n4819 ) ;
  assign n9062 = ( n1521 & n2591 ) | ( n1521 & ~n9061 ) | ( n2591 & ~n9061 ) ;
  assign n9065 = n9064 ^ n9062 ^ n603 ;
  assign n9066 = n4554 ^ n1545 ^ 1'b0 ;
  assign n9067 = n5206 | n9066 ;
  assign n9068 = ( n1114 & n7340 ) | ( n1114 & n9067 ) | ( n7340 & n9067 ) ;
  assign n9069 = n817 & n9068 ;
  assign n9070 = n2092 ^ n780 ^ n249 ;
  assign n9073 = ( n4266 & n5185 ) | ( n4266 & n6591 ) | ( n5185 & n6591 ) ;
  assign n9074 = n5182 & ~n9073 ;
  assign n9075 = n9074 ^ n2457 ^ 1'b0 ;
  assign n9071 = n926 & ~n6885 ;
  assign n9072 = n9071 ^ n6319 ^ 1'b0 ;
  assign n9076 = n9075 ^ n9072 ^ n5544 ;
  assign n9077 = n7255 ^ n6889 ^ n647 ;
  assign n9078 = n1496 & ~n8372 ;
  assign n9079 = n5517 & n9078 ;
  assign n9080 = n1371 & ~n2007 ;
  assign n9081 = n2745 ^ n2143 ^ 1'b0 ;
  assign n9082 = n9080 | n9081 ;
  assign n9083 = ( ~n8375 & n9079 ) | ( ~n8375 & n9082 ) | ( n9079 & n9082 ) ;
  assign n9084 = ( n2795 & n3073 ) | ( n2795 & ~n6664 ) | ( n3073 & ~n6664 ) ;
  assign n9085 = ~n9083 & n9084 ;
  assign n9086 = ~n9077 & n9085 ;
  assign n9087 = n510 & ~n2959 ;
  assign n9088 = ~n8788 & n9087 ;
  assign n9089 = ( n1421 & n5701 ) | ( n1421 & ~n9088 ) | ( n5701 & ~n9088 ) ;
  assign n9090 = n3534 ^ n511 ^ 1'b0 ;
  assign n9091 = ( n505 & n4696 ) | ( n505 & n9090 ) | ( n4696 & n9090 ) ;
  assign n9093 = n3199 ^ n2291 ^ n840 ;
  assign n9092 = ( n811 & n4382 ) | ( n811 & n8647 ) | ( n4382 & n8647 ) ;
  assign n9094 = n9093 ^ n9092 ^ n6225 ;
  assign n9095 = ( n6829 & n9091 ) | ( n6829 & ~n9094 ) | ( n9091 & ~n9094 ) ;
  assign n9096 = n9095 ^ n8049 ^ 1'b0 ;
  assign n9098 = n1570 | n5069 ;
  assign n9099 = n4998 & n9098 ;
  assign n9100 = n9099 ^ n5329 ^ 1'b0 ;
  assign n9097 = n4903 ^ n4487 ^ n4387 ;
  assign n9101 = n9100 ^ n9097 ^ n3812 ;
  assign n9102 = ~n1263 & n8009 ;
  assign n9103 = ~n1191 & n9102 ;
  assign n9104 = ( n2616 & ~n2976 ) | ( n2616 & n3400 ) | ( ~n2976 & n3400 ) ;
  assign n9105 = n9104 ^ n4373 ^ 1'b0 ;
  assign n9106 = ~n1707 & n9105 ;
  assign n9107 = n9106 ^ n3423 ^ 1'b0 ;
  assign n9108 = n6905 & n9107 ;
  assign n9109 = ( n678 & ~n6369 ) | ( n678 & n6454 ) | ( ~n6369 & n6454 ) ;
  assign n9110 = n9109 ^ n8958 ^ n3868 ;
  assign n9111 = n1920 ^ n1125 ^ n579 ;
  assign n9112 = ( n7489 & ~n8254 ) | ( n7489 & n9111 ) | ( ~n8254 & n9111 ) ;
  assign n9113 = ( n4176 & n4417 ) | ( n4176 & ~n6103 ) | ( n4417 & ~n6103 ) ;
  assign n9114 = n9113 ^ n4720 ^ n4202 ;
  assign n9115 = n9114 ^ n9054 ^ n4474 ;
  assign n9116 = n9115 ^ n3877 ^ n1542 ;
  assign n9117 = ( ~n341 & n1369 ) | ( ~n341 & n5882 ) | ( n1369 & n5882 ) ;
  assign n9118 = ( n4102 & ~n8158 ) | ( n4102 & n9117 ) | ( ~n8158 & n9117 ) ;
  assign n9119 = ( n204 & ~n5722 ) | ( n204 & n8143 ) | ( ~n5722 & n8143 ) ;
  assign n9120 = ( n7798 & n7911 ) | ( n7798 & ~n9119 ) | ( n7911 & ~n9119 ) ;
  assign n9121 = n8972 ^ n5707 ^ n3141 ;
  assign n9122 = n9121 ^ n3461 ^ n1518 ;
  assign n9123 = n3852 | n5026 ;
  assign n9124 = n9122 & ~n9123 ;
  assign n9125 = ( ~n3276 & n9120 ) | ( ~n3276 & n9124 ) | ( n9120 & n9124 ) ;
  assign n9126 = ( n7783 & n9118 ) | ( n7783 & n9125 ) | ( n9118 & n9125 ) ;
  assign n9135 = n3916 ^ n256 ^ 1'b0 ;
  assign n9136 = ~n2905 & n9135 ;
  assign n9137 = ~n1894 & n9136 ;
  assign n9138 = n9137 ^ n6234 ^ 1'b0 ;
  assign n9139 = ~n3030 & n9138 ;
  assign n9140 = n5114 | n9139 ;
  assign n9130 = n5082 ^ n2872 ^ 1'b0 ;
  assign n9131 = n5184 & ~n9130 ;
  assign n9132 = n498 | n710 ;
  assign n9133 = n9131 | n9132 ;
  assign n9127 = n780 & ~n1515 ;
  assign n9128 = n3666 ^ n1995 ^ n1050 ;
  assign n9129 = ~n9127 & n9128 ;
  assign n9134 = n9133 ^ n9129 ^ n2835 ;
  assign n9141 = n9140 ^ n9134 ^ 1'b0 ;
  assign n9142 = ~n6358 & n9141 ;
  assign n9143 = n5574 ^ n5090 ^ 1'b0 ;
  assign n9146 = ~n799 & n2739 ;
  assign n9144 = n8234 ^ n3380 ^ 1'b0 ;
  assign n9145 = n9144 ^ n5368 ^ 1'b0 ;
  assign n9147 = n9146 ^ n9145 ^ n4090 ;
  assign n9148 = n5424 ^ n3268 ^ n2726 ;
  assign n9149 = n2799 | n9148 ;
  assign n9150 = n7279 & ~n9149 ;
  assign n9151 = ( n5885 & ~n6922 ) | ( n5885 & n8549 ) | ( ~n6922 & n8549 ) ;
  assign n9152 = ( n4417 & n8170 ) | ( n4417 & ~n9151 ) | ( n8170 & ~n9151 ) ;
  assign n9153 = n2893 ^ n1062 ^ n646 ;
  assign n9154 = n5031 ^ n4966 ^ n1784 ;
  assign n9155 = ~n576 & n2090 ;
  assign n9156 = ~n5254 & n9155 ;
  assign n9157 = n9156 ^ n8382 ^ n6965 ;
  assign n9158 = n9157 ^ n5773 ^ n4199 ;
  assign n9159 = n9154 | n9158 ;
  assign n9160 = ( ~n8489 & n9153 ) | ( ~n8489 & n9159 ) | ( n9153 & n9159 ) ;
  assign n9161 = ( n2118 & n2135 ) | ( n2118 & n5455 ) | ( n2135 & n5455 ) ;
  assign n9163 = n2191 ^ x25 ^ 1'b0 ;
  assign n9164 = n2654 & ~n9163 ;
  assign n9162 = n788 | n4034 ;
  assign n9165 = n9164 ^ n9162 ^ 1'b0 ;
  assign n9166 = ~n2242 & n3486 ;
  assign n9167 = n1178 & n9166 ;
  assign n9168 = ( n3748 & ~n6905 ) | ( n3748 & n9167 ) | ( ~n6905 & n9167 ) ;
  assign n9169 = n2844 ^ n1186 ^ n276 ;
  assign n9170 = n7873 ^ n4691 ^ n2800 ;
  assign n9171 = n9169 | n9170 ;
  assign n9172 = n9171 ^ n4845 ^ 1'b0 ;
  assign n9173 = ~n4318 & n9172 ;
  assign n9174 = ~n1011 & n5218 ;
  assign n9175 = ~n2535 & n9174 ;
  assign n9176 = ( n285 & ~n1872 ) | ( n285 & n8285 ) | ( ~n1872 & n8285 ) ;
  assign n9178 = n7477 ^ n2683 ^ n2586 ;
  assign n9177 = n2734 & n7184 ;
  assign n9179 = n9178 ^ n9177 ^ 1'b0 ;
  assign n9180 = ( n1732 & ~n9176 ) | ( n1732 & n9179 ) | ( ~n9176 & n9179 ) ;
  assign n9181 = ( ~n7618 & n9175 ) | ( ~n7618 & n9180 ) | ( n9175 & n9180 ) ;
  assign n9182 = n9181 ^ n2999 ^ n603 ;
  assign n9183 = n4220 ^ n146 ^ 1'b0 ;
  assign n9184 = ~n628 & n7124 ;
  assign n9185 = n9184 ^ n6303 ^ 1'b0 ;
  assign n9190 = n1391 & ~n4873 ;
  assign n9191 = n9190 ^ n2353 ^ 1'b0 ;
  assign n9186 = n2854 ^ n1438 ^ n727 ;
  assign n9187 = n7203 ^ n1679 ^ 1'b0 ;
  assign n9188 = n9167 | n9187 ;
  assign n9189 = n9186 & ~n9188 ;
  assign n9192 = n9191 ^ n9189 ^ n3114 ;
  assign n9193 = ( ~n9183 & n9185 ) | ( ~n9183 & n9192 ) | ( n9185 & n9192 ) ;
  assign n9202 = ( n1007 & ~n1954 ) | ( n1007 & n2508 ) | ( ~n1954 & n2508 ) ;
  assign n9203 = n9202 ^ n216 ^ 1'b0 ;
  assign n9204 = n9018 | n9203 ;
  assign n9205 = n6390 ^ n4065 ^ n3437 ;
  assign n9206 = n146 | n9205 ;
  assign n9207 = n9204 & ~n9206 ;
  assign n9194 = n7233 ^ n4722 ^ n3397 ;
  assign n9196 = n6170 & n6976 ;
  assign n9197 = n9196 ^ n3231 ^ 1'b0 ;
  assign n9198 = n9197 ^ n2967 ^ n778 ;
  assign n9195 = ( n1044 & n5309 ) | ( n1044 & n6261 ) | ( n5309 & n6261 ) ;
  assign n9199 = n9198 ^ n9195 ^ 1'b0 ;
  assign n9200 = ~n9194 & n9199 ;
  assign n9201 = n7406 & n9200 ;
  assign n9208 = n9207 ^ n9201 ^ 1'b0 ;
  assign n9209 = n8831 ^ n8209 ^ 1'b0 ;
  assign n9210 = n1661 ^ n1117 ^ n465 ;
  assign n9211 = n7415 ^ n3590 ^ 1'b0 ;
  assign n9212 = ~n8538 & n9211 ;
  assign n9213 = ( n6420 & ~n9210 ) | ( n6420 & n9212 ) | ( ~n9210 & n9212 ) ;
  assign n9214 = ( ~x119 & n3693 ) | ( ~x119 & n4011 ) | ( n3693 & n4011 ) ;
  assign n9215 = ( ~n340 & n3144 ) | ( ~n340 & n5060 ) | ( n3144 & n5060 ) ;
  assign n9216 = n2905 ^ n1159 ^ n1095 ;
  assign n9217 = n3835 & ~n9216 ;
  assign n9218 = n9215 & n9217 ;
  assign n9219 = ( n2555 & n3442 ) | ( n2555 & n9218 ) | ( n3442 & n9218 ) ;
  assign n9220 = ( n534 & ~n6407 ) | ( n534 & n9219 ) | ( ~n6407 & n9219 ) ;
  assign n9221 = ( n1721 & n3140 ) | ( n1721 & n6473 ) | ( n3140 & n6473 ) ;
  assign n9222 = n2812 ^ n1419 ^ 1'b0 ;
  assign n9223 = ( n2854 & ~n3458 ) | ( n2854 & n9222 ) | ( ~n3458 & n9222 ) ;
  assign n9224 = ( n2413 & n9221 ) | ( n2413 & ~n9223 ) | ( n9221 & ~n9223 ) ;
  assign n9225 = ( n1479 & n2260 ) | ( n1479 & ~n2499 ) | ( n2260 & ~n2499 ) ;
  assign n9226 = ( n2408 & ~n2724 ) | ( n2408 & n3088 ) | ( ~n2724 & n3088 ) ;
  assign n9227 = ( n2601 & n6672 ) | ( n2601 & n9226 ) | ( n6672 & n9226 ) ;
  assign n9228 = ( n6771 & n9225 ) | ( n6771 & ~n9227 ) | ( n9225 & ~n9227 ) ;
  assign n9229 = ( ~n6293 & n9224 ) | ( ~n6293 & n9228 ) | ( n9224 & n9228 ) ;
  assign n9230 = n9229 ^ n5631 ^ n4471 ;
  assign n9231 = n4148 ^ n1607 ^ 1'b0 ;
  assign n9232 = n9231 ^ n3136 ^ n1308 ;
  assign n9233 = n9232 ^ n8138 ^ n6647 ;
  assign n9234 = n6824 ^ n3236 ^ n3066 ;
  assign n9237 = ( n3372 & n4744 ) | ( n3372 & ~n7980 ) | ( n4744 & ~n7980 ) ;
  assign n9235 = n3946 ^ n2083 ^ 1'b0 ;
  assign n9236 = n3339 | n9235 ;
  assign n9238 = n9237 ^ n9236 ^ n7315 ;
  assign n9239 = n8958 ^ n4465 ^ n1263 ;
  assign n9240 = ( n2106 & n3621 ) | ( n2106 & n8634 ) | ( n3621 & n8634 ) ;
  assign n9241 = n781 ^ n550 ^ 1'b0 ;
  assign n9242 = n6486 ^ x123 ^ 1'b0 ;
  assign n9243 = n1657 & n9242 ;
  assign n9244 = n9243 ^ n6773 ^ n3184 ;
  assign n9245 = n9241 & n9244 ;
  assign n9248 = n3524 ^ n795 ^ 1'b0 ;
  assign n9246 = n2218 & n2742 ;
  assign n9247 = n9246 ^ n7503 ^ 1'b0 ;
  assign n9249 = n9248 ^ n9247 ^ n926 ;
  assign n9250 = n9249 ^ n6209 ^ n4667 ;
  assign n9257 = ( n826 & ~n3222 ) | ( n826 & n5355 ) | ( ~n3222 & n5355 ) ;
  assign n9258 = ( n3872 & n3941 ) | ( n3872 & n9257 ) | ( n3941 & n9257 ) ;
  assign n9261 = ( ~n206 & n1392 ) | ( ~n206 & n1636 ) | ( n1392 & n1636 ) ;
  assign n9259 = n3497 ^ n3352 ^ n541 ;
  assign n9260 = n3188 | n9259 ;
  assign n9262 = n9261 ^ n9260 ^ 1'b0 ;
  assign n9263 = ( n4813 & n9258 ) | ( n4813 & ~n9262 ) | ( n9258 & ~n9262 ) ;
  assign n9251 = n5063 ^ n424 ^ 1'b0 ;
  assign n9252 = n1266 & n3694 ;
  assign n9253 = ( n2846 & ~n5694 ) | ( n2846 & n9252 ) | ( ~n5694 & n9252 ) ;
  assign n9254 = ( n959 & ~n1956 ) | ( n959 & n2587 ) | ( ~n1956 & n2587 ) ;
  assign n9255 = n9253 & n9254 ;
  assign n9256 = ( n8422 & n9251 ) | ( n8422 & ~n9255 ) | ( n9251 & ~n9255 ) ;
  assign n9264 = n9263 ^ n9256 ^ n8938 ;
  assign n9266 = n5279 ^ n1198 ^ n411 ;
  assign n9265 = n3140 ^ n3048 ^ 1'b0 ;
  assign n9267 = n9266 ^ n9265 ^ n3822 ;
  assign n9268 = x103 & n9267 ;
  assign n9269 = n3281 ^ n1965 ^ 1'b0 ;
  assign n9270 = ( n813 & ~n3294 ) | ( n813 & n3543 ) | ( ~n3294 & n3543 ) ;
  assign n9271 = n9270 ^ n182 ^ 1'b0 ;
  assign n9272 = ( n4079 & n7559 ) | ( n4079 & ~n9271 ) | ( n7559 & ~n9271 ) ;
  assign n9273 = ~n5232 & n9272 ;
  assign n9274 = n9269 & n9273 ;
  assign n9280 = n3158 ^ n1799 ^ n1584 ;
  assign n9278 = n1457 ^ n246 ^ 1'b0 ;
  assign n9279 = ( n1555 & ~n2688 ) | ( n1555 & n9278 ) | ( ~n2688 & n9278 ) ;
  assign n9275 = n2047 | n2732 ;
  assign n9276 = n9275 ^ n1918 ^ 1'b0 ;
  assign n9277 = n9276 ^ n5218 ^ n3387 ;
  assign n9281 = n9280 ^ n9279 ^ n9277 ;
  assign n9282 = ( n7864 & n8292 ) | ( n7864 & n8423 ) | ( n8292 & n8423 ) ;
  assign n9283 = n525 & ~n3137 ;
  assign n9284 = n7838 ^ n2168 ^ 1'b0 ;
  assign n9285 = n2496 & n4868 ;
  assign n9286 = n1281 & ~n2697 ;
  assign n9287 = x126 & n9286 ;
  assign n9288 = ~n4722 & n9287 ;
  assign n9289 = n9285 & ~n9288 ;
  assign n9290 = n9289 ^ n4847 ^ 1'b0 ;
  assign n9292 = n2751 ^ n2398 ^ 1'b0 ;
  assign n9293 = n9292 ^ n7354 ^ n1948 ;
  assign n9291 = n4096 | n4810 ;
  assign n9294 = n9293 ^ n9291 ^ n7716 ;
  assign n9303 = ( n584 & n781 ) | ( n584 & ~n1169 ) | ( n781 & ~n1169 ) ;
  assign n9304 = n9303 ^ n6967 ^ n6421 ;
  assign n9301 = ( n1126 & n3603 ) | ( n1126 & n9131 ) | ( n3603 & n9131 ) ;
  assign n9298 = ( n1718 & n1762 ) | ( n1718 & n4133 ) | ( n1762 & n4133 ) ;
  assign n9299 = n2023 & n9298 ;
  assign n9300 = n9299 ^ n4109 ^ 1'b0 ;
  assign n9302 = n9301 ^ n9300 ^ n6806 ;
  assign n9295 = ( ~n833 & n3907 ) | ( ~n833 & n4098 ) | ( n3907 & n4098 ) ;
  assign n9296 = ( ~n867 & n2380 ) | ( ~n867 & n2589 ) | ( n2380 & n2589 ) ;
  assign n9297 = ( n1596 & ~n9295 ) | ( n1596 & n9296 ) | ( ~n9295 & n9296 ) ;
  assign n9305 = n9304 ^ n9302 ^ n9297 ;
  assign n9306 = ( n1257 & n1406 ) | ( n1257 & n3335 ) | ( n1406 & n3335 ) ;
  assign n9307 = n9306 ^ n2591 ^ n1523 ;
  assign n9308 = n9307 ^ n2739 ^ 1'b0 ;
  assign n9320 = n8136 ^ n1623 ^ n1347 ;
  assign n9321 = n9320 ^ n4701 ^ n3464 ;
  assign n9315 = n1557 & ~n2488 ;
  assign n9316 = n9315 ^ n3339 ^ 1'b0 ;
  assign n9317 = n9316 ^ n332 ^ 1'b0 ;
  assign n9318 = ~n7220 & n9317 ;
  assign n9319 = n9318 ^ n681 ^ 1'b0 ;
  assign n9309 = x124 & ~n182 ;
  assign n9310 = n925 ^ n260 ^ 1'b0 ;
  assign n9311 = n5491 | n9310 ;
  assign n9312 = n7016 ^ n6203 ^ 1'b0 ;
  assign n9313 = ~n9311 & n9312 ;
  assign n9314 = ~n9309 & n9313 ;
  assign n9322 = n9321 ^ n9319 ^ n9314 ;
  assign n9323 = ( n8321 & ~n9308 ) | ( n8321 & n9322 ) | ( ~n9308 & n9322 ) ;
  assign n9332 = ( n1471 & n3970 ) | ( n1471 & n4234 ) | ( n3970 & n4234 ) ;
  assign n9333 = n3677 ^ n3082 ^ 1'b0 ;
  assign n9334 = n9333 ^ n160 ^ 1'b0 ;
  assign n9335 = n7541 | n9334 ;
  assign n9336 = n9335 ^ n5216 ^ 1'b0 ;
  assign n9337 = n9332 & ~n9336 ;
  assign n9338 = n9337 ^ n3311 ^ 1'b0 ;
  assign n9326 = n5183 ^ n3528 ^ n2461 ;
  assign n9324 = n6529 ^ n6249 ^ n3709 ;
  assign n9325 = n9324 ^ n6280 ^ n4286 ;
  assign n9327 = n9326 ^ n9325 ^ n1316 ;
  assign n9328 = ( ~n1861 & n3026 ) | ( ~n1861 & n3204 ) | ( n3026 & n3204 ) ;
  assign n9329 = ( n988 & ~n6587 ) | ( n988 & n9328 ) | ( ~n6587 & n9328 ) ;
  assign n9330 = n9329 ^ n4211 ^ n2820 ;
  assign n9331 = ( n8846 & ~n9327 ) | ( n8846 & n9330 ) | ( ~n9327 & n9330 ) ;
  assign n9339 = n9338 ^ n9331 ^ n8884 ;
  assign n9340 = ~n475 & n3944 ;
  assign n9341 = ( n1753 & n5148 ) | ( n1753 & n6137 ) | ( n5148 & n6137 ) ;
  assign n9342 = n9340 | n9341 ;
  assign n9343 = n5341 & ~n9342 ;
  assign n9344 = n6030 ^ n2589 ^ n429 ;
  assign n9345 = ( n2436 & ~n5204 ) | ( n2436 & n9344 ) | ( ~n5204 & n9344 ) ;
  assign n9346 = n709 & n7148 ;
  assign n9347 = n9346 ^ n6849 ^ 1'b0 ;
  assign n9348 = ( ~n3067 & n9345 ) | ( ~n3067 & n9347 ) | ( n9345 & n9347 ) ;
  assign n9349 = n9348 ^ n5659 ^ x0 ;
  assign n9350 = n9349 ^ n8489 ^ 1'b0 ;
  assign n9353 = n216 | n2441 ;
  assign n9354 = n808 | n9353 ;
  assign n9355 = n9354 ^ n7310 ^ 1'b0 ;
  assign n9356 = n5912 & n9355 ;
  assign n9351 = ~n545 & n1097 ;
  assign n9352 = ( n5638 & n6277 ) | ( n5638 & n9351 ) | ( n6277 & n9351 ) ;
  assign n9357 = n9356 ^ n9352 ^ n4459 ;
  assign n9358 = n7963 ^ n2545 ^ n1080 ;
  assign n9359 = ( n3322 & n8113 ) | ( n3322 & n9358 ) | ( n8113 & n9358 ) ;
  assign n9360 = ( n1505 & n9143 ) | ( n1505 & ~n9359 ) | ( n9143 & ~n9359 ) ;
  assign n9361 = ( n2851 & n4458 ) | ( n2851 & n9340 ) | ( n4458 & n9340 ) ;
  assign n9362 = ( ~n2281 & n2588 ) | ( ~n2281 & n8419 ) | ( n2588 & n8419 ) ;
  assign n9363 = n9362 ^ n5836 ^ n3640 ;
  assign n9365 = ~n722 & n5096 ;
  assign n9366 = n1687 & n9365 ;
  assign n9364 = n4778 ^ n1398 ^ 1'b0 ;
  assign n9367 = n9366 ^ n9364 ^ n3213 ;
  assign n9368 = n438 & ~n1674 ;
  assign n9369 = ~n7305 & n9368 ;
  assign n9370 = n9369 ^ n8935 ^ 1'b0 ;
  assign n9371 = n6253 ^ n5943 ^ n1314 ;
  assign n9372 = ( n1799 & ~n7333 ) | ( n1799 & n9371 ) | ( ~n7333 & n9371 ) ;
  assign n9373 = ~n3001 & n9372 ;
  assign n9374 = n9373 ^ n2938 ^ 1'b0 ;
  assign n9375 = ( n1511 & n2307 ) | ( n1511 & n4144 ) | ( n2307 & n4144 ) ;
  assign n9376 = ( n8131 & ~n9374 ) | ( n8131 & n9375 ) | ( ~n9374 & n9375 ) ;
  assign n9379 = n8890 ^ n5858 ^ 1'b0 ;
  assign n9377 = n820 & ~n2379 ;
  assign n9378 = ~n3495 & n9377 ;
  assign n9380 = n9379 ^ n9378 ^ n3210 ;
  assign n9381 = n4734 ^ n2502 ^ 1'b0 ;
  assign n9382 = ~n3487 & n9381 ;
  assign n9383 = n9382 ^ n2839 ^ n1761 ;
  assign n9384 = n9383 ^ n8621 ^ n352 ;
  assign n9385 = n9384 ^ n5271 ^ n1643 ;
  assign n9386 = n8035 ^ n6333 ^ 1'b0 ;
  assign n9387 = n8705 ^ n6773 ^ 1'b0 ;
  assign n9388 = ~n6208 & n9387 ;
  assign n9389 = n6319 | n8006 ;
  assign n9390 = ( n2530 & n3553 ) | ( n2530 & ~n5017 ) | ( n3553 & ~n5017 ) ;
  assign n9391 = ( n5605 & ~n7802 ) | ( n5605 & n9390 ) | ( ~n7802 & n9390 ) ;
  assign n9392 = ( n3048 & ~n7117 ) | ( n3048 & n9391 ) | ( ~n7117 & n9391 ) ;
  assign n9393 = n9392 ^ n2683 ^ 1'b0 ;
  assign n9394 = n8513 & ~n9393 ;
  assign n9398 = n6736 ^ n5912 ^ n784 ;
  assign n9396 = ( n1306 & n2550 ) | ( n1306 & n2799 ) | ( n2550 & n2799 ) ;
  assign n9395 = n1831 ^ n1179 ^ 1'b0 ;
  assign n9397 = n9396 ^ n9395 ^ n6397 ;
  assign n9399 = n9398 ^ n9397 ^ n1438 ;
  assign n9400 = ( ~x113 & n3311 ) | ( ~x113 & n5030 ) | ( n3311 & n5030 ) ;
  assign n9401 = n538 | n9400 ;
  assign n9402 = n9401 ^ n557 ^ 1'b0 ;
  assign n9403 = ( n8924 & ~n9399 ) | ( n8924 & n9402 ) | ( ~n9399 & n9402 ) ;
  assign n9404 = n9403 ^ n6030 ^ n3650 ;
  assign n9405 = ( n289 & n1383 ) | ( n289 & ~n3812 ) | ( n1383 & ~n3812 ) ;
  assign n9406 = n9405 ^ n4623 ^ n2704 ;
  assign n9408 = ( ~n229 & n1597 ) | ( ~n229 & n2377 ) | ( n1597 & n2377 ) ;
  assign n9409 = n9408 ^ n3077 ^ 1'b0 ;
  assign n9410 = n9409 ^ n5725 ^ n796 ;
  assign n9407 = n8385 ^ n2346 ^ n603 ;
  assign n9411 = n9410 ^ n9407 ^ n2326 ;
  assign n9412 = n6677 ^ n1409 ^ 1'b0 ;
  assign n9413 = n4846 ^ n251 ^ 1'b0 ;
  assign n9414 = ( ~n3209 & n9412 ) | ( ~n3209 & n9413 ) | ( n9412 & n9413 ) ;
  assign n9415 = ( ~n5966 & n6573 ) | ( ~n5966 & n9414 ) | ( n6573 & n9414 ) ;
  assign n9417 = n4132 ^ n2719 ^ n1503 ;
  assign n9416 = ( n3505 & n5014 ) | ( n3505 & n6114 ) | ( n5014 & n6114 ) ;
  assign n9418 = n9417 ^ n9416 ^ n5665 ;
  assign n9419 = ~n9415 & n9418 ;
  assign n9420 = n9419 ^ n8818 ^ 1'b0 ;
  assign n9421 = ( n1387 & n3774 ) | ( n1387 & n6789 ) | ( n3774 & n6789 ) ;
  assign n9424 = n1744 ^ n627 ^ n459 ;
  assign n9425 = n5473 | n9424 ;
  assign n9426 = n9425 ^ n5661 ^ 1'b0 ;
  assign n9422 = ~n2836 & n9316 ;
  assign n9423 = n9422 ^ n448 ^ 1'b0 ;
  assign n9427 = n9426 ^ n9423 ^ 1'b0 ;
  assign n9428 = ~n4056 & n9427 ;
  assign n9429 = ( n3493 & n9421 ) | ( n3493 & ~n9428 ) | ( n9421 & ~n9428 ) ;
  assign n9438 = n863 & n1014 ;
  assign n9437 = n8838 ^ n3814 ^ n661 ;
  assign n9439 = n9438 ^ n9437 ^ n4329 ;
  assign n9432 = n2619 ^ n695 ^ 1'b0 ;
  assign n9433 = ~n7862 & n9432 ;
  assign n9434 = ( n2419 & n2806 ) | ( n2419 & ~n9433 ) | ( n2806 & ~n9433 ) ;
  assign n9435 = n9434 ^ n4773 ^ 1'b0 ;
  assign n9436 = ~n1575 & n9435 ;
  assign n9430 = ( ~n826 & n2344 ) | ( ~n826 & n4605 ) | ( n2344 & n4605 ) ;
  assign n9431 = ( n3012 & n8759 ) | ( n3012 & ~n9430 ) | ( n8759 & ~n9430 ) ;
  assign n9440 = n9439 ^ n9436 ^ n9431 ;
  assign n9450 = ( n2705 & n3607 ) | ( n2705 & ~n4876 ) | ( n3607 & ~n4876 ) ;
  assign n9451 = n6038 | n9450 ;
  assign n9441 = n2931 ^ n2335 ^ 1'b0 ;
  assign n9442 = n7104 | n9441 ;
  assign n9443 = n2025 | n9442 ;
  assign n9444 = n3307 ^ n1474 ^ n646 ;
  assign n9445 = n9444 ^ n3021 ^ n442 ;
  assign n9446 = n8731 | n9445 ;
  assign n9447 = n5162 & ~n9446 ;
  assign n9448 = ( n6732 & n8991 ) | ( n6732 & ~n9447 ) | ( n8991 & ~n9447 ) ;
  assign n9449 = ( ~n5924 & n9443 ) | ( ~n5924 & n9448 ) | ( n9443 & n9448 ) ;
  assign n9452 = n9451 ^ n9449 ^ n6038 ;
  assign n9453 = n7593 ^ n5488 ^ n3497 ;
  assign n9458 = n5435 ^ n1617 ^ x5 ;
  assign n9459 = n2733 & n9458 ;
  assign n9454 = ( ~n407 & n6679 ) | ( ~n407 & n7207 ) | ( n6679 & n7207 ) ;
  assign n9455 = ( n2604 & ~n4809 ) | ( n2604 & n7565 ) | ( ~n4809 & n7565 ) ;
  assign n9456 = ( n197 & ~n9454 ) | ( n197 & n9455 ) | ( ~n9454 & n9455 ) ;
  assign n9457 = n9456 ^ n4298 ^ n3252 ;
  assign n9460 = n9459 ^ n9457 ^ 1'b0 ;
  assign n9461 = n9453 | n9460 ;
  assign n9462 = ( n1114 & n7003 ) | ( n1114 & n8337 ) | ( n7003 & n8337 ) ;
  assign n9463 = n7997 ^ n5219 ^ 1'b0 ;
  assign n9464 = n9462 | n9463 ;
  assign n9465 = n3979 | n8440 ;
  assign n9466 = ( n968 & n1449 ) | ( n968 & ~n4792 ) | ( n1449 & ~n4792 ) ;
  assign n9467 = n9466 ^ n2441 ^ 1'b0 ;
  assign n9468 = n4583 | n9467 ;
  assign n9469 = n9468 ^ n6736 ^ n4292 ;
  assign n9470 = n4156 & ~n8638 ;
  assign n9471 = n7203 ^ n2530 ^ 1'b0 ;
  assign n9472 = ~n9470 & n9471 ;
  assign n9473 = n9472 ^ n7958 ^ 1'b0 ;
  assign n9474 = ( ~n7771 & n9469 ) | ( ~n7771 & n9473 ) | ( n9469 & n9473 ) ;
  assign n9475 = ( n3507 & ~n3714 ) | ( n3507 & n5993 ) | ( ~n3714 & n5993 ) ;
  assign n9476 = ( n5708 & n6299 ) | ( n5708 & n9475 ) | ( n6299 & n9475 ) ;
  assign n9477 = n9476 ^ n3599 ^ n206 ;
  assign n9478 = n6972 ^ n5431 ^ n2897 ;
  assign n9479 = n9478 ^ n7629 ^ 1'b0 ;
  assign n9480 = ~n2306 & n9479 ;
  assign n9481 = ~n3355 & n9480 ;
  assign n9482 = n6411 ^ n6363 ^ n1804 ;
  assign n9483 = n3751 & n8475 ;
  assign n9484 = n6838 & n9483 ;
  assign n9485 = ( n362 & ~n9482 ) | ( n362 & n9484 ) | ( ~n9482 & n9484 ) ;
  assign n9486 = ( n7032 & n9204 ) | ( n7032 & ~n9485 ) | ( n9204 & ~n9485 ) ;
  assign n9490 = n2956 ^ n2190 ^ 1'b0 ;
  assign n9491 = n1878 & n9490 ;
  assign n9492 = n8325 & n9491 ;
  assign n9487 = n2902 ^ n2884 ^ n434 ;
  assign n9488 = n239 | n9487 ;
  assign n9489 = n3711 | n9488 ;
  assign n9493 = n9492 ^ n9489 ^ x65 ;
  assign n9494 = n5561 ^ n1413 ^ n374 ;
  assign n9495 = n5097 ^ n3841 ^ n1127 ;
  assign n9496 = n9495 ^ n3616 ^ n2681 ;
  assign n9497 = n9496 ^ n4109 ^ 1'b0 ;
  assign n9498 = n5476 & n9497 ;
  assign n9499 = n1399 & n9498 ;
  assign n9500 = n9499 ^ n4374 ^ 1'b0 ;
  assign n9501 = n4262 ^ n2160 ^ 1'b0 ;
  assign n9502 = ( n939 & n4754 ) | ( n939 & n9501 ) | ( n4754 & n9501 ) ;
  assign n9503 = ( n1159 & n2436 ) | ( n1159 & n8991 ) | ( n2436 & n8991 ) ;
  assign n9504 = n9503 ^ n8610 ^ n5399 ;
  assign n9505 = n192 & ~n2334 ;
  assign n9506 = ~n6226 & n9505 ;
  assign n9507 = n9506 ^ n9152 ^ n231 ;
  assign n9508 = n1612 ^ n1052 ^ 1'b0 ;
  assign n9509 = n5306 & n9508 ;
  assign n9510 = n9509 ^ n8242 ^ n189 ;
  assign n9511 = ~n6884 & n9510 ;
  assign n9512 = n6230 ^ n3420 ^ 1'b0 ;
  assign n9513 = n9511 & ~n9512 ;
  assign n9514 = ~n856 & n1275 ;
  assign n9515 = n9514 ^ n9054 ^ n592 ;
  assign n9516 = ( n702 & n761 ) | ( n702 & n3189 ) | ( n761 & n3189 ) ;
  assign n9517 = n7675 | n9516 ;
  assign n9518 = n9517 ^ n1371 ^ 1'b0 ;
  assign n9519 = n191 | n9518 ;
  assign n9520 = n9519 ^ n4365 ^ 1'b0 ;
  assign n9521 = ( n1038 & ~n2476 ) | ( n1038 & n9520 ) | ( ~n2476 & n9520 ) ;
  assign n9522 = n8708 ^ n4710 ^ 1'b0 ;
  assign n9523 = ( n2876 & n8645 ) | ( n2876 & ~n9522 ) | ( n8645 & ~n9522 ) ;
  assign n9524 = ~n6231 & n6573 ;
  assign n9525 = n3803 | n5280 ;
  assign n9526 = n9525 ^ n2792 ^ 1'b0 ;
  assign n9527 = n9526 ^ n2619 ^ n629 ;
  assign n9528 = ( n9304 & ~n9524 ) | ( n9304 & n9527 ) | ( ~n9524 & n9527 ) ;
  assign n9537 = ( n339 & ~n3355 ) | ( n339 & n3700 ) | ( ~n3355 & n3700 ) ;
  assign n9535 = n5686 ^ n2475 ^ 1'b0 ;
  assign n9536 = ( n763 & ~n4461 ) | ( n763 & n9535 ) | ( ~n4461 & n9535 ) ;
  assign n9529 = n2532 ^ n1835 ^ 1'b0 ;
  assign n9530 = ~n2717 & n9529 ;
  assign n9531 = n9530 ^ n1570 ^ 1'b0 ;
  assign n9532 = ( ~n4403 & n5300 ) | ( ~n4403 & n9531 ) | ( n5300 & n9531 ) ;
  assign n9533 = ~n2854 & n9532 ;
  assign n9534 = n3952 & n9533 ;
  assign n9538 = n9537 ^ n9536 ^ n9534 ;
  assign n9539 = ( n4094 & n6550 ) | ( n4094 & ~n9538 ) | ( n6550 & ~n9538 ) ;
  assign n9540 = n3168 ^ n1713 ^ 1'b0 ;
  assign n9541 = ~n2487 & n9540 ;
  assign n9542 = n4285 ^ n3805 ^ n3597 ;
  assign n9543 = n9542 ^ n958 ^ 1'b0 ;
  assign n9544 = ~n7104 & n9543 ;
  assign n9545 = n9544 ^ n7837 ^ n7146 ;
  assign n9546 = ( n7645 & n9541 ) | ( n7645 & n9545 ) | ( n9541 & n9545 ) ;
  assign n9547 = n3754 | n4486 ;
  assign n9548 = ( x2 & ~n223 ) | ( x2 & n9547 ) | ( ~n223 & n9547 ) ;
  assign n9549 = ( n421 & n9546 ) | ( n421 & ~n9548 ) | ( n9546 & ~n9548 ) ;
  assign n9550 = ( ~n4723 & n5186 ) | ( ~n4723 & n9549 ) | ( n5186 & n9549 ) ;
  assign n9555 = ~n1656 & n3550 ;
  assign n9552 = ( x34 & ~n722 ) | ( x34 & n4346 ) | ( ~n722 & n4346 ) ;
  assign n9553 = ( ~n5361 & n5624 ) | ( ~n5361 & n9552 ) | ( n5624 & n9552 ) ;
  assign n9554 = n2739 & n9553 ;
  assign n9556 = n9555 ^ n9554 ^ 1'b0 ;
  assign n9551 = n6490 ^ n3606 ^ n539 ;
  assign n9557 = n9556 ^ n9551 ^ n7972 ;
  assign n9558 = ~n691 & n9286 ;
  assign n9559 = n9558 ^ n3084 ^ 1'b0 ;
  assign n9560 = n7855 & ~n9559 ;
  assign n9561 = n9560 ^ n9117 ^ n5072 ;
  assign n9562 = n2988 ^ n2322 ^ 1'b0 ;
  assign n9563 = n3072 | n9562 ;
  assign n9564 = ( n7951 & ~n8029 ) | ( n7951 & n9563 ) | ( ~n8029 & n9563 ) ;
  assign n9565 = n9561 | n9564 ;
  assign n9566 = ( n3190 & n5364 ) | ( n3190 & ~n9565 ) | ( n5364 & ~n9565 ) ;
  assign n9567 = n6637 ^ n1466 ^ n452 ;
  assign n9568 = ( x57 & ~n2367 ) | ( x57 & n9567 ) | ( ~n2367 & n9567 ) ;
  assign n9569 = ( ~n413 & n1457 ) | ( ~n413 & n9568 ) | ( n1457 & n9568 ) ;
  assign n9570 = ( ~n1541 & n3059 ) | ( ~n1541 & n9569 ) | ( n3059 & n9569 ) ;
  assign n9571 = n4642 ^ n2654 ^ 1'b0 ;
  assign n9572 = ~n3001 & n3832 ;
  assign n9573 = n9572 ^ n3543 ^ 1'b0 ;
  assign n9574 = ~n1563 & n3007 ;
  assign n9575 = n9574 ^ n5215 ^ 1'b0 ;
  assign n9576 = n1909 & ~n9575 ;
  assign n9577 = n1560 & n9576 ;
  assign n9578 = n9577 ^ n7465 ^ n5951 ;
  assign n9580 = n2140 ^ n1164 ^ 1'b0 ;
  assign n9581 = n2030 | n9580 ;
  assign n9579 = n6863 ^ n6546 ^ n4882 ;
  assign n9582 = n9581 ^ n9579 ^ n452 ;
  assign n9583 = n9582 ^ n8603 ^ n7156 ;
  assign n9584 = ( n4646 & ~n5185 ) | ( n4646 & n5618 ) | ( ~n5185 & n5618 ) ;
  assign n9585 = n9584 ^ n9100 ^ 1'b0 ;
  assign n9587 = n4597 ^ n2222 ^ n299 ;
  assign n9586 = n5076 & n6457 ;
  assign n9588 = n9587 ^ n9586 ^ 1'b0 ;
  assign n9589 = ( n6939 & n9585 ) | ( n6939 & n9588 ) | ( n9585 & n9588 ) ;
  assign n9590 = n978 | n1183 ;
  assign n9591 = n9590 ^ n999 ^ 1'b0 ;
  assign n9592 = n8757 & n9591 ;
  assign n9593 = ( n1400 & ~n2249 ) | ( n1400 & n6527 ) | ( ~n2249 & n6527 ) ;
  assign n9594 = n9382 ^ n903 ^ n197 ;
  assign n9595 = ( n375 & ~n5495 ) | ( n375 & n9594 ) | ( ~n5495 & n9594 ) ;
  assign n9596 = n7340 ^ n5377 ^ n5145 ;
  assign n9597 = n9596 ^ n8034 ^ n2408 ;
  assign n9598 = ( n9593 & ~n9595 ) | ( n9593 & n9597 ) | ( ~n9595 & n9597 ) ;
  assign n9599 = n2413 ^ n207 ^ x83 ;
  assign n9600 = n9599 ^ n6737 ^ 1'b0 ;
  assign n9601 = ~n1731 & n6536 ;
  assign n9602 = n4587 & n9601 ;
  assign n9603 = n9602 ^ n3455 ^ n183 ;
  assign n9604 = n653 & n9603 ;
  assign n9605 = ~n9049 & n9604 ;
  assign n9606 = n8638 ^ n6451 ^ n3701 ;
  assign n9607 = n9606 ^ n5574 ^ n509 ;
  assign n9614 = n3750 ^ n3276 ^ n732 ;
  assign n9611 = n7157 ^ n6415 ^ n3877 ;
  assign n9608 = ( x46 & ~n2118 ) | ( x46 & n3670 ) | ( ~n2118 & n3670 ) ;
  assign n9609 = n1176 & n4918 ;
  assign n9610 = n9608 & n9609 ;
  assign n9612 = n9611 ^ n9610 ^ n1703 ;
  assign n9613 = ( n5808 & ~n7698 ) | ( n5808 & n9612 ) | ( ~n7698 & n9612 ) ;
  assign n9615 = n9614 ^ n9613 ^ 1'b0 ;
  assign n9616 = n9170 ^ n1244 ^ 1'b0 ;
  assign n9617 = n8428 ^ n4946 ^ 1'b0 ;
  assign n9618 = n2609 & n9617 ;
  assign n9619 = n9398 & n9618 ;
  assign n9620 = n5592 & n9619 ;
  assign n9621 = n9620 ^ n3262 ^ x57 ;
  assign n9622 = ( n1189 & ~n4842 ) | ( n1189 & n9621 ) | ( ~n4842 & n9621 ) ;
  assign n9623 = n9622 ^ n6963 ^ n200 ;
  assign n9624 = n3485 & ~n7678 ;
  assign n9625 = n9624 ^ n7528 ^ 1'b0 ;
  assign n9626 = n6456 ^ n2471 ^ n2259 ;
  assign n9627 = ( n815 & ~n5720 ) | ( n815 & n9626 ) | ( ~n5720 & n9626 ) ;
  assign n9628 = n1042 & ~n9627 ;
  assign n9630 = n8489 ^ n5060 ^ n380 ;
  assign n9629 = n3403 ^ n3362 ^ n2129 ;
  assign n9631 = n9630 ^ n9629 ^ n9303 ;
  assign n9632 = n1642 | n5564 ;
  assign n9633 = n2296 ^ n865 ^ 1'b0 ;
  assign n9634 = n9632 & n9633 ;
  assign n9640 = ( n1239 & ~n3101 ) | ( n1239 & n5431 ) | ( ~n3101 & n5431 ) ;
  assign n9641 = n9640 ^ n3990 ^ n2968 ;
  assign n9642 = n9641 ^ n7976 ^ n2318 ;
  assign n9635 = n530 & ~n1381 ;
  assign n9636 = n9635 ^ n3193 ^ 1'b0 ;
  assign n9637 = n6449 ^ n4412 ^ n589 ;
  assign n9638 = ( ~n1308 & n9636 ) | ( ~n1308 & n9637 ) | ( n9636 & n9637 ) ;
  assign n9639 = n9638 ^ n9349 ^ n3012 ;
  assign n9643 = n9642 ^ n9639 ^ n5914 ;
  assign n9644 = n3301 ^ n947 ^ 1'b0 ;
  assign n9645 = n1479 | n9644 ;
  assign n9646 = n4013 ^ n3011 ^ n1886 ;
  assign n9647 = n9646 ^ n9276 ^ n4409 ;
  assign n9648 = ( ~n1731 & n4862 ) | ( ~n1731 & n5759 ) | ( n4862 & n5759 ) ;
  assign n9649 = n2134 ^ n2009 ^ n323 ;
  assign n9650 = ( ~n1356 & n1655 ) | ( ~n1356 & n2207 ) | ( n1655 & n2207 ) ;
  assign n9651 = ~n363 & n3025 ;
  assign n9652 = ~n3419 & n9651 ;
  assign n9653 = ( ~n7671 & n9650 ) | ( ~n7671 & n9652 ) | ( n9650 & n9652 ) ;
  assign n9654 = n9649 & ~n9653 ;
  assign n9655 = n9648 & n9654 ;
  assign n9656 = ( n593 & n7001 ) | ( n593 & n7653 ) | ( n7001 & n7653 ) ;
  assign n9657 = ( n1050 & n1721 ) | ( n1050 & n9656 ) | ( n1721 & n9656 ) ;
  assign n9658 = ( ~n892 & n1890 ) | ( ~n892 & n3569 ) | ( n1890 & n3569 ) ;
  assign n9659 = n8412 | n9658 ;
  assign n9660 = n9657 & ~n9659 ;
  assign n9661 = n9660 ^ n3344 ^ 1'b0 ;
  assign n9662 = ( n496 & n909 ) | ( n496 & n1510 ) | ( n909 & n1510 ) ;
  assign n9663 = n9662 ^ n4777 ^ n737 ;
  assign n9664 = n9663 ^ n5862 ^ n1866 ;
  assign n9670 = ( n472 & n2507 ) | ( n472 & ~n2551 ) | ( n2507 & ~n2551 ) ;
  assign n9668 = n154 | n688 ;
  assign n9669 = n9668 ^ n5590 ^ n3495 ;
  assign n9671 = n9670 ^ n9669 ^ 1'b0 ;
  assign n9666 = n6677 ^ n4549 ^ n940 ;
  assign n9667 = n9666 ^ n5694 ^ n2681 ;
  assign n9665 = ( ~n2715 & n2952 ) | ( ~n2715 & n5295 ) | ( n2952 & n5295 ) ;
  assign n9672 = n9671 ^ n9667 ^ n9665 ;
  assign n9673 = ( n4617 & n4811 ) | ( n4617 & n9672 ) | ( n4811 & n9672 ) ;
  assign n9674 = ( ~n183 & n9664 ) | ( ~n183 & n9673 ) | ( n9664 & n9673 ) ;
  assign n9680 = n2135 & n2435 ;
  assign n9681 = n2338 & n9680 ;
  assign n9677 = ( n1275 & ~n3713 ) | ( n1275 & n7569 ) | ( ~n3713 & n7569 ) ;
  assign n9678 = n9677 ^ n3416 ^ 1'b0 ;
  assign n9679 = ~n4603 & n9678 ;
  assign n9682 = n9681 ^ n9679 ^ n7101 ;
  assign n9683 = n9682 ^ n3691 ^ n2269 ;
  assign n9675 = n569 & n1833 ;
  assign n9676 = n407 & n9675 ;
  assign n9684 = n9683 ^ n9676 ^ 1'b0 ;
  assign n9685 = n3369 | n3841 ;
  assign n9686 = ( n756 & n5525 ) | ( n756 & ~n9685 ) | ( n5525 & ~n9685 ) ;
  assign n9687 = n350 & ~n9686 ;
  assign n9688 = n603 & n9687 ;
  assign n9689 = n224 | n9688 ;
  assign n9690 = ( n5302 & n8419 ) | ( n5302 & ~n8613 ) | ( n8419 & ~n8613 ) ;
  assign n9691 = n5902 ^ n5564 ^ n1733 ;
  assign n9692 = n9691 ^ n4499 ^ 1'b0 ;
  assign n9693 = ~n9441 & n9692 ;
  assign n9694 = n2602 & n4455 ;
  assign n9695 = n9694 ^ n5614 ^ 1'b0 ;
  assign n9696 = ( n445 & n3912 ) | ( n445 & n9695 ) | ( n3912 & n9695 ) ;
  assign n9697 = ~n1694 & n7806 ;
  assign n9698 = n9697 ^ n4882 ^ 1'b0 ;
  assign n9701 = n3180 | n6673 ;
  assign n9702 = n9701 ^ n6869 ^ 1'b0 ;
  assign n9703 = ~n5380 & n9702 ;
  assign n9699 = n4613 & ~n9424 ;
  assign n9700 = ~n7553 & n9699 ;
  assign n9704 = n9703 ^ n9700 ^ 1'b0 ;
  assign n9705 = n6443 ^ n1888 ^ 1'b0 ;
  assign n9706 = n2170 & n4918 ;
  assign n9707 = n9706 ^ n1135 ^ 1'b0 ;
  assign n9708 = ( n7251 & n7452 ) | ( n7251 & ~n9707 ) | ( n7452 & ~n9707 ) ;
  assign n9709 = ( ~n3833 & n8559 ) | ( ~n3833 & n9708 ) | ( n8559 & n9708 ) ;
  assign n9710 = ( n1160 & ~n9705 ) | ( n1160 & n9709 ) | ( ~n9705 & n9709 ) ;
  assign n9711 = n3397 & n9261 ;
  assign n9712 = n1289 & n9711 ;
  assign n9713 = n2754 | n9712 ;
  assign n9714 = n9713 ^ n1319 ^ 1'b0 ;
  assign n9715 = n4056 ^ n1609 ^ n1292 ;
  assign n9716 = n5024 & ~n9715 ;
  assign n9717 = n9714 & n9716 ;
  assign n9718 = n1922 & ~n3156 ;
  assign n9719 = n9718 ^ n4216 ^ 1'b0 ;
  assign n9720 = n8708 | n9719 ;
  assign n9721 = n9717 & ~n9720 ;
  assign n9724 = n7638 ^ n5562 ^ 1'b0 ;
  assign n9725 = n9724 ^ n8972 ^ n5727 ;
  assign n9722 = n5752 ^ n3959 ^ n2636 ;
  assign n9723 = n6621 | n9722 ;
  assign n9726 = n9725 ^ n9723 ^ 1'b0 ;
  assign n9727 = n5412 | n9726 ;
  assign n9728 = ( ~n3153 & n9721 ) | ( ~n3153 & n9727 ) | ( n9721 & n9727 ) ;
  assign n9732 = n8259 ^ n5170 ^ n1614 ;
  assign n9729 = n8606 ^ n7904 ^ n4423 ;
  assign n9730 = n8688 ^ n2953 ^ 1'b0 ;
  assign n9731 = n9729 & n9730 ;
  assign n9733 = n9732 ^ n9731 ^ n7255 ;
  assign n9734 = ( n3188 & n4413 ) | ( n3188 & ~n9430 ) | ( n4413 & ~n9430 ) ;
  assign n9735 = n9734 ^ n3098 ^ n960 ;
  assign n9736 = n9735 ^ n6608 ^ n6401 ;
  assign n9737 = n2102 | n9736 ;
  assign n9738 = ( ~n8067 & n8725 ) | ( ~n8067 & n9737 ) | ( n8725 & n9737 ) ;
  assign n9739 = ( n4723 & n7883 ) | ( n4723 & ~n9738 ) | ( n7883 & ~n9738 ) ;
  assign n9740 = ( n2952 & ~n9733 ) | ( n2952 & n9739 ) | ( ~n9733 & n9739 ) ;
  assign n9745 = ( n911 & n1006 ) | ( n911 & n5368 ) | ( n1006 & n5368 ) ;
  assign n9742 = ~n1606 & n6211 ;
  assign n9743 = ~n2699 & n9742 ;
  assign n9741 = ( n2724 & n5714 ) | ( n2724 & ~n6518 ) | ( n5714 & ~n6518 ) ;
  assign n9744 = n9743 ^ n9741 ^ n4685 ;
  assign n9746 = n9745 ^ n9744 ^ n998 ;
  assign n9747 = ( n1453 & ~n3262 ) | ( n1453 & n4389 ) | ( ~n3262 & n4389 ) ;
  assign n9748 = n9747 ^ n8608 ^ n406 ;
  assign n9749 = n4617 ^ n1559 ^ 1'b0 ;
  assign n9758 = x46 & ~n3396 ;
  assign n9759 = n3712 & n9758 ;
  assign n9753 = ( ~n1289 & n2845 ) | ( ~n1289 & n6526 ) | ( n2845 & n6526 ) ;
  assign n9754 = ( ~n2873 & n3660 ) | ( ~n2873 & n9487 ) | ( n3660 & n9487 ) ;
  assign n9755 = n8647 | n9754 ;
  assign n9756 = n9755 ^ n4321 ^ 1'b0 ;
  assign n9757 = ( n2427 & n9753 ) | ( n2427 & ~n9756 ) | ( n9753 & ~n9756 ) ;
  assign n9750 = n4595 ^ n2128 ^ n1316 ;
  assign n9751 = n9750 ^ n5909 ^ 1'b0 ;
  assign n9752 = n2173 & n9751 ;
  assign n9760 = n9759 ^ n9757 ^ n9752 ;
  assign n9761 = ( ~n680 & n9749 ) | ( ~n680 & n9760 ) | ( n9749 & n9760 ) ;
  assign n9762 = n474 | n1354 ;
  assign n9763 = ( n3203 & n8513 ) | ( n3203 & ~n9762 ) | ( n8513 & ~n9762 ) ;
  assign n9764 = n9645 | n9763 ;
  assign n9765 = n2586 ^ n2175 ^ 1'b0 ;
  assign n9766 = n2424 & n9765 ;
  assign n9767 = n6626 ^ n4613 ^ n1100 ;
  assign n9768 = ( n393 & ~n451 ) | ( n393 & n8417 ) | ( ~n451 & n8417 ) ;
  assign n9769 = ( n1478 & n7820 ) | ( n1478 & n9768 ) | ( n7820 & n9768 ) ;
  assign n9770 = n6536 & ~n9769 ;
  assign n9771 = n9770 ^ n5072 ^ 1'b0 ;
  assign n9772 = n398 & ~n2218 ;
  assign n9773 = n9772 ^ n2008 ^ n1554 ;
  assign n9774 = n9773 ^ n6429 ^ n2161 ;
  assign n9775 = n9774 ^ n4734 ^ n2529 ;
  assign n9776 = n3188 | n9775 ;
  assign n9777 = n9771 | n9776 ;
  assign n9778 = n9777 ^ n4324 ^ x42 ;
  assign n9779 = n9767 | n9778 ;
  assign n9780 = ( n2722 & ~n9766 ) | ( n2722 & n9779 ) | ( ~n9766 & n9779 ) ;
  assign n9781 = x114 & n3899 ;
  assign n9782 = ( x124 & n1847 ) | ( x124 & n3699 ) | ( n1847 & n3699 ) ;
  assign n9783 = ( ~n1550 & n9781 ) | ( ~n1550 & n9782 ) | ( n9781 & n9782 ) ;
  assign n9784 = ( n1853 & ~n7601 ) | ( n1853 & n9783 ) | ( ~n7601 & n9783 ) ;
  assign n9785 = n8549 ^ n2403 ^ 1'b0 ;
  assign n9786 = ~n9092 & n9785 ;
  assign n9787 = n5972 ^ n1898 ^ 1'b0 ;
  assign n9788 = n1392 & n9787 ;
  assign n9789 = ~n3149 & n9788 ;
  assign n9790 = ( n8195 & n8817 ) | ( n8195 & ~n8923 ) | ( n8817 & ~n8923 ) ;
  assign n9791 = n9790 ^ n8010 ^ n3830 ;
  assign n9793 = n3107 & n8479 ;
  assign n9794 = n9793 ^ n6889 ^ 1'b0 ;
  assign n9792 = n5299 ^ n3153 ^ n2291 ;
  assign n9795 = n9794 ^ n9792 ^ n9472 ;
  assign n9796 = n1833 & ~n3422 ;
  assign n9797 = n6204 & n9796 ;
  assign n9798 = ( n349 & n2888 ) | ( n349 & ~n9797 ) | ( n2888 & ~n9797 ) ;
  assign n9799 = n2435 ^ n1342 ^ 1'b0 ;
  assign n9800 = ( ~n2433 & n7607 ) | ( ~n2433 & n9799 ) | ( n7607 & n9799 ) ;
  assign n9801 = ( ~n3748 & n4114 ) | ( ~n3748 & n7272 ) | ( n4114 & n7272 ) ;
  assign n9802 = ( n4829 & ~n8029 ) | ( n4829 & n9801 ) | ( ~n8029 & n9801 ) ;
  assign n9803 = n2851 ^ n1108 ^ n929 ;
  assign n9804 = ( n4001 & ~n4042 ) | ( n4001 & n9803 ) | ( ~n4042 & n9803 ) ;
  assign n9805 = n9804 ^ n8927 ^ n638 ;
  assign n9807 = ( n4038 & ~n4144 ) | ( n4038 & n6052 ) | ( ~n4144 & n6052 ) ;
  assign n9806 = n724 & ~n1203 ;
  assign n9808 = n9807 ^ n9806 ^ n7999 ;
  assign n9809 = n9808 ^ n5915 ^ n1209 ;
  assign n9817 = n4900 ^ n2559 ^ n2145 ;
  assign n9816 = ( n775 & n4861 ) | ( n775 & ~n5517 ) | ( n4861 & ~n5517 ) ;
  assign n9818 = n9817 ^ n9816 ^ 1'b0 ;
  assign n9819 = n3400 | n9818 ;
  assign n9810 = n4864 ^ n3845 ^ 1'b0 ;
  assign n9811 = n8412 ^ n3652 ^ n2897 ;
  assign n9812 = ( n890 & ~n9810 ) | ( n890 & n9811 ) | ( ~n9810 & n9811 ) ;
  assign n9813 = n9812 ^ n4373 ^ n4320 ;
  assign n9814 = ( n2909 & n8606 ) | ( n2909 & n9813 ) | ( n8606 & n9813 ) ;
  assign n9815 = n9814 ^ n1381 ^ 1'b0 ;
  assign n9820 = n9819 ^ n9815 ^ n1458 ;
  assign n9821 = n6528 ^ n5582 ^ n820 ;
  assign n9822 = n9821 ^ n5517 ^ 1'b0 ;
  assign n9823 = n4387 & n4782 ;
  assign n9824 = ~n9822 & n9823 ;
  assign n9825 = n806 & ~n9824 ;
  assign n9826 = n9825 ^ n1244 ^ 1'b0 ;
  assign n9827 = ( n3881 & n5035 ) | ( n3881 & ~n9316 ) | ( n5035 & ~n9316 ) ;
  assign n9828 = n6086 ^ n2732 ^ 1'b0 ;
  assign n9829 = ( n277 & n9827 ) | ( n277 & ~n9828 ) | ( n9827 & ~n9828 ) ;
  assign n9830 = n6592 & ~n9829 ;
  assign n9831 = n5618 ^ n5586 ^ n4636 ;
  assign n9832 = n9831 ^ n6018 ^ n4225 ;
  assign n9833 = ( ~n3538 & n8051 ) | ( ~n3538 & n9832 ) | ( n8051 & n9832 ) ;
  assign n9837 = n5799 ^ x62 ^ x47 ;
  assign n9834 = n9817 ^ n2000 ^ 1'b0 ;
  assign n9835 = ( n1635 & ~n5062 ) | ( n1635 & n9834 ) | ( ~n5062 & n9834 ) ;
  assign n9836 = n9449 | n9835 ;
  assign n9838 = n9837 ^ n9836 ^ n7060 ;
  assign n9839 = ~n935 & n3593 ;
  assign n9840 = n9839 ^ n4543 ^ n975 ;
  assign n9841 = ( n676 & n3567 ) | ( n676 & n9840 ) | ( n3567 & n9840 ) ;
  assign n9842 = ( n3229 & ~n7589 ) | ( n3229 & n9841 ) | ( ~n7589 & n9841 ) ;
  assign n9843 = n841 | n4378 ;
  assign n9844 = n7655 ^ n1088 ^ 1'b0 ;
  assign n9845 = ( n955 & ~n4466 ) | ( n955 & n5704 ) | ( ~n4466 & n5704 ) ;
  assign n9846 = n9845 ^ n6498 ^ n5135 ;
  assign n9847 = ( n238 & n1794 ) | ( n238 & ~n9846 ) | ( n1794 & ~n9846 ) ;
  assign n9848 = n8570 ^ n5350 ^ 1'b0 ;
  assign n9849 = ~n9847 & n9848 ;
  assign n9850 = n3817 ^ n3121 ^ 1'b0 ;
  assign n9851 = ( n796 & n2378 ) | ( n796 & n2982 ) | ( n2378 & n2982 ) ;
  assign n9852 = n9851 ^ n1926 ^ 1'b0 ;
  assign n9853 = n9850 | n9852 ;
  assign n9856 = ( n146 & n310 ) | ( n146 & n3524 ) | ( n310 & n3524 ) ;
  assign n9854 = n3634 | n7134 ;
  assign n9855 = ( n4486 & n6265 ) | ( n4486 & n9854 ) | ( n6265 & n9854 ) ;
  assign n9857 = n9856 ^ n9855 ^ 1'b0 ;
  assign n9858 = n9398 ^ n5584 ^ 1'b0 ;
  assign n9865 = ( ~n5550 & n7326 ) | ( ~n5550 & n8238 ) | ( n7326 & n8238 ) ;
  assign n9866 = ( n284 & n8321 ) | ( n284 & ~n9865 ) | ( n8321 & ~n9865 ) ;
  assign n9859 = n4389 ^ n3415 ^ 1'b0 ;
  assign n9860 = n4020 | n9859 ;
  assign n9861 = ( ~n842 & n5757 ) | ( ~n842 & n7489 ) | ( n5757 & n7489 ) ;
  assign n9862 = ( n1487 & n9860 ) | ( n1487 & ~n9861 ) | ( n9860 & ~n9861 ) ;
  assign n9863 = n4474 ^ n4125 ^ 1'b0 ;
  assign n9864 = ( n754 & n9862 ) | ( n754 & n9863 ) | ( n9862 & n9863 ) ;
  assign n9867 = n9866 ^ n9864 ^ n1903 ;
  assign n9868 = n3367 & n3661 ;
  assign n9869 = n7528 & n9868 ;
  assign n9870 = n9869 ^ n4399 ^ 1'b0 ;
  assign n9871 = ( n4831 & n5926 ) | ( n4831 & n6411 ) | ( n5926 & n6411 ) ;
  assign n9872 = n4277 | n9871 ;
  assign n9873 = n9872 ^ n4264 ^ 1'b0 ;
  assign n9874 = n8844 ^ n7225 ^ n765 ;
  assign n9876 = ( n2569 & ~n4194 ) | ( n2569 & n8411 ) | ( ~n4194 & n8411 ) ;
  assign n9875 = ~n2034 & n6034 ;
  assign n9877 = n9876 ^ n9875 ^ 1'b0 ;
  assign n9883 = n5186 ^ n1820 ^ 1'b0 ;
  assign n9884 = n8175 & n9883 ;
  assign n9885 = ( n6277 & n9093 ) | ( n6277 & n9884 ) | ( n9093 & n9884 ) ;
  assign n9878 = n3359 & ~n8333 ;
  assign n9879 = ~n6697 & n9878 ;
  assign n9880 = n6059 | n6740 ;
  assign n9881 = n9880 ^ n8235 ^ 1'b0 ;
  assign n9882 = ( ~n1827 & n9879 ) | ( ~n1827 & n9881 ) | ( n9879 & n9881 ) ;
  assign n9886 = n9885 ^ n9882 ^ n413 ;
  assign n9887 = n9295 ^ n6661 ^ n5090 ;
  assign n9888 = n9887 ^ n1576 ^ n961 ;
  assign n9889 = ( n2297 & ~n3191 ) | ( n2297 & n8570 ) | ( ~n3191 & n8570 ) ;
  assign n9890 = n4106 & ~n9889 ;
  assign n9891 = n5301 ^ n671 ^ 1'b0 ;
  assign n9892 = n4112 & ~n8296 ;
  assign n9893 = ~n9891 & n9892 ;
  assign n9896 = ~n1797 & n3792 ;
  assign n9897 = n9896 ^ n4471 ^ 1'b0 ;
  assign n9894 = n9399 ^ n6976 ^ n4741 ;
  assign n9895 = n5276 & n9894 ;
  assign n9898 = n9897 ^ n9895 ^ 1'b0 ;
  assign n9899 = ( n4993 & n9893 ) | ( n4993 & n9898 ) | ( n9893 & n9898 ) ;
  assign n9900 = n9879 ^ n4985 ^ n2977 ;
  assign n9902 = n1838 | n7957 ;
  assign n9903 = n9902 ^ n8143 ^ 1'b0 ;
  assign n9901 = n8092 ^ n6843 ^ x41 ;
  assign n9904 = n9903 ^ n9901 ^ n7959 ;
  assign n9905 = n9400 ^ n3949 ^ n2157 ;
  assign n9906 = n9905 ^ n2393 ^ 1'b0 ;
  assign n9907 = n975 & n9906 ;
  assign n9908 = n9907 ^ n7282 ^ x19 ;
  assign n9909 = n9908 ^ n3334 ^ n2802 ;
  assign n9910 = ( n3829 & n6883 ) | ( n3829 & n9367 ) | ( n6883 & n9367 ) ;
  assign n9911 = ( n2737 & n4907 ) | ( n2737 & ~n9167 ) | ( n4907 & ~n9167 ) ;
  assign n9912 = ( n4292 & n4701 ) | ( n4292 & ~n6778 ) | ( n4701 & ~n6778 ) ;
  assign n9913 = n9912 ^ n8475 ^ 1'b0 ;
  assign n9914 = ( n375 & n9911 ) | ( n375 & n9913 ) | ( n9911 & n9913 ) ;
  assign n9922 = n4515 ^ n514 ^ x104 ;
  assign n9923 = n9922 ^ n8034 ^ n2800 ;
  assign n9918 = n360 | n5516 ;
  assign n9919 = n9918 ^ n478 ^ 1'b0 ;
  assign n9920 = ( n3740 & n8185 ) | ( n3740 & n9919 ) | ( n8185 & n9919 ) ;
  assign n9915 = n2405 | n4479 ;
  assign n9916 = n9915 ^ n5988 ^ 1'b0 ;
  assign n9917 = ( ~n1179 & n4645 ) | ( ~n1179 & n9916 ) | ( n4645 & n9916 ) ;
  assign n9921 = n9920 ^ n9917 ^ n323 ;
  assign n9924 = n9923 ^ n9921 ^ n5289 ;
  assign n9939 = n4711 & n6400 ;
  assign n9938 = ( x122 & ~n5218 ) | ( x122 & n5587 ) | ( ~n5218 & n5587 ) ;
  assign n9940 = n9939 ^ n9938 ^ 1'b0 ;
  assign n9926 = n712 & n1270 ;
  assign n9927 = n9926 ^ n5681 ^ 1'b0 ;
  assign n9928 = n9927 ^ n2012 ^ n1041 ;
  assign n9929 = ~n7451 & n9928 ;
  assign n9930 = ( ~n862 & n1792 ) | ( ~n862 & n3664 ) | ( n1792 & n3664 ) ;
  assign n9931 = ( n1371 & ~n1637 ) | ( n1371 & n9930 ) | ( ~n1637 & n9930 ) ;
  assign n9932 = n2517 ^ n1318 ^ n915 ;
  assign n9933 = ( n9774 & ~n9931 ) | ( n9774 & n9932 ) | ( ~n9931 & n9932 ) ;
  assign n9934 = n2375 ^ n2363 ^ n199 ;
  assign n9935 = n9934 ^ n6957 ^ n550 ;
  assign n9936 = ( n838 & ~n9933 ) | ( n838 & n9935 ) | ( ~n9933 & n9935 ) ;
  assign n9937 = n9929 & ~n9936 ;
  assign n9941 = n9940 ^ n9937 ^ 1'b0 ;
  assign n9942 = n9941 ^ n2857 ^ 1'b0 ;
  assign n9943 = n6641 ^ n6326 ^ 1'b0 ;
  assign n9944 = n2229 & n9943 ;
  assign n9945 = ~n7086 & n9944 ;
  assign n9946 = n9945 ^ n8630 ^ n8269 ;
  assign n9947 = ( n287 & n9942 ) | ( n287 & n9946 ) | ( n9942 & n9946 ) ;
  assign n9948 = n9947 ^ n8120 ^ n4869 ;
  assign n9925 = ~n1941 & n3011 ;
  assign n9949 = n9948 ^ n9925 ^ 1'b0 ;
  assign n9950 = ( n711 & n4739 ) | ( n711 & n5624 ) | ( n4739 & n5624 ) ;
  assign n9951 = ( ~n2305 & n3713 ) | ( ~n2305 & n7741 ) | ( n3713 & n7741 ) ;
  assign n9952 = n9951 ^ n7340 ^ n5773 ;
  assign n9953 = n6040 | n9952 ;
  assign n9954 = x119 | n3724 ;
  assign n9955 = n1210 & n6270 ;
  assign n9956 = ( n2915 & ~n9116 ) | ( n2915 & n9955 ) | ( ~n9116 & n9955 ) ;
  assign n9969 = n7692 ^ n3315 ^ n2847 ;
  assign n9964 = n1711 ^ n1552 ^ 1'b0 ;
  assign n9965 = ( n885 & n2662 ) | ( n885 & n3983 ) | ( n2662 & n3983 ) ;
  assign n9966 = ( n3263 & n5317 ) | ( n3263 & n9965 ) | ( n5317 & n9965 ) ;
  assign n9967 = ( n3116 & n9964 ) | ( n3116 & ~n9966 ) | ( n9964 & ~n9966 ) ;
  assign n9961 = ( x37 & ~n1112 ) | ( x37 & n1231 ) | ( ~n1112 & n1231 ) ;
  assign n9962 = n8239 ^ n4240 ^ 1'b0 ;
  assign n9963 = n9961 & ~n9962 ;
  assign n9968 = n9967 ^ n9963 ^ n5426 ;
  assign n9957 = ~n1448 & n2380 ;
  assign n9958 = ( n2286 & n4626 ) | ( n2286 & ~n8069 ) | ( n4626 & ~n8069 ) ;
  assign n9959 = n9958 ^ n8984 ^ n4657 ;
  assign n9960 = ( n171 & ~n9957 ) | ( n171 & n9959 ) | ( ~n9957 & n9959 ) ;
  assign n9970 = n9969 ^ n9968 ^ n9960 ;
  assign n9976 = n846 | n9053 ;
  assign n9977 = n3623 & ~n9976 ;
  assign n9971 = n1865 & n8428 ;
  assign n9972 = n3905 & n9971 ;
  assign n9973 = n9972 ^ n8881 ^ n3728 ;
  assign n9974 = ( ~n7565 & n7631 ) | ( ~n7565 & n9973 ) | ( n7631 & n9973 ) ;
  assign n9975 = ~n4248 & n9974 ;
  assign n9978 = n9977 ^ n9975 ^ n5408 ;
  assign n9979 = n2873 | n8649 ;
  assign n9980 = n9979 ^ n483 ^ 1'b0 ;
  assign n9981 = n4278 ^ n2651 ^ n1723 ;
  assign n9982 = ( n4905 & n9980 ) | ( n4905 & ~n9981 ) | ( n9980 & ~n9981 ) ;
  assign n9983 = n9982 ^ n7380 ^ 1'b0 ;
  assign n9986 = ( n1203 & ~n2066 ) | ( n1203 & n2371 ) | ( ~n2066 & n2371 ) ;
  assign n9984 = n8087 ^ n4700 ^ 1'b0 ;
  assign n9985 = n721 | n9984 ;
  assign n9987 = n9986 ^ n9985 ^ n5031 ;
  assign n9988 = n9987 ^ n4437 ^ n3634 ;
  assign n9989 = n9988 ^ n9433 ^ n4183 ;
  assign n9990 = n2489 | n9989 ;
  assign n9991 = n5183 & ~n9990 ;
  assign n9992 = n9602 ^ n2991 ^ 1'b0 ;
  assign n9993 = n343 & n9992 ;
  assign n9994 = ( n3559 & n3875 ) | ( n3559 & ~n4793 ) | ( n3875 & ~n4793 ) ;
  assign n9995 = n9994 ^ n2012 ^ n823 ;
  assign n9996 = n6779 ^ n1660 ^ 1'b0 ;
  assign n9997 = n9995 & n9996 ;
  assign n9998 = n9997 ^ n6440 ^ n1326 ;
  assign n9999 = ~n2199 & n2869 ;
  assign n10000 = n4331 ^ n1539 ^ n1227 ;
  assign n10001 = n5200 ^ n2761 ^ n1555 ;
  assign n10002 = n10001 ^ n4868 ^ n216 ;
  assign n10003 = ~n4134 & n10002 ;
  assign n10004 = ~n10000 & n10003 ;
  assign n10005 = ( n9998 & ~n9999 ) | ( n9998 & n10004 ) | ( ~n9999 & n10004 ) ;
  assign n10006 = ~n548 & n5113 ;
  assign n10007 = n6104 ^ n5448 ^ n1542 ;
  assign n10008 = n9434 ^ n4235 ^ 1'b0 ;
  assign n10009 = ( n1081 & n3619 ) | ( n1081 & n10008 ) | ( n3619 & n10008 ) ;
  assign n10010 = n10009 ^ n7932 ^ n5630 ;
  assign n10011 = n7859 ^ n5437 ^ 1'b0 ;
  assign n10012 = n4155 & n10011 ;
  assign n10013 = n10012 ^ n5176 ^ n2196 ;
  assign n10014 = ( ~n7617 & n10010 ) | ( ~n7617 & n10013 ) | ( n10010 & n10013 ) ;
  assign n10015 = n7194 ^ n6653 ^ 1'b0 ;
  assign n10016 = n10001 ^ n7222 ^ 1'b0 ;
  assign n10017 = n10016 ^ n3313 ^ n1207 ;
  assign n10018 = ( n3526 & ~n7498 ) | ( n3526 & n10017 ) | ( ~n7498 & n10017 ) ;
  assign n10019 = n7636 ^ n7625 ^ 1'b0 ;
  assign n10020 = n8449 & ~n10019 ;
  assign n10021 = x63 & ~n7936 ;
  assign n10022 = ( n1352 & ~n1678 ) | ( n1352 & n8171 ) | ( ~n1678 & n8171 ) ;
  assign n10023 = ( n1548 & n3073 ) | ( n1548 & ~n7042 ) | ( n3073 & ~n7042 ) ;
  assign n10030 = ~n2583 & n4667 ;
  assign n10031 = n7352 & ~n10030 ;
  assign n10024 = n3139 ^ n1436 ^ 1'b0 ;
  assign n10025 = n10024 ^ n7715 ^ n3046 ;
  assign n10026 = n10025 ^ x98 ^ 1'b0 ;
  assign n10027 = ~n1428 & n10026 ;
  assign n10028 = n5779 ^ n2687 ^ 1'b0 ;
  assign n10029 = ( ~n5221 & n10027 ) | ( ~n5221 & n10028 ) | ( n10027 & n10028 ) ;
  assign n10032 = n10031 ^ n10029 ^ n5912 ;
  assign n10033 = n4850 ^ n4535 ^ n1570 ;
  assign n10034 = n10033 ^ n6941 ^ n159 ;
  assign n10035 = n5712 ^ n4741 ^ n2095 ;
  assign n10036 = n10035 ^ n4494 ^ 1'b0 ;
  assign n10037 = n10036 ^ n8963 ^ n2268 ;
  assign n10038 = n6287 ^ n283 ^ 1'b0 ;
  assign n10039 = n1782 & ~n7554 ;
  assign n10040 = ( ~n841 & n2034 ) | ( ~n841 & n10039 ) | ( n2034 & n10039 ) ;
  assign n10041 = n2828 ^ n2699 ^ 1'b0 ;
  assign n10042 = ~n2249 & n10041 ;
  assign n10043 = n10040 & n10042 ;
  assign n10044 = n10043 ^ n6391 ^ n582 ;
  assign n10048 = n3516 ^ n2069 ^ n1792 ;
  assign n10047 = n1392 & ~n2208 ;
  assign n10049 = n10048 ^ n10047 ^ 1'b0 ;
  assign n10045 = n5023 & ~n5799 ;
  assign n10046 = ~n795 & n10045 ;
  assign n10050 = n10049 ^ n10046 ^ n456 ;
  assign n10051 = n5145 ^ n1328 ^ 1'b0 ;
  assign n10052 = n1991 | n10051 ;
  assign n10053 = n1580 & ~n10052 ;
  assign n10054 = n10053 ^ n9080 ^ n6808 ;
  assign n10055 = n9546 ^ n7182 ^ n3789 ;
  assign n10056 = ( n888 & ~n10054 ) | ( n888 & n10055 ) | ( ~n10054 & n10055 ) ;
  assign n10059 = n2726 ^ n1798 ^ 1'b0 ;
  assign n10057 = n3268 ^ n486 ^ 1'b0 ;
  assign n10058 = n10057 ^ n5982 ^ n4507 ;
  assign n10060 = n10059 ^ n10058 ^ n6059 ;
  assign n10061 = ( n5572 & n8288 ) | ( n5572 & n10060 ) | ( n8288 & n10060 ) ;
  assign n10062 = ( ~n3344 & n3515 ) | ( ~n3344 & n3563 ) | ( n3515 & n3563 ) ;
  assign n10063 = n4812 ^ n2341 ^ 1'b0 ;
  assign n10064 = ~n3122 & n10063 ;
  assign n10065 = n10064 ^ n5919 ^ n4013 ;
  assign n10066 = n10065 ^ n4565 ^ n4434 ;
  assign n10067 = ( ~n6593 & n10062 ) | ( ~n6593 & n10066 ) | ( n10062 & n10066 ) ;
  assign n10068 = ~n6884 & n10067 ;
  assign n10069 = n10068 ^ n5752 ^ 1'b0 ;
  assign n10070 = n7518 ^ n200 ^ 1'b0 ;
  assign n10071 = ~n747 & n4549 ;
  assign n10072 = n10071 ^ n8149 ^ n2077 ;
  assign n10073 = n7266 ^ n2098 ^ n2049 ;
  assign n10074 = n2953 ^ n2311 ^ n1469 ;
  assign n10075 = n5296 & n10074 ;
  assign n10076 = n10073 & n10075 ;
  assign n10079 = ~n2666 & n7579 ;
  assign n10077 = n9943 ^ n1893 ^ 1'b0 ;
  assign n10078 = n1740 & ~n10077 ;
  assign n10080 = n10079 ^ n10078 ^ 1'b0 ;
  assign n10081 = ( ~n934 & n2591 ) | ( ~n934 & n2741 ) | ( n2591 & n2741 ) ;
  assign n10083 = n5956 ^ n3081 ^ 1'b0 ;
  assign n10082 = ( n1062 & ~n1921 ) | ( n1062 & n3030 ) | ( ~n1921 & n3030 ) ;
  assign n10084 = n10083 ^ n10082 ^ n4999 ;
  assign n10085 = ( n1309 & n5058 ) | ( n1309 & n10084 ) | ( n5058 & n10084 ) ;
  assign n10086 = n5643 ^ n3526 ^ x66 ;
  assign n10087 = ( n10081 & ~n10085 ) | ( n10081 & n10086 ) | ( ~n10085 & n10086 ) ;
  assign n10088 = n8392 ^ n1679 ^ 1'b0 ;
  assign n10092 = n8213 ^ n423 ^ 1'b0 ;
  assign n10093 = n4162 | n10092 ;
  assign n10090 = ( n3278 & ~n3626 ) | ( n3278 & n6058 ) | ( ~n3626 & n6058 ) ;
  assign n10089 = ( n1865 & n6234 ) | ( n1865 & n8687 ) | ( n6234 & n8687 ) ;
  assign n10091 = n10090 ^ n10089 ^ n6796 ;
  assign n10094 = n10093 ^ n10091 ^ n2523 ;
  assign n10100 = n2378 ^ n1266 ^ n1263 ;
  assign n10101 = ( n2257 & n5468 ) | ( n2257 & n10100 ) | ( n5468 & n10100 ) ;
  assign n10098 = ~n5526 & n7295 ;
  assign n10099 = n10098 ^ n4087 ^ 1'b0 ;
  assign n10096 = ( ~n736 & n3238 ) | ( ~n736 & n4407 ) | ( n3238 & n4407 ) ;
  assign n10097 = n10096 ^ n4584 ^ n3965 ;
  assign n10102 = n10101 ^ n10099 ^ n10097 ;
  assign n10095 = n673 & ~n7746 ;
  assign n10103 = n10102 ^ n10095 ^ 1'b0 ;
  assign n10106 = n8067 ^ n6778 ^ n2852 ;
  assign n10104 = n9855 ^ n5664 ^ n1113 ;
  assign n10105 = ( ~n3216 & n4890 ) | ( ~n3216 & n10104 ) | ( n4890 & n10104 ) ;
  assign n10107 = n10106 ^ n10105 ^ 1'b0 ;
  assign n10108 = n2727 ^ n2487 ^ n2352 ;
  assign n10109 = n10108 ^ n6915 ^ n1911 ;
  assign n10110 = ~n5945 & n10109 ;
  assign n10112 = n9243 ^ n7264 ^ 1'b0 ;
  assign n10111 = n1627 | n6234 ;
  assign n10113 = n10112 ^ n10111 ^ 1'b0 ;
  assign n10129 = ~n3177 & n8430 ;
  assign n10130 = n8422 & n10129 ;
  assign n10126 = ( n1513 & n2766 ) | ( n1513 & ~n7002 ) | ( n2766 & ~n7002 ) ;
  assign n10127 = n4852 & n5873 ;
  assign n10128 = ( ~n4193 & n10126 ) | ( ~n4193 & n10127 ) | ( n10126 & n10127 ) ;
  assign n10131 = n10130 ^ n10128 ^ n5061 ;
  assign n10114 = n4880 ^ n4001 ^ n798 ;
  assign n10115 = n10114 ^ n2619 ^ n1501 ;
  assign n10116 = x13 & ~n3993 ;
  assign n10117 = n4851 & n10116 ;
  assign n10118 = n4985 & n10117 ;
  assign n10119 = n1116 & n10118 ;
  assign n10120 = n10119 ^ n8449 ^ n4885 ;
  assign n10121 = ( n2279 & n6358 ) | ( n2279 & n10120 ) | ( n6358 & n10120 ) ;
  assign n10122 = ( ~n2129 & n10115 ) | ( ~n2129 & n10121 ) | ( n10115 & n10121 ) ;
  assign n10123 = n4425 & ~n6294 ;
  assign n10124 = n10123 ^ n7377 ^ 1'b0 ;
  assign n10125 = ( ~n2249 & n10122 ) | ( ~n2249 & n10124 ) | ( n10122 & n10124 ) ;
  assign n10132 = n10131 ^ n10125 ^ n1941 ;
  assign n10133 = ( ~n2353 & n6114 ) | ( ~n2353 & n6712 ) | ( n6114 & n6712 ) ;
  assign n10134 = n10133 ^ n3686 ^ n2691 ;
  assign n10135 = n10134 ^ n3806 ^ n397 ;
  assign n10136 = n9020 ^ n3129 ^ 1'b0 ;
  assign n10137 = ( ~x56 & n168 ) | ( ~x56 & n10136 ) | ( n168 & n10136 ) ;
  assign n10138 = n10137 ^ n7812 ^ 1'b0 ;
  assign n10139 = n195 | n10138 ;
  assign n10140 = ( ~n2076 & n4196 ) | ( ~n2076 & n9662 ) | ( n4196 & n9662 ) ;
  assign n10141 = n3975 & n10140 ;
  assign n10142 = ~n3177 & n7788 ;
  assign n10143 = ( n3001 & n7023 ) | ( n3001 & ~n10142 ) | ( n7023 & ~n10142 ) ;
  assign n10144 = ~n6373 & n10143 ;
  assign n10153 = n8357 ^ n4729 ^ 1'b0 ;
  assign n10154 = n6249 & n10153 ;
  assign n10155 = n10154 ^ n7219 ^ n439 ;
  assign n10145 = n8469 ^ n4666 ^ n3082 ;
  assign n10146 = n6489 & n10145 ;
  assign n10147 = n1167 & n2229 ;
  assign n10148 = n10147 ^ n1918 ^ 1'b0 ;
  assign n10149 = ( ~n2599 & n6261 ) | ( ~n2599 & n10148 ) | ( n6261 & n10148 ) ;
  assign n10150 = n2193 & n10149 ;
  assign n10151 = n10150 ^ n6865 ^ n5276 ;
  assign n10152 = n10146 | n10151 ;
  assign n10156 = n10155 ^ n10152 ^ 1'b0 ;
  assign n10157 = n879 & ~n2383 ;
  assign n10158 = ( ~n2562 & n6030 ) | ( ~n2562 & n7207 ) | ( n6030 & n7207 ) ;
  assign n10159 = ~n2157 & n5482 ;
  assign n10160 = n10159 ^ n1351 ^ 1'b0 ;
  assign n10161 = n10158 | n10160 ;
  assign n10162 = ( n4806 & n10157 ) | ( n4806 & ~n10161 ) | ( n10157 & ~n10161 ) ;
  assign n10163 = n10162 ^ n5047 ^ n205 ;
  assign n10164 = n4553 | n6032 ;
  assign n10165 = n4303 ^ n3372 ^ 1'b0 ;
  assign n10166 = n2548 & ~n10165 ;
  assign n10167 = n10166 ^ n4480 ^ n3103 ;
  assign n10168 = ( x68 & n10164 ) | ( x68 & ~n10167 ) | ( n10164 & ~n10167 ) ;
  assign n10169 = n659 & n2127 ;
  assign n10170 = n8080 ^ n7041 ^ n5299 ;
  assign n10171 = ( n4979 & ~n5318 ) | ( n4979 & n10170 ) | ( ~n5318 & n10170 ) ;
  assign n10172 = n10171 ^ n8716 ^ 1'b0 ;
  assign n10173 = ~n3530 & n10172 ;
  assign n10174 = n7281 & n10173 ;
  assign n10175 = ( n822 & ~n7639 ) | ( n822 & n8545 ) | ( ~n7639 & n8545 ) ;
  assign n10176 = n277 & n8307 ;
  assign n10177 = n10176 ^ n4156 ^ 1'b0 ;
  assign n10178 = ~n4601 & n4801 ;
  assign n10179 = n10178 ^ n1588 ^ 1'b0 ;
  assign n10180 = ( n1530 & ~n10177 ) | ( n1530 & n10179 ) | ( ~n10177 & n10179 ) ;
  assign n10181 = n9005 ^ n3221 ^ n2702 ;
  assign n10182 = n10181 ^ n2629 ^ n901 ;
  assign n10183 = n5020 | n10182 ;
  assign n10184 = n8349 & ~n10183 ;
  assign n10190 = n8039 ^ n3281 ^ n817 ;
  assign n10189 = ( n1360 & n2260 ) | ( n1360 & n8709 ) | ( n2260 & n8709 ) ;
  assign n10185 = n3971 | n5548 ;
  assign n10186 = ~n5600 & n10185 ;
  assign n10187 = n2991 & n10186 ;
  assign n10188 = n10187 ^ n9413 ^ n1656 ;
  assign n10191 = n10190 ^ n10189 ^ n10188 ;
  assign n10192 = ( n1285 & n7034 ) | ( n1285 & n10191 ) | ( n7034 & n10191 ) ;
  assign n10193 = ( ~n6887 & n9168 ) | ( ~n6887 & n10192 ) | ( n9168 & n10192 ) ;
  assign n10194 = ( ~n5153 & n7516 ) | ( ~n5153 & n9042 ) | ( n7516 & n9042 ) ;
  assign n10195 = n6414 ^ n1312 ^ 1'b0 ;
  assign n10196 = n10195 ^ n6117 ^ n4931 ;
  assign n10197 = n9277 ^ n8236 ^ n2077 ;
  assign n10198 = ( n8172 & ~n8417 ) | ( n8172 & n10197 ) | ( ~n8417 & n10197 ) ;
  assign n10199 = ( n590 & n6350 ) | ( n590 & n10198 ) | ( n6350 & n10198 ) ;
  assign n10200 = n10199 ^ n5415 ^ n4547 ;
  assign n10201 = n5619 ^ n1203 ^ n162 ;
  assign n10202 = n10201 ^ n3478 ^ n3432 ;
  assign n10203 = n10202 ^ n5616 ^ n3016 ;
  assign n10204 = n1296 & n3256 ;
  assign n10205 = n10204 ^ n5013 ^ 1'b0 ;
  assign n10206 = ~n4568 & n10205 ;
  assign n10207 = ~n5425 & n10206 ;
  assign n10208 = n936 & ~n7147 ;
  assign n10209 = n10207 & n10208 ;
  assign n10210 = n5313 ^ n4918 ^ n1551 ;
  assign n10211 = n232 | n10210 ;
  assign n10212 = n10209 & ~n10211 ;
  assign n10213 = n6670 ^ n1277 ^ n956 ;
  assign n10214 = n10213 ^ n10080 ^ n3226 ;
  assign n10215 = ( n908 & ~n2855 ) | ( n908 & n3087 ) | ( ~n2855 & n3087 ) ;
  assign n10216 = ( n424 & ~n1863 ) | ( n424 & n8725 ) | ( ~n1863 & n8725 ) ;
  assign n10217 = ( ~n4389 & n5670 ) | ( ~n4389 & n9542 ) | ( n5670 & n9542 ) ;
  assign n10218 = ( n635 & n1295 ) | ( n635 & n10217 ) | ( n1295 & n10217 ) ;
  assign n10219 = n10216 | n10218 ;
  assign n10220 = n10219 ^ n6220 ^ 1'b0 ;
  assign n10221 = ( ~n9630 & n10215 ) | ( ~n9630 & n10220 ) | ( n10215 & n10220 ) ;
  assign n10222 = ( ~n302 & n2193 ) | ( ~n302 & n10221 ) | ( n2193 & n10221 ) ;
  assign n10223 = ( ~n187 & n1741 ) | ( ~n187 & n2759 ) | ( n1741 & n2759 ) ;
  assign n10224 = n4128 & ~n4891 ;
  assign n10225 = ~n547 & n10224 ;
  assign n10226 = n10223 & ~n10225 ;
  assign n10227 = n2232 & n8873 ;
  assign n10228 = n10226 & n10227 ;
  assign n10234 = ( n1072 & ~n2032 ) | ( n1072 & n2914 ) | ( ~n2032 & n2914 ) ;
  assign n10235 = n10234 ^ n6730 ^ n6422 ;
  assign n10229 = n6297 ^ n3470 ^ x88 ;
  assign n10230 = ~n3451 & n5512 ;
  assign n10231 = n10230 ^ n4961 ^ 1'b0 ;
  assign n10232 = n10231 ^ n174 ^ 1'b0 ;
  assign n10233 = ~n10229 & n10232 ;
  assign n10236 = n10235 ^ n10233 ^ n6318 ;
  assign n10237 = ( x114 & n396 ) | ( x114 & n4362 ) | ( n396 & n4362 ) ;
  assign n10238 = ( ~n362 & n6944 ) | ( ~n362 & n9569 ) | ( n6944 & n9569 ) ;
  assign n10240 = n9804 ^ n6592 ^ 1'b0 ;
  assign n10241 = n3532 & ~n10240 ;
  assign n10242 = n10241 ^ n5058 ^ n858 ;
  assign n10239 = n5365 ^ n2643 ^ n2224 ;
  assign n10243 = n10242 ^ n10239 ^ n3054 ;
  assign n10244 = ( n10237 & n10238 ) | ( n10237 & ~n10243 ) | ( n10238 & ~n10243 ) ;
  assign n10245 = n3974 & ~n10187 ;
  assign n10246 = n10245 ^ n5644 ^ 1'b0 ;
  assign n10247 = n9936 ^ n5065 ^ n3301 ;
  assign n10251 = ( ~n1717 & n3862 ) | ( ~n1717 & n9974 ) | ( n3862 & n9974 ) ;
  assign n10252 = n10251 ^ n7272 ^ n3880 ;
  assign n10248 = n3907 & ~n9344 ;
  assign n10249 = ~n7511 & n10248 ;
  assign n10250 = ( x47 & n7445 ) | ( x47 & n10249 ) | ( n7445 & n10249 ) ;
  assign n10253 = n10252 ^ n10250 ^ n7930 ;
  assign n10254 = n10253 ^ n6891 ^ 1'b0 ;
  assign n10255 = n10247 & n10254 ;
  assign n10256 = n8087 ^ n3103 ^ n2358 ;
  assign n10257 = ( n3262 & ~n8986 ) | ( n3262 & n10256 ) | ( ~n8986 & n10256 ) ;
  assign n10258 = ( n4247 & ~n7148 ) | ( n4247 & n9178 ) | ( ~n7148 & n9178 ) ;
  assign n10263 = n1205 & n4896 ;
  assign n10264 = n10263 ^ n9050 ^ 1'b0 ;
  assign n10265 = ( ~n7006 & n7644 ) | ( ~n7006 & n10264 ) | ( n7644 & n10264 ) ;
  assign n10266 = ( n5756 & n9773 ) | ( n5756 & ~n10265 ) | ( n9773 & ~n10265 ) ;
  assign n10260 = ( n1745 & n3589 ) | ( n1745 & ~n3860 ) | ( n3589 & ~n3860 ) ;
  assign n10259 = n550 | n6713 ;
  assign n10261 = n10260 ^ n10259 ^ 1'b0 ;
  assign n10262 = ( n2443 & ~n3981 ) | ( n2443 & n10261 ) | ( ~n3981 & n10261 ) ;
  assign n10267 = n10266 ^ n10262 ^ n7549 ;
  assign n10269 = n5087 ^ n2095 ^ n777 ;
  assign n10268 = n8328 ^ n6341 ^ n1320 ;
  assign n10270 = n10269 ^ n10268 ^ n4533 ;
  assign n10271 = n10270 ^ n9936 ^ 1'b0 ;
  assign n10274 = ( n3518 & n4350 ) | ( n3518 & ~n4405 ) | ( n4350 & ~n4405 ) ;
  assign n10272 = n253 & ~n7516 ;
  assign n10273 = n2841 & n10272 ;
  assign n10275 = n10274 ^ n10273 ^ n392 ;
  assign n10276 = n9281 ^ n5366 ^ 1'b0 ;
  assign n10277 = n8711 & n10276 ;
  assign n10278 = n2783 ^ n1329 ^ 1'b0 ;
  assign n10279 = ~n152 & n10278 ;
  assign n10280 = ( n2615 & ~n2909 ) | ( n2615 & n10279 ) | ( ~n2909 & n10279 ) ;
  assign n10281 = ( n4691 & n5875 ) | ( n4691 & n10280 ) | ( n5875 & n10280 ) ;
  assign n10282 = n9568 ^ n5410 ^ n220 ;
  assign n10283 = ( n2027 & n7609 ) | ( n2027 & ~n10282 ) | ( n7609 & ~n10282 ) ;
  assign n10284 = n9144 | n10283 ;
  assign n10285 = n10284 ^ n9649 ^ 1'b0 ;
  assign n10286 = n8009 & ~n8790 ;
  assign n10288 = n1453 & n1982 ;
  assign n10289 = n10288 ^ n4104 ^ 1'b0 ;
  assign n10291 = n6653 ^ n1528 ^ 1'b0 ;
  assign n10292 = ( ~n1378 & n9685 ) | ( ~n1378 & n10291 ) | ( n9685 & n10291 ) ;
  assign n10290 = n3727 | n9871 ;
  assign n10293 = n10292 ^ n10290 ^ 1'b0 ;
  assign n10294 = ( ~n3316 & n10289 ) | ( ~n3316 & n10293 ) | ( n10289 & n10293 ) ;
  assign n10295 = n10294 ^ n582 ^ n480 ;
  assign n10296 = ~n4811 & n10295 ;
  assign n10287 = n9034 ^ n7985 ^ 1'b0 ;
  assign n10297 = n10296 ^ n10287 ^ n5386 ;
  assign n10298 = n2566 | n5953 ;
  assign n10299 = n1249 | n10298 ;
  assign n10300 = n10299 ^ n2160 ^ 1'b0 ;
  assign n10301 = n4623 & n10300 ;
  assign n10302 = n10301 ^ n8666 ^ n428 ;
  assign n10303 = n6920 & ~n9509 ;
  assign n10304 = n10303 ^ n3053 ^ n1169 ;
  assign n10305 = n6645 ^ n6132 ^ 1'b0 ;
  assign n10306 = n10305 ^ n6226 ^ n545 ;
  assign n10307 = ( n873 & n1603 ) | ( n873 & n6576 ) | ( n1603 & n6576 ) ;
  assign n10308 = n10307 ^ n2311 ^ 1'b0 ;
  assign n10309 = ( n693 & n4372 ) | ( n693 & n7923 ) | ( n4372 & n7923 ) ;
  assign n10310 = n10309 ^ n4372 ^ n1437 ;
  assign n10311 = ~n985 & n3152 ;
  assign n10312 = n10311 ^ n2862 ^ 1'b0 ;
  assign n10313 = n570 & ~n4714 ;
  assign n10314 = ~n10312 & n10313 ;
  assign n10315 = n3759 | n10314 ;
  assign n10316 = ( n1700 & n4370 ) | ( n1700 & n7271 ) | ( n4370 & n7271 ) ;
  assign n10317 = n10315 | n10316 ;
  assign n10318 = n10317 ^ x103 ^ 1'b0 ;
  assign n10319 = ( n769 & n771 ) | ( n769 & n3976 ) | ( n771 & n3976 ) ;
  assign n10320 = ( n4013 & n7617 ) | ( n4013 & ~n10319 ) | ( n7617 & ~n10319 ) ;
  assign n10321 = ( n4798 & n10318 ) | ( n4798 & ~n10320 ) | ( n10318 & ~n10320 ) ;
  assign n10322 = n3777 ^ n2940 ^ 1'b0 ;
  assign n10323 = n10322 ^ n4760 ^ n2023 ;
  assign n10324 = n1930 | n8119 ;
  assign n10325 = ( n5625 & n6022 ) | ( n5625 & ~n10324 ) | ( n6022 & ~n10324 ) ;
  assign n10330 = n6658 & n9466 ;
  assign n10331 = ( n5859 & n10319 ) | ( n5859 & n10330 ) | ( n10319 & n10330 ) ;
  assign n10332 = n1134 ^ n472 ^ 1'b0 ;
  assign n10333 = n10332 ^ n7839 ^ x44 ;
  assign n10334 = ( n1848 & n10331 ) | ( n1848 & ~n10333 ) | ( n10331 & ~n10333 ) ;
  assign n10328 = n1601 ^ x75 ^ x59 ;
  assign n10329 = n10328 ^ n5573 ^ n391 ;
  assign n10326 = n3635 ^ n3273 ^ 1'b0 ;
  assign n10327 = ~n4494 & n10326 ;
  assign n10335 = n10334 ^ n10329 ^ n10327 ;
  assign n10336 = ( n1032 & n3492 ) | ( n1032 & ~n10335 ) | ( n3492 & ~n10335 ) ;
  assign n10337 = n2601 ^ n329 ^ x84 ;
  assign n10338 = ~n4575 & n10337 ;
  assign n10339 = n10338 ^ n5718 ^ 1'b0 ;
  assign n10340 = n2326 ^ n1303 ^ 1'b0 ;
  assign n10341 = n10339 & ~n10340 ;
  assign n10342 = ( ~n1091 & n1225 ) | ( ~n1091 & n5429 ) | ( n1225 & n5429 ) ;
  assign n10343 = ( n5423 & n5498 ) | ( n5423 & n10342 ) | ( n5498 & n10342 ) ;
  assign n10344 = ( n1756 & ~n2411 ) | ( n1756 & n10343 ) | ( ~n2411 & n10343 ) ;
  assign n10345 = ( n5154 & ~n7958 ) | ( n5154 & n10344 ) | ( ~n7958 & n10344 ) ;
  assign n10346 = ( n8164 & n8956 ) | ( n8164 & ~n9054 ) | ( n8956 & ~n9054 ) ;
  assign n10347 = n10346 ^ n2326 ^ 1'b0 ;
  assign n10348 = ( n2146 & n4855 ) | ( n2146 & n10347 ) | ( n4855 & n10347 ) ;
  assign n10349 = n10348 ^ n6508 ^ n5865 ;
  assign n10350 = ~n778 & n4365 ;
  assign n10351 = n10350 ^ n8866 ^ n2613 ;
  assign n10352 = ( ~n3263 & n9812 ) | ( ~n3263 & n10351 ) | ( n9812 & n10351 ) ;
  assign n10353 = ( n1108 & n2856 ) | ( n1108 & n10352 ) | ( n2856 & n10352 ) ;
  assign n10354 = x68 & ~n775 ;
  assign n10355 = ~n3707 & n10354 ;
  assign n10356 = ( ~n643 & n2750 ) | ( ~n643 & n10355 ) | ( n2750 & n10355 ) ;
  assign n10357 = n10104 ^ n6099 ^ n424 ;
  assign n10358 = ( n317 & n4268 ) | ( n317 & n5274 ) | ( n4268 & n5274 ) ;
  assign n10359 = n10358 ^ n5407 ^ x81 ;
  assign n10360 = n10359 ^ n2964 ^ n2112 ;
  assign n10361 = n10189 ^ n2348 ^ 1'b0 ;
  assign n10362 = n7041 | n10361 ;
  assign n10363 = ( n958 & ~n2547 ) | ( n958 & n10362 ) | ( ~n2547 & n10362 ) ;
  assign n10364 = n8333 | n10363 ;
  assign n10365 = ( ~n1220 & n2512 ) | ( ~n1220 & n5903 ) | ( n2512 & n5903 ) ;
  assign n10366 = n10365 ^ n2731 ^ 1'b0 ;
  assign n10367 = ~n823 & n10366 ;
  assign n10368 = ( ~n1699 & n3133 ) | ( ~n1699 & n4965 ) | ( n3133 & n4965 ) ;
  assign n10369 = n10368 ^ n7874 ^ n605 ;
  assign n10371 = ~n258 & n3210 ;
  assign n10370 = n2449 & n7295 ;
  assign n10372 = n10371 ^ n10370 ^ 1'b0 ;
  assign n10382 = ( n1112 & n2012 ) | ( n1112 & ~n3897 ) | ( n2012 & ~n3897 ) ;
  assign n10383 = n10382 ^ n1393 ^ n234 ;
  assign n10379 = n3260 ^ n693 ^ 1'b0 ;
  assign n10380 = n10379 ^ n9468 ^ 1'b0 ;
  assign n10375 = n723 | n3220 ;
  assign n10376 = n10375 ^ n887 ^ 1'b0 ;
  assign n10377 = n10376 ^ n3492 ^ 1'b0 ;
  assign n10373 = n5925 ^ n4502 ^ 1'b0 ;
  assign n10374 = n3444 | n10373 ;
  assign n10378 = n10377 ^ n10374 ^ 1'b0 ;
  assign n10381 = n10380 ^ n10378 ^ n130 ;
  assign n10384 = n10383 ^ n10381 ^ n10109 ;
  assign n10386 = ( n911 & ~n2495 ) | ( n911 & n9285 ) | ( ~n2495 & n9285 ) ;
  assign n10385 = n4362 ^ n2312 ^ n1636 ;
  assign n10387 = n10386 ^ n10385 ^ n5147 ;
  assign n10388 = n9884 ^ n7352 ^ n5650 ;
  assign n10389 = n10388 ^ n2049 ^ 1'b0 ;
  assign n10390 = ( n6146 & n9450 ) | ( n6146 & n9734 ) | ( n9450 & n9734 ) ;
  assign n10391 = x7 & ~n10390 ;
  assign n10392 = ~n3741 & n10391 ;
  assign n10401 = n1165 ^ n1161 ^ n546 ;
  assign n10398 = ( n3380 & ~n4565 ) | ( n3380 & n8847 ) | ( ~n4565 & n8847 ) ;
  assign n10393 = ~n2200 & n8006 ;
  assign n10394 = ~n4668 & n10393 ;
  assign n10395 = n8976 & ~n10394 ;
  assign n10396 = n549 & n10395 ;
  assign n10397 = ( n3601 & ~n5468 ) | ( n3601 & n10396 ) | ( ~n5468 & n10396 ) ;
  assign n10399 = n10398 ^ n10397 ^ n10131 ;
  assign n10400 = ~n7818 & n10399 ;
  assign n10402 = n10401 ^ n10400 ^ 1'b0 ;
  assign n10403 = ( n10389 & n10392 ) | ( n10389 & ~n10402 ) | ( n10392 & ~n10402 ) ;
  assign n10404 = ( ~n864 & n2528 ) | ( ~n864 & n3562 ) | ( n2528 & n3562 ) ;
  assign n10405 = n10404 ^ n8932 ^ n7493 ;
  assign n10406 = n6667 ^ n2118 ^ n2115 ;
  assign n10407 = ~n8552 & n10406 ;
  assign n10408 = ~n9613 & n10407 ;
  assign n10409 = n7139 ^ n4946 ^ n2910 ;
  assign n10410 = n4107 & ~n4493 ;
  assign n10411 = ~n2039 & n10410 ;
  assign n10412 = n10409 & n10411 ;
  assign n10413 = n10412 ^ n10384 ^ n10320 ;
  assign n10414 = n4871 ^ n4345 ^ 1'b0 ;
  assign n10415 = n4630 & ~n10414 ;
  assign n10416 = n5795 ^ n4085 ^ 1'b0 ;
  assign n10417 = n4045 ^ n2432 ^ n367 ;
  assign n10418 = n10417 ^ n2235 ^ 1'b0 ;
  assign n10419 = n10416 | n10418 ;
  assign n10420 = ( n1766 & n3798 ) | ( n1766 & n4497 ) | ( n3798 & n4497 ) ;
  assign n10421 = ( n1987 & n5359 ) | ( n1987 & ~n5429 ) | ( n5359 & ~n5429 ) ;
  assign n10422 = ( ~n1360 & n10420 ) | ( ~n1360 & n10421 ) | ( n10420 & n10421 ) ;
  assign n10423 = n10422 ^ n1582 ^ 1'b0 ;
  assign n10424 = ~n10419 & n10423 ;
  assign n10425 = ( n6219 & n10415 ) | ( n6219 & ~n10424 ) | ( n10415 & ~n10424 ) ;
  assign n10426 = ( n200 & n693 ) | ( n200 & ~n1515 ) | ( n693 & ~n1515 ) ;
  assign n10427 = ( n3613 & n5554 ) | ( n3613 & ~n10426 ) | ( n5554 & ~n10426 ) ;
  assign n10428 = n10427 ^ n7566 ^ 1'b0 ;
  assign n10429 = n4078 | n10428 ;
  assign n10430 = n9888 & ~n10429 ;
  assign n10431 = n10430 ^ n9216 ^ 1'b0 ;
  assign n10432 = n1928 ^ n1457 ^ n844 ;
  assign n10433 = ~n3129 & n10432 ;
  assign n10434 = ~n538 & n5049 ;
  assign n10435 = n3933 & n10434 ;
  assign n10436 = n3502 | n10435 ;
  assign n10438 = ( n4376 & n4920 ) | ( n4376 & ~n6275 ) | ( n4920 & ~n6275 ) ;
  assign n10439 = ( n6511 & n9011 ) | ( n6511 & ~n10438 ) | ( n9011 & ~n10438 ) ;
  assign n10437 = n7063 & n8950 ;
  assign n10440 = n10439 ^ n10437 ^ 1'b0 ;
  assign n10444 = n6611 ^ n2982 ^ 1'b0 ;
  assign n10441 = x5 | n3200 ;
  assign n10442 = n10441 ^ n3592 ^ n575 ;
  assign n10443 = n7736 & n10442 ;
  assign n10445 = n10444 ^ n10443 ^ 1'b0 ;
  assign n10446 = ( n4507 & n5326 ) | ( n4507 & n6701 ) | ( n5326 & n6701 ) ;
  assign n10447 = n10446 ^ n7379 ^ n2970 ;
  assign n10448 = n2789 ^ n2004 ^ 1'b0 ;
  assign n10449 = x65 & ~n5440 ;
  assign n10450 = n10449 ^ n4917 ^ n291 ;
  assign n10451 = n924 | n9231 ;
  assign n10452 = n10451 ^ n141 ^ 1'b0 ;
  assign n10453 = n1910 ^ n1723 ^ 1'b0 ;
  assign n10454 = n10452 & ~n10453 ;
  assign n10455 = ( n5187 & n10100 ) | ( n5187 & n10454 ) | ( n10100 & n10454 ) ;
  assign n10456 = n2377 ^ n1874 ^ n1825 ;
  assign n10457 = n10456 ^ n8827 ^ n2375 ;
  assign n10458 = n3815 ^ n1492 ^ n532 ;
  assign n10459 = n1095 & n10458 ;
  assign n10460 = n7848 & ~n10459 ;
  assign n10461 = n8924 ^ n6976 ^ n4821 ;
  assign n10462 = n8588 ^ n6823 ^ n6156 ;
  assign n10466 = ( n6337 & n6716 ) | ( n6337 & n8047 ) | ( n6716 & n8047 ) ;
  assign n10464 = n2262 ^ n520 ^ 1'b0 ;
  assign n10463 = ( n831 & n1416 ) | ( n831 & ~n1922 ) | ( n1416 & ~n1922 ) ;
  assign n10465 = n10464 ^ n10463 ^ n712 ;
  assign n10467 = n10466 ^ n10465 ^ n8737 ;
  assign n10468 = n10462 & ~n10467 ;
  assign n10469 = n10468 ^ n5928 ^ 1'b0 ;
  assign n10470 = ( ~n1892 & n5184 ) | ( ~n1892 & n5341 ) | ( n5184 & n5341 ) ;
  assign n10471 = n5715 ^ n5282 ^ 1'b0 ;
  assign n10472 = n411 | n10471 ;
  assign n10473 = n8866 | n10472 ;
  assign n10474 = n10473 ^ n8713 ^ 1'b0 ;
  assign n10476 = n1006 & ~n4552 ;
  assign n10477 = n10476 ^ n3997 ^ n1718 ;
  assign n10475 = n2207 & n4651 ;
  assign n10478 = n10477 ^ n10475 ^ n1480 ;
  assign n10479 = ( n882 & ~n2147 ) | ( n882 & n8054 ) | ( ~n2147 & n8054 ) ;
  assign n10480 = n10479 ^ n171 ^ 1'b0 ;
  assign n10481 = n9433 ^ n8054 ^ n2876 ;
  assign n10482 = n10481 ^ n4417 ^ 1'b0 ;
  assign n10483 = n7564 & n10482 ;
  assign n10484 = n8560 ^ n2445 ^ 1'b0 ;
  assign n10485 = n7222 | n10484 ;
  assign n10486 = n9281 ^ n6571 ^ 1'b0 ;
  assign n10487 = ( ~n10483 & n10485 ) | ( ~n10483 & n10486 ) | ( n10485 & n10486 ) ;
  assign n10495 = ~n1145 & n1959 ;
  assign n10496 = n3605 & n10495 ;
  assign n10488 = ~n3815 & n7433 ;
  assign n10489 = ( n6749 & ~n9641 ) | ( n6749 & n10488 ) | ( ~n9641 & n10488 ) ;
  assign n10490 = ( ~x47 & n3345 ) | ( ~x47 & n10489 ) | ( n3345 & n10489 ) ;
  assign n10491 = n10490 ^ n4271 ^ n413 ;
  assign n10492 = n5894 ^ n4233 ^ 1'b0 ;
  assign n10493 = n10491 & ~n10492 ;
  assign n10494 = n3151 & n10493 ;
  assign n10497 = n10496 ^ n10494 ^ n1667 ;
  assign n10498 = ( n2534 & n3714 ) | ( n2534 & n7191 ) | ( n3714 & n7191 ) ;
  assign n10499 = n10498 ^ n7490 ^ n436 ;
  assign n10500 = n10499 ^ n3959 ^ 1'b0 ;
  assign n10501 = ( ~n2540 & n7063 ) | ( ~n2540 & n9269 ) | ( n7063 & n9269 ) ;
  assign n10506 = n3353 | n4952 ;
  assign n10507 = n166 & ~n10506 ;
  assign n10508 = ( n2929 & n6331 ) | ( n2929 & ~n10507 ) | ( n6331 & ~n10507 ) ;
  assign n10502 = n9994 ^ n1958 ^ n1645 ;
  assign n10503 = n7111 ^ n7049 ^ n724 ;
  assign n10504 = n10503 ^ n9223 ^ n4613 ;
  assign n10505 = ( n580 & n10502 ) | ( n580 & ~n10504 ) | ( n10502 & ~n10504 ) ;
  assign n10509 = n10508 ^ n10505 ^ n1307 ;
  assign n10510 = n7319 ^ n4053 ^ 1'b0 ;
  assign n10514 = ~n1786 & n8307 ;
  assign n10515 = n1631 & n2189 ;
  assign n10516 = n10515 ^ n4463 ^ 1'b0 ;
  assign n10517 = ( ~n894 & n3873 ) | ( ~n894 & n7451 ) | ( n3873 & n7451 ) ;
  assign n10518 = ( n1347 & n10516 ) | ( n1347 & n10517 ) | ( n10516 & n10517 ) ;
  assign n10519 = ( n3661 & ~n10514 ) | ( n3661 & n10518 ) | ( ~n10514 & n10518 ) ;
  assign n10520 = n5319 & ~n6138 ;
  assign n10521 = ~n4090 & n10520 ;
  assign n10522 = n10521 ^ n6277 ^ x43 ;
  assign n10523 = n10522 ^ n1379 ^ 1'b0 ;
  assign n10524 = n10519 & n10523 ;
  assign n10511 = n2230 ^ n732 ^ 1'b0 ;
  assign n10512 = n10511 ^ n7753 ^ 1'b0 ;
  assign n10513 = n10512 ^ n5080 ^ 1'b0 ;
  assign n10525 = n10524 ^ n10513 ^ n5193 ;
  assign n10529 = n8809 ^ n8556 ^ n5256 ;
  assign n10527 = ( n1614 & n3267 ) | ( n1614 & n7579 ) | ( n3267 & n7579 ) ;
  assign n10526 = n2371 ^ n2102 ^ 1'b0 ;
  assign n10528 = n10527 ^ n10526 ^ n4883 ;
  assign n10530 = n10529 ^ n10528 ^ n409 ;
  assign n10531 = n1115 | n7299 ;
  assign n10532 = n4331 ^ n2277 ^ 1'b0 ;
  assign n10533 = n10532 ^ n6069 ^ n1731 ;
  assign n10534 = n10533 ^ n3423 ^ n1858 ;
  assign n10535 = n6695 ^ n6249 ^ n5658 ;
  assign n10536 = n10535 ^ n6992 ^ n1588 ;
  assign n10537 = ( ~n2175 & n10534 ) | ( ~n2175 & n10536 ) | ( n10534 & n10536 ) ;
  assign n10538 = ( ~n3229 & n4948 ) | ( ~n3229 & n6119 ) | ( n4948 & n6119 ) ;
  assign n10539 = ( n1364 & n9097 ) | ( n1364 & ~n9831 ) | ( n9097 & ~n9831 ) ;
  assign n10543 = n7148 ^ n6204 ^ n5608 ;
  assign n10541 = ( n2778 & n4217 ) | ( n2778 & n4671 ) | ( n4217 & n4671 ) ;
  assign n10542 = ( n1151 & ~n6157 ) | ( n1151 & n10541 ) | ( ~n6157 & n10541 ) ;
  assign n10544 = n10543 ^ n10542 ^ n773 ;
  assign n10540 = n7471 ^ n2640 ^ 1'b0 ;
  assign n10545 = n10544 ^ n10540 ^ n4116 ;
  assign n10546 = n1180 ^ n1015 ^ n223 ;
  assign n10547 = ~n2023 & n10546 ;
  assign n10548 = ~n10546 & n10547 ;
  assign n10549 = n5019 ^ n952 ^ 1'b0 ;
  assign n10550 = ~n4292 & n10549 ;
  assign n10551 = n10550 ^ n3846 ^ n665 ;
  assign n10552 = n4246 ^ n3867 ^ n2532 ;
  assign n10553 = n10551 & n10552 ;
  assign n10554 = n10553 ^ n5977 ^ n2426 ;
  assign n10555 = n10554 ^ n9158 ^ n1007 ;
  assign n10556 = ( ~n168 & n1507 ) | ( ~n168 & n2889 ) | ( n1507 & n2889 ) ;
  assign n10558 = n4719 ^ n1718 ^ 1'b0 ;
  assign n10559 = x119 & ~n10558 ;
  assign n10557 = ~n798 & n2812 ;
  assign n10560 = n10559 ^ n10557 ^ 1'b0 ;
  assign n10561 = ( n1853 & ~n10556 ) | ( n1853 & n10560 ) | ( ~n10556 & n10560 ) ;
  assign n10564 = ( ~n2241 & n5450 ) | ( ~n2241 & n8213 ) | ( n5450 & n8213 ) ;
  assign n10562 = ( n2613 & n2746 ) | ( n2613 & n4876 ) | ( n2746 & n4876 ) ;
  assign n10563 = n10562 ^ n7873 ^ n6630 ;
  assign n10565 = n10564 ^ n10563 ^ 1'b0 ;
  assign n10566 = ~n4541 & n10565 ;
  assign n10567 = n10566 ^ n10499 ^ 1'b0 ;
  assign n10568 = ( n567 & ~n6948 ) | ( n567 & n8906 ) | ( ~n6948 & n8906 ) ;
  assign n10569 = ( ~n2041 & n3272 ) | ( ~n2041 & n7936 ) | ( n3272 & n7936 ) ;
  assign n10570 = ( ~n2593 & n9670 ) | ( ~n2593 & n10569 ) | ( n9670 & n10569 ) ;
  assign n10571 = n1343 | n7309 ;
  assign n10572 = n10570 & ~n10571 ;
  assign n10574 = ~n4557 & n5250 ;
  assign n10575 = ( n1789 & ~n3852 ) | ( n1789 & n10574 ) | ( ~n3852 & n10574 ) ;
  assign n10576 = n2690 ^ n1284 ^ n1124 ;
  assign n10577 = n10576 ^ n8613 ^ n5056 ;
  assign n10578 = n1716 | n10577 ;
  assign n10579 = n10575 | n10578 ;
  assign n10573 = n5090 | n8556 ;
  assign n10580 = n10579 ^ n10573 ^ 1'b0 ;
  assign n10581 = ( n6577 & n10036 ) | ( n6577 & n10580 ) | ( n10036 & n10580 ) ;
  assign n10582 = ( n10568 & ~n10572 ) | ( n10568 & n10581 ) | ( ~n10572 & n10581 ) ;
  assign n10583 = n7422 ^ n2164 ^ 1'b0 ;
  assign n10584 = ( x34 & n2995 ) | ( x34 & n10583 ) | ( n2995 & n10583 ) ;
  assign n10585 = ( ~n2009 & n9648 ) | ( ~n2009 & n10584 ) | ( n9648 & n10584 ) ;
  assign n10586 = ~n1059 & n6951 ;
  assign n10587 = n10586 ^ n2544 ^ 1'b0 ;
  assign n10588 = n10587 ^ n9544 ^ 1'b0 ;
  assign n10589 = n3190 & n10588 ;
  assign n10590 = n10589 ^ n1661 ^ 1'b0 ;
  assign n10591 = n4571 | n10590 ;
  assign n10592 = ( n3059 & ~n6988 ) | ( n3059 & n10591 ) | ( ~n6988 & n10591 ) ;
  assign n10594 = n4139 & n6829 ;
  assign n10595 = n7498 ^ n4641 ^ n3041 ;
  assign n10596 = ( n955 & ~n7549 ) | ( n955 & n10595 ) | ( ~n7549 & n10595 ) ;
  assign n10597 = ( n9176 & n10594 ) | ( n9176 & n10596 ) | ( n10594 & n10596 ) ;
  assign n10598 = n10597 ^ n4191 ^ n3822 ;
  assign n10593 = n4881 ^ n4588 ^ 1'b0 ;
  assign n10599 = n10598 ^ n10593 ^ 1'b0 ;
  assign n10600 = n3620 | n10599 ;
  assign n10601 = n10378 ^ n5402 ^ n4213 ;
  assign n10602 = ( n436 & ~n2714 ) | ( n436 & n10601 ) | ( ~n2714 & n10601 ) ;
  assign n10603 = n7248 ^ n1440 ^ n728 ;
  assign n10604 = n4292 ^ n1335 ^ 1'b0 ;
  assign n10605 = ~n3596 & n10604 ;
  assign n10606 = n10605 ^ n9057 ^ n7162 ;
  assign n10607 = n10606 ^ n2391 ^ 1'b0 ;
  assign n10608 = ~n10603 & n10607 ;
  assign n10614 = n2725 ^ n2630 ^ n1513 ;
  assign n10615 = n10614 ^ n1790 ^ 1'b0 ;
  assign n10609 = n905 & n966 ;
  assign n10610 = ( n219 & ~n1895 ) | ( n219 & n10609 ) | ( ~n1895 & n10609 ) ;
  assign n10611 = ( ~n3923 & n9669 ) | ( ~n3923 & n10610 ) | ( n9669 & n10610 ) ;
  assign n10612 = n10611 ^ n9737 ^ n5549 ;
  assign n10613 = ( n144 & ~n9495 ) | ( n144 & n10612 ) | ( ~n9495 & n10612 ) ;
  assign n10616 = n10615 ^ n10613 ^ n2236 ;
  assign n10617 = n10616 ^ n6384 ^ n736 ;
  assign n10618 = ( n406 & n3269 ) | ( n406 & ~n10322 ) | ( n3269 & ~n10322 ) ;
  assign n10619 = n6456 | n10618 ;
  assign n10620 = ~n574 & n3549 ;
  assign n10621 = ~n5489 & n10620 ;
  assign n10622 = ( n1104 & n1717 ) | ( n1104 & n10621 ) | ( n1717 & n10621 ) ;
  assign n10623 = ( n5915 & ~n6785 ) | ( n5915 & n10622 ) | ( ~n6785 & n10622 ) ;
  assign n10624 = n10623 ^ n7904 ^ n6517 ;
  assign n10625 = ( n2656 & n2973 ) | ( n2656 & ~n6291 ) | ( n2973 & ~n6291 ) ;
  assign n10626 = ~n1469 & n2974 ;
  assign n10627 = n3863 & ~n10626 ;
  assign n10628 = n3614 & n10627 ;
  assign n10629 = n6742 ^ n5388 ^ 1'b0 ;
  assign n10630 = ( n9151 & ~n10628 ) | ( n9151 & n10629 ) | ( ~n10628 & n10629 ) ;
  assign n10631 = ( n3172 & ~n10625 ) | ( n3172 & n10630 ) | ( ~n10625 & n10630 ) ;
  assign n10632 = ( n3459 & n7266 ) | ( n3459 & n7371 ) | ( n7266 & n7371 ) ;
  assign n10633 = ( n263 & n1858 ) | ( n263 & ~n2322 ) | ( n1858 & ~n2322 ) ;
  assign n10634 = ( ~n450 & n5065 ) | ( ~n450 & n10633 ) | ( n5065 & n10633 ) ;
  assign n10635 = n10634 ^ n3852 ^ n523 ;
  assign n10636 = ( n4723 & ~n8169 ) | ( n4723 & n10635 ) | ( ~n8169 & n10635 ) ;
  assign n10637 = ( n2181 & n10632 ) | ( n2181 & ~n10636 ) | ( n10632 & ~n10636 ) ;
  assign n10639 = n1982 & ~n7644 ;
  assign n10640 = n10639 ^ n9518 ^ 1'b0 ;
  assign n10638 = n9235 & n10226 ;
  assign n10641 = n10640 ^ n10638 ^ n1979 ;
  assign n10642 = ( ~n4369 & n7605 ) | ( ~n4369 & n10641 ) | ( n7605 & n10641 ) ;
  assign n10644 = ( n2679 & n3359 ) | ( n2679 & n5001 ) | ( n3359 & n5001 ) ;
  assign n10643 = ( ~n786 & n2997 ) | ( ~n786 & n3009 ) | ( n2997 & n3009 ) ;
  assign n10645 = n10644 ^ n10643 ^ n3158 ;
  assign n10646 = ( n395 & ~n9526 ) | ( n395 & n10645 ) | ( ~n9526 & n10645 ) ;
  assign n10647 = n7009 | n10646 ;
  assign n10648 = n10647 ^ n823 ^ 1'b0 ;
  assign n10656 = n3483 ^ n2526 ^ 1'b0 ;
  assign n10657 = n3873 & ~n10656 ;
  assign n10658 = ( n1233 & ~n4123 ) | ( n1233 & n10657 ) | ( ~n4123 & n10657 ) ;
  assign n10649 = ( n153 & n444 ) | ( n153 & ~n805 ) | ( n444 & ~n805 ) ;
  assign n10650 = n10649 ^ n4522 ^ n810 ;
  assign n10651 = n10650 ^ n4874 ^ n299 ;
  assign n10652 = ~n251 & n1903 ;
  assign n10653 = n10652 ^ n10559 ^ n3859 ;
  assign n10654 = ~n3936 & n10653 ;
  assign n10655 = ~n10651 & n10654 ;
  assign n10659 = n10658 ^ n10655 ^ n4678 ;
  assign n10660 = n748 & n1196 ;
  assign n10661 = ~n3004 & n10660 ;
  assign n10662 = n6747 | n10661 ;
  assign n10663 = ( ~n1027 & n1281 ) | ( ~n1027 & n10662 ) | ( n1281 & n10662 ) ;
  assign n10664 = ( n377 & n2890 ) | ( n377 & ~n8158 ) | ( n2890 & ~n8158 ) ;
  assign n10665 = n966 & n10664 ;
  assign n10666 = ( ~x76 & n3799 ) | ( ~x76 & n10665 ) | ( n3799 & n10665 ) ;
  assign n10667 = n5226 ^ n3941 ^ n3724 ;
  assign n10668 = n10667 ^ n5440 ^ 1'b0 ;
  assign n10669 = ~n6949 & n10668 ;
  assign n10670 = n10669 ^ n7987 ^ n3594 ;
  assign n10671 = n5921 | n7698 ;
  assign n10672 = ~n9450 & n10671 ;
  assign n10673 = n10670 & n10672 ;
  assign n10674 = n10609 ^ n3767 ^ 1'b0 ;
  assign n10675 = n1121 & ~n10674 ;
  assign n10676 = ( n2773 & n5650 ) | ( n2773 & n10675 ) | ( n5650 & n10675 ) ;
  assign n10677 = ~n1027 & n10676 ;
  assign n10678 = n10677 ^ n6804 ^ 1'b0 ;
  assign n10679 = n10190 ^ n2355 ^ n1329 ;
  assign n10680 = n4108 ^ n3224 ^ 1'b0 ;
  assign n10681 = n247 & n10680 ;
  assign n10682 = n10681 ^ n1051 ^ 1'b0 ;
  assign n10683 = n2054 | n10682 ;
  assign n10684 = n10683 ^ n8893 ^ 1'b0 ;
  assign n10685 = n10684 ^ n3821 ^ n2256 ;
  assign n10686 = ( n545 & ~n607 ) | ( n545 & n2579 ) | ( ~n607 & n2579 ) ;
  assign n10687 = ( n1161 & ~n8201 ) | ( n1161 & n10686 ) | ( ~n8201 & n10686 ) ;
  assign n10688 = n901 & n10687 ;
  assign n10689 = ( n6598 & ~n10685 ) | ( n6598 & n10688 ) | ( ~n10685 & n10688 ) ;
  assign n10690 = n4661 & ~n7868 ;
  assign n10693 = n6870 ^ n6819 ^ n6406 ;
  assign n10691 = n1342 ^ n1146 ^ n1009 ;
  assign n10692 = ~n2610 & n10691 ;
  assign n10694 = n10693 ^ n10692 ^ 1'b0 ;
  assign n10695 = n10694 ^ n5529 ^ n3332 ;
  assign n10696 = n10695 ^ n9728 ^ 1'b0 ;
  assign n10697 = n10086 & n10696 ;
  assign n10698 = n9447 ^ n6067 ^ n914 ;
  assign n10701 = n5209 ^ n3511 ^ n1354 ;
  assign n10702 = ( n4781 & n9856 ) | ( n4781 & ~n10701 ) | ( n9856 & ~n10701 ) ;
  assign n10703 = n10702 ^ n9963 ^ n4558 ;
  assign n10704 = n10703 ^ n4422 ^ n1531 ;
  assign n10700 = n1336 & n7577 ;
  assign n10705 = n10704 ^ n10700 ^ 1'b0 ;
  assign n10699 = ( n676 & n2004 ) | ( n676 & n7775 ) | ( n2004 & n7775 ) ;
  assign n10706 = n10705 ^ n10699 ^ 1'b0 ;
  assign n10707 = ( n1801 & n9390 ) | ( n1801 & n10706 ) | ( n9390 & n10706 ) ;
  assign n10715 = ( n421 & n1835 ) | ( n421 & n3050 ) | ( n1835 & n3050 ) ;
  assign n10712 = n5973 ^ n4817 ^ n2714 ;
  assign n10713 = ( n1685 & ~n5896 ) | ( n1685 & n10712 ) | ( ~n5896 & n10712 ) ;
  assign n10714 = n7862 & ~n10713 ;
  assign n10709 = n1144 & n10185 ;
  assign n10710 = n3286 & n10709 ;
  assign n10708 = n9154 ^ n4660 ^ n868 ;
  assign n10711 = n10710 ^ n10708 ^ n7411 ;
  assign n10716 = n10715 ^ n10714 ^ n10711 ;
  assign n10717 = ( x34 & ~n294 ) | ( x34 & n7365 ) | ( ~n294 & n7365 ) ;
  assign n10718 = n5022 ^ n470 ^ 1'b0 ;
  assign n10719 = n8513 & ~n10718 ;
  assign n10720 = n10719 ^ n2823 ^ n1412 ;
  assign n10721 = ~n1359 & n1686 ;
  assign n10722 = n804 & n10721 ;
  assign n10723 = ~n10720 & n10722 ;
  assign n10724 = ~n6593 & n7387 ;
  assign n10725 = n2444 & ~n4553 ;
  assign n10726 = ~n1880 & n10725 ;
  assign n10728 = n4419 ^ n3600 ^ n800 ;
  assign n10729 = n10728 ^ n10715 ^ n465 ;
  assign n10730 = n5373 & ~n10729 ;
  assign n10731 = n10730 ^ n3808 ^ 1'b0 ;
  assign n10727 = n6070 ^ n1675 ^ n746 ;
  assign n10732 = n10731 ^ n10727 ^ n8703 ;
  assign n10736 = x55 & n2328 ;
  assign n10737 = n5972 | n10736 ;
  assign n10738 = n3315 & ~n10737 ;
  assign n10733 = n3225 & ~n7328 ;
  assign n10734 = n10733 ^ n4194 ^ n3649 ;
  assign n10735 = ( n2011 & n2718 ) | ( n2011 & n10734 ) | ( n2718 & n10734 ) ;
  assign n10739 = n10738 ^ n10735 ^ n8970 ;
  assign n10740 = n2365 & n2482 ;
  assign n10741 = n1333 & ~n3369 ;
  assign n10742 = ~n8838 & n10741 ;
  assign n10743 = n5334 ^ n5020 ^ 1'b0 ;
  assign n10744 = ~n10742 & n10743 ;
  assign n10745 = ( n10469 & n10740 ) | ( n10469 & n10744 ) | ( n10740 & n10744 ) ;
  assign n10746 = n6804 ^ n4052 ^ n3323 ;
  assign n10747 = n1403 & n2120 ;
  assign n10748 = ( n7177 & ~n8621 ) | ( n7177 & n10747 ) | ( ~n8621 & n10747 ) ;
  assign n10749 = n10748 ^ n6672 ^ n2032 ;
  assign n10750 = n3161 & n10749 ;
  assign n10751 = n10746 & n10750 ;
  assign n10752 = n10262 ^ n6210 ^ 1'b0 ;
  assign n10753 = ( n799 & n2789 ) | ( n799 & ~n10752 ) | ( n2789 & ~n10752 ) ;
  assign n10754 = n10753 ^ n2188 ^ 1'b0 ;
  assign n10755 = n7581 ^ n6978 ^ 1'b0 ;
  assign n10756 = n10755 ^ n9958 ^ n2754 ;
  assign n10757 = ( n2502 & n3336 ) | ( n2502 & n3427 ) | ( n3336 & n3427 ) ;
  assign n10758 = n4955 ^ n2004 ^ 1'b0 ;
  assign n10759 = n9469 ^ n6541 ^ n1371 ;
  assign n10760 = n3201 ^ n2487 ^ n2296 ;
  assign n10761 = n903 & ~n10760 ;
  assign n10762 = ( n5393 & n10759 ) | ( n5393 & ~n10761 ) | ( n10759 & ~n10761 ) ;
  assign n10763 = ( ~n10757 & n10758 ) | ( ~n10757 & n10762 ) | ( n10758 & n10762 ) ;
  assign n10764 = n3954 ^ n1333 ^ n1195 ;
  assign n10765 = ( n414 & n1234 ) | ( n414 & ~n3376 ) | ( n1234 & ~n3376 ) ;
  assign n10766 = n10765 ^ n10292 ^ n2167 ;
  assign n10767 = ( n1042 & ~n10764 ) | ( n1042 & n10766 ) | ( ~n10764 & n10766 ) ;
  assign n10768 = x86 & n4769 ;
  assign n10774 = n7671 ^ n5726 ^ n1258 ;
  assign n10769 = n10594 ^ n9169 ^ n166 ;
  assign n10770 = n1799 & ~n6133 ;
  assign n10771 = n10770 ^ n4365 ^ n3685 ;
  assign n10772 = ( ~n149 & n10769 ) | ( ~n149 & n10771 ) | ( n10769 & n10771 ) ;
  assign n10773 = ~n1050 & n10772 ;
  assign n10775 = n10774 ^ n10773 ^ 1'b0 ;
  assign n10776 = ( n1842 & n2199 ) | ( n1842 & ~n7445 ) | ( n2199 & ~n7445 ) ;
  assign n10777 = ( ~n553 & n903 ) | ( ~n553 & n5729 ) | ( n903 & n5729 ) ;
  assign n10778 = n10777 ^ n5876 ^ n1144 ;
  assign n10779 = ( n1499 & n2635 ) | ( n1499 & n4086 ) | ( n2635 & n4086 ) ;
  assign n10780 = n7165 | n10779 ;
  assign n10781 = n10778 & ~n10780 ;
  assign n10782 = n4956 & ~n7192 ;
  assign n10783 = ( ~n10776 & n10781 ) | ( ~n10776 & n10782 ) | ( n10781 & n10782 ) ;
  assign n10784 = n3583 | n10783 ;
  assign n10785 = ( x123 & ~n1160 ) | ( x123 & n4691 ) | ( ~n1160 & n4691 ) ;
  assign n10786 = n1999 | n10785 ;
  assign n10787 = ( x112 & n9053 ) | ( x112 & n10577 ) | ( n9053 & n10577 ) ;
  assign n10788 = ( x90 & n1400 ) | ( x90 & ~n10787 ) | ( n1400 & ~n10787 ) ;
  assign n10789 = ( n5701 & n10786 ) | ( n5701 & n10788 ) | ( n10786 & n10788 ) ;
  assign n10790 = ( n1971 & n2060 ) | ( n1971 & ~n5572 ) | ( n2060 & ~n5572 ) ;
  assign n10791 = n4677 & n10790 ;
  assign n10792 = n10791 ^ n3001 ^ 1'b0 ;
  assign n10797 = n3248 & ~n4418 ;
  assign n10798 = ~n453 & n10797 ;
  assign n10799 = ( n4958 & n9077 ) | ( n4958 & n10798 ) | ( n9077 & n10798 ) ;
  assign n10793 = n6764 ^ n5581 ^ n3496 ;
  assign n10794 = n2561 & n10793 ;
  assign n10795 = ~n5096 & n10794 ;
  assign n10796 = n10795 ^ n9158 ^ n3742 ;
  assign n10800 = n10799 ^ n10796 ^ n6923 ;
  assign n10801 = ( ~n3810 & n10792 ) | ( ~n3810 & n10800 ) | ( n10792 & n10800 ) ;
  assign n10802 = ( n258 & n5004 ) | ( n258 & n7582 ) | ( n5004 & n7582 ) ;
  assign n10803 = ( ~n3052 & n7499 ) | ( ~n3052 & n10802 ) | ( n7499 & n10802 ) ;
  assign n10804 = n10803 ^ n5522 ^ n1258 ;
  assign n10805 = n10804 ^ n8124 ^ n6985 ;
  assign n10806 = n7914 ^ n7593 ^ n5920 ;
  assign n10807 = ( n5082 & ~n8642 ) | ( n5082 & n10247 ) | ( ~n8642 & n10247 ) ;
  assign n10808 = n7167 & ~n7592 ;
  assign n10810 = n10722 ^ n8502 ^ n4326 ;
  assign n10809 = n7474 ^ n3760 ^ n960 ;
  assign n10811 = n10810 ^ n10809 ^ 1'b0 ;
  assign n10812 = n10808 & ~n10811 ;
  assign n10813 = n8402 & n8576 ;
  assign n10814 = n6275 ^ n937 ^ n379 ;
  assign n10815 = n10814 ^ n7842 ^ 1'b0 ;
  assign n10816 = n4604 ^ n1182 ^ 1'b0 ;
  assign n10817 = n4407 & ~n10816 ;
  assign n10818 = n10817 ^ n1386 ^ n384 ;
  assign n10819 = n10818 ^ n2240 ^ n1237 ;
  assign n10820 = ~n4840 & n10819 ;
  assign n10821 = n10815 & n10820 ;
  assign n10822 = n10821 ^ n7661 ^ n3691 ;
  assign n10823 = ( x99 & n6681 ) | ( x99 & ~n8334 ) | ( n6681 & ~n8334 ) ;
  assign n10824 = ( n4322 & n5221 ) | ( n4322 & ~n10823 ) | ( n5221 & ~n10823 ) ;
  assign n10832 = n2296 ^ n1879 ^ 1'b0 ;
  assign n10826 = n3214 & ~n6241 ;
  assign n10827 = ~n2632 & n10826 ;
  assign n10828 = n2851 ^ n394 ^ 1'b0 ;
  assign n10829 = n9544 ^ n4032 ^ n2995 ;
  assign n10830 = ( n10827 & n10828 ) | ( n10827 & n10829 ) | ( n10828 & n10829 ) ;
  assign n10825 = n7083 ^ n4571 ^ n3726 ;
  assign n10831 = n10830 ^ n10825 ^ n3093 ;
  assign n10833 = n10832 ^ n10831 ^ n5550 ;
  assign n10834 = ( ~n2079 & n6829 ) | ( ~n2079 & n8412 ) | ( n6829 & n8412 ) ;
  assign n10835 = ( n6843 & n10833 ) | ( n6843 & ~n10834 ) | ( n10833 & ~n10834 ) ;
  assign n10836 = n8884 ^ n2861 ^ x36 ;
  assign n10837 = n10191 ^ n3629 ^ 1'b0 ;
  assign n10844 = n7541 ^ n5522 ^ n1664 ;
  assign n10842 = n1584 | n3017 ;
  assign n10843 = n4281 | n10842 ;
  assign n10838 = n7049 ^ n1484 ^ n381 ;
  assign n10839 = ( ~n2082 & n2845 ) | ( ~n2082 & n6471 ) | ( n2845 & n6471 ) ;
  assign n10840 = ( n5283 & n5328 ) | ( n5283 & n10839 ) | ( n5328 & n10839 ) ;
  assign n10841 = n10838 & ~n10840 ;
  assign n10845 = n10844 ^ n10843 ^ n10841 ;
  assign n10846 = ( n7988 & n10837 ) | ( n7988 & ~n10845 ) | ( n10837 & ~n10845 ) ;
  assign n10847 = n10846 ^ n4729 ^ 1'b0 ;
  assign n10848 = n3320 | n4473 ;
  assign n10849 = n2449 | n10848 ;
  assign n10850 = n8087 ^ n4100 ^ n272 ;
  assign n10851 = ( n439 & n10849 ) | ( n439 & n10850 ) | ( n10849 & n10850 ) ;
  assign n10852 = ( ~n2692 & n5166 ) | ( ~n2692 & n5328 ) | ( n5166 & n5328 ) ;
  assign n10853 = n10852 ^ n5498 ^ n3137 ;
  assign n10854 = n7163 & n7896 ;
  assign n10855 = n7675 & n10854 ;
  assign n10856 = ( n676 & n1765 ) | ( n676 & n10740 ) | ( n1765 & n10740 ) ;
  assign n10857 = ( n7202 & n10459 ) | ( n7202 & ~n10856 ) | ( n10459 & ~n10856 ) ;
  assign n10858 = ( n761 & ~n4320 ) | ( n761 & n6591 ) | ( ~n4320 & n6591 ) ;
  assign n10859 = n2087 | n10858 ;
  assign n10860 = n10859 ^ n2923 ^ 1'b0 ;
  assign n10861 = ( ~n2878 & n3361 ) | ( ~n2878 & n10860 ) | ( n3361 & n10860 ) ;
  assign n10862 = n9699 & n10861 ;
  assign n10864 = n9667 ^ n8852 ^ n5945 ;
  assign n10863 = ( n238 & ~n1872 ) | ( n238 & n2247 ) | ( ~n1872 & n2247 ) ;
  assign n10865 = n10864 ^ n10863 ^ n6272 ;
  assign n10869 = ( n205 & n1079 ) | ( n205 & n3303 ) | ( n1079 & n3303 ) ;
  assign n10868 = ( n4280 & n5619 ) | ( n4280 & ~n10502 ) | ( n5619 & ~n10502 ) ;
  assign n10866 = ( n1359 & ~n7973 ) | ( n1359 & n8014 ) | ( ~n7973 & n8014 ) ;
  assign n10867 = n10866 ^ n2440 ^ n619 ;
  assign n10870 = n10869 ^ n10868 ^ n10867 ;
  assign n10871 = n539 & ~n1601 ;
  assign n10872 = ~n4778 & n10871 ;
  assign n10873 = n8922 ^ n1672 ^ 1'b0 ;
  assign n10874 = ~n10872 & n10873 ;
  assign n10877 = n426 & n10543 ;
  assign n10878 = ( ~n1546 & n4541 ) | ( ~n1546 & n10877 ) | ( n4541 & n10877 ) ;
  assign n10875 = n7314 ^ n4890 ^ 1'b0 ;
  assign n10876 = ~n1634 & n10875 ;
  assign n10879 = n10878 ^ n10876 ^ x15 ;
  assign n10880 = n5723 ^ n2142 ^ 1'b0 ;
  assign n10881 = n9773 & n10880 ;
  assign n10882 = ( n3936 & ~n4132 ) | ( n3936 & n10881 ) | ( ~n4132 & n10881 ) ;
  assign n10883 = ( n488 & n3116 ) | ( n488 & n9919 ) | ( n3116 & n9919 ) ;
  assign n10884 = n8531 ^ n5958 ^ n3775 ;
  assign n10885 = ( n1788 & n2905 ) | ( n1788 & ~n5507 ) | ( n2905 & ~n5507 ) ;
  assign n10886 = n10885 ^ n10650 ^ 1'b0 ;
  assign n10887 = n10884 | n10886 ;
  assign n10888 = n10887 ^ n8187 ^ n1329 ;
  assign n10889 = ( n7142 & ~n10883 ) | ( n7142 & n10888 ) | ( ~n10883 & n10888 ) ;
  assign n10890 = n10889 ^ n5929 ^ n4653 ;
  assign n10891 = n6138 ^ n4451 ^ n354 ;
  assign n10892 = n10891 ^ n4013 ^ n662 ;
  assign n10893 = n10892 ^ n8176 ^ n4812 ;
  assign n10894 = n6380 ^ n5610 ^ n1927 ;
  assign n10895 = n5990 ^ n5468 ^ 1'b0 ;
  assign n10896 = n10894 | n10895 ;
  assign n10897 = n4295 ^ n400 ^ 1'b0 ;
  assign n10898 = n10610 ^ n7613 ^ n2967 ;
  assign n10899 = n4201 ^ n2279 ^ n949 ;
  assign n10900 = n10899 ^ n3643 ^ n1340 ;
  assign n10901 = n10900 ^ n9595 ^ n4178 ;
  assign n10902 = n3426 | n10901 ;
  assign n10903 = n2968 | n4709 ;
  assign n10904 = n10903 ^ n207 ^ 1'b0 ;
  assign n10905 = n10904 ^ n6532 ^ 1'b0 ;
  assign n10906 = n858 & ~n10905 ;
  assign n10907 = ( ~n1925 & n7554 ) | ( ~n1925 & n8665 ) | ( n7554 & n8665 ) ;
  assign n10908 = n10907 ^ n6218 ^ 1'b0 ;
  assign n10909 = n10908 ^ n9487 ^ 1'b0 ;
  assign n10910 = n10906 & ~n10909 ;
  assign n10911 = ( n4266 & n5893 ) | ( n4266 & ~n9344 ) | ( n5893 & ~n9344 ) ;
  assign n10912 = ( ~n277 & n4929 ) | ( ~n277 & n5851 ) | ( n4929 & n5851 ) ;
  assign n10913 = n10912 ^ n4092 ^ 1'b0 ;
  assign n10914 = ( n9218 & n10911 ) | ( n9218 & ~n10913 ) | ( n10911 & ~n10913 ) ;
  assign n10915 = n7653 | n10914 ;
  assign n10916 = ( ~n4187 & n4876 ) | ( ~n4187 & n10915 ) | ( n4876 & n10915 ) ;
  assign n10917 = n3739 & ~n10916 ;
  assign n10918 = ~n10910 & n10917 ;
  assign n10919 = n4414 & ~n7476 ;
  assign n10920 = n10919 ^ n7011 ^ 1'b0 ;
  assign n10921 = n10920 ^ n10074 ^ n7153 ;
  assign n10922 = n9964 ^ n4963 ^ n855 ;
  assign n10923 = n10922 ^ n2631 ^ n338 ;
  assign n10924 = ( n2930 & n9873 ) | ( n2930 & n10923 ) | ( n9873 & n10923 ) ;
  assign n10925 = n5866 ^ n3642 ^ n348 ;
  assign n10926 = n9077 ^ n3432 ^ n1348 ;
  assign n10927 = n8113 ^ n3241 ^ n2379 ;
  assign n10928 = n2732 | n9846 ;
  assign n10929 = n10927 | n10928 ;
  assign n10930 = ( ~x112 & n1600 ) | ( ~x112 & n10929 ) | ( n1600 & n10929 ) ;
  assign n10931 = n3835 ^ n2618 ^ n574 ;
  assign n10932 = n10931 ^ n9359 ^ n3562 ;
  assign n10937 = n10376 ^ n1416 ^ 1'b0 ;
  assign n10938 = n246 | n10937 ;
  assign n10939 = n10938 ^ n5148 ^ n4597 ;
  assign n10933 = n4211 ^ n605 ^ n510 ;
  assign n10934 = n10933 ^ n4413 ^ n1748 ;
  assign n10935 = n10934 ^ n1264 ^ n1251 ;
  assign n10936 = ( n6365 & n6486 ) | ( n6365 & n10935 ) | ( n6486 & n10935 ) ;
  assign n10940 = n10939 ^ n10936 ^ 1'b0 ;
  assign n10941 = n373 ^ n350 ^ 1'b0 ;
  assign n10942 = n2271 & ~n10941 ;
  assign n10943 = n10942 ^ n7660 ^ n5959 ;
  assign n10948 = n7297 ^ n5972 ^ n4195 ;
  assign n10944 = ( n3257 & ~n3307 ) | ( n3257 & n5642 ) | ( ~n3307 & n5642 ) ;
  assign n10945 = ( n389 & ~n1647 ) | ( n389 & n10828 ) | ( ~n1647 & n10828 ) ;
  assign n10946 = n10945 ^ n5341 ^ n737 ;
  assign n10947 = n10944 | n10946 ;
  assign n10949 = n10948 ^ n10947 ^ n3967 ;
  assign n10950 = ( ~x27 & n3213 ) | ( ~x27 & n9285 ) | ( n3213 & n9285 ) ;
  assign n10951 = n8893 ^ n8591 ^ 1'b0 ;
  assign n10952 = ~n4081 & n10951 ;
  assign n10953 = ( n10931 & n10950 ) | ( n10931 & n10952 ) | ( n10950 & n10952 ) ;
  assign n10954 = n10953 ^ n3664 ^ 1'b0 ;
  assign n10955 = n7315 & ~n7805 ;
  assign n10956 = ~n6535 & n10955 ;
  assign n10964 = n10906 ^ n5320 ^ n1124 ;
  assign n10961 = n3981 | n6315 ;
  assign n10962 = n10961 ^ n10933 ^ 1'b0 ;
  assign n10957 = ( n2441 & ~n2909 ) | ( n2441 & n3230 ) | ( ~n2909 & n3230 ) ;
  assign n10958 = ( n4496 & n5142 ) | ( n4496 & ~n10957 ) | ( n5142 & ~n10957 ) ;
  assign n10959 = n10958 ^ n7046 ^ 1'b0 ;
  assign n10960 = x16 & n10959 ;
  assign n10963 = n10962 ^ n10960 ^ 1'b0 ;
  assign n10965 = n10964 ^ n10963 ^ x109 ;
  assign n10966 = ( n2560 & n6986 ) | ( n2560 & n9337 ) | ( n6986 & n9337 ) ;
  assign n10967 = n10966 ^ n1458 ^ 1'b0 ;
  assign n10968 = ( n869 & n3384 ) | ( n869 & n3489 ) | ( n3384 & n3489 ) ;
  assign n10969 = ( n3693 & n8063 ) | ( n3693 & ~n10968 ) | ( n8063 & ~n10968 ) ;
  assign n10970 = ( n8578 & n10634 ) | ( n8578 & n10969 ) | ( n10634 & n10969 ) ;
  assign n10971 = n4384 ^ n319 ^ 1'b0 ;
  assign n10972 = ~n4069 & n10971 ;
  assign n10973 = n10972 ^ n829 ^ 1'b0 ;
  assign n10974 = n9615 & ~n10973 ;
  assign n10975 = ( n1703 & ~n10970 ) | ( n1703 & n10974 ) | ( ~n10970 & n10974 ) ;
  assign n10976 = n4425 ^ n2196 ^ n150 ;
  assign n10977 = ( n4408 & ~n4463 ) | ( n4408 & n10976 ) | ( ~n4463 & n10976 ) ;
  assign n10978 = ( ~n855 & n2236 ) | ( ~n855 & n10977 ) | ( n2236 & n10977 ) ;
  assign n10979 = ( n993 & ~n4883 ) | ( n993 & n9007 ) | ( ~n4883 & n9007 ) ;
  assign n10985 = n6045 ^ n5213 ^ n1790 ;
  assign n10984 = ( n293 & n2561 ) | ( n293 & n10872 ) | ( n2561 & n10872 ) ;
  assign n10986 = n10985 ^ n10984 ^ n10001 ;
  assign n10980 = ~n964 & n1979 ;
  assign n10981 = n10980 ^ n4549 ^ 1'b0 ;
  assign n10982 = n10981 ^ n3589 ^ 1'b0 ;
  assign n10983 = n6361 & ~n10982 ;
  assign n10987 = n10986 ^ n10983 ^ 1'b0 ;
  assign n10988 = ( x17 & ~n10979 ) | ( x17 & n10987 ) | ( ~n10979 & n10987 ) ;
  assign n10989 = n1465 ^ n656 ^ n194 ;
  assign n10990 = n2788 ^ n561 ^ n520 ;
  assign n10991 = ( n3216 & ~n10989 ) | ( n3216 & n10990 ) | ( ~n10989 & n10990 ) ;
  assign n10993 = ( n1655 & ~n5800 ) | ( n1655 & n10373 ) | ( ~n5800 & n10373 ) ;
  assign n10992 = n5896 ^ n5051 ^ x48 ;
  assign n10994 = n10993 ^ n10992 ^ n8039 ;
  assign n10995 = n10888 ^ n7994 ^ 1'b0 ;
  assign n10996 = ( n3442 & ~n9510 ) | ( n3442 & n10223 ) | ( ~n9510 & n10223 ) ;
  assign n10997 = ( n2861 & n7999 ) | ( n2861 & ~n10996 ) | ( n7999 & ~n10996 ) ;
  assign n10998 = n5592 ^ n3135 ^ n582 ;
  assign n10999 = n9681 ^ n6713 ^ 1'b0 ;
  assign n11000 = n10998 & n10999 ;
  assign n11001 = n11000 ^ n4357 ^ n3064 ;
  assign n11002 = n11001 ^ n3226 ^ n1653 ;
  assign n11004 = n1690 & n4617 ;
  assign n11005 = ~n3373 & n11004 ;
  assign n11006 = n11005 ^ n4441 ^ x68 ;
  assign n11003 = n9652 ^ n7273 ^ n2412 ;
  assign n11007 = n11006 ^ n11003 ^ 1'b0 ;
  assign n11008 = n11002 | n11007 ;
  assign n11009 = n7878 ^ n3884 ^ n2667 ;
  assign n11010 = n988 ^ n207 ^ 1'b0 ;
  assign n11011 = n11010 ^ n7183 ^ n737 ;
  assign n11012 = n11011 ^ n8687 ^ 1'b0 ;
  assign n11013 = n340 | n11012 ;
  assign n11014 = n11013 ^ n9253 ^ n4983 ;
  assign n11015 = n2022 & ~n3106 ;
  assign n11016 = n11015 ^ n4764 ^ n1930 ;
  assign n11017 = ( n499 & n9602 ) | ( n499 & n11016 ) | ( n9602 & n11016 ) ;
  assign n11018 = n301 & n1200 ;
  assign n11019 = ( ~n886 & n3304 ) | ( ~n886 & n11018 ) | ( n3304 & n11018 ) ;
  assign n11020 = ( n2906 & n4116 ) | ( n2906 & ~n11019 ) | ( n4116 & ~n11019 ) ;
  assign n11021 = ( x35 & n1772 ) | ( x35 & ~n2343 ) | ( n1772 & ~n2343 ) ;
  assign n11022 = ( n9222 & n11020 ) | ( n9222 & ~n11021 ) | ( n11020 & ~n11021 ) ;
  assign n11023 = n11022 ^ n10830 ^ n1760 ;
  assign n11024 = ~n1363 & n10339 ;
  assign n11025 = ~n11023 & n11024 ;
  assign n11026 = ( n2061 & ~n5836 ) | ( n2061 & n10622 ) | ( ~n5836 & n10622 ) ;
  assign n11027 = ~n3062 & n3616 ;
  assign n11028 = n6354 ^ n3570 ^ n2047 ;
  assign n11029 = ( n4291 & n4578 ) | ( n4291 & n7881 ) | ( n4578 & n7881 ) ;
  assign n11030 = n470 | n3984 ;
  assign n11031 = n11030 ^ n2665 ^ 1'b0 ;
  assign n11032 = n11031 ^ n8524 ^ n1161 ;
  assign n11035 = n5208 ^ n394 ^ n138 ;
  assign n11033 = ( x95 & ~n304 ) | ( x95 & n1354 ) | ( ~n304 & n1354 ) ;
  assign n11034 = ( n8925 & n9560 ) | ( n8925 & n11033 ) | ( n9560 & n11033 ) ;
  assign n11036 = n11035 ^ n11034 ^ 1'b0 ;
  assign n11037 = ~n7238 & n11036 ;
  assign n11038 = n11037 ^ n398 ^ 1'b0 ;
  assign n11039 = n11032 & n11038 ;
  assign n11040 = n11029 & n11039 ;
  assign n11043 = ( n447 & n1694 ) | ( n447 & n8242 ) | ( n1694 & n8242 ) ;
  assign n11041 = n7791 ^ n4195 ^ n1708 ;
  assign n11042 = n8753 & n11041 ;
  assign n11044 = n11043 ^ n11042 ^ 1'b0 ;
  assign n11046 = ( n280 & n501 ) | ( n280 & ~n1273 ) | ( n501 & ~n1273 ) ;
  assign n11047 = n11046 ^ x14 ^ 1'b0 ;
  assign n11048 = ~n4280 & n11047 ;
  assign n11045 = n8897 ^ n8402 ^ n2383 ;
  assign n11049 = n11048 ^ n11045 ^ 1'b0 ;
  assign n11050 = n1299 | n11049 ;
  assign n11051 = ( n799 & ~n1525 ) | ( n799 & n8463 ) | ( ~n1525 & n8463 ) ;
  assign n11052 = n10652 ^ n4616 ^ n1241 ;
  assign n11053 = n11052 ^ n5356 ^ n5181 ;
  assign n11058 = ( n234 & n3458 ) | ( n234 & n4160 ) | ( n3458 & n4160 ) ;
  assign n11059 = n11058 ^ n7403 ^ n3261 ;
  assign n11060 = n11059 ^ n10759 ^ n8412 ;
  assign n11054 = ( n3466 & n8336 ) | ( n3466 & n9276 ) | ( n8336 & n9276 ) ;
  assign n11055 = ( ~n699 & n5055 ) | ( ~n699 & n11054 ) | ( n5055 & n11054 ) ;
  assign n11056 = n11055 ^ n5489 ^ 1'b0 ;
  assign n11057 = ( n4177 & n6851 ) | ( n4177 & ~n11056 ) | ( n6851 & ~n11056 ) ;
  assign n11061 = n11060 ^ n11057 ^ n5782 ;
  assign n11062 = ( ~n804 & n1448 ) | ( ~n804 & n5902 ) | ( n1448 & n5902 ) ;
  assign n11063 = ( n1317 & n1878 ) | ( n1317 & n2737 ) | ( n1878 & n2737 ) ;
  assign n11064 = ( n2615 & ~n5529 ) | ( n2615 & n11063 ) | ( ~n5529 & n11063 ) ;
  assign n11065 = n11064 ^ n10270 ^ n7713 ;
  assign n11066 = ( ~n699 & n3541 ) | ( ~n699 & n5467 ) | ( n3541 & n5467 ) ;
  assign n11067 = n9248 ^ n830 ^ 1'b0 ;
  assign n11068 = n8757 & n11067 ;
  assign n11069 = ~n11066 & n11068 ;
  assign n11071 = ( n672 & n1114 ) | ( n672 & n4819 ) | ( n1114 & n4819 ) ;
  assign n11070 = n2847 ^ n2220 ^ n2100 ;
  assign n11072 = n11071 ^ n11070 ^ n4342 ;
  assign n11073 = n5295 ^ n4176 ^ n515 ;
  assign n11074 = ~n2795 & n11073 ;
  assign n11075 = n6043 ^ n3127 ^ n2445 ;
  assign n11076 = ( n5029 & n7039 ) | ( n5029 & n11075 ) | ( n7039 & n11075 ) ;
  assign n11077 = n11076 ^ n5055 ^ n2853 ;
  assign n11078 = n701 & ~n11077 ;
  assign n11079 = n11074 & n11078 ;
  assign n11080 = ( n2815 & ~n3032 ) | ( n2815 & n10733 ) | ( ~n3032 & n10733 ) ;
  assign n11081 = n11080 ^ n9384 ^ n6197 ;
  assign n11082 = ( n1956 & n11079 ) | ( n1956 & n11081 ) | ( n11079 & n11081 ) ;
  assign n11083 = ( x117 & n4329 ) | ( x117 & ~n7762 ) | ( n4329 & ~n7762 ) ;
  assign n11084 = n11083 ^ n2940 ^ 1'b0 ;
  assign n11085 = ( n7951 & n10402 ) | ( n7951 & ~n11084 ) | ( n10402 & ~n11084 ) ;
  assign n11086 = ( ~n4143 & n6220 ) | ( ~n4143 & n11085 ) | ( n6220 & n11085 ) ;
  assign n11087 = n4909 & ~n5455 ;
  assign n11088 = n11087 ^ n7813 ^ 1'b0 ;
  assign n11089 = ( n3659 & n7578 ) | ( n3659 & ~n11088 ) | ( n7578 & ~n11088 ) ;
  assign n11090 = n5773 ^ n3624 ^ n2217 ;
  assign n11091 = ~n341 & n11090 ;
  assign n11092 = n4793 ^ n3068 ^ n638 ;
  assign n11093 = ( n2581 & n5681 ) | ( n2581 & n11092 ) | ( n5681 & n11092 ) ;
  assign n11094 = ( n268 & ~n10358 ) | ( n268 & n11093 ) | ( ~n10358 & n11093 ) ;
  assign n11095 = ( ~n3423 & n10301 ) | ( ~n3423 & n11094 ) | ( n10301 & n11094 ) ;
  assign n11096 = ~n319 & n10641 ;
  assign n11097 = n11096 ^ n3305 ^ n1926 ;
  assign n11098 = ~n7515 & n9364 ;
  assign n11099 = n896 ^ n570 ^ n211 ;
  assign n11100 = ( n6960 & n9514 ) | ( n6960 & n11099 ) | ( n9514 & n11099 ) ;
  assign n11101 = n11100 ^ n6450 ^ n4077 ;
  assign n11102 = ( ~n3367 & n8637 ) | ( ~n3367 & n11101 ) | ( n8637 & n11101 ) ;
  assign n11103 = ( n799 & ~n2997 ) | ( n799 & n4757 ) | ( ~n2997 & n4757 ) ;
  assign n11104 = ( n1495 & ~n6657 ) | ( n1495 & n11103 ) | ( ~n6657 & n11103 ) ;
  assign n11105 = n4092 ^ n706 ^ 1'b0 ;
  assign n11106 = n2054 ^ n428 ^ 1'b0 ;
  assign n11107 = ( n177 & n2336 ) | ( n177 & ~n11106 ) | ( n2336 & ~n11106 ) ;
  assign n11108 = ( n5014 & n6062 ) | ( n5014 & n11107 ) | ( n6062 & n11107 ) ;
  assign n11109 = ( n11034 & n11105 ) | ( n11034 & ~n11108 ) | ( n11105 & ~n11108 ) ;
  assign n11110 = n7325 & ~n11109 ;
  assign n11111 = n11110 ^ n9524 ^ 1'b0 ;
  assign n11117 = n8144 ^ n2808 ^ n2100 ;
  assign n11112 = n7634 ^ n7409 ^ n163 ;
  assign n11113 = n3722 ^ n1215 ^ n337 ;
  assign n11114 = ( ~n2139 & n3028 ) | ( ~n2139 & n7513 ) | ( n3028 & n7513 ) ;
  assign n11115 = ( n293 & ~n3769 ) | ( n293 & n11114 ) | ( ~n3769 & n11114 ) ;
  assign n11116 = ( ~n11112 & n11113 ) | ( ~n11112 & n11115 ) | ( n11113 & n11115 ) ;
  assign n11118 = n11117 ^ n11116 ^ n9965 ;
  assign n11130 = ( n1873 & n2882 ) | ( n1873 & ~n3564 ) | ( n2882 & ~n3564 ) ;
  assign n11128 = ( n1336 & n1857 ) | ( n1336 & n7272 ) | ( n1857 & n7272 ) ;
  assign n11129 = n11128 ^ n5247 ^ n1296 ;
  assign n11119 = ~n353 & n1686 ;
  assign n11120 = ~n4011 & n11119 ;
  assign n11121 = ( n1775 & n1849 ) | ( n1775 & n5747 ) | ( n1849 & n5747 ) ;
  assign n11122 = n6365 ^ n3191 ^ n1365 ;
  assign n11123 = n11121 & ~n11122 ;
  assign n11124 = ( n3419 & ~n11120 ) | ( n3419 & n11123 ) | ( ~n11120 & n11123 ) ;
  assign n11125 = ( n2489 & n2551 ) | ( n2489 & ~n6647 ) | ( n2551 & ~n6647 ) ;
  assign n11126 = n6345 & ~n11125 ;
  assign n11127 = ~n11124 & n11126 ;
  assign n11131 = n11130 ^ n11129 ^ n11127 ;
  assign n11132 = ( ~n3636 & n4913 ) | ( ~n3636 & n6303 ) | ( n4913 & n6303 ) ;
  assign n11133 = ~n7267 & n11132 ;
  assign n11134 = ~n4387 & n11133 ;
  assign n11135 = ( ~n5761 & n11131 ) | ( ~n5761 & n11134 ) | ( n11131 & n11134 ) ;
  assign n11136 = n2981 ^ n2869 ^ x67 ;
  assign n11137 = n11136 ^ n10380 ^ 1'b0 ;
  assign n11138 = ( ~n3241 & n7436 ) | ( ~n3241 & n10190 ) | ( n7436 & n10190 ) ;
  assign n11139 = ~n8447 & n11138 ;
  assign n11140 = n11139 ^ n1241 ^ 1'b0 ;
  assign n11141 = n8242 & ~n11140 ;
  assign n11142 = n11137 & n11141 ;
  assign n11143 = n2527 & n6510 ;
  assign n11144 = n11143 ^ n5892 ^ 1'b0 ;
  assign n11145 = ( x71 & ~n8456 ) | ( x71 & n11144 ) | ( ~n8456 & n11144 ) ;
  assign n11146 = ~n10846 & n11145 ;
  assign n11150 = n10839 ^ n8404 ^ n3060 ;
  assign n11147 = n5305 ^ n2356 ^ 1'b0 ;
  assign n11148 = n5439 & n11147 ;
  assign n11149 = ( ~n776 & n3971 ) | ( ~n776 & n11148 ) | ( n3971 & n11148 ) ;
  assign n11151 = n11150 ^ n11149 ^ n7164 ;
  assign n11152 = n2190 ^ n2055 ^ 1'b0 ;
  assign n11153 = n11152 ^ n7563 ^ n6609 ;
  assign n11154 = ( ~n9662 & n10429 ) | ( ~n9662 & n11153 ) | ( n10429 & n11153 ) ;
  assign n11165 = n7424 ^ n7268 ^ n4619 ;
  assign n11161 = ( n724 & n835 ) | ( n724 & n2452 ) | ( n835 & n2452 ) ;
  assign n11160 = n2619 & ~n5281 ;
  assign n11162 = n11161 ^ n11160 ^ 1'b0 ;
  assign n11163 = n11162 ^ n10757 ^ 1'b0 ;
  assign n11164 = n6007 | n11163 ;
  assign n11166 = n11165 ^ n11164 ^ n3339 ;
  assign n11158 = n5871 ^ n4383 ^ n2042 ;
  assign n11156 = n5443 ^ n2544 ^ 1'b0 ;
  assign n11157 = ( n1864 & n10000 ) | ( n1864 & ~n11156 ) | ( n10000 & ~n11156 ) ;
  assign n11159 = n11158 ^ n11157 ^ n6808 ;
  assign n11155 = ( n1960 & n6384 ) | ( n1960 & n6637 ) | ( n6384 & n6637 ) ;
  assign n11167 = n11166 ^ n11159 ^ n11155 ;
  assign n11168 = ( n623 & ~n4246 ) | ( n623 & n7155 ) | ( ~n4246 & n7155 ) ;
  assign n11169 = ~n3603 & n11168 ;
  assign n11170 = n3306 & n11169 ;
  assign n11171 = ( n133 & n10002 ) | ( n133 & n11170 ) | ( n10002 & n11170 ) ;
  assign n11172 = n5012 ^ n2483 ^ 1'b0 ;
  assign n11173 = n838 | n11172 ;
  assign n11174 = ( ~n1670 & n3605 ) | ( ~n1670 & n11173 ) | ( n3605 & n11173 ) ;
  assign n11175 = ( n2230 & n5636 ) | ( n2230 & n11174 ) | ( n5636 & n11174 ) ;
  assign n11176 = n11175 ^ n1674 ^ n1272 ;
  assign n11177 = n11176 ^ n8418 ^ 1'b0 ;
  assign n11178 = ( n3639 & ~n3716 ) | ( n3639 & n4651 ) | ( ~n3716 & n4651 ) ;
  assign n11179 = ( ~n2893 & n6267 ) | ( ~n2893 & n11178 ) | ( n6267 & n11178 ) ;
  assign n11180 = n3392 & n9328 ;
  assign n11181 = ~n4604 & n11180 ;
  assign n11182 = ( n777 & n1448 ) | ( n777 & ~n11181 ) | ( n1448 & ~n11181 ) ;
  assign n11183 = n1121 & n11182 ;
  assign n11184 = ~n11179 & n11183 ;
  assign n11185 = ( n163 & n4973 ) | ( n163 & n5697 ) | ( n4973 & n5697 ) ;
  assign n11186 = n9468 ^ n4755 ^ 1'b0 ;
  assign n11187 = n11185 | n11186 ;
  assign n11188 = ( n366 & ~n1196 ) | ( n366 & n3637 ) | ( ~n1196 & n3637 ) ;
  assign n11189 = n8787 ^ n5942 ^ n2976 ;
  assign n11190 = n11189 ^ n2883 ^ n198 ;
  assign n11191 = ~n1787 & n11190 ;
  assign n11192 = n11188 & n11191 ;
  assign n11193 = n2164 & ~n5118 ;
  assign n11194 = n11193 ^ n5975 ^ 1'b0 ;
  assign n11195 = n11194 ^ n6557 ^ n4674 ;
  assign n11196 = n11195 ^ n2968 ^ n935 ;
  assign n11197 = n4747 ^ n2851 ^ 1'b0 ;
  assign n11198 = n9966 | n11197 ;
  assign n11199 = n6471 ^ n6470 ^ n404 ;
  assign n11200 = ( n983 & n1237 ) | ( n983 & n3690 ) | ( n1237 & n3690 ) ;
  assign n11201 = n323 | n11200 ;
  assign n11202 = ~n11199 & n11201 ;
  assign n11203 = n11198 & n11202 ;
  assign n11204 = n2336 & ~n4697 ;
  assign n11205 = n5473 & n11204 ;
  assign n11206 = ~n3288 & n10770 ;
  assign n11207 = n6033 | n6523 ;
  assign n11208 = ( n7665 & n7908 ) | ( n7665 & n11207 ) | ( n7908 & n11207 ) ;
  assign n11209 = n11179 ^ n2671 ^ n810 ;
  assign n11210 = n11209 ^ n10333 ^ 1'b0 ;
  assign n11211 = n3873 ^ n1449 ^ 1'b0 ;
  assign n11212 = ~n7458 & n11211 ;
  assign n11213 = ( n3336 & n4597 ) | ( n3336 & n11212 ) | ( n4597 & n11212 ) ;
  assign n11214 = n11213 ^ n5458 ^ n3184 ;
  assign n11215 = n11214 ^ n3199 ^ n588 ;
  assign n11216 = n4425 ^ n4382 ^ 1'b0 ;
  assign n11217 = n11216 ^ n10729 ^ n4383 ;
  assign n11218 = ( n2497 & n11215 ) | ( n2497 & ~n11217 ) | ( n11215 & ~n11217 ) ;
  assign n11219 = ( ~n538 & n1406 ) | ( ~n538 & n2033 ) | ( n1406 & n2033 ) ;
  assign n11220 = n11219 ^ n2415 ^ n1365 ;
  assign n11221 = n11220 ^ n10105 ^ n2008 ;
  assign n11222 = ( n2592 & n3779 ) | ( n2592 & ~n4121 ) | ( n3779 & ~n4121 ) ;
  assign n11223 = ~n9092 & n11222 ;
  assign n11224 = n10351 ^ n6225 ^ n6094 ;
  assign n11225 = n11224 ^ n1329 ^ 1'b0 ;
  assign n11226 = ( n4500 & n8603 ) | ( n4500 & ~n11225 ) | ( n8603 & ~n11225 ) ;
  assign n11230 = n9856 ^ n8683 ^ n5282 ;
  assign n11231 = ~n4100 & n6770 ;
  assign n11232 = n3966 & n11231 ;
  assign n11233 = n11232 ^ n4181 ^ 1'b0 ;
  assign n11234 = n11230 & n11233 ;
  assign n11227 = n1903 ^ n561 ^ 1'b0 ;
  assign n11228 = n2356 | n4585 ;
  assign n11229 = n11227 | n11228 ;
  assign n11235 = n11234 ^ n11229 ^ n8352 ;
  assign n11236 = ( n1957 & n2016 ) | ( n1957 & n4248 ) | ( n2016 & n4248 ) ;
  assign n11237 = n4599 & ~n8333 ;
  assign n11238 = n11237 ^ n9450 ^ 1'b0 ;
  assign n11239 = n11236 & n11238 ;
  assign n11240 = ( n7123 & n7410 ) | ( n7123 & n8552 ) | ( n7410 & n8552 ) ;
  assign n11241 = n7541 | n11240 ;
  assign n11242 = n3061 | n11241 ;
  assign n11243 = ~n1154 & n4362 ;
  assign n11244 = n3767 & n11243 ;
  assign n11245 = n11244 ^ n986 ^ 1'b0 ;
  assign n11246 = n4956 | n11245 ;
  assign n11247 = n11246 ^ n10322 ^ n3220 ;
  assign n11248 = n2660 ^ n451 ^ 1'b0 ;
  assign n11249 = ~n3425 & n11248 ;
  assign n11250 = n11249 ^ n254 ^ n163 ;
  assign n11251 = n11250 ^ n2434 ^ n1912 ;
  assign n11252 = n11251 ^ n6659 ^ 1'b0 ;
  assign n11253 = n11247 | n11252 ;
  assign n11254 = n4302 ^ n2850 ^ n2723 ;
  assign n11255 = ( n3324 & n5660 ) | ( n3324 & ~n8186 ) | ( n5660 & ~n8186 ) ;
  assign n11256 = ( n10562 & n11254 ) | ( n10562 & n11255 ) | ( n11254 & n11255 ) ;
  assign n11257 = ( ~n6302 & n10378 ) | ( ~n6302 & n10398 ) | ( n10378 & n10398 ) ;
  assign n11259 = ( n6835 & n7371 ) | ( n6835 & n8092 ) | ( n7371 & n8092 ) ;
  assign n11258 = ( n3748 & n7380 ) | ( n3748 & n8414 ) | ( n7380 & n8414 ) ;
  assign n11260 = n11259 ^ n11258 ^ n7601 ;
  assign n11261 = ( n1374 & n6707 ) | ( n1374 & n11260 ) | ( n6707 & n11260 ) ;
  assign n11262 = n5241 & ~n7621 ;
  assign n11263 = n3203 & n11262 ;
  assign n11264 = n7403 ^ n7007 ^ n2051 ;
  assign n11265 = n11263 & n11264 ;
  assign n11266 = ( n1432 & n2962 ) | ( n1432 & ~n5408 ) | ( n2962 & ~n5408 ) ;
  assign n11267 = n8479 ^ n3773 ^ n3315 ;
  assign n11268 = n3349 & n11267 ;
  assign n11269 = n11268 ^ n9064 ^ 1'b0 ;
  assign n11270 = ( ~n2967 & n11266 ) | ( ~n2967 & n11269 ) | ( n11266 & n11269 ) ;
  assign n11271 = ( n4120 & n7703 ) | ( n4120 & n11270 ) | ( n7703 & n11270 ) ;
  assign n11272 = n3097 | n11271 ;
  assign n11273 = x106 & n3325 ;
  assign n11274 = n2806 & n11273 ;
  assign n11275 = n4272 & n11274 ;
  assign n11276 = ( n2293 & ~n4824 ) | ( n2293 & n11275 ) | ( ~n4824 & n11275 ) ;
  assign n11277 = n9862 ^ n9503 ^ n7682 ;
  assign n11278 = n8840 ^ n5672 ^ n1558 ;
  assign n11279 = ( n717 & n2640 ) | ( n717 & ~n4068 ) | ( n2640 & ~n4068 ) ;
  assign n11280 = ( n3285 & ~n7967 ) | ( n3285 & n11279 ) | ( ~n7967 & n11279 ) ;
  assign n11281 = ( n7274 & ~n7876 ) | ( n7274 & n11280 ) | ( ~n7876 & n11280 ) ;
  assign n11282 = n11278 & n11281 ;
  assign n11283 = ~n2921 & n5159 ;
  assign n11284 = n11283 ^ n2093 ^ 1'b0 ;
  assign n11285 = ( n6204 & ~n9104 ) | ( n6204 & n11284 ) | ( ~n9104 & n11284 ) ;
  assign n11286 = n803 & n11242 ;
  assign n11287 = n11285 & n11286 ;
  assign n11288 = n2576 ^ n1215 ^ 1'b0 ;
  assign n11291 = n354 | n8296 ;
  assign n11292 = n2376 & ~n11291 ;
  assign n11293 = n10957 | n11292 ;
  assign n11294 = n10074 & ~n11293 ;
  assign n11289 = n1232 ^ n1222 ^ 1'b0 ;
  assign n11290 = n9030 | n11289 ;
  assign n11295 = n11294 ^ n11290 ^ n8003 ;
  assign n11296 = ( n235 & ~n7191 ) | ( n235 & n7202 ) | ( ~n7191 & n7202 ) ;
  assign n11297 = ( n4606 & n4870 ) | ( n4606 & ~n5489 ) | ( n4870 & ~n5489 ) ;
  assign n11298 = ( n5413 & n9567 ) | ( n5413 & ~n11297 ) | ( n9567 & ~n11297 ) ;
  assign n11299 = n2529 & ~n7644 ;
  assign n11300 = n11299 ^ n4295 ^ 1'b0 ;
  assign n11303 = n5799 ^ n1484 ^ 1'b0 ;
  assign n11304 = n4064 & ~n11303 ;
  assign n11305 = n11304 ^ n147 ^ 1'b0 ;
  assign n11306 = n2925 & ~n11305 ;
  assign n11301 = n2242 ^ n2018 ^ 1'b0 ;
  assign n11302 = n1310 & ~n11301 ;
  assign n11307 = n11306 ^ n11302 ^ 1'b0 ;
  assign n11308 = n5794 & ~n11307 ;
  assign n11309 = n11082 ^ n7128 ^ n1618 ;
  assign n11310 = n7841 ^ n3356 ^ n2839 ;
  assign n11312 = n653 ^ n429 ^ n208 ;
  assign n11311 = ~n3622 & n7673 ;
  assign n11313 = n11312 ^ n11311 ^ n2854 ;
  assign n11314 = ( ~n3532 & n8769 ) | ( ~n3532 & n10210 ) | ( n8769 & n10210 ) ;
  assign n11315 = ( n1893 & ~n4831 ) | ( n1893 & n8902 ) | ( ~n4831 & n8902 ) ;
  assign n11316 = n1477 & n11315 ;
  assign n11317 = ~n2742 & n11316 ;
  assign n11318 = n1227 | n6489 ;
  assign n11319 = n11318 ^ n8140 ^ 1'b0 ;
  assign n11321 = ~n841 & n6156 ;
  assign n11320 = n6935 ^ n3374 ^ n2979 ;
  assign n11322 = n11321 ^ n11320 ^ n6953 ;
  assign n11323 = ( ~n1914 & n2338 ) | ( ~n1914 & n11322 ) | ( n2338 & n11322 ) ;
  assign n11324 = n7831 | n10730 ;
  assign n11325 = n11324 ^ n6630 ^ 1'b0 ;
  assign n11326 = n2892 & n7133 ;
  assign n11327 = ~n7588 & n11326 ;
  assign n11328 = n11327 ^ n6022 ^ n2190 ;
  assign n11329 = ( ~n3279 & n11325 ) | ( ~n3279 & n11328 ) | ( n11325 & n11328 ) ;
  assign n11330 = ( n1438 & n1894 ) | ( n1438 & n2186 ) | ( n1894 & n2186 ) ;
  assign n11331 = n11330 ^ n4428 ^ n586 ;
  assign n11332 = n4890 ^ n3152 ^ 1'b0 ;
  assign n11333 = n673 & ~n11332 ;
  assign n11334 = n7254 ^ n6540 ^ n432 ;
  assign n11335 = ( ~n7849 & n10533 ) | ( ~n7849 & n11334 ) | ( n10533 & n11334 ) ;
  assign n11336 = ( ~n11331 & n11333 ) | ( ~n11331 & n11335 ) | ( n11333 & n11335 ) ;
  assign n11337 = ( n1481 & n2730 ) | ( n1481 & ~n3185 ) | ( n2730 & ~n3185 ) ;
  assign n11338 = ( n3683 & n4173 ) | ( n3683 & ~n11337 ) | ( n4173 & ~n11337 ) ;
  assign n11339 = ( n2599 & n10024 ) | ( n2599 & ~n11338 ) | ( n10024 & ~n11338 ) ;
  assign n11340 = n5862 ^ n2373 ^ n249 ;
  assign n11344 = n10201 ^ n4613 ^ 1'b0 ;
  assign n11345 = n5919 & ~n11344 ;
  assign n11341 = n3760 ^ n2225 ^ n833 ;
  assign n11342 = ( ~n995 & n3579 ) | ( ~n995 & n11341 ) | ( n3579 & n11341 ) ;
  assign n11343 = ( n5388 & ~n7832 ) | ( n5388 & n11342 ) | ( ~n7832 & n11342 ) ;
  assign n11346 = n11345 ^ n11343 ^ n3489 ;
  assign n11347 = ( n2189 & n3683 ) | ( n2189 & n8104 ) | ( n3683 & n8104 ) ;
  assign n11348 = ( n2988 & n8372 ) | ( n2988 & ~n11347 ) | ( n8372 & ~n11347 ) ;
  assign n11349 = n9662 ^ n6575 ^ 1'b0 ;
  assign n11350 = n5885 & ~n11349 ;
  assign n11351 = n1942 ^ n352 ^ x81 ;
  assign n11357 = ( n3320 & n4691 ) | ( n3320 & n7830 ) | ( n4691 & n7830 ) ;
  assign n11354 = n8922 ^ n8338 ^ n3669 ;
  assign n11355 = ( n3116 & n10122 ) | ( n3116 & ~n11354 ) | ( n10122 & ~n11354 ) ;
  assign n11352 = n4828 | n5692 ;
  assign n11353 = x106 | n11352 ;
  assign n11356 = n11355 ^ n11353 ^ n990 ;
  assign n11358 = n11357 ^ n11356 ^ n4190 ;
  assign n11359 = ( n3831 & ~n4008 ) | ( n3831 & n8087 ) | ( ~n4008 & n8087 ) ;
  assign n11360 = n11359 ^ n6621 ^ 1'b0 ;
  assign n11361 = n10404 & ~n11360 ;
  assign n11362 = n4507 | n7909 ;
  assign n11363 = n1469 & ~n11362 ;
  assign n11364 = ( n1957 & ~n11361 ) | ( n1957 & n11363 ) | ( ~n11361 & n11363 ) ;
  assign n11381 = n9593 ^ n3692 ^ 1'b0 ;
  assign n11382 = n5216 & ~n11381 ;
  assign n11378 = n3865 ^ n2475 ^ 1'b0 ;
  assign n11379 = ~n5671 & n11378 ;
  assign n11367 = n2050 ^ n1196 ^ 1'b0 ;
  assign n11368 = n3084 & n11367 ;
  assign n11369 = ( n2748 & n6204 ) | ( n2748 & ~n11368 ) | ( n6204 & ~n11368 ) ;
  assign n11371 = ~n1941 & n6087 ;
  assign n11372 = n11371 ^ n2666 ^ 1'b0 ;
  assign n11370 = ( n1598 & n2028 ) | ( n1598 & ~n3633 ) | ( n2028 & ~n3633 ) ;
  assign n11373 = n11372 ^ n11370 ^ n864 ;
  assign n11374 = n3350 & n11373 ;
  assign n11375 = n11374 ^ n3047 ^ 1'b0 ;
  assign n11376 = ( n7104 & n11369 ) | ( n7104 & n11375 ) | ( n11369 & n11375 ) ;
  assign n11377 = ( n5397 & n9129 ) | ( n5397 & ~n11376 ) | ( n9129 & ~n11376 ) ;
  assign n11365 = n612 & n7765 ;
  assign n11366 = n3063 & n11365 ;
  assign n11380 = n11379 ^ n11377 ^ n11366 ;
  assign n11383 = n11382 ^ n11380 ^ 1'b0 ;
  assign n11384 = n11364 | n11383 ;
  assign n11385 = ( ~n7935 & n11232 ) | ( ~n7935 & n11384 ) | ( n11232 & n11384 ) ;
  assign n11386 = ( n578 & n1883 ) | ( n578 & n6658 ) | ( n1883 & n6658 ) ;
  assign n11387 = n8623 ^ n3050 ^ n809 ;
  assign n11388 = ( n362 & ~n1424 ) | ( n362 & n2599 ) | ( ~n1424 & n2599 ) ;
  assign n11389 = n11388 ^ n3357 ^ 1'b0 ;
  assign n11390 = n11387 | n11389 ;
  assign n11391 = ( x88 & ~n692 ) | ( x88 & n6073 ) | ( ~n692 & n6073 ) ;
  assign n11392 = n11391 ^ n8690 ^ n426 ;
  assign n11393 = n5264 ^ n2982 ^ n1135 ;
  assign n11397 = n2128 ^ n1538 ^ n309 ;
  assign n11394 = ( n2857 & n7065 ) | ( n2857 & n7760 ) | ( n7065 & n7760 ) ;
  assign n11395 = x45 & ~n11394 ;
  assign n11396 = n11395 ^ n380 ^ 1'b0 ;
  assign n11398 = n11397 ^ n11396 ^ n4588 ;
  assign n11399 = ( n9616 & n9890 ) | ( n9616 & n11398 ) | ( n9890 & n11398 ) ;
  assign n11400 = n7943 | n11399 ;
  assign n11401 = n3607 & ~n11400 ;
  assign n11402 = n2981 ^ n2528 ^ n2135 ;
  assign n11403 = n11402 ^ n2550 ^ n627 ;
  assign n11405 = n5165 & n10643 ;
  assign n11404 = n8192 ^ n6796 ^ n3581 ;
  assign n11406 = n11405 ^ n11404 ^ n4098 ;
  assign n11407 = n2311 ^ n2268 ^ x119 ;
  assign n11408 = n10819 | n11407 ;
  assign n11411 = n10576 ^ n6075 ^ n1637 ;
  assign n11410 = n10059 ^ n9271 ^ 1'b0 ;
  assign n11409 = n10828 ^ n8295 ^ n2776 ;
  assign n11412 = n11411 ^ n11410 ^ n11409 ;
  assign n11413 = ( n2990 & n5080 ) | ( n2990 & n8881 ) | ( n5080 & n8881 ) ;
  assign n11414 = n388 | n421 ;
  assign n11415 = n11414 ^ n1303 ^ 1'b0 ;
  assign n11416 = n11415 ^ n2006 ^ 1'b0 ;
  assign n11417 = n11416 ^ n5109 ^ n1005 ;
  assign n11418 = n11413 | n11417 ;
  assign n11419 = n11418 ^ n8897 ^ 1'b0 ;
  assign n11420 = n11419 ^ n2648 ^ 1'b0 ;
  assign n11421 = n11420 ^ n9331 ^ n6493 ;
  assign n11422 = n9744 ^ n8217 ^ 1'b0 ;
  assign n11423 = ~n6325 & n11422 ;
  assign n11431 = n3595 & ~n4161 ;
  assign n11432 = ~x11 & n11431 ;
  assign n11433 = ( n354 & n7566 ) | ( n354 & ~n11432 ) | ( n7566 & ~n11432 ) ;
  assign n11428 = ( n2955 & n4994 ) | ( n2955 & ~n7543 ) | ( n4994 & ~n7543 ) ;
  assign n11429 = n11428 ^ n11092 ^ n6835 ;
  assign n11424 = ( n2493 & n2858 ) | ( n2493 & n6976 ) | ( n2858 & n6976 ) ;
  assign n11425 = ( n191 & ~n376 ) | ( n191 & n1909 ) | ( ~n376 & n1909 ) ;
  assign n11426 = n11425 ^ n7518 ^ n2216 ;
  assign n11427 = n11424 & ~n11426 ;
  assign n11430 = n11429 ^ n11427 ^ 1'b0 ;
  assign n11434 = n11433 ^ n11430 ^ 1'b0 ;
  assign n11435 = ( n159 & n1084 ) | ( n159 & n4444 ) | ( n1084 & n4444 ) ;
  assign n11436 = ( n661 & n10452 ) | ( n661 & ~n11435 ) | ( n10452 & ~n11435 ) ;
  assign n11437 = n11436 ^ n5772 ^ n4604 ;
  assign n11438 = n10064 ^ n9482 ^ n4278 ;
  assign n11439 = n4106 & ~n9433 ;
  assign n11440 = ( ~n7168 & n11438 ) | ( ~n7168 & n11439 ) | ( n11438 & n11439 ) ;
  assign n11441 = ( ~n4663 & n11437 ) | ( ~n4663 & n11440 ) | ( n11437 & n11440 ) ;
  assign n11442 = n11441 ^ n9879 ^ 1'b0 ;
  assign n11443 = n9230 | n11442 ;
  assign n11445 = ~n900 & n2153 ;
  assign n11446 = n2959 & n11445 ;
  assign n11447 = n2089 & n11446 ;
  assign n11444 = ( x39 & n3129 ) | ( x39 & ~n6389 ) | ( n3129 & ~n6389 ) ;
  assign n11448 = n11447 ^ n11444 ^ 1'b0 ;
  assign n11449 = n7532 & ~n11448 ;
  assign n11450 = n2587 ^ n867 ^ n331 ;
  assign n11451 = ( ~n832 & n6646 ) | ( ~n832 & n11450 ) | ( n6646 & n11450 ) ;
  assign n11452 = n11451 ^ n4644 ^ 1'b0 ;
  assign n11453 = ~n7344 & n11452 ;
  assign n11454 = ( n1126 & ~n4346 ) | ( n1126 & n6557 ) | ( ~n4346 & n6557 ) ;
  assign n11455 = n5583 ^ n3901 ^ n133 ;
  assign n11456 = ( n280 & ~n3152 ) | ( n280 & n5260 ) | ( ~n3152 & n5260 ) ;
  assign n11457 = ( n7959 & n11455 ) | ( n7959 & ~n11456 ) | ( n11455 & ~n11456 ) ;
  assign n11458 = ( n6883 & n8844 ) | ( n6883 & n11457 ) | ( n8844 & n11457 ) ;
  assign n11459 = ( ~n3881 & n6515 ) | ( ~n3881 & n10502 ) | ( n6515 & n10502 ) ;
  assign n11460 = ( n3442 & ~n9316 ) | ( n3442 & n11459 ) | ( ~n9316 & n11459 ) ;
  assign n11461 = n5774 | n11460 ;
  assign n11462 = n1344 | n11461 ;
  assign n11463 = n11462 ^ n4851 ^ n620 ;
  assign n11464 = n8451 ^ n4895 ^ n2776 ;
  assign n11465 = n10332 ^ n1852 ^ n888 ;
  assign n11466 = ( n3355 & n5443 ) | ( n3355 & n7608 ) | ( n5443 & n7608 ) ;
  assign n11467 = n5529 ^ n578 ^ 1'b0 ;
  assign n11468 = ( n11465 & n11466 ) | ( n11465 & n11467 ) | ( n11466 & n11467 ) ;
  assign n11469 = n6971 & n9212 ;
  assign n11470 = n2249 ^ n2178 ^ n567 ;
  assign n11471 = n11470 ^ n3581 ^ 1'b0 ;
  assign n11472 = n11469 | n11471 ;
  assign n11474 = n4888 ^ n3434 ^ n373 ;
  assign n11473 = n4045 & ~n5348 ;
  assign n11475 = n11474 ^ n11473 ^ 1'b0 ;
  assign n11476 = ~n2781 & n11475 ;
  assign n11480 = n7487 ^ n6325 ^ n1786 ;
  assign n11478 = ( n790 & n5076 ) | ( n790 & n7960 ) | ( n5076 & n7960 ) ;
  assign n11477 = ( n3153 & n8072 ) | ( n3153 & ~n10511 ) | ( n8072 & ~n10511 ) ;
  assign n11479 = n11478 ^ n11477 ^ n7575 ;
  assign n11481 = n11480 ^ n11479 ^ n8749 ;
  assign n11482 = n9320 ^ n7365 ^ 1'b0 ;
  assign n11484 = n2140 ^ n1887 ^ n1285 ;
  assign n11485 = ~n505 & n11484 ;
  assign n11483 = n3000 & ~n4545 ;
  assign n11486 = n11485 ^ n11483 ^ 1'b0 ;
  assign n11487 = ( ~x114 & n1000 ) | ( ~x114 & n4366 ) | ( n1000 & n4366 ) ;
  assign n11488 = n5422 & n11487 ;
  assign n11489 = n3485 & n10089 ;
  assign n11490 = n10892 ^ n5326 ^ n5178 ;
  assign n11491 = ( n1282 & n3485 ) | ( n1282 & n3924 ) | ( n3485 & n3924 ) ;
  assign n11492 = ( n5951 & n9450 ) | ( n5951 & ~n11491 ) | ( n9450 & ~n11491 ) ;
  assign n11493 = n11490 | n11492 ;
  assign n11494 = n11489 & ~n11493 ;
  assign n11495 = ( n7338 & n11488 ) | ( n7338 & ~n11494 ) | ( n11488 & ~n11494 ) ;
  assign n11496 = n8740 ^ n3289 ^ n2297 ;
  assign n11497 = ~n319 & n1407 ;
  assign n11498 = n11497 ^ n2068 ^ 1'b0 ;
  assign n11499 = n11498 ^ n9932 ^ 1'b0 ;
  assign n11500 = ~n11496 & n11499 ;
  assign n11503 = n3668 ^ n3409 ^ n2069 ;
  assign n11504 = n11503 ^ n2244 ^ n885 ;
  assign n11505 = ( n2883 & n5618 ) | ( n2883 & n11504 ) | ( n5618 & n11504 ) ;
  assign n11501 = ~n1534 & n6534 ;
  assign n11502 = n11501 ^ n6480 ^ n541 ;
  assign n11506 = n11505 ^ n11502 ^ 1'b0 ;
  assign n11507 = n11500 & n11506 ;
  assign n11508 = ( n6668 & ~n7585 ) | ( n6668 & n8012 ) | ( ~n7585 & n8012 ) ;
  assign n11509 = n1165 & ~n8923 ;
  assign n11510 = n11508 & n11509 ;
  assign n11511 = n11510 ^ n1639 ^ n1257 ;
  assign n11512 = ( n2405 & n3689 ) | ( n2405 & n11511 ) | ( n3689 & n11511 ) ;
  assign n11514 = n8787 ^ n8399 ^ n1215 ;
  assign n11513 = ( n906 & n1263 ) | ( n906 & ~n4295 ) | ( n1263 & ~n4295 ) ;
  assign n11515 = n11514 ^ n11513 ^ n906 ;
  assign n11516 = n11515 ^ n2306 ^ 1'b0 ;
  assign n11517 = n11516 ^ n8085 ^ 1'b0 ;
  assign n11518 = n1437 & n2654 ;
  assign n11519 = ~n10771 & n11518 ;
  assign n11520 = ( n1987 & ~n6978 ) | ( n1987 & n8693 ) | ( ~n6978 & n8693 ) ;
  assign n11521 = ( ~n8597 & n11519 ) | ( ~n8597 & n11520 ) | ( n11519 & n11520 ) ;
  assign n11526 = n10191 ^ n2758 ^ 1'b0 ;
  assign n11522 = n2947 | n8368 ;
  assign n11523 = n5987 & ~n11522 ;
  assign n11524 = n11523 ^ n4401 ^ 1'b0 ;
  assign n11525 = n6464 | n11524 ;
  assign n11527 = n11526 ^ n11525 ^ n2297 ;
  assign n11528 = n8461 ^ n4202 ^ n475 ;
  assign n11529 = n11528 ^ n8129 ^ n6950 ;
  assign n11530 = n1632 & ~n4060 ;
  assign n11531 = n6547 & n11530 ;
  assign n11535 = n5307 & ~n8336 ;
  assign n11536 = ( ~n804 & n6736 ) | ( ~n804 & n11535 ) | ( n6736 & n11535 ) ;
  assign n11533 = n9951 ^ n1151 ^ 1'b0 ;
  assign n11534 = ~n138 & n11533 ;
  assign n11532 = n11090 ^ n5756 ^ n5352 ;
  assign n11537 = n11536 ^ n11534 ^ n11532 ;
  assign n11538 = n6123 ^ n3691 ^ n1264 ;
  assign n11539 = ( ~n4558 & n5809 ) | ( ~n4558 & n11538 ) | ( n5809 & n11538 ) ;
  assign n11540 = n9125 ^ n4281 ^ 1'b0 ;
  assign n11541 = ~n9537 & n11540 ;
  assign n11542 = ~n3542 & n6697 ;
  assign n11543 = n381 & n11542 ;
  assign n11544 = n11543 ^ n7867 ^ n1925 ;
  assign n11545 = n11544 ^ n5065 ^ n3179 ;
  assign n11546 = ( n7839 & n8414 ) | ( n7839 & n11545 ) | ( n8414 & n11545 ) ;
  assign n11547 = n10114 ^ n1170 ^ n941 ;
  assign n11548 = ~n992 & n1634 ;
  assign n11549 = n11548 ^ n3124 ^ 1'b0 ;
  assign n11550 = n2797 ^ n1037 ^ n243 ;
  assign n11551 = n11549 | n11550 ;
  assign n11552 = n5517 & ~n11551 ;
  assign n11553 = n4480 & ~n11552 ;
  assign n11554 = ~n11547 & n11553 ;
  assign n11555 = n11554 ^ n10307 ^ n143 ;
  assign n11556 = n11555 ^ x63 ^ 1'b0 ;
  assign n11557 = ( ~x93 & n193 ) | ( ~x93 & n3980 ) | ( n193 & n3980 ) ;
  assign n11558 = n9762 ^ n9506 ^ n7173 ;
  assign n11559 = n11558 ^ n4605 ^ n3697 ;
  assign n11560 = n11557 & n11559 ;
  assign n11561 = n2470 | n3182 ;
  assign n11562 = n4840 ^ n3954 ^ n511 ;
  assign n11563 = n11562 ^ n3518 ^ n2896 ;
  assign n11564 = n9010 & n11563 ;
  assign n11565 = ( n226 & n1184 ) | ( n226 & n5090 ) | ( n1184 & n5090 ) ;
  assign n11566 = ~n776 & n3832 ;
  assign n11567 = n11566 ^ n4559 ^ n2066 ;
  assign n11568 = ( ~n1005 & n11565 ) | ( ~n1005 & n11567 ) | ( n11565 & n11567 ) ;
  assign n11569 = n11568 ^ n9546 ^ n4017 ;
  assign n11570 = n3833 & n11569 ;
  assign n11571 = ~n11564 & n11570 ;
  assign n11572 = n5740 & ~n11571 ;
  assign n11573 = n1478 & n11572 ;
  assign n11574 = ( n4819 & n11561 ) | ( n4819 & n11573 ) | ( n11561 & n11573 ) ;
  assign n11578 = ( n1973 & n5229 ) | ( n1973 & n9272 ) | ( n5229 & n9272 ) ;
  assign n11575 = n6177 ^ n3691 ^ n1922 ;
  assign n11576 = ( ~n1449 & n3261 ) | ( ~n1449 & n3972 ) | ( n3261 & n3972 ) ;
  assign n11577 = ( n10554 & n11575 ) | ( n10554 & ~n11576 ) | ( n11575 & ~n11576 ) ;
  assign n11579 = n11578 ^ n11577 ^ n656 ;
  assign n11580 = ( n4364 & ~n5167 ) | ( n4364 & n9496 ) | ( ~n5167 & n9496 ) ;
  assign n11581 = n8789 ^ n4003 ^ n2256 ;
  assign n11582 = ( n905 & n5511 ) | ( n905 & n7203 ) | ( n5511 & n7203 ) ;
  assign n11584 = n1861 ^ n598 ^ n213 ;
  assign n11583 = n3327 & ~n10786 ;
  assign n11585 = n11584 ^ n11583 ^ n8704 ;
  assign n11586 = n7644 ^ n6843 ^ x112 ;
  assign n11587 = n8156 & ~n9827 ;
  assign n11588 = n1211 & n11587 ;
  assign n11589 = n1865 ^ n819 ^ n751 ;
  assign n11590 = n11589 ^ n2355 ^ n389 ;
  assign n11591 = n685 | n10878 ;
  assign n11592 = n11591 ^ n1588 ^ 1'b0 ;
  assign n11593 = n11592 ^ n9157 ^ n3753 ;
  assign n11594 = n6527 ^ n1644 ^ n648 ;
  assign n11595 = ( n364 & n4965 ) | ( n364 & n9679 ) | ( n4965 & n9679 ) ;
  assign n11596 = n11595 ^ n5649 ^ n4950 ;
  assign n11597 = ( ~n5368 & n11594 ) | ( ~n5368 & n11596 ) | ( n11594 & n11596 ) ;
  assign n11598 = n8174 & n11597 ;
  assign n11599 = n10356 ^ n9302 ^ n7152 ;
  assign n11600 = n1706 & ~n2891 ;
  assign n11601 = ~n5231 & n11600 ;
  assign n11604 = n302 & n4731 ;
  assign n11605 = ( n4285 & n10969 ) | ( n4285 & n11604 ) | ( n10969 & n11604 ) ;
  assign n11602 = n6054 ^ n5023 ^ 1'b0 ;
  assign n11603 = n7557 | n11602 ;
  assign n11606 = n11605 ^ n11603 ^ n2642 ;
  assign n11607 = ( n1977 & n11601 ) | ( n1977 & n11606 ) | ( n11601 & n11606 ) ;
  assign n11608 = n9276 ^ n591 ^ 1'b0 ;
  assign n11617 = ( n1350 & ~n1631 ) | ( n1350 & n1923 ) | ( ~n1631 & n1923 ) ;
  assign n11618 = n10933 ^ n4641 ^ n829 ;
  assign n11619 = ( n4435 & n11617 ) | ( n4435 & ~n11618 ) | ( n11617 & ~n11618 ) ;
  assign n11614 = ~n1973 & n3168 ;
  assign n11615 = n11614 ^ n426 ^ 1'b0 ;
  assign n11613 = ( n1652 & n8950 ) | ( n1652 & n11274 ) | ( n8950 & n11274 ) ;
  assign n11611 = n5763 ^ n3573 ^ n2114 ;
  assign n11612 = n11611 ^ n3757 ^ n1313 ;
  assign n11616 = n11615 ^ n11613 ^ n11612 ;
  assign n11620 = n11619 ^ n11616 ^ n2983 ;
  assign n11609 = ( ~n1201 & n4717 ) | ( ~n1201 & n6923 ) | ( n4717 & n6923 ) ;
  assign n11610 = n846 | n11609 ;
  assign n11621 = n11620 ^ n11610 ^ 1'b0 ;
  assign n11622 = n7079 ^ n6688 ^ n3716 ;
  assign n11623 = n4091 ^ n994 ^ n327 ;
  assign n11624 = n1777 & n11623 ;
  assign n11625 = n7145 | n11624 ;
  assign n11626 = n8970 | n11625 ;
  assign n11633 = ( ~n964 & n2331 ) | ( ~n964 & n3479 ) | ( n2331 & n3479 ) ;
  assign n11631 = n5903 ^ n355 ^ 1'b0 ;
  assign n11632 = n11631 ^ n4079 ^ n1994 ;
  assign n11634 = n11633 ^ n11632 ^ 1'b0 ;
  assign n11627 = ( n610 & ~n3349 ) | ( n610 & n3633 ) | ( ~n3349 & n3633 ) ;
  assign n11628 = n8570 ^ n5849 ^ n3447 ;
  assign n11629 = n11628 ^ n9589 ^ 1'b0 ;
  assign n11630 = n11627 | n11629 ;
  assign n11635 = n11634 ^ n11630 ^ n7264 ;
  assign n11636 = ( n2552 & n3843 ) | ( n2552 & n4824 ) | ( n3843 & n4824 ) ;
  assign n11637 = ~n11416 & n11636 ;
  assign n11647 = ( ~n1675 & n4078 ) | ( ~n1675 & n4921 ) | ( n4078 & n4921 ) ;
  assign n11648 = n11647 ^ n5954 ^ n2879 ;
  assign n11640 = n1662 ^ n1058 ^ n952 ;
  assign n11641 = n11640 ^ n1453 ^ n248 ;
  assign n11642 = n11641 ^ n10426 ^ 1'b0 ;
  assign n11643 = n9998 & n11642 ;
  assign n11644 = ~n4065 & n11643 ;
  assign n11645 = n11644 ^ n6158 ^ 1'b0 ;
  assign n11646 = n11645 ^ n2391 ^ 1'b0 ;
  assign n11638 = n6844 ^ n2079 ^ n1687 ;
  assign n11639 = n11638 ^ n2312 ^ n507 ;
  assign n11649 = n11648 ^ n11646 ^ n11639 ;
  assign n11656 = ( n988 & n4471 ) | ( n988 & ~n7034 ) | ( n4471 & ~n7034 ) ;
  assign n11650 = n1009 & n4382 ;
  assign n11651 = n9035 ^ n1896 ^ n198 ;
  assign n11652 = n11650 | n11651 ;
  assign n11653 = n11652 ^ n4471 ^ 1'b0 ;
  assign n11654 = ( ~n1425 & n3775 ) | ( ~n1425 & n11653 ) | ( n3775 & n11653 ) ;
  assign n11655 = n11654 ^ n4232 ^ 1'b0 ;
  assign n11657 = n11656 ^ n11655 ^ 1'b0 ;
  assign n11658 = n11657 ^ n7909 ^ n5008 ;
  assign n11659 = ( n3372 & n7602 ) | ( n3372 & ~n11658 ) | ( n7602 & ~n11658 ) ;
  assign n11662 = ( ~n935 & n2644 ) | ( ~n935 & n4662 ) | ( n2644 & n4662 ) ;
  assign n11661 = ( n1219 & ~n4203 ) | ( n1219 & n11508 ) | ( ~n4203 & n11508 ) ;
  assign n11663 = n11662 ^ n11661 ^ n3876 ;
  assign n11664 = n11663 ^ n4955 ^ n2891 ;
  assign n11660 = ~n1285 & n3066 ;
  assign n11665 = n11664 ^ n11660 ^ 1'b0 ;
  assign n11666 = n7164 ^ n2405 ^ n1849 ;
  assign n11667 = n11666 ^ n7422 ^ 1'b0 ;
  assign n11668 = n11667 ^ n11207 ^ n5125 ;
  assign n11671 = n3307 & n7885 ;
  assign n11672 = n11671 ^ n1009 ^ n161 ;
  assign n11670 = n4137 ^ n1057 ^ 1'b0 ;
  assign n11669 = n3283 ^ n2037 ^ n1518 ;
  assign n11673 = n11672 ^ n11670 ^ n11669 ;
  assign n11676 = n3409 ^ n452 ^ 1'b0 ;
  assign n11677 = n556 | n11676 ;
  assign n11675 = ~n730 & n869 ;
  assign n11678 = n11677 ^ n11675 ^ n9817 ;
  assign n11674 = n1883 & ~n4562 ;
  assign n11679 = n11678 ^ n11674 ^ n1660 ;
  assign n11680 = n1678 & n2895 ;
  assign n11681 = n11680 ^ n5189 ^ 1'b0 ;
  assign n11682 = n11681 ^ n3615 ^ n318 ;
  assign n11683 = n11682 ^ n9428 ^ n4586 ;
  assign n11685 = n9390 ^ n3758 ^ n2734 ;
  assign n11686 = ( n2801 & n3063 ) | ( n2801 & n11685 ) | ( n3063 & n11685 ) ;
  assign n11684 = n138 | n1105 ;
  assign n11687 = n11686 ^ n11684 ^ 1'b0 ;
  assign n11688 = x39 & ~n7794 ;
  assign n11689 = n11688 ^ n4568 ^ 1'b0 ;
  assign n11690 = ~n541 & n8068 ;
  assign n11691 = n11690 ^ n7446 ^ 1'b0 ;
  assign n11692 = n9886 | n11691 ;
  assign n11693 = n6062 | n11692 ;
  assign n11696 = ( n893 & n1217 ) | ( n893 & ~n10091 ) | ( n1217 & ~n10091 ) ;
  assign n11694 = ( n6294 & n8237 ) | ( n6294 & ~n8690 ) | ( n8237 & ~n8690 ) ;
  assign n11695 = ( n4195 & n7688 ) | ( n4195 & n11694 ) | ( n7688 & n11694 ) ;
  assign n11697 = n11696 ^ n11695 ^ n3357 ;
  assign n11704 = ~n6802 & n11019 ;
  assign n11705 = ( n2634 & ~n7975 ) | ( n2634 & n11704 ) | ( ~n7975 & n11704 ) ;
  assign n11699 = ( n2585 & ~n4331 ) | ( n2585 & n6987 ) | ( ~n4331 & n6987 ) ;
  assign n11700 = n868 & ~n11699 ;
  assign n11701 = ( n523 & n6382 ) | ( n523 & ~n7775 ) | ( n6382 & ~n7775 ) ;
  assign n11702 = ( n6065 & n11700 ) | ( n6065 & ~n11701 ) | ( n11700 & ~n11701 ) ;
  assign n11698 = n3699 & ~n5703 ;
  assign n11703 = n11702 ^ n11698 ^ 1'b0 ;
  assign n11706 = n11705 ^ n11703 ^ n612 ;
  assign n11707 = ( ~n382 & n964 ) | ( ~n382 & n1252 ) | ( n964 & n1252 ) ;
  assign n11708 = n6413 & n11707 ;
  assign n11709 = n11708 ^ n2828 ^ 1'b0 ;
  assign n11710 = ( n7599 & n11706 ) | ( n7599 & n11709 ) | ( n11706 & n11709 ) ;
  assign n11711 = ( n2589 & n7369 ) | ( n2589 & ~n10243 ) | ( n7369 & ~n10243 ) ;
  assign n11718 = n746 ^ n445 ^ 1'b0 ;
  assign n11719 = n11718 ^ n254 ^ 1'b0 ;
  assign n11720 = n2105 & n11719 ;
  assign n11717 = ( x125 & n363 ) | ( x125 & ~n8182 ) | ( n363 & ~n8182 ) ;
  assign n11712 = n4115 ^ n1656 ^ n289 ;
  assign n11713 = n5797 & n9046 ;
  assign n11714 = n11713 ^ n1865 ^ 1'b0 ;
  assign n11715 = ~n1766 & n11714 ;
  assign n11716 = ( n3070 & ~n11712 ) | ( n3070 & n11715 ) | ( ~n11712 & n11715 ) ;
  assign n11721 = n11720 ^ n11717 ^ n11716 ;
  assign n11722 = ( n739 & ~n3557 ) | ( n739 & n5207 ) | ( ~n3557 & n5207 ) ;
  assign n11724 = n3952 | n5451 ;
  assign n11725 = n11724 ^ n2883 ^ 1'b0 ;
  assign n11726 = n11725 ^ n5630 ^ n3656 ;
  assign n11723 = n1495 & ~n11164 ;
  assign n11727 = n11726 ^ n11723 ^ 1'b0 ;
  assign n11728 = ( ~n2630 & n9882 ) | ( ~n2630 & n11727 ) | ( n9882 & n11727 ) ;
  assign n11729 = n7629 | n11728 ;
  assign n11730 = n11722 | n11729 ;
  assign n11731 = ~n3943 & n6727 ;
  assign n11732 = n1705 & n11731 ;
  assign n11733 = n11732 ^ n3277 ^ 1'b0 ;
  assign n11734 = n4382 & ~n11733 ;
  assign n11735 = n9325 & n11734 ;
  assign n11736 = n3200 ^ n1265 ^ x92 ;
  assign n11737 = n11736 ^ n11292 ^ n3652 ;
  assign n11738 = n11737 ^ n6981 ^ n6344 ;
  assign n11739 = ( ~n162 & n11735 ) | ( ~n162 & n11738 ) | ( n11735 & n11738 ) ;
  assign n11740 = ~n1912 & n4345 ;
  assign n11741 = n1373 & n11740 ;
  assign n11742 = n11544 ^ n7195 ^ n1856 ;
  assign n11743 = n453 & n8716 ;
  assign n11744 = n11743 ^ n6095 ^ 1'b0 ;
  assign n11745 = n11742 & ~n11744 ;
  assign n11746 = n11745 ^ n6532 ^ 1'b0 ;
  assign n11747 = n11741 | n11746 ;
  assign n11748 = n3832 ^ n2554 ^ 1'b0 ;
  assign n11749 = n11748 ^ n4115 ^ n3122 ;
  assign n11750 = ( n873 & ~n2408 ) | ( n873 & n6227 ) | ( ~n2408 & n6227 ) ;
  assign n11751 = n11750 ^ n10137 ^ n3528 ;
  assign n11752 = ( ~n3921 & n10645 ) | ( ~n3921 & n11751 ) | ( n10645 & n11751 ) ;
  assign n11753 = n11752 ^ x34 ^ 1'b0 ;
  assign n11760 = ( n969 & ~n1163 ) | ( n969 & n2536 ) | ( ~n1163 & n2536 ) ;
  assign n11758 = n11132 ^ n1272 ^ n822 ;
  assign n11759 = ( ~n3989 & n6469 ) | ( ~n3989 & n11758 ) | ( n6469 & n11758 ) ;
  assign n11761 = n11760 ^ n11759 ^ n2232 ;
  assign n11756 = n3103 & ~n10394 ;
  assign n11754 = n3155 & n3580 ;
  assign n11755 = n6133 | n11754 ;
  assign n11757 = n11756 ^ n11755 ^ n1086 ;
  assign n11762 = n11761 ^ n11757 ^ n10422 ;
  assign n11763 = ( ~n1040 & n1504 ) | ( ~n1040 & n4445 ) | ( n1504 & n4445 ) ;
  assign n11764 = n10693 ^ n6642 ^ n2086 ;
  assign n11765 = ( n10390 & n11001 ) | ( n10390 & n11764 ) | ( n11001 & n11764 ) ;
  assign n11766 = n11765 ^ n8815 ^ n8017 ;
  assign n11767 = n11745 ^ n10518 ^ n4660 ;
  assign n11768 = n11767 ^ n8288 ^ n4236 ;
  assign n11769 = n11768 ^ n9266 ^ n5838 ;
  assign n11772 = ( n1369 & n1422 ) | ( n1369 & ~n7898 ) | ( n1422 & ~n7898 ) ;
  assign n11773 = ( ~n4076 & n4639 ) | ( ~n4076 & n11772 ) | ( n4639 & n11772 ) ;
  assign n11770 = n4541 ^ n877 ^ 1'b0 ;
  assign n11771 = n11770 ^ n10498 ^ n3760 ;
  assign n11774 = n11773 ^ n11771 ^ 1'b0 ;
  assign n11775 = ( ~n6046 & n11769 ) | ( ~n6046 & n11774 ) | ( n11769 & n11774 ) ;
  assign n11776 = ~n3398 & n9809 ;
  assign n11777 = ~n1057 & n11776 ;
  assign n11780 = ( n1339 & n1794 ) | ( n1339 & ~n4795 ) | ( n1794 & ~n4795 ) ;
  assign n11781 = ( ~n3604 & n4092 ) | ( ~n3604 & n7059 ) | ( n4092 & n7059 ) ;
  assign n11782 = ( n9266 & n11780 ) | ( n9266 & ~n11781 ) | ( n11780 & ~n11781 ) ;
  assign n11778 = ( ~n3435 & n3579 ) | ( ~n3435 & n6076 ) | ( n3579 & n6076 ) ;
  assign n11779 = n11778 ^ n4659 ^ n1243 ;
  assign n11783 = n11782 ^ n11779 ^ n5155 ;
  assign n11784 = n2220 ^ x55 ^ 1'b0 ;
  assign n11785 = ( n426 & ~n2292 ) | ( n426 & n11550 ) | ( ~n2292 & n11550 ) ;
  assign n11786 = n11785 ^ n7201 ^ n636 ;
  assign n11787 = ( ~n4085 & n5639 ) | ( ~n4085 & n11786 ) | ( n5639 & n11786 ) ;
  assign n11788 = ( n1572 & n11784 ) | ( n1572 & n11787 ) | ( n11784 & n11787 ) ;
  assign n11789 = ( n8006 & ~n10787 ) | ( n8006 & n10945 ) | ( ~n10787 & n10945 ) ;
  assign n11799 = n5979 ^ n3001 ^ n223 ;
  assign n11790 = n8422 ^ n3570 ^ n2744 ;
  assign n11791 = n11790 ^ n1251 ^ 1'b0 ;
  assign n11792 = n787 & ~n11791 ;
  assign n11793 = n11173 ^ n5134 ^ 1'b0 ;
  assign n11794 = n6528 & n11793 ;
  assign n11795 = ( n3683 & n7654 ) | ( n3683 & n11794 ) | ( n7654 & n11794 ) ;
  assign n11796 = ( n1001 & ~n2577 ) | ( n1001 & n2929 ) | ( ~n2577 & n2929 ) ;
  assign n11797 = n11796 ^ n10463 ^ n3361 ;
  assign n11798 = ( n11792 & n11795 ) | ( n11792 & n11797 ) | ( n11795 & n11797 ) ;
  assign n11800 = n11799 ^ n11798 ^ n337 ;
  assign n11801 = ( n1151 & n5207 ) | ( n1151 & ~n11093 ) | ( n5207 & ~n11093 ) ;
  assign n11802 = n11801 ^ n4173 ^ 1'b0 ;
  assign n11803 = ( n2012 & n10268 ) | ( n2012 & ~n11802 ) | ( n10268 & ~n11802 ) ;
  assign n11804 = ( n5713 & ~n6150 ) | ( n5713 & n11803 ) | ( ~n6150 & n11803 ) ;
  assign n11805 = ( n591 & ~n4756 ) | ( n591 & n10213 ) | ( ~n4756 & n10213 ) ;
  assign n11806 = ( n4458 & n4925 ) | ( n4458 & n7597 ) | ( n4925 & n7597 ) ;
  assign n11807 = ( n638 & n4913 ) | ( n638 & ~n10396 ) | ( n4913 & ~n10396 ) ;
  assign n11808 = n11807 ^ n6590 ^ n2086 ;
  assign n11809 = ( n3365 & n11806 ) | ( n3365 & ~n11808 ) | ( n11806 & ~n11808 ) ;
  assign n11810 = n8923 ^ n6818 ^ 1'b0 ;
  assign n11811 = n11584 ^ n7174 ^ n4400 ;
  assign n11812 = ( n11809 & ~n11810 ) | ( n11809 & n11811 ) | ( ~n11810 & n11811 ) ;
  assign n11813 = n8296 ^ n8051 ^ n2297 ;
  assign n11814 = ( x9 & ~n1183 ) | ( x9 & n11813 ) | ( ~n1183 & n11813 ) ;
  assign n11815 = n11814 ^ n5979 ^ n3122 ;
  assign n11816 = ( n892 & ~n9736 ) | ( n892 & n11815 ) | ( ~n9736 & n11815 ) ;
  assign n11825 = n2679 ^ n787 ^ 1'b0 ;
  assign n11823 = n5513 ^ n3742 ^ n2545 ;
  assign n11824 = n11823 ^ n936 ^ n783 ;
  assign n11826 = n11825 ^ n11824 ^ n1122 ;
  assign n11820 = ( n1141 & ~n1964 ) | ( n1141 & n3911 ) | ( ~n1964 & n3911 ) ;
  assign n11821 = n8568 ^ n900 ^ 1'b0 ;
  assign n11822 = ~n11820 & n11821 ;
  assign n11827 = n11826 ^ n11822 ^ n1907 ;
  assign n11828 = ~n9717 & n10802 ;
  assign n11829 = n11828 ^ n9893 ^ 1'b0 ;
  assign n11830 = ( n3695 & n11827 ) | ( n3695 & n11829 ) | ( n11827 & n11829 ) ;
  assign n11817 = n3405 & n11604 ;
  assign n11818 = n3684 & ~n11817 ;
  assign n11819 = ~n3484 & n11818 ;
  assign n11831 = n11830 ^ n11819 ^ n489 ;
  assign n11832 = n5960 ^ n2445 ^ n1649 ;
  assign n11833 = n11832 ^ n10621 ^ n5082 ;
  assign n11834 = n1282 & ~n4473 ;
  assign n11835 = n2205 | n2716 ;
  assign n11836 = n1469 & ~n11835 ;
  assign n11837 = n11834 & n11836 ;
  assign n11838 = n8626 ^ n5935 ^ n3888 ;
  assign n11839 = n8920 ^ n7505 ^ n5485 ;
  assign n11840 = ( ~n966 & n5196 ) | ( ~n966 & n10507 ) | ( n5196 & n10507 ) ;
  assign n11841 = n11840 ^ n8984 ^ 1'b0 ;
  assign n11842 = n11778 & n11841 ;
  assign n11843 = n1303 | n2494 ;
  assign n11844 = n916 & ~n11843 ;
  assign n11845 = n4921 & n9005 ;
  assign n11846 = n10502 | n11845 ;
  assign n11847 = n11844 & ~n11846 ;
  assign n11848 = n10598 ^ n1458 ^ n487 ;
  assign n11849 = ( n8773 & n11742 ) | ( n8773 & ~n11848 ) | ( n11742 & ~n11848 ) ;
  assign n11850 = ( n4430 & n7103 ) | ( n4430 & n11372 ) | ( n7103 & n11372 ) ;
  assign n11851 = ~n1165 & n11850 ;
  assign n11852 = ( n1375 & n4306 ) | ( n1375 & ~n4351 ) | ( n4306 & ~n4351 ) ;
  assign n11853 = n11852 ^ n4791 ^ n1144 ;
  assign n11854 = n11853 ^ n10746 ^ n4508 ;
  assign n11860 = n4935 & ~n11055 ;
  assign n11861 = n3088 & n11860 ;
  assign n11855 = ( n1879 & ~n2128 ) | ( n1879 & n4731 ) | ( ~n2128 & n4731 ) ;
  assign n11856 = ( n6775 & n7015 ) | ( n6775 & n11855 ) | ( n7015 & n11855 ) ;
  assign n11857 = n11856 ^ n10838 ^ n8130 ;
  assign n11858 = n11857 ^ n1633 ^ x27 ;
  assign n11859 = ~n10957 & n11858 ;
  assign n11862 = n11861 ^ n11859 ^ 1'b0 ;
  assign n11863 = n11112 ^ n5328 ^ n4414 ;
  assign n11864 = ( ~n2472 & n2826 ) | ( ~n2472 & n11863 ) | ( n2826 & n11863 ) ;
  assign n11865 = ( n5727 & n7029 ) | ( n5727 & ~n11864 ) | ( n7029 & ~n11864 ) ;
  assign n11866 = n11862 & ~n11865 ;
  assign n11867 = ~n7963 & n11866 ;
  assign n11870 = n305 & ~n6280 ;
  assign n11871 = ~n570 & n11870 ;
  assign n11872 = ( n495 & n678 ) | ( n495 & ~n3546 ) | ( n678 & ~n3546 ) ;
  assign n11873 = n11872 ^ n5002 ^ n3352 ;
  assign n11874 = ( n3580 & n11871 ) | ( n3580 & n11873 ) | ( n11871 & n11873 ) ;
  assign n11868 = n5342 | n5519 ;
  assign n11869 = n5805 | n11868 ;
  assign n11875 = n11874 ^ n11869 ^ n2625 ;
  assign n11876 = n11767 ^ n9579 ^ n5573 ;
  assign n11877 = n4331 ^ n2613 ^ n2018 ;
  assign n11878 = n4127 & ~n11877 ;
  assign n11879 = n4058 & n11878 ;
  assign n11880 = n4104 & ~n11879 ;
  assign n11881 = n4590 ^ n1126 ^ 1'b0 ;
  assign n11882 = ( n4430 & n11880 ) | ( n4430 & ~n11881 ) | ( n11880 & ~n11881 ) ;
  assign n11883 = ( n2737 & ~n8716 ) | ( n2737 & n8784 ) | ( ~n8716 & n8784 ) ;
  assign n11884 = n11883 ^ n4889 ^ 1'b0 ;
  assign n11885 = n3359 ^ n1653 ^ n614 ;
  assign n11886 = n750 & n11885 ;
  assign n11887 = ~n11884 & n11886 ;
  assign n11888 = n9259 ^ n5830 ^ 1'b0 ;
  assign n11889 = n9507 ^ n635 ^ 1'b0 ;
  assign n11890 = n10560 ^ n8503 ^ n7342 ;
  assign n11897 = ~n212 & n2105 ;
  assign n11898 = ~n1229 & n11897 ;
  assign n11891 = n8238 ^ n3313 ^ n2291 ;
  assign n11892 = ( n1460 & n2816 ) | ( n1460 & ~n7847 ) | ( n2816 & ~n7847 ) ;
  assign n11893 = n11892 ^ n10519 ^ 1'b0 ;
  assign n11894 = n1699 & n11893 ;
  assign n11895 = n11891 & ~n11894 ;
  assign n11896 = n11895 ^ n3733 ^ n1289 ;
  assign n11899 = n11898 ^ n11896 ^ n11429 ;
  assign n11905 = ( n1234 & ~n3345 ) | ( n1234 & n4603 ) | ( ~n3345 & n4603 ) ;
  assign n11900 = n6075 ^ n2767 ^ n512 ;
  assign n11901 = n4646 ^ n3281 ^ 1'b0 ;
  assign n11902 = ( ~n3356 & n8839 ) | ( ~n3356 & n11901 ) | ( n8839 & n11901 ) ;
  assign n11903 = n4208 | n11902 ;
  assign n11904 = n11900 & ~n11903 ;
  assign n11906 = n11905 ^ n11904 ^ 1'b0 ;
  assign n11907 = n3205 & n4645 ;
  assign n11908 = n11907 ^ n1460 ^ 1'b0 ;
  assign n11909 = ~n1063 & n5710 ;
  assign n11910 = n11909 ^ n6228 ^ 1'b0 ;
  assign n11911 = n2234 & ~n4057 ;
  assign n11912 = ( n325 & n1346 ) | ( n325 & n11911 ) | ( n1346 & n11911 ) ;
  assign n11913 = ( n3220 & n11910 ) | ( n3220 & ~n11912 ) | ( n11910 & ~n11912 ) ;
  assign n11914 = n4488 & n10198 ;
  assign n11915 = ( ~n3453 & n10739 ) | ( ~n3453 & n11914 ) | ( n10739 & n11914 ) ;
  assign n11916 = n10261 ^ n6096 ^ n5975 ;
  assign n11917 = n11216 & n11916 ;
  assign n11918 = ~n6169 & n11917 ;
  assign n11919 = n11918 ^ n6962 ^ n5329 ;
  assign n11920 = ( n510 & n2272 ) | ( n510 & ~n4560 ) | ( n2272 & ~n4560 ) ;
  assign n11921 = ( ~n8811 & n9773 ) | ( ~n8811 & n11920 ) | ( n9773 & n11920 ) ;
  assign n11922 = n2727 | n11921 ;
  assign n11923 = n8753 & ~n11922 ;
  assign n11924 = n11923 ^ n11413 ^ 1'b0 ;
  assign n11925 = n7465 ^ n6026 ^ n1277 ;
  assign n11926 = n3045 | n11925 ;
  assign n11927 = n11926 ^ n4538 ^ 1'b0 ;
  assign n11928 = n11927 ^ n11411 ^ n9522 ;
  assign n11929 = n11928 ^ n4497 ^ n1733 ;
  assign n11930 = n205 | n6673 ;
  assign n11931 = n11929 & ~n11930 ;
  assign n11932 = n3423 ^ n2987 ^ 1'b0 ;
  assign n11933 = n10922 & ~n11932 ;
  assign n11934 = n11933 ^ n9509 ^ 1'b0 ;
  assign n11935 = ( n3582 & n3619 ) | ( n3582 & n3989 ) | ( n3619 & n3989 ) ;
  assign n11936 = n11935 ^ n2750 ^ n2313 ;
  assign n11937 = ( ~n1518 & n6139 ) | ( ~n1518 & n6184 ) | ( n6139 & n6184 ) ;
  assign n11938 = n11936 & n11937 ;
  assign n11939 = ~n8420 & n11938 ;
  assign n11940 = ( n5866 & n9134 ) | ( n5866 & n11939 ) | ( n9134 & n11939 ) ;
  assign n11941 = n3666 | n11940 ;
  assign n11942 = n11941 ^ n10698 ^ n226 ;
  assign n11943 = n2152 ^ n498 ^ 1'b0 ;
  assign n11944 = n2826 & n11943 ;
  assign n11945 = ( n3371 & ~n6323 ) | ( n3371 & n11944 ) | ( ~n6323 & n11944 ) ;
  assign n11946 = n11945 ^ n7232 ^ n3233 ;
  assign n11947 = n11946 ^ n9374 ^ n3828 ;
  assign n11949 = ( n697 & ~n763 ) | ( n697 & n4560 ) | ( ~n763 & n4560 ) ;
  assign n11948 = n11662 ^ n4418 ^ n3496 ;
  assign n11950 = n11949 ^ n11948 ^ n2151 ;
  assign n11951 = n4902 ^ n1777 ^ n1740 ;
  assign n11952 = ( n5953 & n10008 ) | ( n5953 & n11951 ) | ( n10008 & n11951 ) ;
  assign n11953 = ( ~n3833 & n11092 ) | ( ~n3833 & n11952 ) | ( n11092 & n11952 ) ;
  assign n11954 = n3700 ^ n3176 ^ n2345 ;
  assign n11955 = ( n3096 & n4626 ) | ( n3096 & ~n11954 ) | ( n4626 & ~n11954 ) ;
  assign n11971 = n10126 ^ n8703 ^ n7852 ;
  assign n11956 = ( n1224 & ~n5446 ) | ( n1224 & n8184 ) | ( ~n5446 & n8184 ) ;
  assign n11957 = ~n1470 & n11956 ;
  assign n11958 = ~n645 & n11957 ;
  assign n11959 = n9336 ^ n7486 ^ x121 ;
  assign n11960 = n3765 | n11959 ;
  assign n11961 = n11958 & ~n11960 ;
  assign n11962 = n4486 ^ n465 ^ 1'b0 ;
  assign n11963 = n5489 & ~n11962 ;
  assign n11964 = ~n1927 & n11963 ;
  assign n11965 = n2130 & n11964 ;
  assign n11966 = x59 & ~n3868 ;
  assign n11967 = n11966 ^ n459 ^ 1'b0 ;
  assign n11968 = ( ~n2138 & n3096 ) | ( ~n2138 & n11967 ) | ( n3096 & n11967 ) ;
  assign n11969 = ( n7558 & ~n11965 ) | ( n7558 & n11968 ) | ( ~n11965 & n11968 ) ;
  assign n11970 = ( n439 & ~n11961 ) | ( n439 & n11969 ) | ( ~n11961 & n11969 ) ;
  assign n11972 = n11971 ^ n11970 ^ n4075 ;
  assign n11973 = n8406 ^ n3536 ^ n2378 ;
  assign n11974 = ( n4253 & ~n10572 ) | ( n4253 & n11973 ) | ( ~n10572 & n11973 ) ;
  assign n11975 = ( n724 & n1435 ) | ( n724 & ~n4646 ) | ( n1435 & ~n4646 ) ;
  assign n11976 = ~n3375 & n7671 ;
  assign n11977 = n11975 & n11976 ;
  assign n11987 = ( n1914 & n4031 ) | ( n1914 & n9891 ) | ( n4031 & n9891 ) ;
  assign n11983 = n10472 ^ n7184 ^ 1'b0 ;
  assign n11984 = n1580 & ~n11983 ;
  assign n11985 = n11984 ^ n10904 ^ n7116 ;
  assign n11986 = ( n4121 & n4211 ) | ( n4121 & n11985 ) | ( n4211 & n11985 ) ;
  assign n11981 = n11491 ^ n2610 ^ 1'b0 ;
  assign n11978 = n3829 ^ x91 ^ 1'b0 ;
  assign n11979 = ~n9514 & n11978 ;
  assign n11980 = n11979 ^ n3962 ^ n846 ;
  assign n11982 = n11981 ^ n11980 ^ n2350 ;
  assign n11988 = n11987 ^ n11986 ^ n11982 ;
  assign n11989 = ( ~n707 & n879 ) | ( ~n707 & n4550 ) | ( n879 & n4550 ) ;
  assign n11990 = ( n2890 & ~n8683 ) | ( n2890 & n9395 ) | ( ~n8683 & n9395 ) ;
  assign n11991 = n11990 ^ n4078 ^ 1'b0 ;
  assign n11992 = n7554 & n11991 ;
  assign n11993 = n898 & n4610 ;
  assign n11994 = ~n577 & n11993 ;
  assign n11995 = n11994 ^ n7394 ^ 1'b0 ;
  assign n11996 = ( ~n1591 & n11992 ) | ( ~n1591 & n11995 ) | ( n11992 & n11995 ) ;
  assign n12007 = n7335 ^ n1189 ^ n1084 ;
  assign n11997 = ( ~n3597 & n6471 ) | ( ~n3597 & n7685 ) | ( n6471 & n7685 ) ;
  assign n11998 = n11997 ^ n11832 ^ n2677 ;
  assign n11999 = ( n5734 & n11402 ) | ( n5734 & n11998 ) | ( n11402 & n11998 ) ;
  assign n12000 = n1636 ^ n159 ^ 1'b0 ;
  assign n12002 = ( n3531 & n5031 ) | ( n3531 & ~n9400 ) | ( n5031 & ~n9400 ) ;
  assign n12001 = n6427 ^ n4685 ^ 1'b0 ;
  assign n12003 = n12002 ^ n12001 ^ n2721 ;
  assign n12004 = ~n12000 & n12003 ;
  assign n12005 = n12004 ^ n2435 ^ 1'b0 ;
  assign n12006 = n11999 & ~n12005 ;
  assign n12008 = n12007 ^ n12006 ^ 1'b0 ;
  assign n12009 = ( n3442 & n8340 ) | ( n3442 & ~n10875 ) | ( n8340 & ~n10875 ) ;
  assign n12010 = ( n2663 & ~n8708 ) | ( n2663 & n8921 ) | ( ~n8708 & n8921 ) ;
  assign n12011 = n484 ^ n270 ^ 1'b0 ;
  assign n12012 = n4384 ^ n4011 ^ n1695 ;
  assign n12013 = ( n11814 & n12011 ) | ( n11814 & ~n12012 ) | ( n12011 & ~n12012 ) ;
  assign n12014 = ( ~n4018 & n5726 ) | ( ~n4018 & n12013 ) | ( n5726 & n12013 ) ;
  assign n12015 = n2023 & ~n4882 ;
  assign n12016 = n12015 ^ n7472 ^ 1'b0 ;
  assign n12017 = n3691 & n5166 ;
  assign n12018 = n147 & n1583 ;
  assign n12019 = n12018 ^ n9797 ^ n4358 ;
  assign n12020 = n12017 & ~n12019 ;
  assign n12021 = ~n12016 & n12020 ;
  assign n12022 = n1969 ^ n1496 ^ n1168 ;
  assign n12023 = n5100 & n12022 ;
  assign n12024 = n12023 ^ n5422 ^ n677 ;
  assign n12031 = ( n2437 & n4508 ) | ( n2437 & ~n8056 ) | ( n4508 & ~n8056 ) ;
  assign n12025 = n5825 ^ n732 ^ 1'b0 ;
  assign n12026 = n12025 ^ n3665 ^ n1695 ;
  assign n12027 = ( n3667 & n6792 ) | ( n3667 & ~n12026 ) | ( n6792 & ~n12026 ) ;
  assign n12028 = n1689 ^ n1521 ^ 1'b0 ;
  assign n12029 = ~n12027 & n12028 ;
  assign n12030 = n12029 ^ n3062 ^ 1'b0 ;
  assign n12032 = n12031 ^ n12030 ^ n8098 ;
  assign n12033 = n1919 & ~n3453 ;
  assign n12034 = n3732 & ~n12033 ;
  assign n12035 = n6513 & n6520 ;
  assign n12036 = ~n12034 & n12035 ;
  assign n12037 = n11213 ^ n9379 ^ 1'b0 ;
  assign n12038 = n12036 | n12037 ;
  assign n12039 = ( n2561 & n9544 ) | ( n2561 & n10894 ) | ( n9544 & n10894 ) ;
  assign n12040 = x3 & n12039 ;
  assign n12041 = ( n10971 & n11850 ) | ( n10971 & ~n12040 ) | ( n11850 & ~n12040 ) ;
  assign n12042 = ~n1889 & n4991 ;
  assign n12043 = n2962 & ~n3705 ;
  assign n12044 = n10686 ^ n8436 ^ n1088 ;
  assign n12045 = ~n4979 & n12044 ;
  assign n12046 = ~n6540 & n12045 ;
  assign n12051 = ( n1217 & ~n3599 ) | ( n1217 & n4770 ) | ( ~n3599 & n4770 ) ;
  assign n12052 = n12051 ^ n1194 ^ n1191 ;
  assign n12049 = ( n1576 & ~n2296 ) | ( n1576 & n9320 ) | ( ~n2296 & n9320 ) ;
  assign n12050 = ( n4942 & n10161 ) | ( n4942 & ~n12049 ) | ( n10161 & ~n12049 ) ;
  assign n12047 = n1271 & n1906 ;
  assign n12048 = n3870 & n12047 ;
  assign n12053 = n12052 ^ n12050 ^ n12048 ;
  assign n12054 = n2758 ^ n1413 ^ 1'b0 ;
  assign n12055 = ( n391 & n9400 ) | ( n391 & n12054 ) | ( n9400 & n12054 ) ;
  assign n12056 = ( n8670 & n12053 ) | ( n8670 & n12055 ) | ( n12053 & n12055 ) ;
  assign n12057 = n12056 ^ n9686 ^ n2224 ;
  assign n12058 = n5082 ^ n1322 ^ n722 ;
  assign n12059 = ( ~n1474 & n2604 ) | ( ~n1474 & n3458 ) | ( n2604 & n3458 ) ;
  assign n12060 = ( x87 & n775 ) | ( x87 & n12059 ) | ( n775 & n12059 ) ;
  assign n12061 = n6662 ^ n3011 ^ n1588 ;
  assign n12062 = ( n12058 & n12060 ) | ( n12058 & ~n12061 ) | ( n12060 & ~n12061 ) ;
  assign n12063 = n3098 ^ n1672 ^ 1'b0 ;
  assign n12064 = ( n1679 & n6980 ) | ( n1679 & n9977 ) | ( n6980 & n9977 ) ;
  assign n12065 = n12064 ^ n10770 ^ 1'b0 ;
  assign n12066 = ~n12063 & n12065 ;
  assign n12067 = n6562 ^ n1712 ^ 1'b0 ;
  assign n12068 = ~n3441 & n12067 ;
  assign n12069 = ( n1980 & ~n11207 ) | ( n1980 & n12068 ) | ( ~n11207 & n12068 ) ;
  assign n12070 = n4810 & n8402 ;
  assign n12071 = n12070 ^ n2691 ^ n1526 ;
  assign n12072 = n4409 ^ n3377 ^ n1980 ;
  assign n12073 = n7810 ^ n2739 ^ 1'b0 ;
  assign n12075 = ( ~n1395 & n5332 ) | ( ~n1395 & n6614 ) | ( n5332 & n6614 ) ;
  assign n12076 = ( n2651 & n5340 ) | ( n2651 & n12075 ) | ( n5340 & n12075 ) ;
  assign n12074 = ( n5366 & n8186 ) | ( n5366 & ~n9332 ) | ( n8186 & ~n9332 ) ;
  assign n12077 = n12076 ^ n12074 ^ n7614 ;
  assign n12081 = n6188 & n8337 ;
  assign n12082 = n12081 ^ n8993 ^ 1'b0 ;
  assign n12078 = ~n6291 & n6393 ;
  assign n12079 = n7940 & n12078 ;
  assign n12080 = n4324 | n12079 ;
  assign n12083 = n12082 ^ n12080 ^ 1'b0 ;
  assign n12087 = n1767 ^ n918 ^ n284 ;
  assign n12084 = n5270 ^ n2821 ^ n665 ;
  assign n12085 = n12084 ^ n1772 ^ n1254 ;
  assign n12086 = n12085 ^ n6794 ^ n4921 ;
  assign n12088 = n12087 ^ n12086 ^ n1062 ;
  assign n12089 = n12088 ^ n2021 ^ 1'b0 ;
  assign n12090 = n12083 & ~n12089 ;
  assign n12091 = n7049 ^ n2193 ^ n541 ;
  assign n12092 = n12091 ^ n8422 ^ n8309 ;
  assign n12095 = ~n527 & n3616 ;
  assign n12093 = n2397 ^ n1686 ^ n1184 ;
  assign n12094 = n12093 ^ n6189 ^ n1966 ;
  assign n12096 = n12095 ^ n12094 ^ n8963 ;
  assign n12097 = ( ~n11970 & n12092 ) | ( ~n11970 & n12096 ) | ( n12092 & n12096 ) ;
  assign n12098 = ( ~n1919 & n5301 ) | ( ~n1919 & n11601 ) | ( n5301 & n11601 ) ;
  assign n12099 = n10532 | n12098 ;
  assign n12100 = n4451 | n12099 ;
  assign n12101 = ( n657 & n2902 ) | ( n657 & n4895 ) | ( n2902 & n4895 ) ;
  assign n12102 = n7045 ^ n1922 ^ n556 ;
  assign n12103 = ( ~n2468 & n6486 ) | ( ~n2468 & n12102 ) | ( n6486 & n12102 ) ;
  assign n12104 = ( ~n9527 & n12101 ) | ( ~n9527 & n12103 ) | ( n12101 & n12103 ) ;
  assign n12107 = n3084 ^ n972 ^ 1'b0 ;
  assign n12105 = n9879 ^ n5705 ^ n5601 ;
  assign n12106 = ~n1189 & n12105 ;
  assign n12108 = n12107 ^ n12106 ^ n8020 ;
  assign n12121 = ( n822 & n2220 ) | ( n822 & ~n4972 ) | ( n2220 & ~n4972 ) ;
  assign n12119 = ~n7678 & n11450 ;
  assign n12118 = n11823 ^ n1713 ^ x97 ;
  assign n12120 = n12119 ^ n12118 ^ n6907 ;
  assign n12109 = n3799 ^ n668 ^ 1'b0 ;
  assign n12110 = n766 & n12109 ;
  assign n12111 = n1893 & n5964 ;
  assign n12112 = n12111 ^ n2609 ^ 1'b0 ;
  assign n12113 = ( n1428 & n8035 ) | ( n1428 & n10394 ) | ( n8035 & n10394 ) ;
  assign n12114 = n12113 ^ n4403 ^ n631 ;
  assign n12115 = ( n1249 & ~n12112 ) | ( n1249 & n12114 ) | ( ~n12112 & n12114 ) ;
  assign n12116 = ( n7424 & ~n10790 ) | ( n7424 & n12115 ) | ( ~n10790 & n12115 ) ;
  assign n12117 = ( ~n7117 & n12110 ) | ( ~n7117 & n12116 ) | ( n12110 & n12116 ) ;
  assign n12122 = n12121 ^ n12120 ^ n12117 ;
  assign n12123 = n6386 ^ n3067 ^ n2174 ;
  assign n12124 = n12123 ^ n10429 ^ n7058 ;
  assign n12126 = ( x99 & n4966 ) | ( x99 & n7103 ) | ( n4966 & n7103 ) ;
  assign n12127 = n12126 ^ n1690 ^ 1'b0 ;
  assign n12128 = n511 & n12127 ;
  assign n12125 = ( n985 & n4006 ) | ( n985 & ~n5619 ) | ( n4006 & ~n5619 ) ;
  assign n12129 = n12128 ^ n12125 ^ n5893 ;
  assign n12130 = n7495 ^ n6173 ^ 1'b0 ;
  assign n12131 = x86 & ~n12130 ;
  assign n12132 = n816 | n5533 ;
  assign n12133 = n12132 ^ n11855 ^ 1'b0 ;
  assign n12134 = n12133 ^ n8041 ^ n5044 ;
  assign n12135 = n2228 & ~n12134 ;
  assign n12136 = n1687 | n4710 ;
  assign n12137 = n4644 | n12136 ;
  assign n12138 = n5963 ^ n1384 ^ 1'b0 ;
  assign n12139 = ( n7773 & n10009 ) | ( n7773 & ~n12138 ) | ( n10009 & ~n12138 ) ;
  assign n12140 = ( n4832 & n12137 ) | ( n4832 & n12139 ) | ( n12137 & n12139 ) ;
  assign n12141 = n6640 ^ n5583 ^ n3424 ;
  assign n12142 = n11601 ^ n3789 ^ 1'b0 ;
  assign n12143 = n12141 & n12142 ;
  assign n12144 = ( ~n1636 & n8111 ) | ( ~n1636 & n12143 ) | ( n8111 & n12143 ) ;
  assign n12145 = n6223 ^ n1701 ^ 1'b0 ;
  assign n12146 = ( n1544 & ~n2241 ) | ( n1544 & n5231 ) | ( ~n2241 & n5231 ) ;
  assign n12147 = n12146 ^ n4744 ^ 1'b0 ;
  assign n12148 = n12145 & n12147 ;
  assign n12149 = n3596 ^ n2336 ^ n209 ;
  assign n12150 = ~n5785 & n12149 ;
  assign n12151 = ~n381 & n12150 ;
  assign n12152 = ( n3406 & n12148 ) | ( n3406 & n12151 ) | ( n12148 & n12151 ) ;
  assign n12153 = ( ~n9566 & n11796 ) | ( ~n9566 & n12152 ) | ( n11796 & n12152 ) ;
  assign n12154 = n4884 & ~n12153 ;
  assign n12160 = n9371 ^ x60 ^ x36 ;
  assign n12159 = ( ~n4083 & n7257 ) | ( ~n4083 & n7476 ) | ( n7257 & n7476 ) ;
  assign n12157 = ( n321 & ~n593 ) | ( n321 & n1050 ) | ( ~n593 & n1050 ) ;
  assign n12155 = n4000 & n6413 ;
  assign n12156 = ~n6976 & n12155 ;
  assign n12158 = n12157 ^ n12156 ^ n10280 ;
  assign n12161 = n12160 ^ n12159 ^ n12158 ;
  assign n12163 = n1778 ^ n1667 ^ x18 ;
  assign n12164 = n12163 ^ n2375 ^ n1193 ;
  assign n12162 = n2280 ^ n1440 ^ n1272 ;
  assign n12165 = n12164 ^ n12162 ^ n8047 ;
  assign n12166 = ~n6363 & n11173 ;
  assign n12167 = n6079 ^ n1235 ^ n495 ;
  assign n12172 = n9058 | n9767 ;
  assign n12168 = ( ~n2494 & n4924 ) | ( ~n2494 & n5162 ) | ( n4924 & n5162 ) ;
  assign n12169 = ~n7513 & n12168 ;
  assign n12170 = n12169 ^ n4238 ^ 1'b0 ;
  assign n12171 = ( ~n424 & n6159 ) | ( ~n424 & n12170 ) | ( n6159 & n12170 ) ;
  assign n12173 = n12172 ^ n12171 ^ n8428 ;
  assign n12174 = n12173 ^ n5147 ^ n4828 ;
  assign n12175 = ( ~n6706 & n12167 ) | ( ~n6706 & n12174 ) | ( n12167 & n12174 ) ;
  assign n12176 = ( ~n4447 & n12166 ) | ( ~n4447 & n12175 ) | ( n12166 & n12175 ) ;
  assign n12177 = ( ~n1456 & n3983 ) | ( ~n1456 & n5905 ) | ( n3983 & n5905 ) ;
  assign n12178 = ( n947 & n10452 ) | ( n947 & n12177 ) | ( n10452 & n12177 ) ;
  assign n12179 = n10852 | n12178 ;
  assign n12180 = ( ~n988 & n1437 ) | ( ~n988 & n7011 ) | ( n1437 & n7011 ) ;
  assign n12181 = ( n5281 & n7053 ) | ( n5281 & n12180 ) | ( n7053 & n12180 ) ;
  assign n12182 = ( n8460 & ~n10891 ) | ( n8460 & n12181 ) | ( ~n10891 & n12181 ) ;
  assign n12183 = n7511 & n8254 ;
  assign n12184 = ( ~n4532 & n4987 ) | ( ~n4532 & n9257 ) | ( n4987 & n9257 ) ;
  assign n12185 = n6636 ^ n1175 ^ n929 ;
  assign n12186 = n333 | n1326 ;
  assign n12187 = n12186 ^ n2716 ^ 1'b0 ;
  assign n12188 = n1110 & ~n5056 ;
  assign n12189 = ( n2376 & n12187 ) | ( n2376 & n12188 ) | ( n12187 & n12188 ) ;
  assign n12190 = ( ~n12094 & n12185 ) | ( ~n12094 & n12189 ) | ( n12185 & n12189 ) ;
  assign n12196 = n497 & ~n9750 ;
  assign n12191 = ( ~n1365 & n4595 ) | ( ~n1365 & n8233 ) | ( n4595 & n8233 ) ;
  assign n12192 = n12191 ^ n3791 ^ n3581 ;
  assign n12193 = ( n11330 & ~n11822 ) | ( n11330 & n12192 ) | ( ~n11822 & n12192 ) ;
  assign n12194 = n12193 ^ n2419 ^ 1'b0 ;
  assign n12195 = ~n1324 & n12194 ;
  assign n12197 = n12196 ^ n12195 ^ n3205 ;
  assign n12198 = n404 | n6570 ;
  assign n12199 = n12198 ^ n2470 ^ n503 ;
  assign n12200 = ~n2698 & n11066 ;
  assign n12201 = n12200 ^ n292 ^ 1'b0 ;
  assign n12202 = ~n11466 & n12201 ;
  assign n12203 = n11970 ^ n6915 ^ 1'b0 ;
  assign n12204 = n6928 ^ n5495 ^ n1545 ;
  assign n12205 = n1056 & n12204 ;
  assign n12206 = n12205 ^ n10410 ^ x7 ;
  assign n12207 = ( ~n2073 & n2511 ) | ( ~n2073 & n12206 ) | ( n2511 & n12206 ) ;
  assign n12208 = ( n820 & n2820 ) | ( n820 & ~n5018 ) | ( n2820 & ~n5018 ) ;
  assign n12209 = n12208 ^ n2886 ^ 1'b0 ;
  assign n12230 = n5504 ^ n3000 ^ 1'b0 ;
  assign n12227 = ( n2729 & ~n3907 ) | ( n2729 & n6268 ) | ( ~n3907 & n6268 ) ;
  assign n12216 = ( n1555 & n2487 ) | ( n1555 & n8354 ) | ( n2487 & n8354 ) ;
  assign n12223 = n10652 ^ n3059 ^ 1'b0 ;
  assign n12220 = n5178 ^ n2697 ^ 1'b0 ;
  assign n12221 = n4613 & n12220 ;
  assign n12217 = ( x111 & n5836 ) | ( x111 & ~n11717 ) | ( n5836 & ~n11717 ) ;
  assign n12218 = ( ~n3422 & n9106 ) | ( ~n3422 & n11601 ) | ( n9106 & n11601 ) ;
  assign n12219 = ~n12217 & n12218 ;
  assign n12222 = n12221 ^ n12219 ^ 1'b0 ;
  assign n12224 = n12223 ^ n12222 ^ n9067 ;
  assign n12225 = n2664 & ~n12224 ;
  assign n12226 = n12216 & n12225 ;
  assign n12228 = n12227 ^ n12226 ^ n470 ;
  assign n12215 = n1564 | n2806 ;
  assign n12229 = n12228 ^ n12215 ^ 1'b0 ;
  assign n12231 = n12230 ^ n12229 ^ 1'b0 ;
  assign n12210 = x43 & ~n5230 ;
  assign n12211 = n12210 ^ n5458 ^ 1'b0 ;
  assign n12212 = ( n1436 & n7538 ) | ( n1436 & n12211 ) | ( n7538 & n12211 ) ;
  assign n12213 = n12212 ^ n8451 ^ n3882 ;
  assign n12214 = n2869 & ~n12213 ;
  assign n12232 = n12231 ^ n12214 ^ 1'b0 ;
  assign n12233 = n4505 & n7233 ;
  assign n12234 = ( n397 & n869 ) | ( n397 & ~n12233 ) | ( n869 & ~n12233 ) ;
  assign n12235 = ( n656 & n7674 ) | ( n656 & ~n9530 ) | ( n7674 & ~n9530 ) ;
  assign n12236 = n8009 ^ n7585 ^ n7165 ;
  assign n12237 = ( n3489 & n5858 ) | ( n3489 & ~n12236 ) | ( n5858 & ~n12236 ) ;
  assign n12240 = n11662 ^ n9819 ^ n1337 ;
  assign n12238 = ( n359 & n548 ) | ( n359 & ~n3509 ) | ( n548 & ~n3509 ) ;
  assign n12239 = ( n4194 & n5892 ) | ( n4194 & ~n12238 ) | ( n5892 & ~n12238 ) ;
  assign n12241 = n12240 ^ n12239 ^ 1'b0 ;
  assign n12242 = ~n10466 & n12241 ;
  assign n12243 = n12242 ^ n12116 ^ n3851 ;
  assign n12244 = ~n12237 & n12243 ;
  assign n12245 = n11935 ^ n11647 ^ n6626 ;
  assign n12246 = ( ~n6372 & n9666 ) | ( ~n6372 & n12245 ) | ( n9666 & n12245 ) ;
  assign n12251 = ( n362 & ~n4471 ) | ( n362 & n5148 ) | ( ~n4471 & n5148 ) ;
  assign n12252 = n7171 | n12251 ;
  assign n12253 = n12252 ^ n6673 ^ 1'b0 ;
  assign n12249 = n8050 ^ n1136 ^ 1'b0 ;
  assign n12247 = x59 & ~n4759 ;
  assign n12248 = n2371 & n12247 ;
  assign n12250 = n12249 ^ n12248 ^ n11128 ;
  assign n12254 = n12253 ^ n12250 ^ n3683 ;
  assign n12255 = n7859 ^ n4527 ^ n641 ;
  assign n12256 = ( ~n6302 & n7848 ) | ( ~n6302 & n12255 ) | ( n7848 & n12255 ) ;
  assign n12257 = ~n5171 & n12256 ;
  assign n12258 = ( n4647 & n8457 ) | ( n4647 & ~n12257 ) | ( n8457 & ~n12257 ) ;
  assign n12259 = n7692 ^ n5718 ^ n3255 ;
  assign n12260 = ( n1472 & n4115 ) | ( n1472 & n5310 ) | ( n4115 & n5310 ) ;
  assign n12261 = ~n3998 & n12260 ;
  assign n12262 = n12261 ^ n937 ^ 1'b0 ;
  assign n12267 = n3799 ^ n3413 ^ 1'b0 ;
  assign n12268 = ( ~n1976 & n2396 ) | ( ~n1976 & n4677 ) | ( n2396 & n4677 ) ;
  assign n12269 = n12268 ^ n10990 ^ 1'b0 ;
  assign n12270 = n12267 & ~n12269 ;
  assign n12265 = n3302 ^ n3117 ^ 1'b0 ;
  assign n12263 = n5967 | n7863 ;
  assign n12264 = n12263 ^ n5088 ^ n5073 ;
  assign n12266 = n12265 ^ n12264 ^ 1'b0 ;
  assign n12271 = n12270 ^ n12266 ^ n1266 ;
  assign n12272 = ( n586 & ~n5360 ) | ( n586 & n11832 ) | ( ~n5360 & n11832 ) ;
  assign n12274 = n2993 | n3285 ;
  assign n12273 = n4059 | n9549 ;
  assign n12275 = n12274 ^ n12273 ^ 1'b0 ;
  assign n12276 = ( n1886 & n6177 ) | ( n1886 & ~n12275 ) | ( n6177 & ~n12275 ) ;
  assign n12277 = n3522 ^ n252 ^ 1'b0 ;
  assign n12278 = ( n444 & n1224 ) | ( n444 & ~n12277 ) | ( n1224 & ~n12277 ) ;
  assign n12279 = n5606 | n12278 ;
  assign n12280 = n12276 & ~n12279 ;
  assign n12281 = n12280 ^ n8849 ^ n4659 ;
  assign n12282 = ( n2858 & ~n3610 ) | ( n2858 & n10195 ) | ( ~n3610 & n10195 ) ;
  assign n12283 = n11082 ^ n524 ^ 1'b0 ;
  assign n12284 = n2989 | n12283 ;
  assign n12285 = ( ~n2137 & n12083 ) | ( ~n2137 & n12284 ) | ( n12083 & n12284 ) ;
  assign n12286 = ( n597 & ~n1527 ) | ( n597 & n6473 ) | ( ~n1527 & n6473 ) ;
  assign n12287 = n12286 ^ n7137 ^ n2411 ;
  assign n12288 = n12287 ^ n11259 ^ 1'b0 ;
  assign n12289 = n2750 & n12288 ;
  assign n12290 = n3522 ^ n153 ^ 1'b0 ;
  assign n12291 = ( n4094 & n7152 ) | ( n4094 & n12290 ) | ( n7152 & n12290 ) ;
  assign n12292 = n1822 ^ n251 ^ 1'b0 ;
  assign n12293 = n4556 & ~n12292 ;
  assign n12294 = ~n3748 & n12293 ;
  assign n12295 = ( ~n512 & n5164 ) | ( ~n512 & n10049 ) | ( n5164 & n10049 ) ;
  assign n12296 = ( n7631 & n9337 ) | ( n7631 & ~n12295 ) | ( n9337 & ~n12295 ) ;
  assign n12297 = x89 & ~n4740 ;
  assign n12298 = ( n12294 & n12296 ) | ( n12294 & n12297 ) | ( n12296 & n12297 ) ;
  assign n12299 = ~n4465 & n7996 ;
  assign n12300 = n9610 ^ n3436 ^ 1'b0 ;
  assign n12301 = n12299 | n12300 ;
  assign n12302 = ( n1639 & n3786 ) | ( n1639 & n12301 ) | ( n3786 & n12301 ) ;
  assign n12303 = n12270 ^ n6709 ^ n4847 ;
  assign n12304 = ( n1073 & n2276 ) | ( n1073 & n8642 ) | ( n2276 & n8642 ) ;
  assign n12307 = ( n194 & n1874 ) | ( n194 & n4764 ) | ( n1874 & n4764 ) ;
  assign n12308 = ( n2875 & ~n5686 ) | ( n2875 & n8538 ) | ( ~n5686 & n8538 ) ;
  assign n12309 = n12307 & ~n12308 ;
  assign n12310 = n12309 ^ n1051 ^ 1'b0 ;
  assign n12305 = n4298 ^ n1510 ^ 1'b0 ;
  assign n12306 = n12305 ^ n8014 ^ n7249 ;
  assign n12311 = n12310 ^ n12306 ^ n9181 ;
  assign n12316 = n6152 ^ n5687 ^ n282 ;
  assign n12312 = n6459 ^ n1620 ^ n1245 ;
  assign n12313 = n3225 & ~n12312 ;
  assign n12314 = n8644 & ~n12313 ;
  assign n12315 = n12314 ^ n1035 ^ 1'b0 ;
  assign n12317 = n12316 ^ n12315 ^ n8983 ;
  assign n12318 = ( n7142 & ~n9936 ) | ( n7142 & n10939 ) | ( ~n9936 & n10939 ) ;
  assign n12319 = n1715 & n5427 ;
  assign n12320 = n4858 & n12319 ;
  assign n12321 = ( ~n2769 & n3009 ) | ( ~n2769 & n12320 ) | ( n3009 & n12320 ) ;
  assign n12322 = n6313 ^ n4476 ^ n2727 ;
  assign n12323 = ( n4200 & n7472 ) | ( n4200 & n12322 ) | ( n7472 & n12322 ) ;
  assign n12324 = n12323 ^ n2417 ^ n1417 ;
  assign n12325 = n12324 ^ n10017 ^ n2422 ;
  assign n12326 = ( ~n2720 & n3617 ) | ( ~n2720 & n7963 ) | ( n3617 & n7963 ) ;
  assign n12327 = ( ~n1677 & n4291 ) | ( ~n1677 & n12326 ) | ( n4291 & n12326 ) ;
  assign n12328 = n10827 ^ n4270 ^ 1'b0 ;
  assign n12329 = n1978 ^ n136 ^ 1'b0 ;
  assign n12330 = n3161 & n12329 ;
  assign n12331 = ( n357 & n3138 ) | ( n357 & n12052 ) | ( n3138 & n12052 ) ;
  assign n12332 = ( n609 & n10796 ) | ( n609 & ~n12331 ) | ( n10796 & ~n12331 ) ;
  assign n12334 = n3217 ^ n2020 ^ n788 ;
  assign n12333 = n9861 ^ n2616 ^ n440 ;
  assign n12335 = n12334 ^ n12333 ^ n9077 ;
  assign n12342 = ( x69 & n4910 ) | ( x69 & n5657 ) | ( n4910 & n5657 ) ;
  assign n12336 = n7020 ^ n243 ^ 1'b0 ;
  assign n12337 = ( n7257 & n7644 ) | ( n7257 & n12336 ) | ( n7644 & n12336 ) ;
  assign n12338 = ( n232 & n2535 ) | ( n232 & n7979 ) | ( n2535 & n7979 ) ;
  assign n12339 = n12338 ^ n1949 ^ 1'b0 ;
  assign n12340 = n6617 & ~n12339 ;
  assign n12341 = ( n5736 & ~n12337 ) | ( n5736 & n12340 ) | ( ~n12337 & n12340 ) ;
  assign n12343 = n12342 ^ n12341 ^ n1705 ;
  assign n12344 = ( x68 & n2665 ) | ( x68 & ~n5185 ) | ( n2665 & ~n5185 ) ;
  assign n12345 = n10521 ^ n2439 ^ 1'b0 ;
  assign n12346 = ~n12344 & n12345 ;
  assign n12347 = n2555 | n5287 ;
  assign n12348 = ( n6701 & n7175 ) | ( n6701 & ~n12347 ) | ( n7175 & ~n12347 ) ;
  assign n12349 = ~n12346 & n12348 ;
  assign n12350 = ~n396 & n6655 ;
  assign n12351 = n12350 ^ n11138 ^ 1'b0 ;
  assign n12355 = ~n2745 & n3952 ;
  assign n12352 = n7326 ^ n3168 ^ 1'b0 ;
  assign n12353 = ~n8131 & n12352 ;
  assign n12354 = ( n953 & n2132 ) | ( n953 & n12353 ) | ( n2132 & n12353 ) ;
  assign n12356 = n12355 ^ n12354 ^ n9244 ;
  assign n12357 = ( n3434 & n6223 ) | ( n3434 & n7422 ) | ( n6223 & n7422 ) ;
  assign n12358 = n12357 ^ n673 ^ 1'b0 ;
  assign n12359 = ~n7395 & n12358 ;
  assign n12360 = n12359 ^ n12113 ^ 1'b0 ;
  assign n12361 = ( n3420 & ~n8562 ) | ( n3420 & n12360 ) | ( ~n8562 & n12360 ) ;
  assign n12362 = ( n2751 & n3543 ) | ( n2751 & n5287 ) | ( n3543 & n5287 ) ;
  assign n12363 = n12362 ^ n8425 ^ n3235 ;
  assign n12364 = n7979 ^ n7933 ^ n3952 ;
  assign n12365 = ~n5400 & n7655 ;
  assign n12366 = n4221 & n12365 ;
  assign n12367 = ( n2862 & n3291 ) | ( n2862 & ~n9575 ) | ( n3291 & ~n9575 ) ;
  assign n12368 = ( ~n1160 & n12366 ) | ( ~n1160 & n12367 ) | ( n12366 & n12367 ) ;
  assign n12369 = ( ~n6007 & n6643 ) | ( ~n6007 & n12368 ) | ( n6643 & n12368 ) ;
  assign n12370 = ( ~n11528 & n12364 ) | ( ~n11528 & n12369 ) | ( n12364 & n12369 ) ;
  assign n12371 = ~n500 & n1475 ;
  assign n12372 = n12371 ^ n5581 ^ 1'b0 ;
  assign n12373 = ~n3581 & n8010 ;
  assign n12374 = ~n4303 & n12373 ;
  assign n12375 = n12374 ^ n8721 ^ 1'b0 ;
  assign n12376 = ~n12372 & n12375 ;
  assign n12377 = ( n1969 & ~n5683 ) | ( n1969 & n8380 ) | ( ~n5683 & n8380 ) ;
  assign n12378 = n10127 & ~n12377 ;
  assign n12379 = ~n856 & n12378 ;
  assign n12380 = n3935 ^ n3317 ^ 1'b0 ;
  assign n12381 = n12380 ^ n9929 ^ n8078 ;
  assign n12382 = n3510 ^ n3363 ^ n287 ;
  assign n12383 = ( n1985 & n4786 ) | ( n1985 & ~n12382 ) | ( n4786 & ~n12382 ) ;
  assign n12388 = ~n1781 & n2664 ;
  assign n12389 = n12388 ^ n2688 ^ 1'b0 ;
  assign n12390 = n12389 ^ n4196 ^ n292 ;
  assign n12391 = ( ~n383 & n4041 ) | ( ~n383 & n12390 ) | ( n4041 & n12390 ) ;
  assign n12384 = n5296 ^ n1164 ^ 1'b0 ;
  assign n12385 = n2884 | n12384 ;
  assign n12386 = n6241 | n12385 ;
  assign n12387 = n7059 | n12386 ;
  assign n12392 = n12391 ^ n12387 ^ 1'b0 ;
  assign n12393 = ~n3642 & n6980 ;
  assign n12394 = ~n4773 & n12393 ;
  assign n12395 = ~x28 & n12394 ;
  assign n12396 = n12395 ^ n2530 ^ x2 ;
  assign n12397 = n9072 ^ n5375 ^ n5367 ;
  assign n12398 = ( n3189 & n5080 ) | ( n3189 & ~n7429 ) | ( n5080 & ~n7429 ) ;
  assign n12401 = ( ~n251 & n2337 ) | ( ~n251 & n9662 ) | ( n2337 & n9662 ) ;
  assign n12399 = n9197 ^ n1385 ^ 1'b0 ;
  assign n12400 = n7867 & ~n12399 ;
  assign n12402 = n12401 ^ n12400 ^ n6886 ;
  assign n12403 = ( n10792 & n12398 ) | ( n10792 & n12402 ) | ( n12398 & n12402 ) ;
  assign n12404 = ( n3910 & n6499 ) | ( n3910 & n7467 ) | ( n6499 & n7467 ) ;
  assign n12405 = n12404 ^ n5161 ^ n1243 ;
  assign n12406 = n473 | n4239 ;
  assign n12407 = n3983 & ~n12406 ;
  assign n12408 = n12407 ^ n3966 ^ 1'b0 ;
  assign n12409 = n12408 ^ n8028 ^ n4566 ;
  assign n12410 = ( n4987 & n8726 ) | ( n4987 & ~n9131 ) | ( n8726 & ~n9131 ) ;
  assign n12411 = ( ~n6238 & n8241 ) | ( ~n6238 & n12410 ) | ( n8241 & n12410 ) ;
  assign n12412 = ( n4155 & ~n4447 ) | ( n4155 & n12411 ) | ( ~n4447 & n12411 ) ;
  assign n12413 = n9067 ^ n8841 ^ 1'b0 ;
  assign n12416 = n6858 & ~n10938 ;
  assign n12417 = ~n10442 & n12416 ;
  assign n12414 = n4514 ^ n1239 ^ n248 ;
  assign n12415 = n2152 | n12414 ;
  assign n12418 = n12417 ^ n12415 ^ 1'b0 ;
  assign n12427 = ( n3349 & n5027 ) | ( n3349 & n7204 ) | ( n5027 & n7204 ) ;
  assign n12422 = n5578 ^ n2630 ^ 1'b0 ;
  assign n12423 = ~n1627 & n12422 ;
  assign n12419 = n1160 | n8296 ;
  assign n12420 = n4828 & ~n12419 ;
  assign n12421 = n6021 | n12420 ;
  assign n12424 = n12423 ^ n12421 ^ n2842 ;
  assign n12425 = ~n10273 & n12424 ;
  assign n12426 = n12425 ^ n11433 ^ 1'b0 ;
  assign n12428 = n12427 ^ n12426 ^ 1'b0 ;
  assign n12429 = ( n2879 & n6761 ) | ( n2879 & n10720 ) | ( n6761 & n10720 ) ;
  assign n12430 = ( n7564 & n7593 ) | ( n7564 & n12429 ) | ( n7593 & n12429 ) ;
  assign n12431 = n12430 ^ n10823 ^ n10762 ;
  assign n12432 = n7446 & n10713 ;
  assign n12433 = n2906 ^ n2352 ^ 1'b0 ;
  assign n12434 = ~n6562 & n9559 ;
  assign n12435 = n12200 ^ n7979 ^ n3877 ;
  assign n12440 = n10008 ^ n4401 ^ n4244 ;
  assign n12441 = n649 & ~n12440 ;
  assign n12439 = n3141 ^ n1693 ^ 1'b0 ;
  assign n12442 = n12441 ^ n12439 ^ 1'b0 ;
  assign n12436 = ~n4536 & n8976 ;
  assign n12437 = ~n2073 & n12436 ;
  assign n12438 = n12437 ^ n4826 ^ n3979 ;
  assign n12443 = n12442 ^ n12438 ^ 1'b0 ;
  assign n12444 = n12435 & ~n12443 ;
  assign n12445 = n12444 ^ n11749 ^ n7560 ;
  assign n12447 = n8465 ^ n7191 ^ n272 ;
  assign n12446 = ( n3048 & n4764 ) | ( n3048 & n4895 ) | ( n4764 & n4895 ) ;
  assign n12448 = n12447 ^ n12446 ^ 1'b0 ;
  assign n12449 = n1184 & ~n12448 ;
  assign n12450 = n2428 | n12449 ;
  assign n12451 = n5382 ^ n1665 ^ 1'b0 ;
  assign n12452 = n10377 ^ n10226 ^ 1'b0 ;
  assign n12455 = ( ~n4120 & n5298 ) | ( ~n4120 & n5736 ) | ( n5298 & n5736 ) ;
  assign n12453 = ( n1166 & n1878 ) | ( n1166 & n6336 ) | ( n1878 & n6336 ) ;
  assign n12454 = n6013 & n12453 ;
  assign n12456 = n12455 ^ n12454 ^ 1'b0 ;
  assign n12457 = ~n2142 & n12456 ;
  assign n12458 = n12457 ^ n3931 ^ 1'b0 ;
  assign n12459 = ( n7443 & n9397 ) | ( n7443 & ~n12458 ) | ( n9397 & ~n12458 ) ;
  assign n12460 = n10900 ^ n4822 ^ n1466 ;
  assign n12461 = ( n3382 & ~n6393 ) | ( n3382 & n12460 ) | ( ~n6393 & n12460 ) ;
  assign n12462 = ( n200 & ~n4997 ) | ( n200 & n6435 ) | ( ~n4997 & n6435 ) ;
  assign n12463 = n12462 ^ n11415 ^ 1'b0 ;
  assign n12464 = n3585 ^ n2081 ^ 1'b0 ;
  assign n12465 = ( n2255 & n12463 ) | ( n2255 & ~n12464 ) | ( n12463 & ~n12464 ) ;
  assign n12466 = n1735 | n2929 ;
  assign n12467 = n12466 ^ n5881 ^ n5370 ;
  assign n12475 = n11480 ^ n9763 ^ x60 ;
  assign n12468 = n11307 ^ n5050 ^ 1'b0 ;
  assign n12469 = n7972 ^ n6515 ^ n2258 ;
  assign n12470 = ( n6094 & n12016 ) | ( n6094 & n12469 ) | ( n12016 & n12469 ) ;
  assign n12471 = ~n9348 & n12470 ;
  assign n12472 = n12471 ^ x73 ^ 1'b0 ;
  assign n12473 = ~n12468 & n12472 ;
  assign n12474 = n12473 ^ n8611 ^ 1'b0 ;
  assign n12476 = n12475 ^ n12474 ^ n1983 ;
  assign n12477 = ( n6883 & n7198 ) | ( n6883 & n11965 ) | ( n7198 & n11965 ) ;
  assign n12478 = n12477 ^ n7276 ^ n496 ;
  assign n12479 = n12478 ^ n4476 ^ 1'b0 ;
  assign n12483 = n10358 ^ n7781 ^ n3673 ;
  assign n12484 = n12483 ^ n8124 ^ n4940 ;
  assign n12485 = ( n9831 & n12098 ) | ( n9831 & n12484 ) | ( n12098 & n12484 ) ;
  assign n12480 = n5242 ^ n1226 ^ n1150 ;
  assign n12481 = ( n1731 & n4770 ) | ( n1731 & ~n12480 ) | ( n4770 & ~n12480 ) ;
  assign n12482 = ( n2732 & n8680 ) | ( n2732 & n12481 ) | ( n8680 & n12481 ) ;
  assign n12486 = n12485 ^ n12482 ^ n2372 ;
  assign n12487 = n12486 ^ n3455 ^ n1095 ;
  assign n12492 = n696 ^ x52 ^ 1'b0 ;
  assign n12493 = ( n6934 & n11785 ) | ( n6934 & n12492 ) | ( n11785 & n12492 ) ;
  assign n12490 = ~n6969 & n10382 ;
  assign n12491 = n12490 ^ n11237 ^ 1'b0 ;
  assign n12488 = n11855 ^ n9961 ^ n7070 ;
  assign n12489 = n12488 ^ n1774 ^ 1'b0 ;
  assign n12494 = n12493 ^ n12491 ^ n12489 ;
  assign n12495 = n9568 ^ n3518 ^ 1'b0 ;
  assign n12503 = n3218 & ~n9681 ;
  assign n12504 = n12503 ^ n1320 ^ 1'b0 ;
  assign n12502 = n4562 ^ n4111 ^ n2047 ;
  assign n12505 = n12504 ^ n12502 ^ 1'b0 ;
  assign n12496 = n10025 ^ n8588 ^ n2902 ;
  assign n12498 = n1563 ^ n749 ^ 1'b0 ;
  assign n12497 = ( n1418 & n2531 ) | ( n1418 & ~n7806 ) | ( n2531 & ~n7806 ) ;
  assign n12499 = n12498 ^ n12497 ^ n8412 ;
  assign n12500 = ( n1504 & n8821 ) | ( n1504 & n12499 ) | ( n8821 & n12499 ) ;
  assign n12501 = n12496 & ~n12500 ;
  assign n12506 = n12505 ^ n12501 ^ 1'b0 ;
  assign n12507 = ( ~n2696 & n7356 ) | ( ~n2696 & n7699 ) | ( n7356 & n7699 ) ;
  assign n12513 = ( n4379 & n5815 ) | ( n4379 & n6932 ) | ( n5815 & n6932 ) ;
  assign n12511 = ( n3678 & n5773 ) | ( n3678 & ~n11526 ) | ( n5773 & ~n11526 ) ;
  assign n12512 = ( ~n4249 & n11817 ) | ( ~n4249 & n12511 ) | ( n11817 & n12511 ) ;
  assign n12509 = ~n649 & n8972 ;
  assign n12508 = n11284 ^ n6103 ^ n3515 ;
  assign n12510 = n12509 ^ n12508 ^ n5293 ;
  assign n12514 = n12513 ^ n12512 ^ n12510 ;
  assign n12515 = ( n4520 & n4685 ) | ( n4520 & n10711 ) | ( n4685 & n10711 ) ;
  assign n12516 = ~n11988 & n12515 ;
  assign n12517 = ( n1045 & n3197 ) | ( n1045 & n3249 ) | ( n3197 & n3249 ) ;
  assign n12518 = n12517 ^ n6582 ^ n4474 ;
  assign n12519 = n8217 ^ n603 ^ n340 ;
  assign n12520 = n4018 & ~n4125 ;
  assign n12521 = ~n2374 & n4689 ;
  assign n12522 = n12521 ^ n10752 ^ 1'b0 ;
  assign n12523 = n6657 & ~n12522 ;
  assign n12524 = ( n5756 & n9224 ) | ( n5756 & n12523 ) | ( n9224 & n12523 ) ;
  assign n12525 = ( n12519 & n12520 ) | ( n12519 & n12524 ) | ( n12520 & n12524 ) ;
  assign n12531 = n10066 ^ n9008 ^ n8856 ;
  assign n12526 = ~n268 & n5419 ;
  assign n12527 = n12526 ^ n5937 ^ 1'b0 ;
  assign n12528 = n12527 ^ n4121 ^ n2642 ;
  assign n12529 = ( n3299 & ~n8582 ) | ( n3299 & n12528 ) | ( ~n8582 & n12528 ) ;
  assign n12530 = n11921 | n12529 ;
  assign n12532 = n12531 ^ n12530 ^ 1'b0 ;
  assign n12533 = ( ~n10939 & n12025 ) | ( ~n10939 & n12532 ) | ( n12025 & n12532 ) ;
  assign n12534 = n6032 ^ n2061 ^ n951 ;
  assign n12535 = ( ~n1138 & n3033 ) | ( ~n1138 & n12401 ) | ( n3033 & n12401 ) ;
  assign n12536 = n4020 & n4527 ;
  assign n12537 = ( n3215 & n7450 ) | ( n3215 & n12536 ) | ( n7450 & n12536 ) ;
  assign n12538 = n7486 | n12537 ;
  assign n12539 = n12538 ^ n11736 ^ 1'b0 ;
  assign n12540 = ( n12534 & ~n12535 ) | ( n12534 & n12539 ) | ( ~n12535 & n12539 ) ;
  assign n12543 = n7342 ^ n142 ^ 1'b0 ;
  assign n12544 = n12543 ^ n4513 ^ n1271 ;
  assign n12541 = n499 | n6470 ;
  assign n12542 = n12541 ^ n9977 ^ n2642 ;
  assign n12545 = n12544 ^ n12542 ^ n499 ;
  assign n12546 = ( ~n2598 & n3380 ) | ( ~n2598 & n3870 ) | ( n3380 & n3870 ) ;
  assign n12547 = n1635 & ~n12546 ;
  assign n12548 = n7479 & n12547 ;
  assign n12549 = ~n12030 & n12548 ;
  assign n12550 = ( n312 & ~n1020 ) | ( n312 & n1220 ) | ( ~n1020 & n1220 ) ;
  assign n12552 = n840 & ~n9325 ;
  assign n12553 = n8844 & n12552 ;
  assign n12551 = n8577 & n10850 ;
  assign n12554 = n12553 ^ n12551 ^ n5182 ;
  assign n12555 = ( ~n3322 & n12550 ) | ( ~n3322 & n12554 ) | ( n12550 & n12554 ) ;
  assign n12556 = n12555 ^ n7103 ^ 1'b0 ;
  assign n12557 = n2706 & ~n6636 ;
  assign n12558 = ( n1477 & n8502 ) | ( n1477 & n12557 ) | ( n8502 & n12557 ) ;
  assign n12559 = ( n1887 & n3639 ) | ( n1887 & ~n10541 ) | ( n3639 & ~n10541 ) ;
  assign n12560 = n12559 ^ n4878 ^ n4822 ;
  assign n12562 = n7849 ^ n6382 ^ n323 ;
  assign n12563 = n12562 ^ n2043 ^ n1920 ;
  assign n12561 = n2062 & ~n7120 ;
  assign n12564 = n12563 ^ n12561 ^ 1'b0 ;
  assign n12565 = ( n4189 & ~n4575 ) | ( n4189 & n4769 ) | ( ~n4575 & n4769 ) ;
  assign n12566 = ~n3857 & n12565 ;
  assign n12567 = n12529 & n12566 ;
  assign n12568 = n12567 ^ n7911 ^ n1920 ;
  assign n12569 = n5336 ^ n5313 ^ 1'b0 ;
  assign n12571 = n1526 ^ n1186 ^ x11 ;
  assign n12572 = n12571 ^ n9819 ^ n5568 ;
  assign n12573 = ( x58 & ~n906 ) | ( x58 & n12572 ) | ( ~n906 & n12572 ) ;
  assign n12570 = ( n6292 & n7865 ) | ( n6292 & n10368 ) | ( n7865 & n10368 ) ;
  assign n12574 = n12573 ^ n12570 ^ n6182 ;
  assign n12575 = ~n500 & n2376 ;
  assign n12579 = n10479 ^ n3923 ^ n578 ;
  assign n12578 = n10404 ^ n7414 ^ n3283 ;
  assign n12576 = n4352 & n12505 ;
  assign n12577 = n12576 ^ n7290 ^ 1'b0 ;
  assign n12580 = n12579 ^ n12578 ^ n12577 ;
  assign n12581 = n10968 ^ n7377 ^ n4131 ;
  assign n12582 = ( ~n12575 & n12580 ) | ( ~n12575 & n12581 ) | ( n12580 & n12581 ) ;
  assign n12583 = ( ~x93 & n718 ) | ( ~x93 & n1485 ) | ( n718 & n1485 ) ;
  assign n12584 = n2260 | n6024 ;
  assign n12585 = n12583 | n12584 ;
  assign n12586 = ( ~n1406 & n2792 ) | ( ~n1406 & n4439 ) | ( n2792 & n4439 ) ;
  assign n12587 = n7840 & ~n12586 ;
  assign n12588 = n6557 ^ n4333 ^ 1'b0 ;
  assign n12589 = ~n3032 & n7062 ;
  assign n12590 = ~n5106 & n12589 ;
  assign n12591 = n10860 ^ n6261 ^ n5982 ;
  assign n12592 = n7928 ^ n3342 ^ n2183 ;
  assign n12593 = n4982 | n12592 ;
  assign n12594 = n8722 ^ n8043 ^ n6414 ;
  assign n12595 = ( ~n4826 & n12455 ) | ( ~n4826 & n12594 ) | ( n12455 & n12594 ) ;
  assign n12596 = n12595 ^ n236 ^ 1'b0 ;
  assign n12597 = n2830 | n12596 ;
  assign n12598 = ( n2060 & ~n6268 ) | ( n2060 & n6639 ) | ( ~n6268 & n6639 ) ;
  assign n12599 = n10189 ^ n5018 ^ n923 ;
  assign n12600 = ( n1861 & ~n6107 ) | ( n1861 & n12599 ) | ( ~n6107 & n12599 ) ;
  assign n12601 = ( n11781 & n12598 ) | ( n11781 & n12600 ) | ( n12598 & n12600 ) ;
  assign n12602 = n9931 ^ n3807 ^ n1917 ;
  assign n12603 = n12602 ^ n10420 ^ n8077 ;
  assign n12604 = ~n12099 & n12603 ;
  assign n12605 = n6024 ^ n4664 ^ n1507 ;
  assign n12606 = n10479 ^ n5408 ^ n890 ;
  assign n12607 = n5708 & n12606 ;
  assign n12608 = ~n4203 & n12607 ;
  assign n12609 = n6447 ^ n5296 ^ n3000 ;
  assign n12610 = ~n12608 & n12609 ;
  assign n12611 = ~n5906 & n12610 ;
  assign n12612 = ( n749 & ~n12605 ) | ( n749 & n12611 ) | ( ~n12605 & n12611 ) ;
  assign n12613 = n9153 ^ n2852 ^ 1'b0 ;
  assign n12614 = ~n12113 & n12613 ;
  assign n12615 = ( n482 & n662 ) | ( n482 & n980 ) | ( n662 & n980 ) ;
  assign n12616 = ( n1731 & n12307 ) | ( n1731 & ~n12615 ) | ( n12307 & ~n12615 ) ;
  assign n12617 = ( ~n5657 & n12614 ) | ( ~n5657 & n12616 ) | ( n12614 & n12616 ) ;
  assign n12618 = n12617 ^ n2122 ^ 1'b0 ;
  assign n12619 = n2345 & n12618 ;
  assign n12621 = ( x7 & n885 ) | ( x7 & ~n11388 ) | ( n885 & ~n11388 ) ;
  assign n12620 = n1145 | n8407 ;
  assign n12622 = n12621 ^ n12620 ^ 1'b0 ;
  assign n12623 = n12622 ^ n9104 ^ n6943 ;
  assign n12626 = n7862 ^ n6603 ^ n850 ;
  assign n12624 = n4127 & ~n8457 ;
  assign n12625 = ~n326 & n12624 ;
  assign n12627 = n12626 ^ n12625 ^ 1'b0 ;
  assign n12628 = n12623 | n12627 ;
  assign n12629 = ( n3567 & ~n4841 ) | ( n3567 & n6437 ) | ( ~n4841 & n6437 ) ;
  assign n12630 = ( n1116 & ~n4064 ) | ( n1116 & n4078 ) | ( ~n4064 & n4078 ) ;
  assign n12631 = n12630 ^ n2957 ^ n2858 ;
  assign n12632 = n12631 ^ n3895 ^ n2444 ;
  assign n12633 = n12632 ^ n3557 ^ n1980 ;
  assign n12634 = n12633 ^ n11467 ^ n9288 ;
  assign n12635 = n5803 ^ n5799 ^ 1'b0 ;
  assign n12636 = ~n1875 & n12635 ;
  assign n12637 = n12636 ^ n7072 ^ 1'b0 ;
  assign n12638 = n4905 | n12637 ;
  assign n12639 = n8120 ^ n4465 ^ n995 ;
  assign n12640 = ( n136 & ~n3640 ) | ( n136 & n8658 ) | ( ~n3640 & n8658 ) ;
  assign n12641 = n12640 ^ n9881 ^ n5786 ;
  assign n12642 = n11927 ^ n5727 ^ 1'b0 ;
  assign n12643 = ( n928 & n1008 ) | ( n928 & ~n2283 ) | ( n1008 & ~n2283 ) ;
  assign n12644 = ( n3157 & n12642 ) | ( n3157 & n12643 ) | ( n12642 & n12643 ) ;
  assign n12645 = ( n1625 & ~n6471 ) | ( n1625 & n11115 ) | ( ~n6471 & n11115 ) ;
  assign n12648 = n8446 ^ n2241 ^ n1006 ;
  assign n12646 = n6926 ^ n3108 ^ n2047 ;
  assign n12647 = n12646 ^ n11836 ^ n529 ;
  assign n12649 = n12648 ^ n12647 ^ n7571 ;
  assign n12650 = n12649 ^ n6899 ^ n3594 ;
  assign n12651 = n12650 ^ n4118 ^ 1'b0 ;
  assign n12652 = ( n769 & n12357 ) | ( n769 & n12651 ) | ( n12357 & n12651 ) ;
  assign n12653 = ( n2599 & ~n4036 ) | ( n2599 & n4639 ) | ( ~n4036 & n4639 ) ;
  assign n12654 = ( n4224 & ~n7049 ) | ( n4224 & n12653 ) | ( ~n7049 & n12653 ) ;
  assign n12655 = n12654 ^ n11043 ^ n1412 ;
  assign n12656 = n4395 ^ n665 ^ n475 ;
  assign n12657 = n12656 ^ n5763 ^ n3998 ;
  assign n12658 = n12657 ^ n8452 ^ n6685 ;
  assign n12659 = n12658 ^ n5577 ^ n1001 ;
  assign n12660 = n7632 ^ n5718 ^ n4842 ;
  assign n12661 = ( n868 & ~n7847 ) | ( n868 & n12660 ) | ( ~n7847 & n12660 ) ;
  assign n12662 = n1926 ^ x54 ^ 1'b0 ;
  assign n12663 = n2121 | n12662 ;
  assign n12664 = n3665 & n12663 ;
  assign n12665 = ( n758 & n12661 ) | ( n758 & n12664 ) | ( n12661 & n12664 ) ;
  assign n12666 = ( n7207 & ~n12659 ) | ( n7207 & n12665 ) | ( ~n12659 & n12665 ) ;
  assign n12667 = n12666 ^ n4530 ^ 1'b0 ;
  assign n12668 = n11439 & n12667 ;
  assign n12669 = n8293 ^ n4046 ^ n3880 ;
  assign n12670 = ( ~n3149 & n4011 ) | ( ~n3149 & n5464 ) | ( n4011 & n5464 ) ;
  assign n12671 = ( n1051 & n11038 ) | ( n1051 & ~n12670 ) | ( n11038 & ~n12670 ) ;
  assign n12672 = n8296 ^ n3102 ^ n616 ;
  assign n12673 = n12672 ^ n4331 ^ 1'b0 ;
  assign n12674 = n4366 & n12673 ;
  assign n12675 = ( ~n5650 & n6042 ) | ( ~n5650 & n12674 ) | ( n6042 & n12674 ) ;
  assign n12676 = n3521 & n6653 ;
  assign n12679 = ( ~x65 & n4765 ) | ( ~x65 & n5486 ) | ( n4765 & n5486 ) ;
  assign n12677 = ~n3398 & n12221 ;
  assign n12678 = n12677 ^ n1244 ^ 1'b0 ;
  assign n12680 = n12679 ^ n12678 ^ n2762 ;
  assign n12681 = n4728 ^ n3246 ^ 1'b0 ;
  assign n12682 = ~n4100 & n12681 ;
  assign n12683 = n12682 ^ n3450 ^ n3302 ;
  assign n12684 = n12683 ^ n8713 ^ n6098 ;
  assign n12685 = n12684 ^ n10498 ^ n2262 ;
  assign n12686 = ~n1361 & n1962 ;
  assign n12687 = n12686 ^ x112 ^ 1'b0 ;
  assign n12689 = n377 & ~n3020 ;
  assign n12688 = ( n890 & n8124 ) | ( n890 & n11357 ) | ( n8124 & n11357 ) ;
  assign n12690 = n12689 ^ n12688 ^ n883 ;
  assign n12691 = ( n5429 & ~n12687 ) | ( n5429 & n12690 ) | ( ~n12687 & n12690 ) ;
  assign n12692 = n1997 | n12691 ;
  assign n12693 = n12692 ^ n12453 ^ 1'b0 ;
  assign n12694 = ( n626 & ~n1677 ) | ( n626 & n1823 ) | ( ~n1677 & n1823 ) ;
  assign n12695 = n12694 ^ n9568 ^ n2220 ;
  assign n12696 = ( n396 & n5840 ) | ( n396 & n12695 ) | ( n5840 & n12695 ) ;
  assign n12697 = n7424 ^ n4891 ^ x64 ;
  assign n12698 = n5565 ^ n479 ^ 1'b0 ;
  assign n12699 = ~n12697 & n12698 ;
  assign n12700 = n603 & n12699 ;
  assign n12701 = ( n1751 & n12696 ) | ( n1751 & ~n12700 ) | ( n12696 & ~n12700 ) ;
  assign n12702 = n12257 ^ n12133 ^ n5563 ;
  assign n12704 = ~n2639 & n9495 ;
  assign n12705 = n12704 ^ n5757 ^ 1'b0 ;
  assign n12703 = n2190 | n7047 ;
  assign n12706 = n12705 ^ n12703 ^ 1'b0 ;
  assign n12707 = n7585 & ~n8124 ;
  assign n12708 = ( ~n2652 & n6047 ) | ( ~n2652 & n12707 ) | ( n6047 & n12707 ) ;
  assign n12709 = n10212 ^ n9153 ^ 1'b0 ;
  assign n12710 = n4519 & ~n12709 ;
  assign n12711 = n209 & ~n4703 ;
  assign n12712 = n6997 & ~n12711 ;
  assign n12713 = n8135 ^ n2755 ^ 1'b0 ;
  assign n12714 = n12712 & ~n12713 ;
  assign n12715 = ( n12708 & n12710 ) | ( n12708 & n12714 ) | ( n12710 & n12714 ) ;
  assign n12718 = n2831 & n3507 ;
  assign n12719 = n871 & n12718 ;
  assign n12720 = n7514 | n12719 ;
  assign n12716 = n6232 & ~n9050 ;
  assign n12717 = n12716 ^ n9270 ^ 1'b0 ;
  assign n12721 = n12720 ^ n12717 ^ 1'b0 ;
  assign n12722 = n8858 ^ n2183 ^ 1'b0 ;
  assign n12723 = n8169 ^ n5552 ^ 1'b0 ;
  assign n12724 = n12723 ^ n1833 ^ n869 ;
  assign n12725 = ( ~n5601 & n12722 ) | ( ~n5601 & n12724 ) | ( n12722 & n12724 ) ;
  assign n12726 = n5196 ^ n830 ^ n207 ;
  assign n12727 = ( n1206 & ~n4915 ) | ( n1206 & n12726 ) | ( ~n4915 & n12726 ) ;
  assign n12728 = n9194 ^ n6080 ^ n2959 ;
  assign n12729 = ( ~n8844 & n11484 ) | ( ~n8844 & n12728 ) | ( n11484 & n12728 ) ;
  assign n12730 = ( x13 & n5899 ) | ( x13 & n9835 ) | ( n5899 & n9835 ) ;
  assign n12731 = n6027 | n10517 ;
  assign n12732 = n12731 ^ n9292 ^ n2096 ;
  assign n12733 = ( ~n12729 & n12730 ) | ( ~n12729 & n12732 ) | ( n12730 & n12732 ) ;
  assign n12734 = n11214 ^ n9186 ^ n7125 ;
  assign n12735 = n11985 ^ n2591 ^ 1'b0 ;
  assign n12736 = n12734 & n12735 ;
  assign n12737 = n2337 & ~n12133 ;
  assign n12738 = n12737 ^ n10554 ^ 1'b0 ;
  assign n12742 = n7460 ^ n2322 ^ 1'b0 ;
  assign n12743 = ( n659 & n1725 ) | ( n659 & n2200 ) | ( n1725 & n2200 ) ;
  assign n12744 = ( n4071 & n12742 ) | ( n4071 & ~n12743 ) | ( n12742 & ~n12743 ) ;
  assign n12745 = n12744 ^ n7651 ^ n3420 ;
  assign n12741 = n12204 ^ n11285 ^ n4073 ;
  assign n12746 = n12745 ^ n12741 ^ n12414 ;
  assign n12739 = n9271 & ~n9629 ;
  assign n12740 = n12739 ^ n8619 ^ 1'b0 ;
  assign n12747 = n12746 ^ n12740 ^ n10198 ;
  assign n12751 = ( x112 & n1091 ) | ( x112 & n4003 ) | ( n1091 & n4003 ) ;
  assign n12752 = ( ~n855 & n2135 ) | ( ~n855 & n5073 ) | ( n2135 & n5073 ) ;
  assign n12753 = ~n12751 & n12752 ;
  assign n12754 = n12753 ^ n2950 ^ 1'b0 ;
  assign n12748 = ( n1518 & ~n2077 ) | ( n1518 & n7424 ) | ( ~n2077 & n7424 ) ;
  assign n12749 = n7268 & ~n12748 ;
  assign n12750 = ( n4228 & n7017 ) | ( n4228 & n12749 ) | ( n7017 & n12749 ) ;
  assign n12755 = n12754 ^ n12750 ^ n4793 ;
  assign n12756 = ( n696 & ~n2049 ) | ( n696 & n12236 ) | ( ~n2049 & n12236 ) ;
  assign n12757 = n5311 ^ n4109 ^ 1'b0 ;
  assign n12758 = n12757 ^ n3937 ^ 1'b0 ;
  assign n12759 = n7361 & ~n12758 ;
  assign n12762 = n11862 ^ n10365 ^ n8503 ;
  assign n12760 = n10827 ^ n1642 ^ n829 ;
  assign n12761 = ~n912 & n12760 ;
  assign n12763 = n12762 ^ n12761 ^ 1'b0 ;
  assign n12764 = ~n1709 & n12763 ;
  assign n12765 = n12764 ^ n628 ^ 1'b0 ;
  assign n12766 = ( n7602 & ~n10664 ) | ( n7602 & n11440 ) | ( ~n10664 & n11440 ) ;
  assign n12767 = n912 & n2540 ;
  assign n12768 = n12767 ^ n859 ^ 1'b0 ;
  assign n12769 = ( n3563 & n7153 ) | ( n3563 & n10221 ) | ( n7153 & n10221 ) ;
  assign n12770 = ( n2595 & n6279 ) | ( n2595 & n6960 ) | ( n6279 & n6960 ) ;
  assign n12771 = n6884 | n6934 ;
  assign n12772 = n12770 | n12771 ;
  assign n12779 = x119 & ~n2275 ;
  assign n12780 = ~n2279 & n12779 ;
  assign n12778 = n596 & ~n12164 ;
  assign n12781 = n12780 ^ n12778 ^ 1'b0 ;
  assign n12782 = ~n5802 & n12781 ;
  assign n12773 = ( x85 & ~n1122 ) | ( x85 & n4655 ) | ( ~n1122 & n4655 ) ;
  assign n12774 = n9542 & ~n12773 ;
  assign n12775 = n6413 ^ n5966 ^ n388 ;
  assign n12776 = n12775 ^ n9966 ^ n4292 ;
  assign n12777 = n12774 | n12776 ;
  assign n12783 = n12782 ^ n12777 ^ 1'b0 ;
  assign n12784 = ( n464 & n3227 ) | ( n464 & ~n5468 ) | ( n3227 & ~n5468 ) ;
  assign n12785 = n12784 ^ n11561 ^ n4971 ;
  assign n12786 = n12785 ^ n5121 ^ n3994 ;
  assign n12787 = n10761 & ~n12786 ;
  assign n12788 = n10030 ^ n6785 ^ n1455 ;
  assign n12789 = n1284 ^ n327 ^ 1'b0 ;
  assign n12790 = ( ~n1761 & n6291 ) | ( ~n1761 & n12789 ) | ( n6291 & n12789 ) ;
  assign n12791 = ( n4732 & n6874 ) | ( n4732 & n12790 ) | ( n6874 & n12790 ) ;
  assign n12792 = n12791 ^ n3201 ^ 1'b0 ;
  assign n12793 = n946 & ~n2519 ;
  assign n12794 = n12793 ^ n2722 ^ 1'b0 ;
  assign n12795 = n410 & n12794 ;
  assign n12796 = n2979 | n5791 ;
  assign n12797 = n12795 & ~n12796 ;
  assign n12798 = ( ~n2962 & n3855 ) | ( ~n2962 & n4128 ) | ( n3855 & n4128 ) ;
  assign n12799 = n12798 ^ n424 ^ 1'b0 ;
  assign n12800 = ( ~n846 & n6149 ) | ( ~n846 & n6502 ) | ( n6149 & n6502 ) ;
  assign n12801 = n12800 ^ n8863 ^ n4227 ;
  assign n12802 = ( ~n3452 & n12799 ) | ( ~n3452 & n12801 ) | ( n12799 & n12801 ) ;
  assign n12803 = ( n6291 & n12797 ) | ( n6291 & n12802 ) | ( n12797 & n12802 ) ;
  assign n12804 = n12803 ^ n12477 ^ n3858 ;
  assign n12805 = n10420 ^ n8016 ^ n4398 ;
  assign n12806 = n9145 ^ n8725 ^ 1'b0 ;
  assign n12807 = n12805 | n12806 ;
  assign n12809 = ( ~n2644 & n3341 ) | ( ~n2644 & n3400 ) | ( n3341 & n3400 ) ;
  assign n12808 = n12342 ^ n11063 ^ n2688 ;
  assign n12810 = n12809 ^ n12808 ^ n5394 ;
  assign n12813 = n10922 ^ n2955 ^ 1'b0 ;
  assign n12814 = ~n5460 & n12813 ;
  assign n12811 = n4514 ^ n4003 ^ n1713 ;
  assign n12812 = n12811 ^ n5588 ^ n935 ;
  assign n12815 = n12814 ^ n12812 ^ n1629 ;
  assign n12821 = ( ~n2636 & n4942 ) | ( ~n2636 & n11181 ) | ( n4942 & n11181 ) ;
  assign n12816 = n3031 & n9960 ;
  assign n12817 = n3170 ^ n1382 ^ 1'b0 ;
  assign n12818 = n631 & n12817 ;
  assign n12819 = n11505 & n12818 ;
  assign n12820 = n12816 & n12819 ;
  assign n12822 = n12821 ^ n12820 ^ 1'b0 ;
  assign n12823 = n10757 & n12822 ;
  assign n12824 = n8932 ^ n7447 ^ 1'b0 ;
  assign n12825 = ( n9325 & n12351 ) | ( n9325 & n12824 ) | ( n12351 & n12824 ) ;
  assign n12826 = ~n5134 & n7100 ;
  assign n12827 = n12826 ^ n2952 ^ 1'b0 ;
  assign n12831 = ( n611 & ~n6315 ) | ( n611 & n8343 ) | ( ~n6315 & n8343 ) ;
  assign n12830 = ( n4081 & n4700 ) | ( n4081 & ~n9714 ) | ( n4700 & ~n9714 ) ;
  assign n12828 = n2664 & n6977 ;
  assign n12829 = n12828 ^ n10899 ^ 1'b0 ;
  assign n12832 = n12831 ^ n12830 ^ n12829 ;
  assign n12833 = n12294 ^ n6421 ^ n6132 ;
  assign n12834 = ( n12827 & ~n12832 ) | ( n12827 & n12833 ) | ( ~n12832 & n12833 ) ;
  assign n12835 = n6590 ^ n2216 ^ 1'b0 ;
  assign n12836 = n4348 | n8338 ;
  assign n12837 = n12835 | n12836 ;
  assign n12838 = n12837 ^ n8084 ^ n2938 ;
  assign n12839 = n11850 ^ n8195 ^ n358 ;
  assign n12840 = n12839 ^ n8575 ^ n3136 ;
  assign n12841 = ( n7781 & n9955 ) | ( n7781 & ~n12134 ) | ( n9955 & ~n12134 ) ;
  assign n12842 = n4364 ^ n4352 ^ n2678 ;
  assign n12843 = n12842 ^ n5269 ^ 1'b0 ;
  assign n12844 = n6708 ^ n5784 ^ n349 ;
  assign n12845 = ( n3562 & n12843 ) | ( n3562 & ~n12844 ) | ( n12843 & ~n12844 ) ;
  assign n12846 = n12260 ^ n4842 ^ 1'b0 ;
  assign n12847 = n12846 ^ n2144 ^ 1'b0 ;
  assign n12853 = ( n3668 & ~n7052 ) | ( n3668 & n8766 ) | ( ~n7052 & n8766 ) ;
  assign n12848 = n4628 ^ n1453 ^ x6 ;
  assign n12849 = n862 & ~n1065 ;
  assign n12850 = n12849 ^ n141 ^ 1'b0 ;
  assign n12851 = n12850 ^ n3397 ^ 1'b0 ;
  assign n12852 = n12848 & ~n12851 ;
  assign n12854 = n12853 ^ n12852 ^ n4336 ;
  assign n12855 = n12854 ^ n6873 ^ n2050 ;
  assign n12856 = ( n2687 & n5702 ) | ( n2687 & ~n6594 ) | ( n5702 & ~n6594 ) ;
  assign n12857 = n11501 | n12856 ;
  assign n12858 = n12857 ^ n1380 ^ 1'b0 ;
  assign n12859 = ~n6433 & n11795 ;
  assign n12860 = n12859 ^ n4986 ^ 1'b0 ;
  assign n12861 = ( n10048 & ~n12858 ) | ( n10048 & n12860 ) | ( ~n12858 & n12860 ) ;
  assign n12864 = ( ~n3916 & n4032 ) | ( ~n3916 & n8827 ) | ( n4032 & n8827 ) ;
  assign n12865 = ( n3378 & ~n6767 ) | ( n3378 & n12864 ) | ( ~n6767 & n12864 ) ;
  assign n12862 = n9834 ^ n5424 ^ n2699 ;
  assign n12863 = n2880 & n12862 ;
  assign n12866 = n12865 ^ n12863 ^ 1'b0 ;
  assign n12867 = n11714 ^ n2268 ^ 1'b0 ;
  assign n12868 = n5793 & n12867 ;
  assign n12869 = ( ~n7242 & n7907 ) | ( ~n7242 & n12868 ) | ( n7907 & n12868 ) ;
  assign n12870 = ( n2499 & n12866 ) | ( n2499 & n12869 ) | ( n12866 & n12869 ) ;
  assign n12871 = n5410 ^ n4974 ^ n1868 ;
  assign n12872 = ( n2810 & ~n6462 ) | ( n2810 & n12871 ) | ( ~n6462 & n12871 ) ;
  assign n12875 = n7926 ^ n7675 ^ n3111 ;
  assign n12873 = ~n175 & n3686 ;
  assign n12874 = n7187 & n12873 ;
  assign n12876 = n12875 ^ n12874 ^ n8393 ;
  assign n12877 = n6073 ^ n4911 ^ n2289 ;
  assign n12878 = n6673 ^ n3336 ^ n2045 ;
  assign n12879 = n708 & ~n2032 ;
  assign n12880 = n12879 ^ n1726 ^ 1'b0 ;
  assign n12881 = n12880 ^ n10328 ^ n2265 ;
  assign n12882 = n11965 ^ n416 ^ 1'b0 ;
  assign n12883 = ~n10736 & n12882 ;
  assign n12884 = n6951 ^ n1198 ^ 1'b0 ;
  assign n12885 = ~n2808 & n12884 ;
  assign n12886 = ( ~n2699 & n3137 ) | ( ~n2699 & n12885 ) | ( n3137 & n12885 ) ;
  assign n12887 = ( n12881 & n12883 ) | ( n12881 & n12886 ) | ( n12883 & n12886 ) ;
  assign n12888 = ( ~n12877 & n12878 ) | ( ~n12877 & n12887 ) | ( n12878 & n12887 ) ;
  assign n12889 = n12888 ^ n7779 ^ n1008 ;
  assign n12890 = n6143 | n12889 ;
  assign n12891 = n12890 ^ n9214 ^ 1'b0 ;
  assign n12892 = n6312 ^ n3334 ^ n2592 ;
  assign n12893 = ( n525 & n2084 ) | ( n525 & n2733 ) | ( n2084 & n2733 ) ;
  assign n12894 = ( n11813 & n12892 ) | ( n11813 & n12893 ) | ( n12892 & n12893 ) ;
  assign n12895 = n12894 ^ n7922 ^ n4883 ;
  assign n12896 = n883 | n2822 ;
  assign n12897 = n12896 ^ n6241 ^ 1'b0 ;
  assign n12898 = ( n5702 & n12895 ) | ( n5702 & n12897 ) | ( n12895 & n12897 ) ;
  assign n12899 = ( ~n8666 & n9931 ) | ( ~n8666 & n12898 ) | ( n9931 & n12898 ) ;
  assign n12900 = ( n1086 & ~n9414 ) | ( n1086 & n10669 ) | ( ~n9414 & n10669 ) ;
  assign n12901 = n12900 ^ n5244 ^ n3782 ;
  assign n12902 = n7674 ^ n3835 ^ 1'b0 ;
  assign n12903 = n2591 & ~n12902 ;
  assign n12904 = ~n12003 & n12903 ;
  assign n12905 = n859 & ~n2025 ;
  assign n12906 = ( n9337 & n10878 ) | ( n9337 & ~n11709 ) | ( n10878 & ~n11709 ) ;
  assign n12907 = n9891 ^ n4934 ^ x84 ;
  assign n12908 = n12907 ^ n11294 ^ 1'b0 ;
  assign n12911 = n9618 ^ n6479 ^ n2762 ;
  assign n12909 = n318 & ~n6430 ;
  assign n12910 = ~n5142 & n12909 ;
  assign n12912 = n12911 ^ n12910 ^ n9621 ;
  assign n12913 = ( ~n483 & n3488 ) | ( ~n483 & n9964 ) | ( n3488 & n9964 ) ;
  assign n12914 = n12913 ^ n1167 ^ 1'b0 ;
  assign n12915 = n12914 ^ n8649 ^ 1'b0 ;
  assign n12916 = ( n2435 & n9044 ) | ( n2435 & n10120 ) | ( n9044 & n10120 ) ;
  assign n12917 = ( n2958 & ~n3580 ) | ( n2958 & n12916 ) | ( ~n3580 & n12916 ) ;
  assign n12918 = n10071 ^ n9811 ^ n3509 ;
  assign n12919 = n5898 ^ n5350 ^ n1195 ;
  assign n12920 = ( n9224 & ~n12918 ) | ( n9224 & n12919 ) | ( ~n12918 & n12919 ) ;
  assign n12922 = ~n2023 & n3605 ;
  assign n12923 = n12922 ^ n1796 ^ 1'b0 ;
  assign n12924 = n12923 ^ n11823 ^ n3943 ;
  assign n12925 = n12924 ^ n1363 ^ n449 ;
  assign n12921 = n7644 | n8459 ;
  assign n12926 = n12925 ^ n12921 ^ 1'b0 ;
  assign n12927 = ( ~n461 & n4161 ) | ( ~n461 & n11279 ) | ( n4161 & n11279 ) ;
  assign n12929 = x2 | n195 ;
  assign n12928 = ( n1054 & ~n1539 ) | ( n1054 & n7031 ) | ( ~n1539 & n7031 ) ;
  assign n12930 = n12929 ^ n12928 ^ n3844 ;
  assign n12931 = n12930 ^ n9865 ^ n3416 ;
  assign n12932 = n752 | n1898 ;
  assign n12933 = ( n8544 & ~n11792 ) | ( n8544 & n12932 ) | ( ~n11792 & n12932 ) ;
  assign n12934 = n1711 ^ n1433 ^ n1093 ;
  assign n12935 = ( n1810 & ~n4828 ) | ( n1810 & n12934 ) | ( ~n4828 & n12934 ) ;
  assign n12936 = n10195 ^ n8568 ^ n7536 ;
  assign n12937 = n12936 ^ n4729 ^ n1791 ;
  assign n12941 = n1942 ^ n924 ^ 1'b0 ;
  assign n12942 = ~n1527 & n12941 ;
  assign n12943 = n12942 ^ n6767 ^ n4840 ;
  assign n12938 = n1501 | n6029 ;
  assign n12939 = n12938 ^ n4009 ^ 1'b0 ;
  assign n12940 = ( n4742 & n11484 ) | ( n4742 & ~n12939 ) | ( n11484 & ~n12939 ) ;
  assign n12944 = n12943 ^ n12940 ^ 1'b0 ;
  assign n12945 = n5485 ^ n5001 ^ n4560 ;
  assign n12946 = ( ~n2230 & n8948 ) | ( ~n2230 & n11650 ) | ( n8948 & n11650 ) ;
  assign n12947 = ( ~n10446 & n12945 ) | ( ~n10446 & n12946 ) | ( n12945 & n12946 ) ;
  assign n12948 = n1044 & n12296 ;
  assign n12949 = ( n3260 & n12803 ) | ( n3260 & ~n12948 ) | ( n12803 & ~n12948 ) ;
  assign n12950 = ( n12151 & n12947 ) | ( n12151 & ~n12949 ) | ( n12947 & ~n12949 ) ;
  assign n12951 = n12290 ^ n11450 ^ n1361 ;
  assign n12952 = ( n7530 & ~n8578 ) | ( n7530 & n12951 ) | ( ~n8578 & n12951 ) ;
  assign n12953 = n10148 ^ n7979 ^ n1822 ;
  assign n12954 = n12953 ^ n2964 ^ n986 ;
  assign n12959 = ( ~n3500 & n5802 ) | ( ~n3500 & n6657 ) | ( n5802 & n6657 ) ;
  assign n12956 = n12504 ^ n2889 ^ 1'b0 ;
  assign n12957 = ( n3186 & ~n7447 ) | ( n3186 & n7735 ) | ( ~n7447 & n7735 ) ;
  assign n12958 = ( ~n12151 & n12956 ) | ( ~n12151 & n12957 ) | ( n12956 & n12957 ) ;
  assign n12955 = ~x11 & n9632 ;
  assign n12960 = n12959 ^ n12958 ^ n12955 ;
  assign n12961 = n12744 ^ n1448 ^ 1'b0 ;
  assign n12962 = n12961 ^ n4624 ^ n1513 ;
  assign n12963 = n12962 ^ n8156 ^ n1493 ;
  assign n12964 = ( n1135 & n2688 ) | ( n1135 & n12963 ) | ( n2688 & n12963 ) ;
  assign n12967 = n11161 ^ n9226 ^ n185 ;
  assign n12968 = ( n129 & n4043 ) | ( n129 & n12967 ) | ( n4043 & n12967 ) ;
  assign n12965 = ( ~n1016 & n5571 ) | ( ~n1016 & n10048 ) | ( n5571 & n10048 ) ;
  assign n12966 = n12965 ^ n1087 ^ n915 ;
  assign n12969 = n12968 ^ n12966 ^ n6403 ;
  assign n12970 = ( n2257 & ~n4721 ) | ( n2257 & n7635 ) | ( ~n4721 & n7635 ) ;
  assign n12971 = ( n1675 & n4755 ) | ( n1675 & ~n12970 ) | ( n4755 & ~n12970 ) ;
  assign n12972 = ( n460 & ~n4006 ) | ( n460 & n12971 ) | ( ~n4006 & n12971 ) ;
  assign n12973 = n4571 ^ n3294 ^ n1254 ;
  assign n12974 = n7998 ^ n5881 ^ 1'b0 ;
  assign n12975 = n12973 & n12974 ;
  assign n12976 = n4588 | n12975 ;
  assign n12977 = n5581 & n12976 ;
  assign n12978 = n12977 ^ n459 ^ 1'b0 ;
  assign n12979 = n4818 ^ n4717 ^ n2185 ;
  assign n12980 = n6226 & ~n12979 ;
  assign n12981 = n12980 ^ n10499 ^ n9975 ;
  assign n12982 = ( ~n3011 & n6489 ) | ( ~n3011 & n12885 ) | ( n6489 & n12885 ) ;
  assign n12983 = n3190 & n9326 ;
  assign n12984 = n12983 ^ n12880 ^ n10177 ;
  assign n12988 = n10720 ^ n8434 ^ n6839 ;
  assign n12985 = n10452 ^ n7864 ^ n7028 ;
  assign n12986 = n12985 ^ n7849 ^ n2900 ;
  assign n12987 = ~n1393 & n12986 ;
  assign n12989 = n12988 ^ n12987 ^ 1'b0 ;
  assign n12991 = n2062 & ~n3958 ;
  assign n12992 = n4135 & n12991 ;
  assign n12993 = n12992 ^ n8870 ^ n5455 ;
  assign n12990 = n10074 | n11649 ;
  assign n12994 = n12993 ^ n12990 ^ 1'b0 ;
  assign n12995 = n12994 ^ n7563 ^ 1'b0 ;
  assign n12996 = ( n1545 & n1944 ) | ( n1545 & ~n2851 ) | ( n1944 & ~n2851 ) ;
  assign n12997 = ( ~n232 & n7876 ) | ( ~n232 & n12996 ) | ( n7876 & n12996 ) ;
  assign n12998 = ( n5392 & n12931 ) | ( n5392 & ~n12997 ) | ( n12931 & ~n12997 ) ;
  assign n12999 = ( n2428 & n5979 ) | ( n2428 & n12180 ) | ( n5979 & n12180 ) ;
  assign n13000 = ( n4260 & n12193 ) | ( n4260 & ~n12999 ) | ( n12193 & ~n12999 ) ;
  assign n13001 = n573 & n4548 ;
  assign n13002 = n13001 ^ n2713 ^ 1'b0 ;
  assign n13003 = n13002 ^ n11121 ^ n3171 ;
  assign n13004 = n13003 ^ n8869 ^ 1'b0 ;
  assign n13005 = n11137 | n13004 ;
  assign n13006 = n13005 ^ n8970 ^ n7452 ;
  assign n13007 = n13006 ^ n7441 ^ n775 ;
  assign n13008 = n13007 ^ n7296 ^ n3355 ;
  assign n13009 = ( n1244 & n3147 ) | ( n1244 & ~n5024 ) | ( n3147 & ~n5024 ) ;
  assign n13010 = n13009 ^ n10209 ^ n7112 ;
  assign n13011 = n13010 ^ n10658 ^ n7009 ;
  assign n13012 = ( n465 & ~n3585 ) | ( n465 & n8816 ) | ( ~n3585 & n8816 ) ;
  assign n13013 = ( n10187 & n13011 ) | ( n10187 & n13012 ) | ( n13011 & n13012 ) ;
  assign n13014 = n2786 & ~n8710 ;
  assign n13015 = n13014 ^ n3494 ^ n458 ;
  assign n13016 = n4835 & ~n13015 ;
  assign n13017 = n4414 ^ x98 ^ 1'b0 ;
  assign n13018 = n13017 ^ n4697 ^ n3151 ;
  assign n13019 = n8718 ^ n4571 ^ 1'b0 ;
  assign n13020 = n13018 & n13019 ;
  assign n13021 = ( ~n456 & n1821 ) | ( ~n456 & n12025 ) | ( n1821 & n12025 ) ;
  assign n13022 = n13021 ^ n9819 ^ n4003 ;
  assign n13023 = n13022 ^ n4448 ^ n576 ;
  assign n13024 = n7614 ^ n6620 ^ n6396 ;
  assign n13025 = n4539 & n6203 ;
  assign n13026 = n10764 ^ n6414 ^ n3689 ;
  assign n13027 = n11425 ^ n9516 ^ n3579 ;
  assign n13028 = ( n1397 & ~n13026 ) | ( n1397 & n13027 ) | ( ~n13026 & n13027 ) ;
  assign n13029 = ( n12495 & ~n13025 ) | ( n12495 & n13028 ) | ( ~n13025 & n13028 ) ;
  assign n13030 = n12496 ^ n12384 ^ n4418 ;
  assign n13031 = n13030 ^ n3208 ^ 1'b0 ;
  assign n13032 = ( n1904 & n3156 ) | ( n1904 & n13031 ) | ( n3156 & n13031 ) ;
  assign n13033 = n13032 ^ n5733 ^ n1264 ;
  assign n13035 = ( n341 & n4816 ) | ( n341 & ~n5131 ) | ( n4816 & ~n5131 ) ;
  assign n13034 = ( n767 & n1319 ) | ( n767 & ~n2816 ) | ( n1319 & ~n2816 ) ;
  assign n13036 = n13035 ^ n13034 ^ n7240 ;
  assign n13037 = n4920 | n13036 ;
  assign n13038 = n10140 ^ n5134 ^ n257 ;
  assign n13039 = n8096 ^ n7616 ^ 1'b0 ;
  assign n13040 = n13038 & ~n13039 ;
  assign n13041 = n12620 & n13040 ;
  assign n13050 = n11071 ^ n6113 ^ 1'b0 ;
  assign n13051 = ( ~x17 & n7863 ) | ( ~x17 & n13050 ) | ( n7863 & n13050 ) ;
  assign n13047 = ( n1289 & n3753 ) | ( n1289 & n8900 ) | ( n3753 & n8900 ) ;
  assign n13048 = ( ~n2129 & n2497 ) | ( ~n2129 & n13047 ) | ( n2497 & n13047 ) ;
  assign n13049 = n13048 ^ n3732 ^ 1'b0 ;
  assign n13052 = n13051 ^ n13049 ^ n2644 ;
  assign n13042 = n4336 ^ n4190 ^ x62 ;
  assign n13043 = n7671 ^ n6422 ^ 1'b0 ;
  assign n13044 = n13042 | n13043 ;
  assign n13045 = ( n5587 & n7757 ) | ( n5587 & ~n8628 ) | ( n7757 & ~n8628 ) ;
  assign n13046 = n13044 | n13045 ;
  assign n13053 = n13052 ^ n13046 ^ 1'b0 ;
  assign n13054 = n11712 ^ n6148 ^ 1'b0 ;
  assign n13055 = ( n2468 & ~n10976 ) | ( n2468 & n13054 ) | ( ~n10976 & n13054 ) ;
  assign n13056 = n3195 & ~n13055 ;
  assign n13057 = ( ~n2612 & n13053 ) | ( ~n2612 & n13056 ) | ( n13053 & n13056 ) ;
  assign n13058 = n2591 | n6521 ;
  assign n13059 = n13058 ^ n9588 ^ n8983 ;
  assign n13060 = n11320 ^ n1189 ^ 1'b0 ;
  assign n13065 = ~n3335 & n9811 ;
  assign n13066 = n887 & n13065 ;
  assign n13067 = n4280 | n13066 ;
  assign n13061 = n5940 ^ n3035 ^ n1229 ;
  assign n13062 = n11001 ^ n7706 ^ n6920 ;
  assign n13063 = ~n13061 & n13062 ;
  assign n13064 = n2570 & n13063 ;
  assign n13068 = n13067 ^ n13064 ^ n7862 ;
  assign n13069 = n6771 & ~n7207 ;
  assign n13070 = n13069 ^ n2808 ^ 1'b0 ;
  assign n13071 = ~n5675 & n10379 ;
  assign n13072 = n2487 & n13071 ;
  assign n13074 = n3507 ^ n1133 ^ 1'b0 ;
  assign n13073 = n8213 ^ n2588 ^ 1'b0 ;
  assign n13075 = n13074 ^ n13073 ^ n4042 ;
  assign n13076 = n13072 & n13075 ;
  assign n13077 = n12364 ^ n4901 ^ 1'b0 ;
  assign n13078 = n13077 ^ n5008 ^ n1009 ;
  assign n13079 = ( n1886 & n3566 ) | ( n1886 & n5199 ) | ( n3566 & n5199 ) ;
  assign n13080 = n497 & n6769 ;
  assign n13081 = n6337 & n13080 ;
  assign n13082 = n3682 | n13081 ;
  assign n13083 = ( n7561 & n7883 ) | ( n7561 & ~n13082 ) | ( n7883 & ~n13082 ) ;
  assign n13084 = ( n442 & n3030 ) | ( n442 & ~n13083 ) | ( n3030 & ~n13083 ) ;
  assign n13085 = n13084 ^ n3118 ^ n1813 ;
  assign n13086 = ( ~n3423 & n13079 ) | ( ~n3423 & n13085 ) | ( n13079 & n13085 ) ;
  assign n13088 = n10818 ^ n2566 ^ n1576 ;
  assign n13087 = n662 & n11123 ;
  assign n13089 = n13088 ^ n13087 ^ n597 ;
  assign n13090 = n3582 ^ n3568 ^ x22 ;
  assign n13091 = n13090 ^ n4628 ^ 1'b0 ;
  assign n13092 = ( n5129 & n5752 ) | ( n5129 & ~n13091 ) | ( n5752 & ~n13091 ) ;
  assign n13093 = n6013 & n6486 ;
  assign n13094 = ~n5878 & n13093 ;
  assign n13095 = n1225 & ~n8329 ;
  assign n13096 = n11498 & n13095 ;
  assign n13097 = n13096 ^ n8161 ^ n3143 ;
  assign n13098 = ~n9893 & n13097 ;
  assign n13099 = ( ~n11650 & n13094 ) | ( ~n11650 & n13098 ) | ( n13094 & n13098 ) ;
  assign n13100 = n8115 ^ n6293 ^ n6210 ;
  assign n13101 = n4247 & n13100 ;
  assign n13102 = n9669 ^ n1496 ^ n925 ;
  assign n13103 = ( n2536 & n5190 ) | ( n2536 & ~n5595 ) | ( n5190 & ~n5595 ) ;
  assign n13104 = n1499 ^ n809 ^ n163 ;
  assign n13105 = ~n2569 & n13104 ;
  assign n13106 = n13105 ^ n3061 ^ 1'b0 ;
  assign n13107 = ~n1248 & n4460 ;
  assign n13108 = n13106 & n13107 ;
  assign n13109 = n3729 & ~n13108 ;
  assign n13110 = n13109 ^ n2835 ^ 1'b0 ;
  assign n13111 = ( n13102 & ~n13103 ) | ( n13102 & n13110 ) | ( ~n13103 & n13110 ) ;
  assign n13112 = n7494 ^ n4866 ^ n745 ;
  assign n13116 = n2665 ^ n1573 ^ n735 ;
  assign n13117 = ( n4083 & n7322 ) | ( n4083 & ~n13116 ) | ( n7322 & ~n13116 ) ;
  assign n13113 = n6283 ^ n4648 ^ n3137 ;
  assign n13114 = ( n8334 & n10260 ) | ( n8334 & ~n13113 ) | ( n10260 & ~n13113 ) ;
  assign n13115 = ~n6045 & n13114 ;
  assign n13118 = n13117 ^ n13115 ^ 1'b0 ;
  assign n13119 = n11023 ^ n9790 ^ n2076 ;
  assign n13120 = n3728 ^ n1005 ^ n470 ;
  assign n13121 = ( n6299 & n12803 ) | ( n6299 & n13120 ) | ( n12803 & n13120 ) ;
  assign n13122 = n7817 ^ n1473 ^ n477 ;
  assign n13123 = n2769 ^ n186 ^ x38 ;
  assign n13124 = n12946 & ~n13123 ;
  assign n13125 = ~n285 & n13124 ;
  assign n13126 = ( n1406 & ~n7458 ) | ( n1406 & n13125 ) | ( ~n7458 & n13125 ) ;
  assign n13127 = n9750 & ~n13126 ;
  assign n13128 = n13127 ^ n13009 ^ 1'b0 ;
  assign n13129 = n4666 & ~n13128 ;
  assign n13130 = n352 & n13129 ;
  assign n13131 = ( ~n5749 & n7154 ) | ( ~n5749 & n8202 ) | ( n7154 & n8202 ) ;
  assign n13132 = ( n2405 & n5452 ) | ( n2405 & ~n13131 ) | ( n5452 & ~n13131 ) ;
  assign n13133 = n10657 ^ n2551 ^ n875 ;
  assign n13135 = ~n2971 & n4456 ;
  assign n13134 = n1828 | n3338 ;
  assign n13136 = n13135 ^ n13134 ^ 1'b0 ;
  assign n13137 = n13136 ^ n1996 ^ 1'b0 ;
  assign n13138 = n5868 ^ n2609 ^ n448 ;
  assign n13139 = ( n5412 & n12052 ) | ( n5412 & n13138 ) | ( n12052 & n13138 ) ;
  assign n13140 = n13139 ^ n11136 ^ n8134 ;
  assign n13141 = ~n4682 & n8149 ;
  assign n13142 = ( n12760 & n13140 ) | ( n12760 & ~n13141 ) | ( n13140 & ~n13141 ) ;
  assign n13144 = n2074 ^ n1694 ^ 1'b0 ;
  assign n13143 = n4718 ^ n4448 ^ n2801 ;
  assign n13145 = n13144 ^ n13143 ^ n4514 ;
  assign n13147 = n6653 ^ n2344 ^ 1'b0 ;
  assign n13146 = n12795 ^ n929 ^ 1'b0 ;
  assign n13148 = n13147 ^ n13146 ^ n5630 ;
  assign n13149 = n3967 & ~n11871 ;
  assign n13150 = n13149 ^ n1944 ^ 1'b0 ;
  assign n13151 = ( n7951 & ~n12908 ) | ( n7951 & n13150 ) | ( ~n12908 & n13150 ) ;
  assign n13152 = n1492 ^ x47 ^ 1'b0 ;
  assign n13153 = n13152 ^ n7176 ^ n1212 ;
  assign n13154 = n5312 ^ n3519 ^ n1704 ;
  assign n13155 = n13153 | n13154 ;
  assign n13156 = n10878 | n13155 ;
  assign n13157 = n13156 ^ n12565 ^ n1528 ;
  assign n13159 = n2116 & n3263 ;
  assign n13160 = n13159 ^ n2688 ^ 1'b0 ;
  assign n13158 = n3387 & ~n5582 ;
  assign n13161 = n13160 ^ n13158 ^ 1'b0 ;
  assign n13162 = ( n1364 & n5163 ) | ( n1364 & ~n10292 ) | ( n5163 & ~n10292 ) ;
  assign n13163 = n4189 ^ n2445 ^ 1'b0 ;
  assign n13164 = n8603 & ~n13163 ;
  assign n13165 = ( x28 & n3398 ) | ( x28 & ~n13164 ) | ( n3398 & ~n13164 ) ;
  assign n13166 = ( n9356 & n13162 ) | ( n9356 & n13165 ) | ( n13162 & n13165 ) ;
  assign n13167 = n13166 ^ n12496 ^ 1'b0 ;
  assign n13168 = n9170 ^ n4217 ^ 1'b0 ;
  assign n13169 = n13168 ^ n3171 ^ 1'b0 ;
  assign n13170 = ( ~n1580 & n6516 ) | ( ~n1580 & n13169 ) | ( n6516 & n13169 ) ;
  assign n13171 = n13170 ^ n3313 ^ n2326 ;
  assign n13176 = n4494 ^ n3185 ^ n912 ;
  assign n13172 = ( n1458 & n6556 ) | ( n1458 & n10610 ) | ( n6556 & n10610 ) ;
  assign n13173 = ( ~n5372 & n8213 ) | ( ~n5372 & n13172 ) | ( n8213 & n13172 ) ;
  assign n13174 = n13173 ^ n5920 ^ n4587 ;
  assign n13175 = ( n7561 & ~n8260 ) | ( n7561 & n13174 ) | ( ~n8260 & n13174 ) ;
  assign n13177 = n13176 ^ n13175 ^ n6923 ;
  assign n13178 = ( n4080 & n13171 ) | ( n4080 & n13177 ) | ( n13171 & n13177 ) ;
  assign n13179 = ~n5181 & n10971 ;
  assign n13180 = n13179 ^ n3380 ^ 1'b0 ;
  assign n13181 = n13180 ^ n10758 ^ n9841 ;
  assign n13183 = ~n671 & n4053 ;
  assign n13184 = n13183 ^ n4346 ^ n3369 ;
  assign n13182 = n909 | n2971 ;
  assign n13185 = n13184 ^ n13182 ^ n7098 ;
  assign n13186 = n2572 | n4387 ;
  assign n13187 = n13186 ^ n3933 ^ 1'b0 ;
  assign n13188 = n7776 ^ n3569 ^ n2691 ;
  assign n13189 = ( n3327 & n13187 ) | ( n3327 & n13188 ) | ( n13187 & n13188 ) ;
  assign n13191 = n827 & ~n1937 ;
  assign n13190 = n10027 ^ n6495 ^ n2761 ;
  assign n13192 = n13191 ^ n13190 ^ n977 ;
  assign n13193 = n2485 & ~n6078 ;
  assign n13194 = n13193 ^ n9763 ^ 1'b0 ;
  assign n13195 = n13194 ^ n8296 ^ n4961 ;
  assign n13196 = ( n9303 & n13192 ) | ( n9303 & n13195 ) | ( n13192 & n13195 ) ;
  assign n13197 = n13196 ^ n9022 ^ n7375 ;
  assign n13198 = ( n13185 & ~n13189 ) | ( n13185 & n13197 ) | ( ~n13189 & n13197 ) ;
  assign n13199 = ( n3206 & n5298 ) | ( n3206 & n10733 ) | ( n5298 & n10733 ) ;
  assign n13200 = ( n5989 & n6055 ) | ( n5989 & n13199 ) | ( n6055 & n13199 ) ;
  assign n13201 = ( n155 & n6691 ) | ( n155 & ~n13200 ) | ( n6691 & ~n13200 ) ;
  assign n13202 = ( n634 & ~n3138 ) | ( n634 & n12315 ) | ( ~n3138 & n12315 ) ;
  assign n13203 = n5425 ^ n970 ^ 1'b0 ;
  assign n13204 = n6769 & ~n13203 ;
  assign n13205 = n5784 ^ n1882 ^ n869 ;
  assign n13206 = ( n161 & n1759 ) | ( n161 & n13136 ) | ( n1759 & n13136 ) ;
  assign n13207 = ~n13205 & n13206 ;
  assign n13208 = n11712 & n13207 ;
  assign n13210 = ( n5573 & ~n5713 ) | ( n5573 & n8348 ) | ( ~n5713 & n8348 ) ;
  assign n13209 = n10982 ^ n3685 ^ n676 ;
  assign n13211 = n13210 ^ n13209 ^ n3823 ;
  assign n13212 = ( ~n3885 & n9303 ) | ( ~n3885 & n11478 ) | ( n9303 & n11478 ) ;
  assign n13213 = n9812 ^ n9456 ^ n1773 ;
  assign n13214 = ~n143 & n12346 ;
  assign n13215 = ~n13213 & n13214 ;
  assign n13218 = n8532 ^ n6285 ^ n6253 ;
  assign n13217 = n3385 ^ n1279 ^ 1'b0 ;
  assign n13216 = ( n5406 & n6499 ) | ( n5406 & ~n11284 ) | ( n6499 & ~n11284 ) ;
  assign n13219 = n13218 ^ n13217 ^ n13216 ;
  assign n13223 = ( n4502 & n4580 ) | ( n4502 & ~n10985 ) | ( n4580 & ~n10985 ) ;
  assign n13220 = n6689 ^ n4096 ^ n3038 ;
  assign n13221 = n11657 ^ n5356 ^ n337 ;
  assign n13222 = ( n321 & n13220 ) | ( n321 & n13221 ) | ( n13220 & n13221 ) ;
  assign n13224 = n13223 ^ n13222 ^ n1395 ;
  assign n13225 = n9418 & n11857 ;
  assign n13226 = n2346 & n3920 ;
  assign n13227 = n11873 & ~n13226 ;
  assign n13228 = ~x119 & n13227 ;
  assign n13230 = ( n838 & n901 ) | ( n838 & n1401 ) | ( n901 & n1401 ) ;
  assign n13229 = n2484 | n12774 ;
  assign n13231 = n13230 ^ n13229 ^ 1'b0 ;
  assign n13232 = n12729 ^ n8178 ^ n3172 ;
  assign n13233 = ( ~n872 & n6686 ) | ( ~n872 & n13232 ) | ( n6686 & n13232 ) ;
  assign n13234 = n564 | n2413 ;
  assign n13235 = n3799 | n13234 ;
  assign n13236 = ( n533 & n13088 ) | ( n533 & n13235 ) | ( n13088 & n13235 ) ;
  assign n13237 = n13236 ^ n2994 ^ 1'b0 ;
  assign n13238 = n13237 ^ n10229 ^ 1'b0 ;
  assign n13239 = ( n520 & ~n4116 ) | ( n520 & n10957 ) | ( ~n4116 & n10957 ) ;
  assign n13240 = n13239 ^ n8694 ^ 1'b0 ;
  assign n13241 = n12481 ^ n9409 ^ n688 ;
  assign n13242 = n12534 ^ n7204 ^ n4403 ;
  assign n13243 = n13242 ^ n1918 ^ n1765 ;
  assign n13244 = n13243 ^ n10868 ^ n8777 ;
  assign n13245 = n4755 & ~n7328 ;
  assign n13246 = n2164 & ~n6280 ;
  assign n13247 = n13246 ^ n875 ^ 1'b0 ;
  assign n13248 = n2632 & n13247 ;
  assign n13249 = n13248 ^ n11416 ^ 1'b0 ;
  assign n13250 = n13245 & n13249 ;
  assign n13251 = n13250 ^ n8361 ^ 1'b0 ;
  assign n13252 = ( n1853 & n4157 ) | ( n1853 & n4382 ) | ( n4157 & n4382 ) ;
  assign n13253 = n13252 ^ n6951 ^ n142 ;
  assign n13254 = n13253 ^ n8534 ^ 1'b0 ;
  assign n13255 = ~n7690 & n13254 ;
  assign n13256 = ( n5630 & ~n9648 ) | ( n5630 & n11321 ) | ( ~n9648 & n11321 ) ;
  assign n13257 = ( ~x57 & n275 ) | ( ~x57 & n11743 ) | ( n275 & n11743 ) ;
  assign n13258 = ( n2573 & ~n5879 ) | ( n2573 & n6931 ) | ( ~n5879 & n6931 ) ;
  assign n13259 = ( ~n7469 & n10546 ) | ( ~n7469 & n13258 ) | ( n10546 & n13258 ) ;
  assign n13260 = ( n159 & ~n2512 ) | ( n159 & n6670 ) | ( ~n2512 & n6670 ) ;
  assign n13261 = n11615 ^ n5293 ^ n2861 ;
  assign n13262 = n6378 ^ n5005 ^ 1'b0 ;
  assign n13263 = n13261 & n13262 ;
  assign n13264 = ( ~n281 & n12455 ) | ( ~n281 & n13263 ) | ( n12455 & n13263 ) ;
  assign n13265 = n3991 | n13264 ;
  assign n13266 = n13265 ^ n1105 ^ 1'b0 ;
  assign n13267 = n9316 ^ n5437 ^ n3637 ;
  assign n13268 = ( ~n13015 & n13266 ) | ( ~n13015 & n13267 ) | ( n13266 & n13267 ) ;
  assign n13269 = ( n5458 & n7993 ) | ( n5458 & ~n11075 ) | ( n7993 & ~n11075 ) ;
  assign n13275 = n4157 ^ n2515 ^ 1'b0 ;
  assign n13273 = n1387 | n3937 ;
  assign n13272 = n8653 ^ n7192 ^ n382 ;
  assign n13271 = ( n724 & n2711 ) | ( n724 & n10817 ) | ( n2711 & n10817 ) ;
  assign n13274 = n13273 ^ n13272 ^ n13271 ;
  assign n13276 = n13275 ^ n13274 ^ 1'b0 ;
  assign n13270 = n3897 | n13012 ;
  assign n13277 = n13276 ^ n13270 ^ 1'b0 ;
  assign n13278 = n7039 ^ n2346 ^ n179 ;
  assign n13279 = n13278 ^ n11910 ^ n11707 ;
  assign n13280 = ( n9498 & n10249 ) | ( n9498 & n13279 ) | ( n10249 & n13279 ) ;
  assign n13281 = n10628 ^ n6870 ^ 1'b0 ;
  assign n13282 = ~n1896 & n7893 ;
  assign n13283 = n13282 ^ n5989 ^ 1'b0 ;
  assign n13284 = n3949 | n13283 ;
  assign n13285 = ( n2487 & n5425 ) | ( n2487 & n7461 ) | ( n5425 & n7461 ) ;
  assign n13286 = ( n5991 & n11216 ) | ( n5991 & n13285 ) | ( n11216 & n13285 ) ;
  assign n13287 = n13286 ^ n12705 ^ 1'b0 ;
  assign n13288 = ~n1920 & n3766 ;
  assign n13289 = n13288 ^ n9639 ^ 1'b0 ;
  assign n13290 = ( n7278 & n8431 ) | ( n7278 & n13289 ) | ( n8431 & n13289 ) ;
  assign n13291 = n4407 ^ n1120 ^ 1'b0 ;
  assign n13292 = x73 & ~n13291 ;
  assign n13293 = n6948 ^ n3659 ^ n2910 ;
  assign n13294 = ( n3491 & n5060 ) | ( n3491 & n11411 ) | ( n5060 & n11411 ) ;
  assign n13295 = n7204 & ~n13294 ;
  assign n13296 = ( n13292 & ~n13293 ) | ( n13292 & n13295 ) | ( ~n13293 & n13295 ) ;
  assign n13297 = n11450 ^ n6413 ^ 1'b0 ;
  assign n13298 = n6426 ^ n988 ^ 1'b0 ;
  assign n13299 = n3039 | n13298 ;
  assign n13300 = ( n3042 & ~n3150 ) | ( n3042 & n5111 ) | ( ~n3150 & n5111 ) ;
  assign n13301 = ( n8338 & n13194 ) | ( n8338 & ~n13300 ) | ( n13194 & ~n13300 ) ;
  assign n13302 = ( n2958 & ~n13299 ) | ( n2958 & n13301 ) | ( ~n13299 & n13301 ) ;
  assign n13306 = n4025 ^ n3640 ^ 1'b0 ;
  assign n13307 = n13306 ^ n10171 ^ n3324 ;
  assign n13308 = n13307 ^ n4000 ^ n2624 ;
  assign n13303 = n12798 ^ n8018 ^ n732 ;
  assign n13304 = ~n4710 & n9210 ;
  assign n13305 = ~n13303 & n13304 ;
  assign n13309 = n13308 ^ n13305 ^ n10782 ;
  assign n13310 = n13309 ^ n5172 ^ 1'b0 ;
  assign n13311 = n850 | n13310 ;
  assign n13316 = ( n827 & n5360 ) | ( n827 & n5446 ) | ( n5360 & n5446 ) ;
  assign n13317 = ( n6804 & n10985 ) | ( n6804 & n13316 ) | ( n10985 & n13316 ) ;
  assign n13312 = n11864 ^ n7097 ^ 1'b0 ;
  assign n13313 = ( n133 & ~n1231 ) | ( n133 & n1765 ) | ( ~n1231 & n1765 ) ;
  assign n13314 = n13313 ^ n4037 ^ 1'b0 ;
  assign n13315 = n13312 | n13314 ;
  assign n13318 = n13317 ^ n13315 ^ n5769 ;
  assign n13319 = x58 & ~n13318 ;
  assign n13320 = n3143 & n13319 ;
  assign n13321 = n4581 ^ n3074 ^ n1796 ;
  assign n13322 = n13321 ^ n835 ^ 1'b0 ;
  assign n13323 = ~n3033 & n13322 ;
  assign n13324 = n7071 | n11999 ;
  assign n13325 = n2488 | n4950 ;
  assign n13326 = n3886 | n13325 ;
  assign n13327 = ( n1940 & ~n2716 ) | ( n1940 & n3600 ) | ( ~n2716 & n3600 ) ;
  assign n13328 = ( n6103 & ~n9095 ) | ( n6103 & n13327 ) | ( ~n9095 & n13327 ) ;
  assign n13329 = ( ~n6863 & n13326 ) | ( ~n6863 & n13328 ) | ( n13326 & n13328 ) ;
  assign n13330 = ( n13303 & ~n13324 ) | ( n13303 & n13329 ) | ( ~n13324 & n13329 ) ;
  assign n13331 = n5889 ^ n2028 ^ 1'b0 ;
  assign n13332 = ( ~n772 & n1024 ) | ( ~n772 & n11249 ) | ( n1024 & n11249 ) ;
  assign n13333 = n7411 & ~n12572 ;
  assign n13334 = n13333 ^ n5538 ^ 1'b0 ;
  assign n13335 = n13334 ^ n7493 ^ n841 ;
  assign n13336 = n4573 ^ n3210 ^ n2881 ;
  assign n13337 = ( n8966 & ~n9863 ) | ( n8966 & n13336 ) | ( ~n9863 & n13336 ) ;
  assign n13340 = n6789 ^ n5935 ^ n976 ;
  assign n13338 = n6740 ^ n6065 ^ n1174 ;
  assign n13339 = n10990 | n13338 ;
  assign n13341 = n13340 ^ n13339 ^ n1903 ;
  assign n13342 = n13341 ^ n4940 ^ n4371 ;
  assign n13343 = ~n9536 & n13342 ;
  assign n13344 = ( ~n2741 & n13337 ) | ( ~n2741 & n13343 ) | ( n13337 & n13343 ) ;
  assign n13347 = n3111 ^ n1416 ^ n932 ;
  assign n13345 = n12263 ^ n11869 ^ n7610 ;
  assign n13346 = n9436 & n13345 ;
  assign n13348 = n13347 ^ n13346 ^ 1'b0 ;
  assign n13349 = n3457 | n9897 ;
  assign n13350 = n13349 ^ n7320 ^ 1'b0 ;
  assign n13351 = n11601 ^ n8482 ^ n5291 ;
  assign n13352 = n13350 & n13351 ;
  assign n13353 = n13352 ^ n5627 ^ 1'b0 ;
  assign n13354 = ( n5618 & n5929 ) | ( n5618 & n8856 ) | ( n5929 & n8856 ) ;
  assign n13355 = n13354 ^ n12515 ^ n7143 ;
  assign n13356 = n6447 | n11292 ;
  assign n13357 = n13356 ^ n13072 ^ 1'b0 ;
  assign n13358 = n13357 ^ n8550 ^ 1'b0 ;
  assign n13359 = ( n5416 & n6116 ) | ( n5416 & ~n10615 ) | ( n6116 & ~n10615 ) ;
  assign n13360 = n960 & n13359 ;
  assign n13361 = ~n5852 & n13360 ;
  assign n13362 = n790 | n4091 ;
  assign n13363 = n4990 | n13362 ;
  assign n13368 = n892 & ~n3213 ;
  assign n13369 = n13368 ^ n4022 ^ 1'b0 ;
  assign n13364 = n6689 ^ n1398 ^ 1'b0 ;
  assign n13365 = ~n5340 & n13364 ;
  assign n13366 = n295 & n13365 ;
  assign n13367 = ~n11685 & n13366 ;
  assign n13370 = n13369 ^ n13367 ^ n6844 ;
  assign n13371 = n1973 ^ n871 ^ n867 ;
  assign n13372 = n634 | n3174 ;
  assign n13373 = n13371 & ~n13372 ;
  assign n13374 = n13373 ^ n8577 ^ n5000 ;
  assign n13375 = n10279 ^ n8344 ^ 1'b0 ;
  assign n13376 = ( n2630 & ~n13374 ) | ( n2630 & n13375 ) | ( ~n13374 & n13375 ) ;
  assign n13377 = n13376 ^ n10535 ^ n8433 ;
  assign n13378 = n5042 ^ n2876 ^ 1'b0 ;
  assign n13379 = ( n4929 & ~n7837 ) | ( n4929 & n13378 ) | ( ~n7837 & n13378 ) ;
  assign n13380 = ( ~n5153 & n9372 ) | ( ~n5153 & n13379 ) | ( n9372 & n13379 ) ;
  assign n13381 = ( n2943 & n13052 ) | ( n2943 & ~n13380 ) | ( n13052 & ~n13380 ) ;
  assign n13382 = n9712 ^ n2575 ^ n1481 ;
  assign n13383 = n6915 ^ n6400 ^ 1'b0 ;
  assign n13384 = n13383 ^ n3213 ^ n736 ;
  assign n13385 = n13384 ^ n11200 ^ n9514 ;
  assign n13386 = n1678 & n2821 ;
  assign n13387 = n13386 ^ n3150 ^ 1'b0 ;
  assign n13388 = n13387 ^ n5716 ^ n3134 ;
  assign n13389 = n13388 ^ n4562 ^ n4058 ;
  assign n13390 = n1987 & n11270 ;
  assign n13391 = n13389 & ~n13390 ;
  assign n13392 = ( ~n13382 & n13385 ) | ( ~n13382 & n13391 ) | ( n13385 & n13391 ) ;
  assign n13393 = ~n3982 & n7957 ;
  assign n13394 = n7348 ^ n2633 ^ n2036 ;
  assign n13395 = n5506 & n8947 ;
  assign n13396 = n13395 ^ n8940 ^ 1'b0 ;
  assign n13397 = n13396 ^ n8213 ^ 1'b0 ;
  assign n13398 = ( n2039 & ~n13394 ) | ( n2039 & n13397 ) | ( ~n13394 & n13397 ) ;
  assign n13399 = n2033 | n10071 ;
  assign n13400 = n13399 ^ n2472 ^ 1'b0 ;
  assign n13401 = ( n1557 & n5317 ) | ( n1557 & ~n13400 ) | ( n5317 & ~n13400 ) ;
  assign n13402 = n1866 ^ n1180 ^ 1'b0 ;
  assign n13403 = ( n850 & n4016 ) | ( n850 & ~n9390 ) | ( n4016 & ~n9390 ) ;
  assign n13404 = n13402 | n13403 ;
  assign n13405 = ( n3248 & ~n5462 ) | ( n3248 & n6369 ) | ( ~n5462 & n6369 ) ;
  assign n13406 = n10611 ^ n9544 ^ n7761 ;
  assign n13407 = ( n1862 & n13405 ) | ( n1862 & n13406 ) | ( n13405 & n13406 ) ;
  assign n13408 = n13407 ^ n7719 ^ n4978 ;
  assign n13409 = n5826 ^ n374 ^ 1'b0 ;
  assign n13410 = n2885 | n13409 ;
  assign n13411 = n2723 & ~n13410 ;
  assign n13412 = ( ~n1144 & n1472 ) | ( ~n1144 & n3971 ) | ( n1472 & n3971 ) ;
  assign n13413 = n13412 ^ n974 ^ n471 ;
  assign n13414 = n3563 ^ n3339 ^ 1'b0 ;
  assign n13415 = n8626 ^ n1146 ^ n1097 ;
  assign n13416 = ( n4124 & n11236 ) | ( n4124 & n13415 ) | ( n11236 & n13415 ) ;
  assign n13417 = ( n1907 & n9438 ) | ( n1907 & ~n13416 ) | ( n9438 & ~n13416 ) ;
  assign n13418 = n6407 & n6483 ;
  assign n13419 = ~n6513 & n13418 ;
  assign n13422 = n7933 ^ n3928 ^ n3434 ;
  assign n13420 = n12286 ^ n8097 ^ n6223 ;
  assign n13421 = n13420 ^ n1904 ^ x108 ;
  assign n13423 = n13422 ^ n13421 ^ n4844 ;
  assign n13424 = n10048 ^ n7753 ^ n3530 ;
  assign n13425 = n13424 ^ n6747 ^ n3787 ;
  assign n13430 = ( n3886 & n5667 ) | ( n3886 & ~n6951 ) | ( n5667 & ~n6951 ) ;
  assign n13426 = n8467 & n9618 ;
  assign n13427 = n13426 ^ n7849 ^ 1'b0 ;
  assign n13428 = ( n2396 & n10231 ) | ( n2396 & n13427 ) | ( n10231 & n13427 ) ;
  assign n13429 = n10509 | n13428 ;
  assign n13431 = n13430 ^ n13429 ^ 1'b0 ;
  assign n13440 = n6470 ^ n6379 ^ 1'b0 ;
  assign n13432 = n11174 ^ n2726 ^ 1'b0 ;
  assign n13433 = ~n2958 & n13432 ;
  assign n13434 = ( n2852 & ~n11751 ) | ( n2852 & n13433 ) | ( ~n11751 & n13433 ) ;
  assign n13435 = n8722 ^ n1970 ^ 1'b0 ;
  assign n13436 = n11616 ^ n5454 ^ n4098 ;
  assign n13437 = ( n2482 & ~n13435 ) | ( n2482 & n13436 ) | ( ~n13435 & n13436 ) ;
  assign n13438 = n13437 ^ n10693 ^ n9891 ;
  assign n13439 = ( n6696 & ~n13434 ) | ( n6696 & n13438 ) | ( ~n13434 & n13438 ) ;
  assign n13441 = n13440 ^ n13439 ^ n1230 ;
  assign n13449 = n6559 | n9104 ;
  assign n13447 = n7827 ^ x86 ^ 1'b0 ;
  assign n13448 = ~n3634 & n13447 ;
  assign n13442 = ( n2516 & n8985 ) | ( n2516 & ~n9061 ) | ( n8985 & ~n9061 ) ;
  assign n13443 = n13442 ^ n7060 ^ n129 ;
  assign n13444 = n13443 ^ n8561 ^ 1'b0 ;
  assign n13445 = n9610 | n13444 ;
  assign n13446 = ( ~n3176 & n9943 ) | ( ~n3176 & n13445 ) | ( n9943 & n13445 ) ;
  assign n13450 = n13449 ^ n13448 ^ n13446 ;
  assign n13451 = n6949 ^ n3605 ^ n3205 ;
  assign n13452 = ( ~n11385 & n12988 ) | ( ~n11385 & n13451 ) | ( n12988 & n13451 ) ;
  assign n13453 = n11883 ^ n3249 ^ n1108 ;
  assign n13454 = ( n474 & ~n4011 ) | ( n474 & n13453 ) | ( ~n4011 & n13453 ) ;
  assign n13455 = n10494 ^ n5367 ^ n1654 ;
  assign n13456 = n11125 ^ n9686 ^ n5726 ;
  assign n13457 = n12103 ^ n6318 ^ n3884 ;
  assign n13460 = n4494 & ~n4507 ;
  assign n13458 = ( ~n3710 & n4783 ) | ( ~n3710 & n5279 ) | ( n4783 & n5279 ) ;
  assign n13459 = ( n2565 & n12773 ) | ( n2565 & ~n13458 ) | ( n12773 & ~n13458 ) ;
  assign n13461 = n13460 ^ n13459 ^ n4590 ;
  assign n13462 = ( ~n1927 & n7848 ) | ( ~n1927 & n8734 ) | ( n7848 & n8734 ) ;
  assign n13463 = n13462 ^ n11093 ^ n5520 ;
  assign n13464 = ( n742 & n12163 ) | ( n742 & ~n13463 ) | ( n12163 & ~n13463 ) ;
  assign n13467 = n6046 ^ n4569 ^ n975 ;
  assign n13465 = n6188 ^ n5305 ^ 1'b0 ;
  assign n13466 = n2525 & ~n13465 ;
  assign n13468 = n13467 ^ n13466 ^ 1'b0 ;
  assign n13469 = ( n6055 & n9407 ) | ( n6055 & ~n13468 ) | ( n9407 & ~n13468 ) ;
  assign n13470 = n8604 ^ n2479 ^ n484 ;
  assign n13471 = ( n3617 & ~n6507 ) | ( n3617 & n10817 ) | ( ~n6507 & n10817 ) ;
  assign n13472 = ( ~n4530 & n11077 ) | ( ~n4530 & n13471 ) | ( n11077 & n13471 ) ;
  assign n13473 = n12508 ^ n4645 ^ x118 ;
  assign n13474 = n11759 ^ n4235 ^ n178 ;
  assign n13478 = n11456 ^ n9328 ^ n6720 ;
  assign n13475 = n9186 | n10210 ;
  assign n13476 = n7739 | n13475 ;
  assign n13477 = n5556 & n13476 ;
  assign n13479 = n13478 ^ n13477 ^ 1'b0 ;
  assign n13480 = n11557 ^ n2728 ^ n2557 ;
  assign n13481 = ( ~n373 & n5352 ) | ( ~n373 & n13480 ) | ( n5352 & n13480 ) ;
  assign n13482 = ( n1470 & n6220 ) | ( n1470 & n13481 ) | ( n6220 & n13481 ) ;
  assign n13483 = n3118 & n13482 ;
  assign n13487 = n8910 ^ n6241 ^ 1'b0 ;
  assign n13488 = n7526 & n13487 ;
  assign n13489 = ( n727 & n6905 ) | ( n727 & ~n11736 ) | ( n6905 & ~n11736 ) ;
  assign n13490 = n1230 ^ n1172 ^ n448 ;
  assign n13491 = n13490 ^ n12342 ^ n7563 ;
  assign n13492 = n13489 & ~n13491 ;
  assign n13493 = ~n13488 & n13492 ;
  assign n13494 = n966 ^ x104 ^ 1'b0 ;
  assign n13495 = ~n13493 & n13494 ;
  assign n13484 = n11748 ^ n7799 ^ n3879 ;
  assign n13485 = n13484 ^ n7389 ^ 1'b0 ;
  assign n13486 = ~n3659 & n13485 ;
  assign n13496 = n13495 ^ n13486 ^ n10294 ;
  assign n13497 = ( n2375 & n6808 ) | ( n2375 & n13496 ) | ( n6808 & n13496 ) ;
  assign n13498 = ( ~n3634 & n7166 ) | ( ~n3634 & n7531 ) | ( n7166 & n7531 ) ;
  assign n13499 = n13498 ^ n3927 ^ n2103 ;
  assign n13500 = ~n7688 & n13499 ;
  assign n13501 = n5803 ^ n775 ^ 1'b0 ;
  assign n13502 = n13500 | n13501 ;
  assign n13503 = ( n1013 & n10456 ) | ( n1013 & n13502 ) | ( n10456 & n13502 ) ;
  assign n13504 = ( n4508 & ~n4783 ) | ( n4508 & n5479 ) | ( ~n4783 & n5479 ) ;
  assign n13505 = n8149 & ~n13504 ;
  assign n13506 = n13505 ^ n8293 ^ 1'b0 ;
  assign n13507 = n7556 ^ n3469 ^ 1'b0 ;
  assign n13508 = n13507 ^ n3728 ^ n3050 ;
  assign n13509 = ( ~n958 & n2406 ) | ( ~n958 & n2882 ) | ( n2406 & n2882 ) ;
  assign n13510 = n13509 ^ n6558 ^ n4774 ;
  assign n13511 = n13510 ^ n12336 ^ 1'b0 ;
  assign n13512 = ~n1377 & n13511 ;
  assign n13513 = n12164 ^ n3949 ^ n763 ;
  assign n13514 = ( ~n2455 & n4772 ) | ( ~n2455 & n13513 ) | ( n4772 & n13513 ) ;
  assign n13526 = ( n691 & ~n842 ) | ( n691 & n2624 ) | ( ~n842 & n2624 ) ;
  assign n13516 = n6687 ^ n1534 ^ 1'b0 ;
  assign n13517 = n13516 ^ n6175 ^ n3973 ;
  assign n13518 = n6146 ^ n4879 ^ 1'b0 ;
  assign n13519 = n3135 & n13518 ;
  assign n13520 = n5247 & n11106 ;
  assign n13521 = ~n5145 & n13520 ;
  assign n13522 = n13521 ^ n1598 ^ 1'b0 ;
  assign n13523 = n13519 & n13522 ;
  assign n13524 = ( ~n11116 & n13517 ) | ( ~n11116 & n13523 ) | ( n13517 & n13523 ) ;
  assign n13525 = n13524 ^ n12101 ^ n565 ;
  assign n13527 = n13526 ^ n13525 ^ n2739 ;
  assign n13528 = n13527 ^ n13045 ^ n1719 ;
  assign n13515 = n12166 ^ n11827 ^ 1'b0 ;
  assign n13529 = n13528 ^ n13515 ^ n5112 ;
  assign n13530 = ~n5908 & n7154 ;
  assign n13531 = n3485 & n13530 ;
  assign n13532 = n6132 ^ n352 ^ 1'b0 ;
  assign n13533 = n13532 ^ n2922 ^ n2620 ;
  assign n13534 = n9945 ^ n4792 ^ 1'b0 ;
  assign n13536 = ( n6972 & ~n7325 ) | ( n6972 & n12255 ) | ( ~n7325 & n12255 ) ;
  assign n13535 = n1296 & n1581 ;
  assign n13537 = n13536 ^ n13535 ^ 1'b0 ;
  assign n13538 = n13537 ^ n11501 ^ x29 ;
  assign n13539 = ( n13533 & ~n13534 ) | ( n13533 & n13538 ) | ( ~n13534 & n13538 ) ;
  assign n13540 = n9344 ^ n5359 ^ 1'b0 ;
  assign n13541 = n13540 ^ n13403 ^ n5930 ;
  assign n13542 = n1159 & ~n3035 ;
  assign n13543 = n13542 ^ n265 ^ 1'b0 ;
  assign n13544 = n5977 ^ n5101 ^ n243 ;
  assign n13545 = ( ~n5705 & n11694 ) | ( ~n5705 & n13544 ) | ( n11694 & n13544 ) ;
  assign n13546 = n6365 | n9113 ;
  assign n13547 = n6914 ^ n4370 ^ 1'b0 ;
  assign n13548 = n937 & ~n13547 ;
  assign n13549 = n5880 ^ n2843 ^ 1'b0 ;
  assign n13550 = n13548 & n13549 ;
  assign n13551 = ~n3396 & n13550 ;
  assign n13552 = n13551 ^ n209 ^ 1'b0 ;
  assign n13553 = n13552 ^ n6480 ^ n3100 ;
  assign n13554 = ( n813 & n13546 ) | ( n813 & n13553 ) | ( n13546 & n13553 ) ;
  assign n13557 = n1647 & n3496 ;
  assign n13558 = n6420 ^ n195 ^ 1'b0 ;
  assign n13559 = ( ~n4217 & n13557 ) | ( ~n4217 & n13558 ) | ( n13557 & n13558 ) ;
  assign n13555 = ( n1894 & n3136 ) | ( n1894 & n4452 ) | ( n3136 & n4452 ) ;
  assign n13556 = n13555 ^ n1674 ^ 1'b0 ;
  assign n13560 = n13559 ^ n13556 ^ n1973 ;
  assign n13561 = ( n6199 & n9999 ) | ( n6199 & ~n12125 ) | ( n9999 & ~n12125 ) ;
  assign n13562 = n7532 ^ n7313 ^ n4468 ;
  assign n13563 = n381 | n3536 ;
  assign n13564 = n5419 & n7710 ;
  assign n13565 = n13564 ^ n977 ^ 1'b0 ;
  assign n13566 = ( ~n2043 & n2157 ) | ( ~n2043 & n5360 ) | ( n2157 & n5360 ) ;
  assign n13567 = n13566 ^ n3543 ^ n1201 ;
  assign n13568 = n8788 & n10934 ;
  assign n13569 = n13568 ^ n6152 ^ 1'b0 ;
  assign n13570 = ( ~n603 & n3271 ) | ( ~n603 & n7113 ) | ( n3271 & n7113 ) ;
  assign n13571 = n13570 ^ n12362 ^ n3302 ;
  assign n13572 = n7489 & n13571 ;
  assign n13573 = ( n8342 & n11144 ) | ( n8342 & n13572 ) | ( n11144 & n13572 ) ;
  assign n13574 = ( n480 & n4603 ) | ( n480 & ~n13573 ) | ( n4603 & ~n13573 ) ;
  assign n13575 = n10970 ^ n8360 ^ x123 ;
  assign n13576 = n461 & ~n11825 ;
  assign n13577 = n13576 ^ n10987 ^ 1'b0 ;
  assign n13578 = n6518 | n13577 ;
  assign n13579 = n9178 ^ n8532 ^ n5223 ;
  assign n13580 = n13033 ^ n4235 ^ n2573 ;
  assign n13583 = n8305 ^ n3873 ^ 1'b0 ;
  assign n13584 = n4395 & ~n13583 ;
  assign n13581 = n5849 ^ n3667 ^ 1'b0 ;
  assign n13582 = ( n2851 & n7543 ) | ( n2851 & ~n13581 ) | ( n7543 & ~n13581 ) ;
  assign n13585 = n13584 ^ n13582 ^ n1857 ;
  assign n13588 = n10701 ^ n7433 ^ n761 ;
  assign n13586 = n8589 & n9104 ;
  assign n13587 = n13586 ^ n10704 ^ 1'b0 ;
  assign n13589 = n13588 ^ n13587 ^ n780 ;
  assign n13590 = n6384 ^ n5390 ^ n667 ;
  assign n13591 = ( n10477 & ~n10546 ) | ( n10477 & n13590 ) | ( ~n10546 & n13590 ) ;
  assign n13592 = n7092 ^ n5740 ^ n3049 ;
  assign n13593 = n6173 & n13592 ;
  assign n13594 = n13593 ^ n10963 ^ 1'b0 ;
  assign n13595 = n13594 ^ n599 ^ 1'b0 ;
  assign n13596 = ( n272 & n2091 ) | ( n272 & n2139 ) | ( n2091 & n2139 ) ;
  assign n13597 = ( n390 & ~n1934 ) | ( n390 & n13596 ) | ( ~n1934 & n13596 ) ;
  assign n13598 = ~n12055 & n13597 ;
  assign n13599 = ~n302 & n13598 ;
  assign n13600 = n9544 ^ n1808 ^ n1113 ;
  assign n13601 = ( n5925 & ~n11869 ) | ( n5925 & n13600 ) | ( ~n11869 & n13600 ) ;
  assign n13606 = n2374 & ~n4315 ;
  assign n13607 = ( ~n3985 & n9660 ) | ( ~n3985 & n13606 ) | ( n9660 & n13606 ) ;
  assign n13602 = n1021 | n5870 ;
  assign n13603 = n2747 | n13602 ;
  assign n13604 = n13603 ^ n9080 ^ 1'b0 ;
  assign n13605 = ( ~n7070 & n8846 ) | ( ~n7070 & n13604 ) | ( n8846 & n13604 ) ;
  assign n13608 = n13607 ^ n13605 ^ n5479 ;
  assign n13616 = ( n1377 & n2260 ) | ( n1377 & n11631 ) | ( n2260 & n11631 ) ;
  assign n13617 = ( n8690 & n8947 ) | ( n8690 & n13616 ) | ( n8947 & n13616 ) ;
  assign n13618 = n11015 ^ n6102 ^ n5040 ;
  assign n13619 = ( n8447 & n13617 ) | ( n8447 & ~n13618 ) | ( n13617 & ~n13618 ) ;
  assign n13620 = n8900 ^ n3278 ^ n2974 ;
  assign n13621 = n13620 ^ n10491 ^ n3666 ;
  assign n13622 = n13621 ^ n5513 ^ 1'b0 ;
  assign n13623 = n13622 ^ n294 ^ 1'b0 ;
  assign n13624 = ~n13619 & n13623 ;
  assign n13611 = n3017 | n4369 ;
  assign n13612 = n6924 & ~n13611 ;
  assign n13613 = ( n152 & n464 ) | ( n152 & n983 ) | ( n464 & n983 ) ;
  assign n13614 = n13612 | n13613 ;
  assign n13609 = n8540 ^ n7964 ^ n2430 ;
  assign n13610 = ( n3478 & n12414 ) | ( n3478 & ~n13609 ) | ( n12414 & ~n13609 ) ;
  assign n13615 = n13614 ^ n13610 ^ n9255 ;
  assign n13625 = n13624 ^ n13615 ^ n2367 ;
  assign n13627 = n1416 & ~n10059 ;
  assign n13628 = ~n4506 & n13627 ;
  assign n13626 = n2929 ^ n956 ^ n813 ;
  assign n13629 = n13628 ^ n13626 ^ n1688 ;
  assign n13630 = n13629 ^ n11209 ^ 1'b0 ;
  assign n13631 = n13625 | n13630 ;
  assign n13632 = ( n2165 & n11999 ) | ( n2165 & ~n12957 ) | ( n11999 & ~n12957 ) ;
  assign n13634 = n9470 ^ n2042 ^ n1513 ;
  assign n13635 = ~n8827 & n13634 ;
  assign n13636 = ( n4819 & n5732 ) | ( n4819 & n13635 ) | ( n5732 & n13635 ) ;
  assign n13637 = n13636 ^ n12172 ^ n7661 ;
  assign n13633 = n5296 ^ n4058 ^ n2095 ;
  assign n13638 = n13637 ^ n13633 ^ n9443 ;
  assign n13639 = ( n3073 & n12781 ) | ( n3073 & n13638 ) | ( n12781 & n13638 ) ;
  assign n13640 = n13305 ^ n2325 ^ 1'b0 ;
  assign n13641 = n1652 | n13640 ;
  assign n13642 = n9545 ^ n8556 ^ n470 ;
  assign n13643 = ( n1792 & n3142 ) | ( n1792 & n7076 ) | ( n3142 & n7076 ) ;
  assign n13644 = ( ~n8923 & n10815 ) | ( ~n8923 & n13643 ) | ( n10815 & n13643 ) ;
  assign n13645 = n8705 ^ n7788 ^ n6165 ;
  assign n13646 = ( n4185 & n11500 ) | ( n4185 & n13645 ) | ( n11500 & n13645 ) ;
  assign n13653 = ( ~n4786 & n6075 ) | ( ~n4786 & n10736 ) | ( n6075 & n10736 ) ;
  assign n13651 = n2609 ^ n1687 ^ n1239 ;
  assign n13649 = n4190 ^ n2790 ^ n1233 ;
  assign n13650 = ( n409 & n10136 ) | ( n409 & ~n13649 ) | ( n10136 & ~n13649 ) ;
  assign n13652 = n13651 ^ n13650 ^ x54 ;
  assign n13654 = n13653 ^ n13652 ^ n3080 ;
  assign n13647 = n899 | n4913 ;
  assign n13648 = n2701 | n13647 ;
  assign n13655 = n13654 ^ n13648 ^ 1'b0 ;
  assign n13656 = n13646 & ~n13655 ;
  assign n13657 = ( n1801 & n4930 ) | ( n1801 & n11871 ) | ( n4930 & n11871 ) ;
  assign n13658 = n13657 ^ n12914 ^ n11726 ;
  assign n13659 = ( n2956 & n10841 ) | ( n2956 & n13658 ) | ( n10841 & n13658 ) ;
  assign n13660 = n5270 ^ n3661 ^ n3056 ;
  assign n13661 = ( n1107 & n4898 ) | ( n1107 & ~n13660 ) | ( n4898 & ~n13660 ) ;
  assign n13663 = n5027 ^ n3893 ^ n1326 ;
  assign n13664 = n9860 ^ n4271 ^ n2271 ;
  assign n13665 = n13664 ^ n8105 ^ 1'b0 ;
  assign n13666 = ~n13663 & n13665 ;
  assign n13662 = n6763 ^ n2781 ^ n796 ;
  assign n13667 = n13666 ^ n13662 ^ n2715 ;
  assign n13668 = ( n2577 & n13661 ) | ( n2577 & ~n13667 ) | ( n13661 & ~n13667 ) ;
  assign n13669 = n8154 ^ n6587 ^ 1'b0 ;
  assign n13670 = n13669 ^ n7526 ^ n4452 ;
  assign n13674 = ( n2573 & n5600 ) | ( n2573 & ~n6454 ) | ( n5600 & ~n6454 ) ;
  assign n13673 = ( n3684 & n5667 ) | ( n3684 & n8414 ) | ( n5667 & n8414 ) ;
  assign n13671 = n5639 | n12018 ;
  assign n13672 = n2085 | n13671 ;
  assign n13675 = n13674 ^ n13673 ^ n13672 ;
  assign n13676 = ( n181 & n2610 ) | ( n181 & ~n5661 ) | ( n2610 & ~n5661 ) ;
  assign n13677 = ( n9200 & n10628 ) | ( n9200 & n13676 ) | ( n10628 & n13676 ) ;
  assign n13678 = n11306 ^ n10262 ^ n2704 ;
  assign n13679 = n4735 & n13678 ;
  assign n13680 = ( n1909 & n2606 ) | ( n1909 & ~n12016 ) | ( n2606 & ~n12016 ) ;
  assign n13681 = n13680 ^ n2994 ^ 1'b0 ;
  assign n13682 = ( n901 & n8652 ) | ( n901 & n10517 ) | ( n8652 & n10517 ) ;
  assign n13683 = n12741 ^ n3879 ^ 1'b0 ;
  assign n13684 = n5671 ^ n5239 ^ n4471 ;
  assign n13685 = ( n900 & ~n11217 ) | ( n900 & n13684 ) | ( ~n11217 & n13684 ) ;
  assign n13686 = ( n13682 & ~n13683 ) | ( n13682 & n13685 ) | ( ~n13683 & n13685 ) ;
  assign n13687 = n6904 | n13140 ;
  assign n13688 = n6770 ^ n6641 ^ n2754 ;
  assign n13689 = ~n8322 & n11473 ;
  assign n13690 = n5658 ^ n1001 ^ x97 ;
  assign n13691 = n13690 ^ n11369 ^ 1'b0 ;
  assign n13692 = ~n9732 & n13691 ;
  assign n13693 = n6751 & n13692 ;
  assign n13695 = ( n2694 & n7253 ) | ( n2694 & ~n8701 ) | ( n7253 & ~n8701 ) ;
  assign n13694 = n944 | n3623 ;
  assign n13696 = n13695 ^ n13694 ^ 1'b0 ;
  assign n13697 = n13696 ^ n12390 ^ n2236 ;
  assign n13698 = n4735 & ~n7049 ;
  assign n13699 = ~n1802 & n13698 ;
  assign n13703 = n13622 ^ n5074 ^ 1'b0 ;
  assign n13704 = ~n5963 & n13703 ;
  assign n13700 = n7479 ^ n2891 ^ n1246 ;
  assign n13701 = n13700 ^ n9098 ^ 1'b0 ;
  assign n13702 = n10489 & n13701 ;
  assign n13705 = n13704 ^ n13702 ^ 1'b0 ;
  assign n13706 = ( n7824 & n13699 ) | ( n7824 & n13705 ) | ( n13699 & n13705 ) ;
  assign n13707 = ( n6099 & n13697 ) | ( n6099 & n13706 ) | ( n13697 & n13706 ) ;
  assign n13711 = n793 | n9336 ;
  assign n13712 = n13711 ^ n7479 ^ 1'b0 ;
  assign n13713 = n13712 ^ n5337 ^ 1'b0 ;
  assign n13708 = n6218 ^ n4993 ^ n603 ;
  assign n13709 = ( n474 & n8629 ) | ( n474 & ~n8966 ) | ( n8629 & ~n8966 ) ;
  assign n13710 = ( n4334 & n13708 ) | ( n4334 & n13709 ) | ( n13708 & n13709 ) ;
  assign n13714 = n13713 ^ n13710 ^ n1390 ;
  assign n13715 = ( n2420 & ~n9121 ) | ( n2420 & n9897 ) | ( ~n9121 & n9897 ) ;
  assign n13716 = n13715 ^ n12184 ^ n2071 ;
  assign n13717 = n2774 ^ n1415 ^ 1'b0 ;
  assign n13718 = n11571 | n13717 ;
  assign n13719 = n819 & ~n3418 ;
  assign n13720 = n13719 ^ n2096 ^ 1'b0 ;
  assign n13721 = n5432 ^ n226 ^ 1'b0 ;
  assign n13722 = n13721 ^ n7513 ^ n5597 ;
  assign n13723 = ( n3228 & n10852 ) | ( n3228 & ~n13722 ) | ( n10852 & ~n13722 ) ;
  assign n13724 = ( ~n7327 & n10644 ) | ( ~n7327 & n13723 ) | ( n10644 & n13723 ) ;
  assign n13725 = ( n975 & n2504 ) | ( n975 & n13724 ) | ( n2504 & n13724 ) ;
  assign n13726 = ( n2787 & n13720 ) | ( n2787 & n13725 ) | ( n13720 & n13725 ) ;
  assign n13727 = ( n3216 & n5157 ) | ( n3216 & ~n5931 ) | ( n5157 & ~n5931 ) ;
  assign n13728 = n3411 & ~n12648 ;
  assign n13729 = ~n13727 & n13728 ;
  assign n13730 = n9090 & n10853 ;
  assign n13731 = n1386 & n13730 ;
  assign n13732 = ( n247 & ~n13729 ) | ( n247 & n13731 ) | ( ~n13729 & n13731 ) ;
  assign n13733 = ( n3218 & n9722 ) | ( n3218 & n9756 ) | ( n9722 & n9756 ) ;
  assign n13734 = n12885 ^ n7586 ^ n4030 ;
  assign n13735 = n6370 ^ n5841 ^ 1'b0 ;
  assign n13736 = n11995 & ~n13735 ;
  assign n13737 = n12812 & n13736 ;
  assign n13738 = n13734 & n13737 ;
  assign n13739 = n11368 ^ n664 ^ x71 ;
  assign n13740 = ( n859 & n9911 ) | ( n859 & n13739 ) | ( n9911 & n13739 ) ;
  assign n13741 = ( n2323 & ~n7933 ) | ( n2323 & n13740 ) | ( ~n7933 & n13740 ) ;
  assign n13743 = ( n1876 & n2685 ) | ( n1876 & n7461 ) | ( n2685 & n7461 ) ;
  assign n13742 = n6077 | n12722 ;
  assign n13744 = n13743 ^ n13742 ^ 1'b0 ;
  assign n13745 = n13741 & ~n13744 ;
  assign n13746 = n4379 & n13745 ;
  assign n13747 = n5831 ^ n4476 ^ n1995 ;
  assign n13748 = n10420 ^ n8418 ^ n4588 ;
  assign n13749 = n2619 & n7543 ;
  assign n13750 = n13749 ^ n2378 ^ 1'b0 ;
  assign n13751 = n13750 ^ n13106 ^ n3226 ;
  assign n13752 = n9967 ^ n9300 ^ 1'b0 ;
  assign n13753 = n13751 & n13752 ;
  assign n13754 = ~n13748 & n13753 ;
  assign n13755 = n13754 ^ n12141 ^ n4505 ;
  assign n13756 = n10187 ^ n7305 ^ n3724 ;
  assign n13757 = n6258 | n11618 ;
  assign n13758 = n8254 & ~n13757 ;
  assign n13759 = ( ~n3172 & n13756 ) | ( ~n3172 & n13758 ) | ( n13756 & n13758 ) ;
  assign n13760 = n9479 ^ n5190 ^ 1'b0 ;
  assign n13761 = n5157 ^ n4059 ^ n472 ;
  assign n13762 = n12688 ^ n1154 ^ n696 ;
  assign n13763 = ( n1129 & n6693 ) | ( n1129 & ~n13103 ) | ( n6693 & ~n13103 ) ;
  assign n13764 = n13763 ^ n9769 ^ n7396 ;
  assign n13765 = ( n13761 & n13762 ) | ( n13761 & ~n13764 ) | ( n13762 & ~n13764 ) ;
  assign n13766 = ( n1960 & ~n6956 ) | ( n1960 & n10831 ) | ( ~n6956 & n10831 ) ;
  assign n13772 = n7942 ^ n4079 ^ n3296 ;
  assign n13767 = n7657 ^ n1718 ^ 1'b0 ;
  assign n13768 = n11790 | n13767 ;
  assign n13769 = n7951 | n13768 ;
  assign n13770 = n4390 & ~n13769 ;
  assign n13771 = n11259 & ~n13770 ;
  assign n13773 = n13772 ^ n13771 ^ 1'b0 ;
  assign n13779 = n1242 | n4843 ;
  assign n13780 = n13779 ^ n5959 ^ 1'b0 ;
  assign n13781 = ( n9930 & n10490 ) | ( n9930 & n13780 ) | ( n10490 & n13780 ) ;
  assign n13778 = ( n413 & n8137 ) | ( n413 & n11000 ) | ( n8137 & n11000 ) ;
  assign n13782 = n13781 ^ n13778 ^ n6027 ;
  assign n13774 = ( n1934 & n3580 ) | ( n1934 & n4202 ) | ( n3580 & n4202 ) ;
  assign n13775 = n13774 ^ n3756 ^ n2976 ;
  assign n13776 = ( ~n1587 & n7643 ) | ( ~n1587 & n13775 ) | ( n7643 & n13775 ) ;
  assign n13777 = ( n1948 & n11101 ) | ( n1948 & ~n13776 ) | ( n11101 & ~n13776 ) ;
  assign n13783 = n13782 ^ n13777 ^ n6659 ;
  assign n13784 = n13317 | n13783 ;
  assign n13785 = n456 & n11066 ;
  assign n13786 = n1705 | n5022 ;
  assign n13787 = ( ~n740 & n1559 ) | ( ~n740 & n8801 ) | ( n1559 & n8801 ) ;
  assign n13788 = ( ~n10733 & n13786 ) | ( ~n10733 & n13787 ) | ( n13786 & n13787 ) ;
  assign n13791 = ( n826 & ~n3531 ) | ( n826 & n9410 ) | ( ~n3531 & n9410 ) ;
  assign n13792 = n13791 ^ n1432 ^ 1'b0 ;
  assign n13789 = ( n209 & ~n1268 ) | ( n209 & n4619 ) | ( ~n1268 & n4619 ) ;
  assign n13790 = ( n6886 & ~n12656 ) | ( n6886 & n13789 ) | ( ~n12656 & n13789 ) ;
  assign n13793 = n13792 ^ n13790 ^ n10618 ;
  assign n13794 = n8525 ^ n3478 ^ n2139 ;
  assign n13795 = ( n411 & n1413 ) | ( n411 & ~n1803 ) | ( n1413 & ~n1803 ) ;
  assign n13796 = n13795 ^ n3480 ^ n643 ;
  assign n13797 = n5753 | n12856 ;
  assign n13798 = n13796 | n13797 ;
  assign n13799 = ( ~n4481 & n4803 ) | ( ~n4481 & n13798 ) | ( n4803 & n13798 ) ;
  assign n13800 = n8496 ^ n7032 ^ 1'b0 ;
  assign n13801 = ( x47 & ~n5250 ) | ( x47 & n13800 ) | ( ~n5250 & n13800 ) ;
  assign n13802 = ~n13799 & n13801 ;
  assign n13803 = ( n476 & n3840 ) | ( n476 & n13802 ) | ( n3840 & n13802 ) ;
  assign n13804 = n9148 ^ n4544 ^ n1346 ;
  assign n13805 = n13804 ^ n11020 ^ n7838 ;
  assign n13806 = ( n11462 & ~n13125 ) | ( n11462 & n13805 ) | ( ~n13125 & n13805 ) ;
  assign n13807 = n560 & ~n13371 ;
  assign n13808 = n3859 & n13807 ;
  assign n13809 = ( n887 & ~n3424 ) | ( n887 & n10041 ) | ( ~n3424 & n10041 ) ;
  assign n13810 = n4425 ^ n1004 ^ n765 ;
  assign n13811 = ( ~n13808 & n13809 ) | ( ~n13808 & n13810 ) | ( n13809 & n13810 ) ;
  assign n13812 = n13811 ^ n3355 ^ n829 ;
  assign n13813 = n6163 ^ n5215 ^ n4760 ;
  assign n13814 = n12205 ^ n1479 ^ 1'b0 ;
  assign n13815 = n13814 ^ n11498 ^ n6401 ;
  assign n13816 = ( n421 & n13813 ) | ( n421 & n13815 ) | ( n13813 & n13815 ) ;
  assign n13817 = n2151 | n2275 ;
  assign n13818 = n13817 ^ n6475 ^ 1'b0 ;
  assign n13819 = ( n8101 & n13816 ) | ( n8101 & ~n13818 ) | ( n13816 & ~n13818 ) ;
  assign n13820 = n7518 ^ n6723 ^ n3057 ;
  assign n13821 = ~n2874 & n13820 ;
  assign n13823 = ~n3709 & n3973 ;
  assign n13824 = n8511 & n13823 ;
  assign n13825 = n13824 ^ n7670 ^ n6173 ;
  assign n13822 = ( x11 & n3782 ) | ( x11 & n12794 ) | ( n3782 & n12794 ) ;
  assign n13826 = n13825 ^ n13822 ^ 1'b0 ;
  assign n13827 = n10295 & n13826 ;
  assign n13828 = ( n6493 & n9378 ) | ( n6493 & n13827 ) | ( n9378 & n13827 ) ;
  assign n13829 = n8439 ^ n563 ^ 1'b0 ;
  assign n13830 = n4585 ^ n3185 ^ n2989 ;
  assign n13831 = ( n6588 & n7054 ) | ( n6588 & n13830 ) | ( n7054 & n13830 ) ;
  assign n13832 = ~n5709 & n12168 ;
  assign n13833 = ( n1561 & ~n4203 ) | ( n1561 & n13832 ) | ( ~n4203 & n13832 ) ;
  assign n13834 = n13833 ^ n12956 ^ n4732 ;
  assign n13835 = ~n8687 & n8755 ;
  assign n13836 = ~n13834 & n13835 ;
  assign n13837 = n13836 ^ n13295 ^ 1'b0 ;
  assign n13838 = n4481 ^ n2268 ^ 1'b0 ;
  assign n13839 = ( ~n2637 & n8895 ) | ( ~n2637 & n13838 ) | ( n8895 & n13838 ) ;
  assign n13840 = ( n2882 & ~n13521 ) | ( n2882 & n13839 ) | ( ~n13521 & n13839 ) ;
  assign n13841 = n1073 ^ n439 ^ 1'b0 ;
  assign n13842 = ~n5358 & n13841 ;
  assign n13844 = n4175 & n6550 ;
  assign n13843 = n2512 | n11812 ;
  assign n13845 = n13844 ^ n13843 ^ 1'b0 ;
  assign n13846 = n2419 & ~n12223 ;
  assign n13847 = n13846 ^ n4011 ^ n1617 ;
  assign n13848 = n13847 ^ n8349 ^ n1048 ;
  assign n13849 = ( n2449 & n3232 ) | ( n2449 & n4673 ) | ( n3232 & n4673 ) ;
  assign n13850 = ( n5712 & ~n6674 ) | ( n5712 & n13849 ) | ( ~n6674 & n13849 ) ;
  assign n13851 = ~n4691 & n13850 ;
  assign n13858 = n6501 ^ n3241 ^ n2112 ;
  assign n13859 = ( n5100 & n13026 ) | ( n5100 & ~n13858 ) | ( n13026 & ~n13858 ) ;
  assign n13857 = n11797 ^ n2120 ^ n335 ;
  assign n13852 = ( n129 & n672 ) | ( n129 & n2510 ) | ( n672 & n2510 ) ;
  assign n13853 = n13852 ^ n7503 ^ n3091 ;
  assign n13854 = n13853 ^ n4127 ^ 1'b0 ;
  assign n13855 = ( n3367 & ~n8085 ) | ( n3367 & n13854 ) | ( ~n8085 & n13854 ) ;
  assign n13856 = n10496 | n13855 ;
  assign n13860 = n13859 ^ n13857 ^ n13856 ;
  assign n13861 = n8577 & n10735 ;
  assign n13862 = n3398 | n13818 ;
  assign n13863 = n13862 ^ n10488 ^ 1'b0 ;
  assign n13864 = n9668 ^ n6500 ^ 1'b0 ;
  assign n13865 = ( n3779 & ~n10358 ) | ( n3779 & n12606 ) | ( ~n10358 & n12606 ) ;
  assign n13866 = n13865 ^ n801 ^ 1'b0 ;
  assign n13867 = n13864 & ~n13866 ;
  assign n13868 = n13867 ^ n4039 ^ 1'b0 ;
  assign n13869 = n10441 & n13868 ;
  assign n13870 = n10615 ^ n5566 ^ n2350 ;
  assign n13871 = n13870 ^ n10933 ^ n8930 ;
  assign n13876 = ( n294 & n6157 ) | ( n294 & ~n12022 ) | ( n6157 & ~n12022 ) ;
  assign n13875 = n5306 ^ n1093 ^ x14 ;
  assign n13872 = ( ~n1268 & n2970 ) | ( ~n1268 & n3509 ) | ( n2970 & n3509 ) ;
  assign n13873 = n13872 ^ n10864 ^ 1'b0 ;
  assign n13874 = n13873 ^ n9622 ^ n5693 ;
  assign n13877 = n13876 ^ n13875 ^ n13874 ;
  assign n13878 = n12263 ^ n11054 ^ n4009 ;
  assign n13879 = ( n7917 & ~n9002 ) | ( n7917 & n13316 ) | ( ~n9002 & n13316 ) ;
  assign n13880 = ~n9006 & n13879 ;
  assign n13881 = ~n11209 & n13880 ;
  assign n13882 = n2310 ^ n2228 ^ 1'b0 ;
  assign n13883 = ~n2412 & n13882 ;
  assign n13884 = ~n9945 & n13883 ;
  assign n13885 = n13884 ^ n10522 ^ 1'b0 ;
  assign n13886 = ( n294 & ~n484 ) | ( n294 & n13885 ) | ( ~n484 & n13885 ) ;
  assign n13887 = n13886 ^ n1866 ^ n148 ;
  assign n13888 = ( n8895 & n13881 ) | ( n8895 & ~n13887 ) | ( n13881 & ~n13887 ) ;
  assign n13889 = n8531 ^ n7096 ^ n2417 ;
  assign n13890 = n7260 ^ n1174 ^ 1'b0 ;
  assign n13891 = ~n10308 & n13890 ;
  assign n13892 = n7274 ^ n4561 ^ n3865 ;
  assign n13893 = n13892 ^ n9437 ^ 1'b0 ;
  assign n13894 = n6635 | n13893 ;
  assign n13895 = ( n4608 & n5120 ) | ( n4608 & ~n12455 ) | ( n5120 & ~n12455 ) ;
  assign n13896 = ~n6901 & n13895 ;
  assign n13897 = n10648 & n13896 ;
  assign n13898 = n6188 ^ n5874 ^ n2652 ;
  assign n13899 = ( ~n11075 & n12930 ) | ( ~n11075 & n13898 ) | ( n12930 & n13898 ) ;
  assign n13901 = ( x5 & ~n4195 ) | ( x5 & n12635 ) | ( ~n4195 & n12635 ) ;
  assign n13900 = n11207 | n11817 ;
  assign n13902 = n13901 ^ n13900 ^ n4473 ;
  assign n13903 = n5954 ^ n5499 ^ 1'b0 ;
  assign n13904 = n4793 | n13903 ;
  assign n13905 = ( n8694 & n12318 ) | ( n8694 & n13351 ) | ( n12318 & n13351 ) ;
  assign n13906 = ( n5618 & ~n7812 ) | ( n5618 & n12125 ) | ( ~n7812 & n12125 ) ;
  assign n13907 = n8149 ^ n565 ^ 1'b0 ;
  assign n13908 = n13907 ^ n8753 ^ 1'b0 ;
  assign n13909 = x117 & n10589 ;
  assign n13910 = n2640 & n3866 ;
  assign n13911 = ~n13909 & n13910 ;
  assign n13912 = ( n1073 & ~n2446 ) | ( n1073 & n5393 ) | ( ~n2446 & n5393 ) ;
  assign n13913 = n9298 ^ n4310 ^ n946 ;
  assign n13914 = ( ~n2875 & n13912 ) | ( ~n2875 & n13913 ) | ( n13912 & n13913 ) ;
  assign n13916 = n4123 ^ n2504 ^ 1'b0 ;
  assign n13917 = n7013 & n13916 ;
  assign n13915 = n7370 ^ n4424 ^ n3579 ;
  assign n13918 = n13917 ^ n13915 ^ n1676 ;
  assign n13919 = n9743 ^ n7230 ^ n3056 ;
  assign n13920 = n13919 ^ n4119 ^ n1959 ;
  assign n13921 = n13920 ^ n12216 ^ n3235 ;
  assign n13922 = n13921 ^ n4609 ^ 1'b0 ;
  assign n13923 = n13918 & n13922 ;
  assign n13924 = n8182 ^ n5069 ^ n3041 ;
  assign n13925 = n13924 ^ n2749 ^ n1596 ;
  assign n13926 = n13925 ^ n5606 ^ n797 ;
  assign n13927 = n4529 ^ n4163 ^ n1146 ;
  assign n13928 = ( ~n5018 & n11490 ) | ( ~n5018 & n13927 ) | ( n11490 & n13927 ) ;
  assign n13929 = n3372 ^ n3278 ^ n1016 ;
  assign n13931 = n3915 & n7074 ;
  assign n13930 = ( n1207 & n2224 ) | ( n1207 & ~n12878 ) | ( n2224 & ~n12878 ) ;
  assign n13932 = n13931 ^ n13930 ^ 1'b0 ;
  assign n13933 = n4799 & n13932 ;
  assign n13934 = n9121 ^ n4690 ^ 1'b0 ;
  assign n13935 = n9414 & n13934 ;
  assign n13936 = ( ~n13929 & n13933 ) | ( ~n13929 & n13935 ) | ( n13933 & n13935 ) ;
  assign n13939 = n359 & n7704 ;
  assign n13940 = n563 & n13939 ;
  assign n13937 = n2098 | n4659 ;
  assign n13938 = n13937 ^ n9356 ^ 1'b0 ;
  assign n13941 = n13940 ^ n13938 ^ n6433 ;
  assign n13942 = n13373 ^ n12042 ^ n5062 ;
  assign n13943 = ( n2259 & ~n5381 ) | ( n2259 & n7196 ) | ( ~n5381 & n7196 ) ;
  assign n13944 = ~n5115 & n13943 ;
  assign n13945 = n13944 ^ n9443 ^ x83 ;
  assign n13946 = ( n10650 & n11994 ) | ( n10650 & n13945 ) | ( n11994 & n13945 ) ;
  assign n13948 = ( ~n2169 & n2513 ) | ( ~n2169 & n4112 ) | ( n2513 & n4112 ) ;
  assign n13947 = n11411 ^ n1550 ^ 1'b0 ;
  assign n13949 = n13948 ^ n13947 ^ n9383 ;
  assign n13950 = ( n6478 & n13946 ) | ( n6478 & n13949 ) | ( n13946 & n13949 ) ;
  assign n13951 = n13950 ^ n11413 ^ n4513 ;
  assign n13952 = ( n2507 & ~n2535 ) | ( n2507 & n3737 ) | ( ~n2535 & n3737 ) ;
  assign n13953 = ( n7187 & n13626 ) | ( n7187 & n13952 ) | ( n13626 & n13952 ) ;
  assign n13954 = n6535 ^ n4830 ^ n1960 ;
  assign n13955 = n13954 ^ n7622 ^ 1'b0 ;
  assign n13956 = n8769 ^ n4538 ^ 1'b0 ;
  assign n13957 = n4661 ^ n517 ^ 1'b0 ;
  assign n13958 = n7848 | n13957 ;
  assign n13959 = n13138 ^ n5609 ^ 1'b0 ;
  assign n13960 = ( n3538 & ~n10093 ) | ( n3538 & n13959 ) | ( ~n10093 & n13959 ) ;
  assign n13961 = n13960 ^ n12110 ^ n10564 ;
  assign n13962 = n10790 ^ n9079 ^ n669 ;
  assign n13963 = ( ~n688 & n10512 ) | ( ~n688 & n13962 ) | ( n10512 & n13962 ) ;
  assign n13964 = n11535 ^ n10056 ^ n8273 ;
  assign n13965 = n11419 ^ n4637 ^ n2494 ;
  assign n13966 = ( ~n857 & n922 ) | ( ~n857 & n4852 ) | ( n922 & n4852 ) ;
  assign n13967 = n7342 & ~n13966 ;
  assign n13968 = ~n13965 & n13967 ;
  assign n13969 = ( ~n4628 & n9855 ) | ( ~n4628 & n11451 ) | ( n9855 & n11451 ) ;
  assign n13970 = n7841 ^ n4578 ^ n1842 ;
  assign n13971 = n9675 ^ n1670 ^ 1'b0 ;
  assign n13972 = ( n9773 & n11206 ) | ( n9773 & n13971 ) | ( n11206 & n13971 ) ;
  assign n13973 = n13972 ^ n8084 ^ n3219 ;
  assign n13974 = ( n800 & ~n2267 ) | ( n800 & n2886 ) | ( ~n2267 & n2886 ) ;
  assign n13975 = n13306 ^ n11565 ^ n3293 ;
  assign n13976 = ( ~n13872 & n13974 ) | ( ~n13872 & n13975 ) | ( n13974 & n13975 ) ;
  assign n13977 = ( n765 & ~n3693 ) | ( n765 & n13976 ) | ( ~n3693 & n13976 ) ;
  assign n13978 = ( n1285 & ~n3247 ) | ( n1285 & n8114 ) | ( ~n3247 & n8114 ) ;
  assign n13981 = ( ~n1719 & n9469 ) | ( ~n1719 & n13974 ) | ( n9469 & n13974 ) ;
  assign n13982 = n13981 ^ n6943 ^ n1049 ;
  assign n13983 = n10081 ^ n1617 ^ n375 ;
  assign n13984 = n13982 | n13983 ;
  assign n13979 = n4372 & ~n6162 ;
  assign n13980 = n13979 ^ n7309 ^ 1'b0 ;
  assign n13985 = n13984 ^ n13980 ^ n5583 ;
  assign n13986 = ( ~n8058 & n13978 ) | ( ~n8058 & n13985 ) | ( n13978 & n13985 ) ;
  assign n13987 = n12418 ^ n10464 ^ 1'b0 ;
  assign n13988 = ( n3859 & n6062 ) | ( n3859 & n6643 ) | ( n6062 & n6643 ) ;
  assign n13989 = ( n3595 & ~n8637 ) | ( n3595 & n13988 ) | ( ~n8637 & n13988 ) ;
  assign n13991 = ( n5973 & ~n7460 ) | ( n5973 & n8514 ) | ( ~n7460 & n8514 ) ;
  assign n13990 = ~n2721 & n10615 ;
  assign n13992 = n13991 ^ n13990 ^ 1'b0 ;
  assign n13993 = ( n7253 & n13104 ) | ( n7253 & n13992 ) | ( n13104 & n13992 ) ;
  assign n13994 = n2538 ^ n1469 ^ 1'b0 ;
  assign n13995 = x71 & ~n13994 ;
  assign n13996 = ( n4939 & n7257 ) | ( n4939 & n13995 ) | ( n7257 & n13995 ) ;
  assign n13997 = ( ~n4259 & n10142 ) | ( ~n4259 & n10143 ) | ( n10142 & n10143 ) ;
  assign n13998 = ( ~n235 & n8718 ) | ( ~n235 & n13997 ) | ( n8718 & n13997 ) ;
  assign n13999 = ( n765 & ~n1721 ) | ( n765 & n12368 ) | ( ~n1721 & n12368 ) ;
  assign n14009 = n2429 ^ n1367 ^ 1'b0 ;
  assign n14004 = n2286 | n4273 ;
  assign n14005 = n9567 ^ n1966 ^ n764 ;
  assign n14006 = ( n2888 & n13983 ) | ( n2888 & n14005 ) | ( n13983 & n14005 ) ;
  assign n14007 = n14006 ^ n9879 ^ n2998 ;
  assign n14008 = ( n1979 & ~n14004 ) | ( n1979 & n14007 ) | ( ~n14004 & n14007 ) ;
  assign n14010 = n14009 ^ n14008 ^ n1602 ;
  assign n14011 = ( n9679 & n11285 ) | ( n9679 & ~n14010 ) | ( n11285 & ~n14010 ) ;
  assign n14000 = n11251 | n12106 ;
  assign n14001 = n14000 ^ n12404 ^ n6985 ;
  assign n14002 = ( n6677 & n12440 ) | ( n6677 & n13647 ) | ( n12440 & n13647 ) ;
  assign n14003 = n14001 & n14002 ;
  assign n14012 = n14011 ^ n14003 ^ 1'b0 ;
  assign n14013 = n4575 | n14012 ;
  assign n14014 = n13999 | n14013 ;
  assign n14023 = n5261 ^ n3693 ^ n1334 ;
  assign n14024 = n1477 | n14023 ;
  assign n14021 = n1689 ^ n1504 ^ n1245 ;
  assign n14022 = n14021 ^ n9252 ^ n5493 ;
  assign n14019 = n11863 ^ n4020 ^ n2633 ;
  assign n14015 = n13326 ^ n4136 ^ n3808 ;
  assign n14016 = n13519 & n14015 ;
  assign n14017 = ~n6645 & n14016 ;
  assign n14018 = ( n3607 & ~n13094 ) | ( n3607 & n14017 ) | ( ~n13094 & n14017 ) ;
  assign n14020 = n14019 ^ n14018 ^ n1171 ;
  assign n14025 = n14024 ^ n14022 ^ n14020 ;
  assign n14027 = n6008 ^ x27 ^ 1'b0 ;
  assign n14026 = ( n1677 & n2240 ) | ( n1677 & n11552 ) | ( n2240 & n11552 ) ;
  assign n14028 = n14027 ^ n14026 ^ n12865 ;
  assign n14029 = ( n1876 & ~n2286 ) | ( n1876 & n2845 ) | ( ~n2286 & n2845 ) ;
  assign n14030 = n4579 ^ n2142 ^ n366 ;
  assign n14031 = n14030 ^ n10091 ^ n4604 ;
  assign n14034 = ( n382 & ~n2360 ) | ( n382 & n3121 ) | ( ~n2360 & n3121 ) ;
  assign n14032 = n9298 ^ n8199 ^ n7494 ;
  assign n14033 = n213 & ~n14032 ;
  assign n14035 = n14034 ^ n14033 ^ 1'b0 ;
  assign n14036 = n4801 & ~n14035 ;
  assign n14037 = n11456 ^ n10552 ^ 1'b0 ;
  assign n14042 = ( n2472 & n3466 ) | ( n2472 & ~n7886 ) | ( n3466 & ~n7886 ) ;
  assign n14038 = n3711 | n3716 ;
  assign n14039 = n14038 ^ n4280 ^ 1'b0 ;
  assign n14040 = ( n302 & n6054 ) | ( n302 & n14039 ) | ( n6054 & n14039 ) ;
  assign n14041 = n1850 | n14040 ;
  assign n14043 = n14042 ^ n14041 ^ n10841 ;
  assign n14044 = n12224 ^ n4685 ^ n2515 ;
  assign n14045 = ( n2666 & ~n12519 ) | ( n2666 & n14044 ) | ( ~n12519 & n14044 ) ;
  assign n14046 = n6733 & n6734 ;
  assign n14047 = n14046 ^ n7081 ^ n2259 ;
  assign n14048 = ( n14005 & n14045 ) | ( n14005 & ~n14047 ) | ( n14045 & ~n14047 ) ;
  assign n14049 = ( x80 & n4857 ) | ( x80 & ~n10339 ) | ( n4857 & ~n10339 ) ;
  assign n14050 = ( ~n355 & n12442 ) | ( ~n355 & n13723 ) | ( n12442 & n13723 ) ;
  assign n14051 = n9383 ^ n595 ^ 1'b0 ;
  assign n14052 = ( n5934 & n8351 ) | ( n5934 & n14051 ) | ( n8351 & n14051 ) ;
  assign n14053 = n10082 ^ n7840 ^ n7382 ;
  assign n14054 = n6730 ^ n1576 ^ 1'b0 ;
  assign n14055 = n13846 | n14054 ;
  assign n14056 = ( n6671 & n14053 ) | ( n6671 & n14055 ) | ( n14053 & n14055 ) ;
  assign n14057 = n14056 ^ n5244 ^ n2788 ;
  assign n14058 = n6910 & n14057 ;
  assign n14059 = ( ~n4452 & n7212 ) | ( ~n4452 & n10601 ) | ( n7212 & n10601 ) ;
  assign n14060 = n14059 ^ n12168 ^ n4342 ;
  assign n14061 = n3978 ^ n638 ^ 1'b0 ;
  assign n14062 = ~n2511 & n13680 ;
  assign n14063 = n14062 ^ n5822 ^ 1'b0 ;
  assign n14064 = ( ~x127 & n4372 ) | ( ~x127 & n10422 ) | ( n4372 & n10422 ) ;
  assign n14065 = n3082 & n4532 ;
  assign n14066 = n14065 ^ n14007 ^ 1'b0 ;
  assign n14067 = ( n9079 & n12593 ) | ( n9079 & ~n14066 ) | ( n12593 & ~n14066 ) ;
  assign n14070 = n7607 ^ n4544 ^ n1142 ;
  assign n14068 = n8168 & ~n9341 ;
  assign n14069 = n1728 & n14068 ;
  assign n14071 = n14070 ^ n14069 ^ 1'b0 ;
  assign n14072 = n5874 & ~n11116 ;
  assign n14073 = n8368 | n14072 ;
  assign n14074 = n14073 ^ n2196 ^ 1'b0 ;
  assign n14075 = n7406 ^ n5584 ^ 1'b0 ;
  assign n14076 = ( ~n2970 & n3926 ) | ( ~n2970 & n13870 ) | ( n3926 & n13870 ) ;
  assign n14077 = n14076 ^ n11281 ^ n6271 ;
  assign n14078 = n10107 ^ n4345 ^ 1'b0 ;
  assign n14079 = n10644 ^ n8439 ^ n3485 ;
  assign n14080 = n14079 ^ n944 ^ 1'b0 ;
  assign n14081 = n2341 & n14080 ;
  assign n14082 = ( x67 & ~n5665 ) | ( x67 & n11796 ) | ( ~n5665 & n11796 ) ;
  assign n14083 = n14082 ^ n13729 ^ n596 ;
  assign n14084 = ( n496 & ~n5951 ) | ( n496 & n13202 ) | ( ~n5951 & n13202 ) ;
  assign n14085 = n7329 ^ n2236 ^ n243 ;
  assign n14086 = n1325 | n4169 ;
  assign n14087 = n14086 ^ n5962 ^ 1'b0 ;
  assign n14088 = ( ~n3073 & n4160 ) | ( ~n3073 & n14087 ) | ( n4160 & n14087 ) ;
  assign n14089 = n14088 ^ n5983 ^ n2122 ;
  assign n14090 = n14089 ^ n11853 ^ n7555 ;
  assign n14091 = n1340 & n11388 ;
  assign n14092 = n14091 ^ x60 ^ 1'b0 ;
  assign n14093 = ( n953 & n6249 ) | ( n953 & n7615 ) | ( n6249 & n7615 ) ;
  assign n14094 = ( n4651 & n14092 ) | ( n4651 & n14093 ) | ( n14092 & n14093 ) ;
  assign n14095 = ( n4598 & n14090 ) | ( n4598 & n14094 ) | ( n14090 & n14094 ) ;
  assign n14096 = n14095 ^ n13764 ^ 1'b0 ;
  assign n14097 = ( ~n10069 & n14085 ) | ( ~n10069 & n14096 ) | ( n14085 & n14096 ) ;
  assign n14098 = n2724 ^ n2598 ^ 1'b0 ;
  assign n14099 = n13135 & ~n14098 ;
  assign n14109 = n2487 ^ n658 ^ x6 ;
  assign n14106 = n439 | n8319 ;
  assign n14107 = x79 | n14106 ;
  assign n14108 = n14107 ^ n9204 ^ n6257 ;
  assign n14102 = n6614 ^ x73 ^ x16 ;
  assign n14103 = ( n1041 & n8821 ) | ( n1041 & n14102 ) | ( n8821 & n14102 ) ;
  assign n14104 = n14103 ^ x88 ^ 1'b0 ;
  assign n14100 = ~n856 & n2131 ;
  assign n14101 = n6681 | n14100 ;
  assign n14105 = n14104 ^ n14101 ^ n2751 ;
  assign n14110 = n14109 ^ n14108 ^ n14105 ;
  assign n14111 = n1736 ^ n1551 ^ 1'b0 ;
  assign n14112 = n4123 & ~n14111 ;
  assign n14113 = n14112 ^ n12648 ^ 1'b0 ;
  assign n14114 = n6033 & ~n14113 ;
  assign n14117 = ( n1145 & n4641 ) | ( n1145 & ~n7513 ) | ( n4641 & ~n7513 ) ;
  assign n14115 = n12429 ^ n8399 ^ n6035 ;
  assign n14116 = n6077 | n14115 ;
  assign n14118 = n14117 ^ n14116 ^ 1'b0 ;
  assign n14119 = ( n10114 & n14114 ) | ( n10114 & ~n14118 ) | ( n14114 & ~n14118 ) ;
  assign n14120 = ( n4603 & ~n4853 ) | ( n4603 & n12880 ) | ( ~n4853 & n12880 ) ;
  assign n14121 = ( n2694 & n3129 ) | ( n2694 & n14120 ) | ( n3129 & n14120 ) ;
  assign n14122 = n7511 ^ n6380 ^ n2426 ;
  assign n14123 = n14122 ^ n5964 ^ n1167 ;
  assign n14124 = n3459 ^ n421 ^ 1'b0 ;
  assign n14125 = ( n2679 & n3294 ) | ( n2679 & n7236 ) | ( n3294 & n7236 ) ;
  assign n14126 = n1187 & n14125 ;
  assign n14127 = n13236 ^ n4048 ^ n2217 ;
  assign n14128 = ( n3042 & n14126 ) | ( n3042 & n14127 ) | ( n14126 & n14127 ) ;
  assign n14129 = n9951 ^ n4208 ^ 1'b0 ;
  assign n14130 = n12318 & ~n14129 ;
  assign n14131 = ( n1049 & n10125 ) | ( n1049 & ~n11446 ) | ( n10125 & ~n11446 ) ;
  assign n14132 = ( n9018 & n10522 ) | ( n9018 & n12591 ) | ( n10522 & n12591 ) ;
  assign n14133 = ( n2662 & ~n9932 ) | ( n2662 & n10765 ) | ( ~n9932 & n10765 ) ;
  assign n14134 = ( n5490 & n10761 ) | ( n5490 & n14133 ) | ( n10761 & n14133 ) ;
  assign n14135 = n14134 ^ n10086 ^ n7561 ;
  assign n14138 = ( ~n3051 & n5922 ) | ( ~n3051 & n9091 ) | ( n5922 & n9091 ) ;
  assign n14137 = n7227 & n11368 ;
  assign n14136 = n10267 ^ n9869 ^ n6889 ;
  assign n14139 = n14138 ^ n14137 ^ n14136 ;
  assign n14140 = ( n395 & n5285 ) | ( n395 & ~n5481 ) | ( n5285 & ~n5481 ) ;
  assign n14141 = ( ~n4732 & n5799 ) | ( ~n4732 & n14140 ) | ( n5799 & n14140 ) ;
  assign n14142 = ( n3059 & n10122 ) | ( n3059 & n14141 ) | ( n10122 & n14141 ) ;
  assign n14148 = n3753 | n8280 ;
  assign n14149 = n14148 ^ n9891 ^ 1'b0 ;
  assign n14143 = ( n1058 & n1834 ) | ( n1058 & n6773 ) | ( n1834 & n6773 ) ;
  assign n14144 = n14143 ^ n4476 ^ n2904 ;
  assign n14145 = n14144 ^ n12649 ^ n10869 ;
  assign n14146 = ( ~n7148 & n10542 ) | ( ~n7148 & n14145 ) | ( n10542 & n14145 ) ;
  assign n14147 = ~n5056 & n14146 ;
  assign n14150 = n14149 ^ n14147 ^ 1'b0 ;
  assign n14151 = n2340 & ~n9510 ;
  assign n14152 = ~x90 & n14151 ;
  assign n14153 = ( n4056 & n9813 ) | ( n4056 & ~n14152 ) | ( n9813 & ~n14152 ) ;
  assign n14154 = n14153 ^ n11883 ^ n8367 ;
  assign n14155 = n14154 ^ n9274 ^ 1'b0 ;
  assign n14156 = n11364 ^ n7528 ^ 1'b0 ;
  assign n14157 = ~n14155 & n14156 ;
  assign n14159 = n6086 ^ n3686 ^ 1'b0 ;
  assign n14160 = n6358 | n14159 ;
  assign n14158 = n11584 ^ n9642 ^ n994 ;
  assign n14161 = n14160 ^ n14158 ^ n7426 ;
  assign n14162 = n14161 ^ n8560 ^ 1'b0 ;
  assign n14163 = ( n862 & ~n6657 ) | ( n862 & n8346 ) | ( ~n6657 & n8346 ) ;
  assign n14164 = n14163 ^ n11041 ^ n7832 ;
  assign n14169 = ( n3041 & n5511 ) | ( n3041 & n11575 ) | ( n5511 & n11575 ) ;
  assign n14166 = ( n1034 & ~n1797 ) | ( n1034 & n3762 ) | ( ~n1797 & n3762 ) ;
  assign n14167 = n14166 ^ n5337 ^ n1175 ;
  assign n14165 = ( ~n4918 & n5915 ) | ( ~n4918 & n12312 ) | ( n5915 & n12312 ) ;
  assign n14168 = n14167 ^ n14165 ^ n12740 ;
  assign n14170 = n14169 ^ n14168 ^ n1626 ;
  assign n14171 = ~n157 & n1460 ;
  assign n14172 = n14171 ^ n12593 ^ n3585 ;
  assign n14173 = ( n329 & n10397 ) | ( n329 & n11206 ) | ( n10397 & n11206 ) ;
  assign n14174 = ( ~n2606 & n12168 ) | ( ~n2606 & n14173 ) | ( n12168 & n14173 ) ;
  assign n14175 = n3799 ^ n509 ^ 1'b0 ;
  assign n14176 = n149 ^ x30 ^ 1'b0 ;
  assign n14177 = n14176 ^ n11545 ^ n5601 ;
  assign n14178 = ( ~n1360 & n10720 ) | ( ~n1360 & n12496 ) | ( n10720 & n12496 ) ;
  assign n14179 = ( ~n9421 & n14177 ) | ( ~n9421 & n14178 ) | ( n14177 & n14178 ) ;
  assign n14180 = n10415 ^ n3886 ^ 1'b0 ;
  assign n14181 = n5354 ^ n3308 ^ 1'b0 ;
  assign n14182 = n4459 & n14181 ;
  assign n14183 = n2868 & n14182 ;
  assign n14184 = ( n4165 & n7125 ) | ( n4165 & n14183 ) | ( n7125 & n14183 ) ;
  assign n14185 = n14184 ^ n9616 ^ n9358 ;
  assign n14186 = ( ~n3660 & n8375 ) | ( ~n3660 & n12653 ) | ( n8375 & n12653 ) ;
  assign n14187 = n14186 ^ n5010 ^ n2179 ;
  assign n14188 = n14187 ^ n7267 ^ n1179 ;
  assign n14189 = n4298 & n14188 ;
  assign n14190 = n11387 & n14189 ;
  assign n14191 = n13548 ^ n11607 ^ n5062 ;
  assign n14192 = ~n3619 & n6467 ;
  assign n14193 = n14192 ^ n12994 ^ 1'b0 ;
  assign n14194 = ( ~n3782 & n10074 ) | ( ~n3782 & n14193 ) | ( n10074 & n14193 ) ;
  assign n14195 = n3082 & ~n9198 ;
  assign n14196 = n1748 & n14195 ;
  assign n14197 = n13489 ^ n2968 ^ 1'b0 ;
  assign n14198 = n14197 ^ n940 ^ 1'b0 ;
  assign n14199 = ~n14196 & n14198 ;
  assign n14201 = n8042 ^ n2673 ^ 1'b0 ;
  assign n14200 = n7071 | n10192 ;
  assign n14202 = n14201 ^ n14200 ^ 1'b0 ;
  assign n14203 = n14202 ^ n7519 ^ n3514 ;
  assign n14204 = n6141 & ~n7688 ;
  assign n14205 = ( n149 & ~n1670 ) | ( n149 & n5757 ) | ( ~n1670 & n5757 ) ;
  assign n14206 = ~n4169 & n12238 ;
  assign n14207 = n14205 & n14206 ;
  assign n14208 = ( n6366 & ~n12916 ) | ( n6366 & n14207 ) | ( ~n12916 & n14207 ) ;
  assign n14209 = n5858 ^ n1080 ^ n401 ;
  assign n14210 = ( n2391 & n10008 ) | ( n2391 & ~n14209 ) | ( n10008 & ~n14209 ) ;
  assign n14211 = n10479 ^ n486 ^ 1'b0 ;
  assign n14212 = n7349 ^ n3714 ^ n2761 ;
  assign n14213 = ( n8741 & ~n14211 ) | ( n8741 & n14212 ) | ( ~n14211 & n14212 ) ;
  assign n14214 = n11470 ^ n8170 ^ 1'b0 ;
  assign n14215 = n14213 & ~n14214 ;
  assign n14216 = n4613 & ~n12164 ;
  assign n14217 = n14216 ^ n7068 ^ 1'b0 ;
  assign n14218 = ( n8593 & ~n12812 ) | ( n8593 & n14217 ) | ( ~n12812 & n14217 ) ;
  assign n14219 = ( n11808 & ~n11852 ) | ( n11808 & n14218 ) | ( ~n11852 & n14218 ) ;
  assign n14220 = n3150 ^ n2183 ^ 1'b0 ;
  assign n14221 = n1836 | n14220 ;
  assign n14222 = n14221 ^ n9560 ^ n5391 ;
  assign n14223 = ( n1778 & n10337 ) | ( n1778 & n14222 ) | ( n10337 & n14222 ) ;
  assign n14224 = n14223 ^ n1178 ^ 1'b0 ;
  assign n14225 = n2808 | n5481 ;
  assign n14226 = n11122 & ~n14225 ;
  assign n14227 = n3998 ^ n1633 ^ 1'b0 ;
  assign n14228 = ~n781 & n14227 ;
  assign n14229 = n2724 & n14228 ;
  assign n14230 = ( n13106 & n13614 ) | ( n13106 & n14229 ) | ( n13614 & n14229 ) ;
  assign n14231 = n11092 ^ n5237 ^ 1'b0 ;
  assign n14235 = ( n760 & ~n4940 ) | ( n760 & n13347 ) | ( ~n4940 & n13347 ) ;
  assign n14233 = n546 & ~n553 ;
  assign n14234 = n14233 ^ n975 ^ 1'b0 ;
  assign n14232 = ( ~n4863 & n5733 ) | ( ~n4863 & n14006 ) | ( n5733 & n14006 ) ;
  assign n14236 = n14235 ^ n14234 ^ n14232 ;
  assign n14237 = ( ~n2306 & n14231 ) | ( ~n2306 & n14236 ) | ( n14231 & n14236 ) ;
  assign n14238 = n9228 & ~n9803 ;
  assign n14239 = n13153 ^ n11920 ^ n1420 ;
  assign n14240 = ( n4388 & ~n10739 ) | ( n4388 & n14239 ) | ( ~n10739 & n14239 ) ;
  assign n14241 = n7810 ^ n3423 ^ n2066 ;
  assign n14242 = ( n2934 & n6139 ) | ( n2934 & n14241 ) | ( n6139 & n14241 ) ;
  assign n14244 = ( n746 & ~n8856 ) | ( n746 & n13872 ) | ( ~n8856 & n13872 ) ;
  assign n14243 = n10187 ^ n2235 ^ n382 ;
  assign n14245 = n14244 ^ n14243 ^ n3299 ;
  assign n14246 = n5991 ^ n3117 ^ 1'b0 ;
  assign n14247 = n14104 & ~n14246 ;
  assign n14248 = n14247 ^ n10237 ^ n9931 ;
  assign n14249 = n342 | n3385 ;
  assign n14250 = n5650 & ~n14249 ;
  assign n14251 = n2411 ^ n569 ^ 1'b0 ;
  assign n14252 = n9563 | n14251 ;
  assign n14253 = n14252 ^ n8705 ^ 1'b0 ;
  assign n14254 = n11215 ^ n4141 ^ n2561 ;
  assign n14255 = n14254 ^ n11206 ^ n3441 ;
  assign n14256 = ( n10365 & n10651 ) | ( n10365 & ~n13983 ) | ( n10651 & ~n13983 ) ;
  assign n14257 = ~n10331 & n13806 ;
  assign n14258 = n14257 ^ n4872 ^ 1'b0 ;
  assign n14259 = n1994 & n4477 ;
  assign n14260 = n14259 ^ n10262 ^ 1'b0 ;
  assign n14262 = ( x1 & n523 ) | ( x1 & ~n7668 ) | ( n523 & ~n7668 ) ;
  assign n14261 = n4042 & ~n12947 ;
  assign n14263 = n14262 ^ n14261 ^ n6750 ;
  assign n14270 = ( n3878 & ~n6209 ) | ( n3878 & n13490 ) | ( ~n6209 & n13490 ) ;
  assign n14271 = n14270 ^ n194 ^ 1'b0 ;
  assign n14264 = ( ~n1623 & n3110 ) | ( ~n1623 & n10190 ) | ( n3110 & n10190 ) ;
  assign n14265 = n14264 ^ n7859 ^ n3767 ;
  assign n14266 = ( n3008 & n13715 ) | ( n3008 & ~n14265 ) | ( n13715 & ~n14265 ) ;
  assign n14267 = n1084 ^ n890 ^ x13 ;
  assign n14268 = ~n14266 & n14267 ;
  assign n14269 = n6459 & n14268 ;
  assign n14272 = n14271 ^ n14269 ^ n5391 ;
  assign n14273 = ( n9491 & n12091 ) | ( n9491 & ~n14272 ) | ( n12091 & ~n14272 ) ;
  assign n14275 = n14187 ^ n14082 ^ n8823 ;
  assign n14274 = n3705 | n10918 ;
  assign n14276 = n14275 ^ n14274 ^ 1'b0 ;
  assign n14277 = n4644 ^ n3217 ^ n251 ;
  assign n14278 = ( n4757 & ~n10962 ) | ( n4757 & n14277 ) | ( ~n10962 & n14277 ) ;
  assign n14279 = n14278 ^ n10636 ^ n8192 ;
  assign n14280 = ( n9009 & ~n11177 ) | ( n9009 & n14279 ) | ( ~n11177 & n14279 ) ;
  assign n14281 = n7499 ^ n6814 ^ 1'b0 ;
  assign n14282 = n6226 ^ n3177 ^ 1'b0 ;
  assign n14283 = n6292 ^ n2340 ^ 1'b0 ;
  assign n14284 = ( n4000 & n6157 ) | ( n4000 & n8619 ) | ( n6157 & n8619 ) ;
  assign n14285 = ( n2251 & ~n6306 ) | ( n2251 & n7730 ) | ( ~n6306 & n7730 ) ;
  assign n14286 = ( ~n4199 & n14284 ) | ( ~n4199 & n14285 ) | ( n14284 & n14285 ) ;
  assign n14287 = ~n925 & n9005 ;
  assign n14288 = n8576 & n14287 ;
  assign n14289 = ( ~n1466 & n8831 ) | ( ~n1466 & n14288 ) | ( n8831 & n14288 ) ;
  assign n14290 = n14289 ^ n6965 ^ n6343 ;
  assign n14291 = n14286 & ~n14290 ;
  assign n14292 = ( ~x45 & n14283 ) | ( ~x45 & n14291 ) | ( n14283 & n14291 ) ;
  assign n14293 = n8336 ^ n3495 ^ n2908 ;
  assign n14294 = n14293 ^ n13421 ^ n7706 ;
  assign n14295 = ( n10987 & ~n11257 ) | ( n10987 & n13756 ) | ( ~n11257 & n13756 ) ;
  assign n14296 = n7827 ^ n1428 ^ 1'b0 ;
  assign n14297 = n14296 ^ n7329 ^ 1'b0 ;
  assign n14298 = n1770 & n14297 ;
  assign n14299 = n1887 & n3297 ;
  assign n14300 = ~n6173 & n14299 ;
  assign n14301 = n14300 ^ n3998 ^ 1'b0 ;
  assign n14302 = ~n12362 & n14301 ;
  assign n14303 = n14302 ^ n9640 ^ n2257 ;
  assign n14304 = n14303 ^ n6199 ^ n5426 ;
  assign n14305 = n13915 ^ n12881 ^ n8460 ;
  assign n14306 = n1917 & ~n1940 ;
  assign n14307 = n14306 ^ n5779 ^ 1'b0 ;
  assign n14308 = n2151 | n8613 ;
  assign n14309 = n8618 & n14308 ;
  assign n14310 = ~n14307 & n14309 ;
  assign n14311 = n2513 & ~n14310 ;
  assign n14312 = n14305 & n14311 ;
  assign n14313 = ( n5182 & ~n6646 ) | ( n5182 & n11544 ) | ( ~n6646 & n11544 ) ;
  assign n14314 = ( n2720 & ~n8626 ) | ( n2720 & n14313 ) | ( ~n8626 & n14313 ) ;
  assign n14315 = n3149 ^ n2237 ^ n1593 ;
  assign n14316 = n7779 & n14315 ;
  assign n14317 = n14316 ^ n8352 ^ 1'b0 ;
  assign n14318 = n14317 ^ n4791 ^ n4010 ;
  assign n14319 = n14318 ^ n3098 ^ n1377 ;
  assign n14320 = ( n1654 & n11781 ) | ( n1654 & ~n12164 ) | ( n11781 & ~n12164 ) ;
  assign n14321 = n4217 | n12799 ;
  assign n14322 = n14321 ^ n13038 ^ 1'b0 ;
  assign n14323 = n5478 & ~n14322 ;
  assign n14324 = ~n2691 & n14323 ;
  assign n14326 = n7518 ^ n6130 ^ n4884 ;
  assign n14325 = n9067 ^ n4236 ^ n1467 ;
  assign n14327 = n14326 ^ n14325 ^ n364 ;
  assign n14328 = n2501 & ~n13966 ;
  assign n14329 = n14328 ^ n6047 ^ 1'b0 ;
  assign n14330 = n9645 ^ n2976 ^ 1'b0 ;
  assign n14331 = n10456 ^ n5628 ^ 1'b0 ;
  assign n14332 = n1576 & n14331 ;
  assign n14334 = ~n1544 & n1767 ;
  assign n14335 = n14334 ^ n7351 ^ 1'b0 ;
  assign n14336 = n14335 ^ n1911 ^ n212 ;
  assign n14337 = n14336 ^ n3935 ^ n2614 ;
  assign n14333 = ~n2222 & n6657 ;
  assign n14338 = n14337 ^ n14333 ^ 1'b0 ;
  assign n14339 = ( ~n8969 & n14332 ) | ( ~n8969 & n14338 ) | ( n14332 & n14338 ) ;
  assign n14340 = ( n14329 & n14330 ) | ( n14329 & ~n14339 ) | ( n14330 & ~n14339 ) ;
  assign n14341 = n721 | n10257 ;
  assign n14345 = n9768 ^ n5145 ^ 1'b0 ;
  assign n14342 = n9366 ^ n1180 ^ n143 ;
  assign n14343 = n11856 ^ n10353 ^ 1'b0 ;
  assign n14344 = n14342 & ~n14343 ;
  assign n14346 = n14345 ^ n14344 ^ n8104 ;
  assign n14347 = ( n1979 & n2722 ) | ( n1979 & ~n4837 ) | ( n2722 & ~n4837 ) ;
  assign n14348 = ( n8024 & n10118 ) | ( n8024 & n14347 ) | ( n10118 & n14347 ) ;
  assign n14349 = n14348 ^ n7431 ^ n5710 ;
  assign n14350 = n14349 ^ n14081 ^ n8989 ;
  assign n14351 = n9121 ^ n2277 ^ 1'b0 ;
  assign n14352 = n793 | n7284 ;
  assign n14353 = ( ~n6687 & n8647 ) | ( ~n6687 & n14352 ) | ( n8647 & n14352 ) ;
  assign n14354 = ( n550 & n6481 ) | ( n550 & ~n12074 ) | ( n6481 & ~n12074 ) ;
  assign n14355 = ( ~n777 & n14353 ) | ( ~n777 & n14354 ) | ( n14353 & n14354 ) ;
  assign n14356 = n13279 ^ n4119 ^ n1998 ;
  assign n14357 = ( ~n3767 & n6661 ) | ( ~n3767 & n7985 ) | ( n6661 & n7985 ) ;
  assign n14358 = ( ~n1562 & n12098 ) | ( ~n1562 & n14357 ) | ( n12098 & n14357 ) ;
  assign n14359 = ( ~n4147 & n7566 ) | ( ~n4147 & n14358 ) | ( n7566 & n14358 ) ;
  assign n14360 = ( ~n7007 & n8256 ) | ( ~n7007 & n14359 ) | ( n8256 & n14359 ) ;
  assign n14361 = ( n761 & ~n2502 ) | ( n761 & n14360 ) | ( ~n2502 & n14360 ) ;
  assign n14362 = n253 | n9526 ;
  assign n14363 = ( n4481 & n6297 ) | ( n4481 & n14362 ) | ( n6297 & n14362 ) ;
  assign n14364 = ( n2804 & n10852 ) | ( n2804 & n14363 ) | ( n10852 & n14363 ) ;
  assign n14365 = ( n1233 & n4720 ) | ( n1233 & ~n14364 ) | ( n4720 & ~n14364 ) ;
  assign n14367 = n11813 ^ n4255 ^ n3917 ;
  assign n14368 = n14367 ^ n11759 ^ n4146 ;
  assign n14366 = n13597 ^ n10182 ^ 1'b0 ;
  assign n14369 = n14368 ^ n14366 ^ 1'b0 ;
  assign n14370 = n671 & ~n4764 ;
  assign n14371 = n10695 & n14370 ;
  assign n14372 = n10071 ^ n2479 ^ 1'b0 ;
  assign n14373 = ( ~n7788 & n9922 ) | ( ~n7788 & n14372 ) | ( n9922 & n14372 ) ;
  assign n14376 = n12079 ^ n6282 ^ 1'b0 ;
  assign n14377 = n570 & n14376 ;
  assign n14378 = ( n1607 & n12980 ) | ( n1607 & ~n14377 ) | ( n12980 & ~n14377 ) ;
  assign n14374 = n4023 & ~n13787 ;
  assign n14375 = n14374 ^ n5813 ^ 1'b0 ;
  assign n14379 = n14378 ^ n14375 ^ n6798 ;
  assign n14380 = n1669 ^ n1338 ^ 1'b0 ;
  assign n14381 = n596 & n14380 ;
  assign n14382 = n14247 ^ n3067 ^ n2019 ;
  assign n14383 = n7673 & n14382 ;
  assign n14384 = n14383 ^ n13808 ^ 1'b0 ;
  assign n14385 = ( n12696 & n14381 ) | ( n12696 & n14384 ) | ( n14381 & n14384 ) ;
  assign n14386 = n1448 ^ n420 ^ n150 ;
  assign n14387 = n14386 ^ n8240 ^ n342 ;
  assign n14388 = ( ~n2760 & n8027 ) | ( ~n2760 & n14387 ) | ( n8027 & n14387 ) ;
  assign n14389 = n3142 & ~n14388 ;
  assign n14390 = n14319 ^ n13678 ^ n6089 ;
  assign n14391 = n6480 ^ n2751 ^ n2662 ;
  assign n14392 = n14391 ^ n13702 ^ n1153 ;
  assign n14393 = n14392 ^ n3144 ^ 1'b0 ;
  assign n14394 = ( n3017 & n4143 ) | ( n3017 & n6948 ) | ( n4143 & n6948 ) ;
  assign n14395 = ( n5393 & ~n7411 ) | ( n5393 & n12222 ) | ( ~n7411 & n12222 ) ;
  assign n14396 = n14395 ^ n12512 ^ 1'b0 ;
  assign n14397 = n9789 | n12199 ;
  assign n14398 = n14397 ^ n566 ^ 1'b0 ;
  assign n14399 = n644 & ~n8124 ;
  assign n14400 = ( x114 & ~n7116 ) | ( x114 & n11515 ) | ( ~n7116 & n11515 ) ;
  assign n14404 = ( n508 & n519 ) | ( n508 & n7607 ) | ( n519 & n7607 ) ;
  assign n14401 = ( n395 & ~n940 ) | ( n395 & n1181 ) | ( ~n940 & n1181 ) ;
  assign n14402 = n14401 ^ n2341 ^ 1'b0 ;
  assign n14403 = n8875 & n14402 ;
  assign n14405 = n14404 ^ n14403 ^ n6824 ;
  assign n14406 = n1964 ^ n953 ^ n350 ;
  assign n14407 = ( n2713 & n6226 ) | ( n2713 & ~n7408 ) | ( n6226 & ~n7408 ) ;
  assign n14408 = n14407 ^ n1675 ^ 1'b0 ;
  assign n14409 = n14406 | n14408 ;
  assign n14410 = n448 & ~n5348 ;
  assign n14411 = ~n445 & n14410 ;
  assign n14412 = n6925 ^ n2544 ^ n357 ;
  assign n14413 = n5773 & n14412 ;
  assign n14414 = n14413 ^ n4210 ^ 1'b0 ;
  assign n14415 = n14414 ^ n183 ^ 1'b0 ;
  assign n14416 = n14411 | n14415 ;
  assign n14417 = n3353 ^ n2492 ^ x122 ;
  assign n14418 = n7356 | n10634 ;
  assign n14419 = n14417 & ~n14418 ;
  assign n14421 = ( ~n2651 & n4869 ) | ( ~n2651 & n5416 ) | ( n4869 & n5416 ) ;
  assign n14422 = ( ~n2905 & n2972 ) | ( ~n2905 & n14421 ) | ( n2972 & n14421 ) ;
  assign n14423 = n1745 & n14422 ;
  assign n14424 = ~n4061 & n14423 ;
  assign n14420 = ( x121 & ~n774 ) | ( x121 & n5962 ) | ( ~n774 & n5962 ) ;
  assign n14425 = n14424 ^ n14420 ^ n8469 ;
  assign n14426 = n484 & n8115 ;
  assign n14427 = n11967 & n14426 ;
  assign n14428 = ( n6860 & ~n12260 ) | ( n6860 & n12892 ) | ( ~n12260 & n12892 ) ;
  assign n14429 = n14428 ^ n12456 ^ n10237 ;
  assign n14430 = n14429 ^ n1203 ^ 1'b0 ;
  assign n14431 = n644 & ~n1492 ;
  assign n14432 = ( ~n6425 & n10191 ) | ( ~n6425 & n14431 ) | ( n10191 & n14431 ) ;
  assign n14433 = n1213 & ~n12983 ;
  assign n14434 = n14433 ^ n6469 ^ 1'b0 ;
  assign n14435 = n14434 ^ n6119 ^ n3980 ;
  assign n14436 = n6776 ^ n6264 ^ n2457 ;
  assign n14437 = n9214 & n14436 ;
  assign n14438 = ~n14435 & n14437 ;
  assign n14439 = n12385 ^ n3645 ^ n1105 ;
  assign n14440 = n1156 | n14439 ;
  assign n14441 = n14440 ^ n6928 ^ 1'b0 ;
  assign n14442 = ~n1315 & n10217 ;
  assign n14443 = n14442 ^ n242 ^ 1'b0 ;
  assign n14444 = n14443 ^ n2167 ^ n551 ;
  assign n14445 = n13940 ^ n2592 ^ n2310 ;
  assign n14446 = n14444 & ~n14445 ;
  assign n14447 = ~n14441 & n14446 ;
  assign n14451 = n1863 ^ n1381 ^ n256 ;
  assign n14448 = n2663 ^ n1273 ^ 1'b0 ;
  assign n14449 = n3142 & n14448 ;
  assign n14450 = n14449 ^ n4017 ^ n2329 ;
  assign n14452 = n14451 ^ n14450 ^ n2866 ;
  assign n14454 = ( n2619 & n2726 ) | ( n2619 & ~n2998 ) | ( n2726 & ~n2998 ) ;
  assign n14455 = n14454 ^ n12293 ^ n11566 ;
  assign n14456 = ( n6548 & ~n13236 ) | ( n6548 & n14455 ) | ( ~n13236 & n14455 ) ;
  assign n14453 = n8412 ^ n7348 ^ n5271 ;
  assign n14457 = n14456 ^ n14453 ^ n8193 ;
  assign n14458 = ( n2922 & n12334 ) | ( n2922 & n13651 ) | ( n12334 & n13651 ) ;
  assign n14459 = ( n4976 & n9568 ) | ( n4976 & ~n14458 ) | ( n9568 & ~n14458 ) ;
  assign n14460 = n4816 ^ n1641 ^ n1169 ;
  assign n14461 = ( ~n2635 & n14459 ) | ( ~n2635 & n14460 ) | ( n14459 & n14460 ) ;
  assign n14462 = n14461 ^ n7290 ^ n3057 ;
  assign n14463 = ~n7220 & n11411 ;
  assign n14464 = ( n813 & n880 ) | ( n813 & ~n13750 ) | ( n880 & ~n13750 ) ;
  assign n14465 = n14464 ^ n11970 ^ n3540 ;
  assign n14466 = n11301 ^ n11153 ^ n762 ;
  assign n14467 = n1417 & n14466 ;
  assign n14468 = ( n1773 & n6186 ) | ( n1773 & n10922 ) | ( n6186 & n10922 ) ;
  assign n14469 = n14468 ^ n2720 ^ 1'b0 ;
  assign n14470 = n3992 | n9966 ;
  assign n14471 = n5735 & ~n14470 ;
  assign n14472 = ( ~n6792 & n6839 ) | ( ~n6792 & n14032 ) | ( n6839 & n14032 ) ;
  assign n14473 = n423 & ~n6770 ;
  assign n14475 = n9885 | n13713 ;
  assign n14474 = n2721 | n10899 ;
  assign n14476 = n14475 ^ n14474 ^ 1'b0 ;
  assign n14477 = ( n1314 & n3782 ) | ( n1314 & n6291 ) | ( n3782 & n6291 ) ;
  assign n14478 = n14477 ^ n2384 ^ x21 ;
  assign n14479 = n14478 ^ n4341 ^ x82 ;
  assign n14480 = ( n5125 & n5425 ) | ( n5125 & n10876 ) | ( n5425 & n10876 ) ;
  assign n14481 = ( ~n4630 & n6868 ) | ( ~n4630 & n7851 ) | ( n6868 & n7851 ) ;
  assign n14482 = ( ~n364 & n5129 ) | ( ~n364 & n14481 ) | ( n5129 & n14481 ) ;
  assign n14483 = ( ~n167 & n9594 ) | ( ~n167 & n10503 ) | ( n9594 & n10503 ) ;
  assign n14484 = n14483 ^ n4455 ^ n3042 ;
  assign n14485 = n13328 ^ n10360 ^ 1'b0 ;
  assign n14486 = n14484 | n14485 ;
  assign n14491 = n623 | n11001 ;
  assign n14492 = n14491 ^ n3145 ^ 1'b0 ;
  assign n14487 = n2268 | n6761 ;
  assign n14488 = n4660 | n5671 ;
  assign n14489 = n14488 ^ n7251 ^ 1'b0 ;
  assign n14490 = ( n720 & ~n14487 ) | ( n720 & n14489 ) | ( ~n14487 & n14489 ) ;
  assign n14493 = n14492 ^ n14490 ^ n7233 ;
  assign n14494 = n14493 ^ n3928 ^ n3581 ;
  assign n14495 = n1806 | n4160 ;
  assign n14496 = n14495 ^ n4868 ^ 1'b0 ;
  assign n14497 = n3204 | n14496 ;
  assign n14500 = ~n8004 & n13097 ;
  assign n14498 = n3634 ^ n2427 ^ x102 ;
  assign n14499 = ( n788 & n1822 ) | ( n788 & ~n14498 ) | ( n1822 & ~n14498 ) ;
  assign n14501 = n14500 ^ n14499 ^ n3146 ;
  assign n14502 = n14501 ^ n12287 ^ 1'b0 ;
  assign n14503 = n1100 ^ n523 ^ 1'b0 ;
  assign n14504 = n5007 ^ n4612 ^ n346 ;
  assign n14505 = n14504 ^ n7776 ^ n6423 ;
  assign n14506 = n14505 ^ n9640 ^ n968 ;
  assign n14507 = ( n2316 & n14503 ) | ( n2316 & ~n14506 ) | ( n14503 & ~n14506 ) ;
  assign n14508 = ~n13770 & n14507 ;
  assign n14509 = n4671 ^ n1210 ^ 1'b0 ;
  assign n14510 = x120 & n14509 ;
  assign n14511 = n2624 & n14510 ;
  assign n14512 = n14098 ^ x85 ^ 1'b0 ;
  assign n14513 = n14512 ^ n3980 ^ n1539 ;
  assign n14514 = x94 & ~n1674 ;
  assign n14515 = n14514 ^ n1940 ^ 1'b0 ;
  assign n14516 = n14515 ^ n11136 ^ x67 ;
  assign n14517 = ( n4079 & n13606 ) | ( n4079 & ~n14516 ) | ( n13606 & ~n14516 ) ;
  assign n14518 = ( n1371 & ~n2191 ) | ( n1371 & n14517 ) | ( ~n2191 & n14517 ) ;
  assign n14519 = ( n4550 & n14082 ) | ( n4550 & n14518 ) | ( n14082 & n14518 ) ;
  assign n14520 = ( n7721 & n12965 ) | ( n7721 & ~n14125 ) | ( n12965 & ~n14125 ) ;
  assign n14521 = ( n6580 & ~n6655 ) | ( n6580 & n14520 ) | ( ~n6655 & n14520 ) ;
  assign n14522 = n3052 & n3618 ;
  assign n14523 = n14522 ^ n9336 ^ 1'b0 ;
  assign n14524 = ~n419 & n849 ;
  assign n14525 = ( n1933 & n4404 ) | ( n1933 & ~n14524 ) | ( n4404 & ~n14524 ) ;
  assign n14526 = n6913 & ~n14525 ;
  assign n14527 = n14526 ^ n10242 ^ n8358 ;
  assign n14528 = ( n2868 & n7791 ) | ( n2868 & ~n12049 ) | ( n7791 & ~n12049 ) ;
  assign n14529 = ( ~n7675 & n10779 ) | ( ~n7675 & n14528 ) | ( n10779 & n14528 ) ;
  assign n14530 = n12391 ^ n9595 ^ n3933 ;
  assign n14531 = n14530 ^ n8272 ^ n5924 ;
  assign n14532 = n2806 ^ n1055 ^ n1005 ;
  assign n14533 = ( n2235 & ~n6511 ) | ( n2235 & n14532 ) | ( ~n6511 & n14532 ) ;
  assign n14534 = n11778 ^ n4806 ^ 1'b0 ;
  assign n14537 = n3116 & ~n6183 ;
  assign n14538 = ~n3078 & n14537 ;
  assign n14535 = n11855 ^ n10136 ^ n8513 ;
  assign n14536 = n14535 ^ n5904 ^ n2289 ;
  assign n14539 = n14538 ^ n14536 ^ n5803 ;
  assign n14540 = n14534 | n14539 ;
  assign n14541 = n4969 & ~n14540 ;
  assign n14542 = ( ~n6234 & n14533 ) | ( ~n6234 & n14541 ) | ( n14533 & n14541 ) ;
  assign n14543 = n5759 ^ n5171 ^ 1'b0 ;
  assign n14544 = ~n9952 & n14543 ;
  assign n14546 = n1003 & n1225 ;
  assign n14547 = n14546 ^ n1361 ^ 1'b0 ;
  assign n14545 = ( n720 & ~n4681 ) | ( n720 & n7950 ) | ( ~n4681 & n7950 ) ;
  assign n14548 = n14547 ^ n14545 ^ n10609 ;
  assign n14549 = ( n3810 & ~n10273 ) | ( n3810 & n14548 ) | ( ~n10273 & n14548 ) ;
  assign n14551 = ( ~n554 & n3391 ) | ( ~n554 & n6340 ) | ( n3391 & n6340 ) ;
  assign n14552 = n3822 & n14551 ;
  assign n14553 = ( ~n1772 & n2082 ) | ( ~n1772 & n14552 ) | ( n2082 & n14552 ) ;
  assign n14550 = n12256 ^ n9470 ^ n5190 ;
  assign n14554 = n14553 ^ n14550 ^ n382 ;
  assign n14555 = n4508 ^ n1395 ^ 1'b0 ;
  assign n14556 = ( n4281 & n14554 ) | ( n4281 & ~n14555 ) | ( n14554 & ~n14555 ) ;
  assign n14557 = ( n3573 & ~n4925 ) | ( n3573 & n7409 ) | ( ~n4925 & n7409 ) ;
  assign n14558 = ( n3981 & n9762 ) | ( n3981 & n14557 ) | ( n9762 & n14557 ) ;
  assign n14565 = ( x121 & n5980 ) | ( x121 & ~n10518 ) | ( n5980 & ~n10518 ) ;
  assign n14559 = n5721 ^ n2786 ^ n149 ;
  assign n14560 = ( n932 & ~n1644 ) | ( n932 & n8295 ) | ( ~n1644 & n8295 ) ;
  assign n14561 = ( n2331 & n12970 ) | ( n2331 & n14560 ) | ( n12970 & n14560 ) ;
  assign n14562 = ~n8012 & n10188 ;
  assign n14563 = ~n14561 & n14562 ;
  assign n14564 = n14559 & n14563 ;
  assign n14566 = n14565 ^ n14564 ^ n4327 ;
  assign n14569 = n10712 ^ n5173 ^ n1735 ;
  assign n14570 = ( n1334 & n7196 ) | ( n1334 & n7964 ) | ( n7196 & n7964 ) ;
  assign n14571 = ( n1536 & ~n14569 ) | ( n1536 & n14570 ) | ( ~n14569 & n14570 ) ;
  assign n14567 = n772 & ~n8528 ;
  assign n14568 = n3952 | n14567 ;
  assign n14572 = n14571 ^ n14568 ^ n14347 ;
  assign n14573 = n5997 ^ n2383 ^ 1'b0 ;
  assign n14574 = ( n1214 & n8852 ) | ( n1214 & n14506 ) | ( n8852 & n14506 ) ;
  assign n14575 = n1290 ^ n727 ^ 1'b0 ;
  assign n14576 = n14109 & n14575 ;
  assign n14577 = n10463 ^ n7893 ^ x5 ;
  assign n14578 = ~n220 & n14001 ;
  assign n14579 = n1936 & n14578 ;
  assign n14580 = ( n2472 & n14577 ) | ( n2472 & ~n14579 ) | ( n14577 & ~n14579 ) ;
  assign n14581 = n8822 ^ n8729 ^ n1988 ;
  assign n14582 = n14581 ^ n9484 ^ x112 ;
  assign n14583 = n4452 & ~n6107 ;
  assign n14584 = ~n644 & n14583 ;
  assign n14585 = ( n6778 & ~n8044 ) | ( n6778 & n14584 ) | ( ~n8044 & n14584 ) ;
  assign n14586 = n6677 & n14585 ;
  assign n14587 = n2156 | n6942 ;
  assign n14588 = n3158 | n14587 ;
  assign n14596 = n11189 ^ n1829 ^ n881 ;
  assign n14597 = ( n4440 & n7974 ) | ( n4440 & n14596 ) | ( n7974 & n14596 ) ;
  assign n14594 = n12145 ^ n10365 ^ 1'b0 ;
  assign n14590 = n7039 & ~n10133 ;
  assign n14591 = n14590 ^ n6009 ^ 1'b0 ;
  assign n14589 = n11484 ^ n4455 ^ n1863 ;
  assign n14592 = n14591 ^ n14589 ^ n3066 ;
  assign n14593 = ( ~n4331 & n12453 ) | ( ~n4331 & n14592 ) | ( n12453 & n14592 ) ;
  assign n14595 = n14594 ^ n14593 ^ n5014 ;
  assign n14598 = n14597 ^ n14595 ^ n2853 ;
  assign n14599 = n11397 ^ n8708 ^ n7790 ;
  assign n14600 = n14599 ^ n12820 ^ n3829 ;
  assign n14601 = n8920 ^ n4669 ^ n667 ;
  assign n14602 = n4434 ^ n1707 ^ n840 ;
  assign n14603 = ( ~n329 & n9854 ) | ( ~n329 & n14602 ) | ( n9854 & n14602 ) ;
  assign n14604 = ( ~n8317 & n10685 ) | ( ~n8317 & n14603 ) | ( n10685 & n14603 ) ;
  assign n14605 = ~n1357 & n5495 ;
  assign n14606 = n12881 ^ n1235 ^ n529 ;
  assign n14607 = n2105 & ~n9468 ;
  assign n14608 = n14607 ^ n7218 ^ 1'b0 ;
  assign n14609 = ( n584 & n694 ) | ( n584 & ~n14608 ) | ( n694 & ~n14608 ) ;
  assign n14610 = ( ~n11704 & n12799 ) | ( ~n11704 & n14609 ) | ( n12799 & n14609 ) ;
  assign n14611 = ( n4881 & n12268 ) | ( n4881 & n14610 ) | ( n12268 & n14610 ) ;
  assign n14612 = n14611 ^ n14088 ^ n2558 ;
  assign n14613 = ( n8532 & n14606 ) | ( n8532 & n14612 ) | ( n14606 & n14612 ) ;
  assign n14614 = ( n2473 & ~n2822 ) | ( n2473 & n4871 ) | ( ~n2822 & n4871 ) ;
  assign n14615 = n14614 ^ n10164 ^ n3158 ;
  assign n14616 = n14615 ^ n11290 ^ 1'b0 ;
  assign n14617 = ~n13515 & n14616 ;
  assign n14618 = n6383 ^ n3230 ^ 1'b0 ;
  assign n14619 = n13721 ^ n3281 ^ n1061 ;
  assign n14620 = n586 | n14619 ;
  assign n14621 = n7958 ^ n6523 ^ n394 ;
  assign n14622 = ( n1182 & n11170 ) | ( n1182 & n14621 ) | ( n11170 & n14621 ) ;
  assign n14623 = ( n4136 & ~n4597 ) | ( n4136 & n5636 ) | ( ~n4597 & n5636 ) ;
  assign n14624 = n14623 ^ n9251 ^ n2077 ;
  assign n14625 = n14624 ^ n5909 ^ n1375 ;
  assign n14626 = ( n4629 & n6340 ) | ( n4629 & ~n14625 ) | ( n6340 & ~n14625 ) ;
  assign n14627 = n2777 | n3466 ;
  assign n14628 = n5262 ^ n2642 ^ 1'b0 ;
  assign n14629 = n14627 & ~n14628 ;
  assign n14630 = n8313 ^ n5044 ^ 1'b0 ;
  assign n14631 = ( n3103 & n3972 ) | ( n3103 & n6212 ) | ( n3972 & n6212 ) ;
  assign n14632 = ( n11806 & n12277 ) | ( n11806 & n14631 ) | ( n12277 & n14631 ) ;
  assign n14633 = ( ~n2649 & n11220 ) | ( ~n2649 & n14552 ) | ( n11220 & n14552 ) ;
  assign n14634 = n4272 ^ n2947 ^ n404 ;
  assign n14635 = n14634 ^ n9998 ^ n2820 ;
  assign n14636 = ( ~n3020 & n6891 ) | ( ~n3020 & n8922 ) | ( n6891 & n8922 ) ;
  assign n14638 = n2968 ^ n1306 ^ 1'b0 ;
  assign n14637 = n14545 ^ n6131 ^ n4730 ;
  assign n14639 = n14638 ^ n14637 ^ n6507 ;
  assign n14640 = n7898 ^ n7586 ^ n5307 ;
  assign n14641 = n14640 ^ n11883 ^ n2485 ;
  assign n14642 = ( ~x38 & n3721 ) | ( ~x38 & n9575 ) | ( n3721 & n9575 ) ;
  assign n14643 = n14642 ^ n2363 ^ 1'b0 ;
  assign n14644 = ~n10335 & n14643 ;
  assign n14645 = ( n2749 & n9224 ) | ( n2749 & n14644 ) | ( n9224 & n14644 ) ;
  assign n14646 = ( n1417 & n14641 ) | ( n1417 & n14645 ) | ( n14641 & n14645 ) ;
  assign n14647 = ~n8187 & n14646 ;
  assign n14648 = n14639 & n14647 ;
  assign n14649 = ( n1148 & n4189 ) | ( n1148 & n12967 ) | ( n4189 & n12967 ) ;
  assign n14650 = ~n9216 & n14649 ;
  assign n14651 = ~n8682 & n14650 ;
  assign n14652 = n8890 ^ n5701 ^ n5352 ;
  assign n14653 = ( ~n11489 & n13374 ) | ( ~n11489 & n14652 ) | ( n13374 & n14652 ) ;
  assign n14654 = ( n4948 & n7103 ) | ( n4948 & ~n14653 ) | ( n7103 & ~n14653 ) ;
  assign n14655 = ( n7727 & ~n14651 ) | ( n7727 & n14654 ) | ( ~n14651 & n14654 ) ;
  assign n14656 = ( n1064 & ~n3416 ) | ( n1064 & n12584 ) | ( ~n3416 & n12584 ) ;
  assign n14657 = n4663 | n14656 ;
  assign n14658 = n11810 ^ n8982 ^ n849 ;
  assign n14659 = n14004 ^ n12480 ^ n9285 ;
  assign n14660 = n7475 & n14659 ;
  assign n14661 = n811 & n9501 ;
  assign n14662 = n8595 | n14661 ;
  assign n14663 = n14660 | n14662 ;
  assign n14664 = ( n2433 & n5318 ) | ( n2433 & ~n6867 ) | ( n5318 & ~n6867 ) ;
  assign n14665 = n411 & ~n14664 ;
  assign n14666 = n14665 ^ n11937 ^ n11250 ;
  assign n14667 = n11891 ^ n11883 ^ 1'b0 ;
  assign n14668 = n2800 ^ n2348 ^ n1876 ;
  assign n14669 = n14668 ^ n7409 ^ n4136 ;
  assign n14670 = ~n345 & n14669 ;
  assign n14671 = n14670 ^ n6723 ^ n6345 ;
  assign n14672 = n8196 & n14671 ;
  assign n14673 = n3851 & n14672 ;
  assign n14674 = n12614 | n14673 ;
  assign n14677 = n951 ^ n806 ^ x24 ;
  assign n14678 = n7394 | n14677 ;
  assign n14679 = n14678 ^ n9124 ^ 1'b0 ;
  assign n14680 = n14679 ^ n8998 ^ n6075 ;
  assign n14675 = ~n1938 & n9965 ;
  assign n14676 = n14675 ^ n12029 ^ n2688 ;
  assign n14681 = n14680 ^ n14676 ^ 1'b0 ;
  assign n14682 = n4802 & ~n5283 ;
  assign n14683 = n14682 ^ n3950 ^ n2182 ;
  assign n14684 = n11412 ^ n2322 ^ n1818 ;
  assign n14685 = n3115 & n6802 ;
  assign n14686 = n3746 ^ n1091 ^ n670 ;
  assign n14687 = n3792 & ~n10594 ;
  assign n14688 = n14687 ^ n11948 ^ n502 ;
  assign n14689 = ( n6967 & n14686 ) | ( n6967 & n14688 ) | ( n14686 & n14688 ) ;
  assign n14690 = ( n1655 & n2588 ) | ( n1655 & ~n8626 ) | ( n2588 & ~n8626 ) ;
  assign n14691 = ( n3587 & n12688 ) | ( n3587 & ~n14690 ) | ( n12688 & ~n14690 ) ;
  assign n14692 = n14691 ^ n14548 ^ n6413 ;
  assign n14693 = ( n1578 & n4697 ) | ( n1578 & ~n5486 ) | ( n4697 & ~n5486 ) ;
  assign n14694 = ~n2470 & n7468 ;
  assign n14695 = n14693 & n14694 ;
  assign n14696 = ( ~n6315 & n6524 ) | ( ~n6315 & n14695 ) | ( n6524 & n14695 ) ;
  assign n14697 = n14696 ^ n11770 ^ n4791 ;
  assign n14698 = n1490 & ~n4004 ;
  assign n14699 = n374 & n14698 ;
  assign n14700 = ( n8549 & n14359 ) | ( n8549 & ~n14699 ) | ( n14359 & ~n14699 ) ;
  assign n14704 = n11156 ^ n184 ^ 1'b0 ;
  assign n14701 = n6306 ^ n3771 ^ 1'b0 ;
  assign n14702 = n1918 & ~n14701 ;
  assign n14703 = x93 | n14702 ;
  assign n14705 = n14704 ^ n14703 ^ 1'b0 ;
  assign n14706 = n7544 & ~n7930 ;
  assign n14707 = n14706 ^ n6391 ^ 1'b0 ;
  assign n14709 = ( n1092 & n1267 ) | ( n1092 & ~n2004 ) | ( n1267 & ~n2004 ) ;
  assign n14708 = ~n2547 & n13236 ;
  assign n14710 = n14709 ^ n14708 ^ 1'b0 ;
  assign n14715 = n4900 & n9685 ;
  assign n14716 = n14715 ^ n248 ^ 1'b0 ;
  assign n14712 = ( n923 & n2304 ) | ( n923 & ~n11115 ) | ( n2304 & ~n11115 ) ;
  assign n14713 = n14712 ^ n12661 ^ n5701 ;
  assign n14714 = ~n12881 & n14713 ;
  assign n14717 = n14716 ^ n14714 ^ 1'b0 ;
  assign n14711 = n14535 ^ n3535 ^ n256 ;
  assign n14718 = n14717 ^ n14711 ^ n12791 ;
  assign n14719 = n13375 | n14478 ;
  assign n14721 = n3096 ^ n3053 ^ 1'b0 ;
  assign n14722 = ( ~n987 & n5516 ) | ( ~n987 & n14721 ) | ( n5516 & n14721 ) ;
  assign n14720 = n6985 & ~n8602 ;
  assign n14723 = n14722 ^ n14720 ^ 1'b0 ;
  assign n14724 = n8763 ^ n1438 ^ 1'b0 ;
  assign n14725 = n10109 ^ n8755 ^ 1'b0 ;
  assign n14726 = n14725 ^ n14679 ^ 1'b0 ;
  assign n14727 = ( x43 & ~n3048 ) | ( x43 & n4132 ) | ( ~n3048 & n4132 ) ;
  assign n14728 = n8039 ^ n823 ^ n466 ;
  assign n14729 = n14728 ^ n5127 ^ n4092 ;
  assign n14730 = ~n7684 & n13801 ;
  assign n14731 = n14730 ^ n3964 ^ n3666 ;
  assign n14732 = n14731 ^ n7111 ^ 1'b0 ;
  assign n14733 = n14729 & n14732 ;
  assign n14734 = n13308 ^ n11373 ^ n5366 ;
  assign n14735 = n14712 ^ n7171 ^ 1'b0 ;
  assign n14736 = ~n941 & n14735 ;
  assign n14737 = ( n6798 & ~n14734 ) | ( n6798 & n14736 ) | ( ~n14734 & n14736 ) ;
  assign n14743 = n6903 ^ n3500 ^ n2398 ;
  assign n14742 = ( n514 & n5163 ) | ( n514 & n6026 ) | ( n5163 & n6026 ) ;
  assign n14744 = n14743 ^ n14742 ^ 1'b0 ;
  assign n14745 = n2932 & ~n14744 ;
  assign n14740 = ( n1805 & n2055 ) | ( n1805 & n4871 ) | ( n2055 & n4871 ) ;
  assign n14741 = n8836 & ~n14740 ;
  assign n14746 = n14745 ^ n14741 ^ 1'b0 ;
  assign n14738 = ( n1019 & ~n3342 ) | ( n1019 & n4224 ) | ( ~n3342 & n4224 ) ;
  assign n14739 = n6308 & ~n14738 ;
  assign n14747 = n14746 ^ n14739 ^ 1'b0 ;
  assign n14748 = n14747 ^ n11398 ^ 1'b0 ;
  assign n14749 = n14748 ^ n9067 ^ n2908 ;
  assign n14750 = ( x72 & ~n2114 ) | ( x72 & n8531 ) | ( ~n2114 & n8531 ) ;
  assign n14751 = n14750 ^ n3982 ^ 1'b0 ;
  assign n14752 = n13634 & n14751 ;
  assign n14753 = n7974 ^ n1735 ^ 1'b0 ;
  assign n14754 = ( n6169 & n14752 ) | ( n6169 & ~n14753 ) | ( n14752 & ~n14753 ) ;
  assign n14755 = n14754 ^ n8033 ^ 1'b0 ;
  assign n14756 = n14755 ^ n12559 ^ n2408 ;
  assign n14757 = ( n529 & ~n964 ) | ( n529 & n7379 ) | ( ~n964 & n7379 ) ;
  assign n14758 = n14336 ^ n9899 ^ 1'b0 ;
  assign n14759 = ( x19 & ~n2376 ) | ( x19 & n5020 ) | ( ~n2376 & n5020 ) ;
  assign n14760 = ( n3130 & ~n3235 ) | ( n3130 & n14759 ) | ( ~n3235 & n14759 ) ;
  assign n14762 = ( n1999 & n6373 ) | ( n1999 & ~n8382 ) | ( n6373 & ~n8382 ) ;
  assign n14761 = ( x105 & n551 ) | ( x105 & n8032 ) | ( n551 & n8032 ) ;
  assign n14763 = n14762 ^ n14761 ^ n14008 ;
  assign n14764 = n2855 & ~n14763 ;
  assign n14765 = n5641 | n11327 ;
  assign n14766 = n14765 ^ n7802 ^ 1'b0 ;
  assign n14767 = n1820 | n14460 ;
  assign n14769 = ~n1743 & n7129 ;
  assign n14770 = n1942 & n14769 ;
  assign n14768 = n9669 ^ n9172 ^ n4207 ;
  assign n14771 = n14770 ^ n14768 ^ n7762 ;
  assign n14772 = ( ~n1898 & n4058 ) | ( ~n1898 & n6212 ) | ( n4058 & n6212 ) ;
  assign n14773 = n9861 ^ n6545 ^ n2010 ;
  assign n14774 = n10646 ^ n1742 ^ 1'b0 ;
  assign n14776 = n13018 ^ n7052 ^ n4368 ;
  assign n14775 = n1340 & ~n10314 ;
  assign n14777 = n14776 ^ n14775 ^ 1'b0 ;
  assign n14778 = ( n11830 & n14774 ) | ( n11830 & n14777 ) | ( n14774 & n14777 ) ;
  assign n14779 = n4221 | n7104 ;
  assign n14780 = n14517 ^ n3288 ^ n376 ;
  assign n14781 = n14780 ^ n8084 ^ n5208 ;
  assign n14782 = ( ~n8065 & n8849 ) | ( ~n8065 & n9005 ) | ( n8849 & n9005 ) ;
  assign n14783 = n5511 ^ n5413 ^ n4220 ;
  assign n14784 = ~n5103 & n5740 ;
  assign n14785 = ( n1152 & n12265 ) | ( n1152 & n14784 ) | ( n12265 & n14784 ) ;
  assign n14788 = n7023 ^ n3908 ^ n943 ;
  assign n14786 = ( n301 & n2244 ) | ( n301 & ~n4377 ) | ( n2244 & ~n4377 ) ;
  assign n14787 = ( ~n11754 & n11857 ) | ( ~n11754 & n14786 ) | ( n11857 & n14786 ) ;
  assign n14789 = n14788 ^ n14787 ^ n6262 ;
  assign n14790 = n14789 ^ n13725 ^ n9534 ;
  assign n14791 = n9264 ^ n3373 ^ n3129 ;
  assign n14792 = ( n3485 & n5419 ) | ( n3485 & n14791 ) | ( n5419 & n14791 ) ;
  assign n14794 = n489 | n1178 ;
  assign n14795 = n14794 ^ n3980 ^ 1'b0 ;
  assign n14796 = n14795 ^ n1472 ^ n149 ;
  assign n14793 = n13669 ^ n11375 ^ 1'b0 ;
  assign n14797 = n14796 ^ n14793 ^ n8977 ;
  assign n14798 = ( n7091 & n7350 ) | ( n7091 & n13271 ) | ( n7350 & n13271 ) ;
  assign n14799 = ( n1516 & n4504 ) | ( n1516 & n5922 ) | ( n4504 & n5922 ) ;
  assign n14810 = ( n3268 & ~n9797 ) | ( n3268 & n13695 ) | ( ~n9797 & n13695 ) ;
  assign n14809 = n5763 ^ n4399 ^ n3880 ;
  assign n14811 = n14810 ^ n14809 ^ n980 ;
  assign n14802 = n6373 ^ n4895 ^ 1'b0 ;
  assign n14800 = n6921 ^ n1360 ^ n329 ;
  assign n14801 = n14800 ^ n2839 ^ n1876 ;
  assign n14803 = n14802 ^ n14801 ^ n10681 ;
  assign n14804 = n14803 ^ n8671 ^ n6134 ;
  assign n14805 = ( n4460 & n5064 ) | ( n4460 & ~n14545 ) | ( n5064 & ~n14545 ) ;
  assign n14806 = n8223 ^ n3721 ^ n1387 ;
  assign n14807 = ~n14805 & n14806 ;
  assign n14808 = ( n7954 & ~n14804 ) | ( n7954 & n14807 ) | ( ~n14804 & n14807 ) ;
  assign n14812 = n14811 ^ n14808 ^ n13758 ;
  assign n14813 = n8154 ^ n501 ^ x48 ;
  assign n14814 = ( n3485 & ~n6559 ) | ( n3485 & n6568 ) | ( ~n6559 & n6568 ) ;
  assign n14815 = ~n7363 & n14814 ;
  assign n14816 = n14815 ^ n13036 ^ 1'b0 ;
  assign n14817 = n7928 ^ n4089 ^ 1'b0 ;
  assign n14818 = ( n381 & n2681 ) | ( n381 & ~n11877 ) | ( n2681 & ~n11877 ) ;
  assign n14819 = ( n710 & n3610 ) | ( n710 & ~n5253 ) | ( n3610 & ~n5253 ) ;
  assign n14820 = ( n2524 & n8032 ) | ( n2524 & n14819 ) | ( n8032 & n14819 ) ;
  assign n14821 = ( n2792 & ~n11275 ) | ( n2792 & n14820 ) | ( ~n11275 & n14820 ) ;
  assign n14822 = ( ~n2761 & n14818 ) | ( ~n2761 & n14821 ) | ( n14818 & n14821 ) ;
  assign n14823 = ( n13434 & ~n14817 ) | ( n13434 & n14822 ) | ( ~n14817 & n14822 ) ;
  assign n14824 = n5729 ^ x91 ^ 1'b0 ;
  assign n14825 = n14824 ^ n9035 ^ 1'b0 ;
  assign n14826 = n6959 ^ n5520 ^ 1'b0 ;
  assign n14827 = n14826 ^ n5813 ^ 1'b0 ;
  assign n14828 = n14827 ^ n1930 ^ x124 ;
  assign n14829 = n5546 ^ n2880 ^ 1'b0 ;
  assign n14830 = ( n4377 & n10119 ) | ( n4377 & n14829 ) | ( n10119 & n14829 ) ;
  assign n14831 = n14830 ^ n11909 ^ 1'b0 ;
  assign n14833 = n10476 ^ n6365 ^ n1674 ;
  assign n14834 = n14833 ^ n5760 ^ n3204 ;
  assign n14832 = ( n1586 & n7612 ) | ( n1586 & ~n9221 ) | ( n7612 & ~n9221 ) ;
  assign n14835 = n14834 ^ n14832 ^ n10195 ;
  assign n14846 = n2652 ^ n480 ^ 1'b0 ;
  assign n14847 = ~n1265 & n14846 ;
  assign n14848 = n14847 ^ n3915 ^ n3877 ;
  assign n14849 = n5000 | n11735 ;
  assign n14850 = n14849 ^ n6318 ^ 1'b0 ;
  assign n14851 = ( ~n13984 & n14848 ) | ( ~n13984 & n14850 ) | ( n14848 & n14850 ) ;
  assign n14852 = n6536 & ~n14851 ;
  assign n14853 = n14852 ^ n226 ^ 1'b0 ;
  assign n14844 = ( n207 & n3417 ) | ( n207 & ~n6587 ) | ( n3417 & ~n6587 ) ;
  assign n14843 = n6635 | n9537 ;
  assign n14836 = n14402 ^ n12128 ^ n7477 ;
  assign n14837 = n14551 ^ n3382 ^ 1'b0 ;
  assign n14838 = n14836 & ~n14837 ;
  assign n14839 = ( n2872 & ~n13635 ) | ( n2872 & n14838 ) | ( ~n13635 & n14838 ) ;
  assign n14840 = n3835 ^ n3513 ^ n2652 ;
  assign n14841 = ~n2908 & n14840 ;
  assign n14842 = ~n14839 & n14841 ;
  assign n14845 = n14844 ^ n14843 ^ n14842 ;
  assign n14854 = n14853 ^ n14845 ^ n584 ;
  assign n14855 = n3344 & n11284 ;
  assign n14856 = n14855 ^ n1048 ^ n557 ;
  assign n14857 = ~n572 & n6525 ;
  assign n14858 = ~n14856 & n14857 ;
  assign n14861 = n10686 ^ n4497 ^ n3621 ;
  assign n14859 = ( n1856 & ~n5662 ) | ( n1856 & n9965 ) | ( ~n5662 & n9965 ) ;
  assign n14860 = n14859 ^ n601 ^ 1'b0 ;
  assign n14862 = n14861 ^ n14860 ^ 1'b0 ;
  assign n14863 = n3523 ^ n1101 ^ 1'b0 ;
  assign n14864 = ~n2635 & n14863 ;
  assign n14865 = ( n11616 & n12390 ) | ( n11616 & n14864 ) | ( n12390 & n14864 ) ;
  assign n14866 = n14865 ^ n3308 ^ n2405 ;
  assign n14867 = n2871 ^ n1728 ^ 1'b0 ;
  assign n14868 = n5485 & ~n14867 ;
  assign n14869 = n8568 ^ n6573 ^ n5028 ;
  assign n14870 = ~n6603 & n14869 ;
  assign n14871 = ~n7031 & n14870 ;
  assign n14872 = ( n11718 & n14868 ) | ( n11718 & n14871 ) | ( n14868 & n14871 ) ;
  assign n14873 = n13649 ^ n5671 ^ x93 ;
  assign n14874 = ~n11894 & n14873 ;
  assign n14875 = n14788 & n14874 ;
  assign n14876 = ~n1912 & n12534 ;
  assign n14878 = n12382 ^ n1488 ^ n251 ;
  assign n14877 = n1596 ^ n912 ^ x123 ;
  assign n14879 = n14878 ^ n14877 ^ n580 ;
  assign n14880 = ( n2452 & n10651 ) | ( n2452 & n14879 ) | ( n10651 & n14879 ) ;
  assign n14881 = ( n12519 & n14876 ) | ( n12519 & ~n14880 ) | ( n14876 & ~n14880 ) ;
  assign n14882 = ( n2740 & n14875 ) | ( n2740 & n14881 ) | ( n14875 & n14881 ) ;
  assign n14883 = n8997 ^ n7849 ^ n5481 ;
  assign n14884 = ( n1127 & n4777 ) | ( n1127 & ~n14883 ) | ( n4777 & ~n14883 ) ;
  assign n14885 = n14884 ^ n9602 ^ 1'b0 ;
  assign n14888 = ( ~n7116 & n10307 ) | ( ~n7116 & n11077 ) | ( n10307 & n11077 ) ;
  assign n14886 = n5286 ^ n5126 ^ n3830 ;
  assign n14887 = n149 | n14886 ;
  assign n14889 = n14888 ^ n14887 ^ n11916 ;
  assign n14890 = n10605 ^ n3131 ^ n2233 ;
  assign n14891 = n14890 ^ n11799 ^ n4381 ;
  assign n14892 = ( ~n3407 & n6600 ) | ( ~n3407 & n14891 ) | ( n6600 & n14891 ) ;
  assign n14893 = ( ~n2083 & n2771 ) | ( ~n2083 & n5967 ) | ( n2771 & n5967 ) ;
  assign n14894 = ( ~n6268 & n6694 ) | ( ~n6268 & n14893 ) | ( n6694 & n14893 ) ;
  assign n14895 = ( n3158 & ~n14892 ) | ( n3158 & n14894 ) | ( ~n14892 & n14894 ) ;
  assign n14896 = n9169 ^ n4133 ^ n1562 ;
  assign n14897 = ( ~n4214 & n5803 ) | ( ~n4214 & n14896 ) | ( n5803 & n14896 ) ;
  assign n14898 = x66 & n14897 ;
  assign n14899 = n14898 ^ n2249 ^ 1'b0 ;
  assign n14905 = n3121 ^ n1862 ^ n532 ;
  assign n14903 = n885 & ~n12774 ;
  assign n14904 = n14903 ^ n13242 ^ 1'b0 ;
  assign n14906 = n14905 ^ n14904 ^ n5730 ;
  assign n14900 = ~n6261 & n13570 ;
  assign n14901 = n8113 & n14900 ;
  assign n14902 = n988 | n14901 ;
  assign n14907 = n14906 ^ n14902 ^ 1'b0 ;
  assign n14908 = n14907 ^ n11354 ^ n6685 ;
  assign n14914 = ( n3621 & n8370 ) | ( n3621 & ~n12970 ) | ( n8370 & ~n12970 ) ;
  assign n14909 = ( n410 & n5318 ) | ( n410 & n5665 ) | ( n5318 & n5665 ) ;
  assign n14911 = n6411 ^ n1710 ^ n1675 ;
  assign n14910 = ( ~n5224 & n6391 ) | ( ~n5224 & n7557 ) | ( n6391 & n7557 ) ;
  assign n14912 = n14911 ^ n14910 ^ 1'b0 ;
  assign n14913 = n14909 & ~n14912 ;
  assign n14915 = n14914 ^ n14913 ^ n7516 ;
  assign n14916 = n14915 ^ n8349 ^ n1234 ;
  assign n14917 = n11236 ^ n7712 ^ n3038 ;
  assign n14918 = n9187 & n14917 ;
  assign n14919 = n2294 | n11162 ;
  assign n14920 = n12742 & ~n14919 ;
  assign n14921 = ( n1499 & n2872 ) | ( n1499 & n6218 ) | ( n2872 & n6218 ) ;
  assign n14922 = ( n3610 & n14920 ) | ( n3610 & n14921 ) | ( n14920 & n14921 ) ;
  assign n14923 = n6639 ^ n5389 ^ n1205 ;
  assign n14924 = ( x83 & n14444 ) | ( x83 & ~n14923 ) | ( n14444 & ~n14923 ) ;
  assign n14927 = n3855 ^ n804 ^ n153 ;
  assign n14925 = ~n2924 & n5306 ;
  assign n14926 = n14925 ^ n14450 ^ n1158 ;
  assign n14928 = n14927 ^ n14926 ^ n14596 ;
  assign n14929 = n1466 | n4073 ;
  assign n14930 = n14929 ^ n3543 ^ 1'b0 ;
  assign n14931 = ( n6054 & ~n8143 ) | ( n6054 & n11451 ) | ( ~n8143 & n11451 ) ;
  assign n14932 = ( n5024 & ~n8647 ) | ( n5024 & n13612 ) | ( ~n8647 & n13612 ) ;
  assign n14933 = n14640 & n14932 ;
  assign n14934 = n3176 & n14933 ;
  assign n14935 = n14934 ^ n8660 ^ 1'b0 ;
  assign n14936 = n14931 & n14935 ;
  assign n14937 = n14533 ^ n8522 ^ n5196 ;
  assign n14938 = n14937 ^ n14492 ^ n8170 ;
  assign n14939 = ( n4003 & ~n13221 ) | ( n4003 & n14938 ) | ( ~n13221 & n14938 ) ;
  assign n14940 = ( n2279 & n10205 ) | ( n2279 & ~n14939 ) | ( n10205 & ~n14939 ) ;
  assign n14941 = n14901 ^ n2122 ^ n629 ;
  assign n14942 = n3342 | n5566 ;
  assign n14943 = ( n8998 & n14941 ) | ( n8998 & n14942 ) | ( n14941 & n14942 ) ;
  assign n14944 = ( n12496 & ~n14940 ) | ( n12496 & n14943 ) | ( ~n14940 & n14943 ) ;
  assign n14945 = n2220 ^ n1647 ^ n1388 ;
  assign n14946 = n14945 ^ n12550 ^ n10483 ;
  assign n14947 = n478 & ~n4214 ;
  assign n14948 = n14947 ^ n7434 ^ 1'b0 ;
  assign n14949 = n6400 ^ n2977 ^ 1'b0 ;
  assign n14950 = n7730 ^ n3976 ^ n810 ;
  assign n14951 = n1927 | n14950 ;
  assign n14952 = n14951 ^ n9083 ^ 1'b0 ;
  assign n14953 = n14952 ^ n11056 ^ n5381 ;
  assign n14954 = n14953 ^ n14645 ^ n11564 ;
  assign n14955 = n9152 & n14954 ;
  assign n14956 = ~n145 & n14955 ;
  assign n14957 = ( n5259 & ~n8034 ) | ( n5259 & n8354 ) | ( ~n8034 & n8354 ) ;
  assign n14958 = ( n1589 & n5526 ) | ( n1589 & ~n8149 ) | ( n5526 & ~n8149 ) ;
  assign n14959 = ( n4882 & n14957 ) | ( n4882 & ~n14958 ) | ( n14957 & ~n14958 ) ;
  assign n14960 = n14959 ^ n2509 ^ 1'b0 ;
  assign n14961 = x66 & ~n14960 ;
  assign n14962 = n1298 & n4888 ;
  assign n14963 = ~n12943 & n14962 ;
  assign n14964 = n12472 ^ n6770 ^ n6610 ;
  assign n14965 = n12128 ^ n11462 ^ n1611 ;
  assign n14966 = ( n14963 & n14964 ) | ( n14963 & ~n14965 ) | ( n14964 & ~n14965 ) ;
  assign n14967 = ( ~n5599 & n5618 ) | ( ~n5599 & n14966 ) | ( n5618 & n14966 ) ;
  assign n14968 = ( n6007 & ~n12918 ) | ( n6007 & n13751 ) | ( ~n12918 & n13751 ) ;
  assign n14969 = n14968 ^ n13476 ^ n11820 ;
  assign n14970 = n12648 ^ n3860 ^ n1699 ;
  assign n14971 = n8913 ^ n3520 ^ n1485 ;
  assign n14972 = n12946 & n14971 ;
  assign n14973 = n11868 ^ n9042 ^ n6766 ;
  assign n14974 = n11444 ^ n4587 ^ n3567 ;
  assign n14975 = ( n13839 & n14559 ) | ( n13839 & n14974 ) | ( n14559 & n14974 ) ;
  assign n14981 = n2002 ^ n471 ^ n257 ;
  assign n14976 = n10899 ^ n9767 ^ n2822 ;
  assign n14977 = ( n5836 & ~n5854 ) | ( n5836 & n14976 ) | ( ~n5854 & n14976 ) ;
  assign n14978 = ( ~n5610 & n6630 ) | ( ~n5610 & n14977 ) | ( n6630 & n14977 ) ;
  assign n14979 = n14978 ^ n2023 ^ 1'b0 ;
  assign n14980 = ~n13526 & n14979 ;
  assign n14982 = n14981 ^ n14980 ^ n3193 ;
  assign n14983 = n7381 & n14702 ;
  assign n14984 = n14983 ^ n7979 ^ 1'b0 ;
  assign n14985 = n4321 & n14984 ;
  assign n14986 = ( ~n6218 & n9023 ) | ( ~n6218 & n14985 ) | ( n9023 & n14985 ) ;
  assign n14987 = n7950 ^ n5839 ^ n2446 ;
  assign n14988 = ( n7805 & n8296 ) | ( n7805 & n14987 ) | ( n8296 & n14987 ) ;
  assign n14989 = ( n10417 & n14112 ) | ( n10417 & ~n14988 ) | ( n14112 & ~n14988 ) ;
  assign n14990 = ( n2747 & ~n5435 ) | ( n2747 & n14989 ) | ( ~n5435 & n14989 ) ;
  assign n14991 = n11780 ^ n8130 ^ n4762 ;
  assign n14992 = n3609 ^ n364 ^ x57 ;
  assign n14993 = ( n4681 & n9251 ) | ( n4681 & n14992 ) | ( n9251 & n14992 ) ;
  assign n14994 = n14993 ^ n185 ^ 1'b0 ;
  assign n14995 = ( n832 & n14991 ) | ( n832 & n14994 ) | ( n14991 & n14994 ) ;
  assign n14996 = ( n3956 & n4693 ) | ( n3956 & n11515 ) | ( n4693 & n11515 ) ;
  assign n14997 = n6008 ^ n2575 ^ n2236 ;
  assign n14998 = n14997 ^ n12429 ^ n12007 ;
  assign n14999 = ( n14995 & n14996 ) | ( n14995 & ~n14998 ) | ( n14996 & ~n14998 ) ;
  assign n15000 = ( ~n5625 & n6366 ) | ( ~n5625 & n9705 ) | ( n6366 & n9705 ) ;
  assign n15001 = n4266 ^ n3020 ^ 1'b0 ;
  assign n15002 = ~n1687 & n15001 ;
  assign n15003 = ~n10081 & n15002 ;
  assign n15004 = ~n612 & n15003 ;
  assign n15005 = ( n4428 & n15000 ) | ( n4428 & ~n15004 ) | ( n15000 & ~n15004 ) ;
  assign n15008 = n6046 ^ n5785 ^ n2139 ;
  assign n15006 = ( n5736 & n6931 ) | ( n5736 & n9514 ) | ( n6931 & n9514 ) ;
  assign n15007 = n15006 ^ n648 ^ n493 ;
  assign n15009 = n15008 ^ n15007 ^ n12318 ;
  assign n15010 = n13663 ^ n6396 ^ n6079 ;
  assign n15011 = n767 | n2573 ;
  assign n15012 = n15011 ^ n1178 ^ 1'b0 ;
  assign n15013 = ( ~n768 & n4548 ) | ( ~n768 & n15012 ) | ( n4548 & n15012 ) ;
  assign n15014 = n3232 | n15013 ;
  assign n15015 = ( n2455 & n8759 ) | ( n2455 & n9255 ) | ( n8759 & n9255 ) ;
  assign n15016 = ( n2783 & ~n3524 ) | ( n2783 & n15015 ) | ( ~n3524 & n15015 ) ;
  assign n15017 = ( n10989 & n15014 ) | ( n10989 & ~n15016 ) | ( n15014 & ~n15016 ) ;
  assign n15019 = ( n1542 & n2344 ) | ( n1542 & ~n2550 ) | ( n2344 & ~n2550 ) ;
  assign n15018 = n10885 ^ n2784 ^ n2719 ;
  assign n15020 = n15019 ^ n15018 ^ n10328 ;
  assign n15021 = n8710 ^ n5391 ^ 1'b0 ;
  assign n15022 = ~n1784 & n15013 ;
  assign n15023 = n1465 & ~n6915 ;
  assign n15024 = n15022 & n15023 ;
  assign n15025 = n6896 | n10077 ;
  assign n15026 = n15025 ^ n8092 ^ 1'b0 ;
  assign n15027 = n332 & ~n2741 ;
  assign n15028 = n15027 ^ n12211 ^ 1'b0 ;
  assign n15029 = n15028 ^ n1395 ^ 1'b0 ;
  assign n15030 = n15029 ^ n10565 ^ n6868 ;
  assign n15031 = ( n9418 & n15026 ) | ( n9418 & ~n15030 ) | ( n15026 & ~n15030 ) ;
  assign n15032 = ( ~n7157 & n15024 ) | ( ~n7157 & n15031 ) | ( n15024 & n15031 ) ;
  assign n15033 = ( ~n3396 & n3659 ) | ( ~n3396 & n9663 ) | ( n3659 & n9663 ) ;
  assign n15034 = n15033 ^ n12481 ^ n2038 ;
  assign n15041 = ( ~n346 & n2577 ) | ( ~n346 & n7458 ) | ( n2577 & n7458 ) ;
  assign n15035 = n1348 | n6500 ;
  assign n15036 = n7919 & ~n15035 ;
  assign n15037 = n6250 ^ n597 ^ 1'b0 ;
  assign n15038 = ~n15036 & n15037 ;
  assign n15039 = ~n8986 & n15038 ;
  assign n15040 = ~n10671 & n15039 ;
  assign n15042 = n15041 ^ n15040 ^ n14596 ;
  assign n15043 = n15042 ^ n8382 ^ 1'b0 ;
  assign n15044 = ( n477 & ~n1406 ) | ( n477 & n14591 ) | ( ~n1406 & n14591 ) ;
  assign n15045 = n13438 ^ n2821 ^ 1'b0 ;
  assign n15046 = ( n13680 & n15044 ) | ( n13680 & ~n15045 ) | ( n15044 & ~n15045 ) ;
  assign n15047 = n10735 ^ n8970 ^ n4238 ;
  assign n15048 = n237 & n1455 ;
  assign n15049 = ~n12123 & n15048 ;
  assign n15050 = ( n4861 & n11778 ) | ( n4861 & ~n15049 ) | ( n11778 & ~n15049 ) ;
  assign n15051 = n4529 ^ n4157 ^ 1'b0 ;
  assign n15052 = n1690 & n15051 ;
  assign n15053 = n15052 ^ n12286 ^ n2168 ;
  assign n15054 = n14585 ^ n1855 ^ 1'b0 ;
  assign n15055 = ~n10061 & n15054 ;
  assign n15056 = n15053 & n15055 ;
  assign n15058 = n5964 ^ n2558 ^ 1'b0 ;
  assign n15059 = n15058 ^ n4345 ^ n1715 ;
  assign n15057 = n10025 & n10125 ;
  assign n15060 = n15059 ^ n15057 ^ 1'b0 ;
  assign n15061 = n15060 ^ n10405 ^ n5749 ;
  assign n15062 = ( ~n1116 & n3896 ) | ( ~n1116 & n4220 ) | ( n3896 & n4220 ) ;
  assign n15064 = n12600 ^ n5773 ^ 1'b0 ;
  assign n15065 = ~n598 & n15064 ;
  assign n15066 = ~n8665 & n15065 ;
  assign n15067 = n15066 ^ n7894 ^ 1'b0 ;
  assign n15063 = n5242 ^ n3595 ^ n2486 ;
  assign n15068 = n15067 ^ n15063 ^ n5482 ;
  assign n15069 = n9170 ^ n6487 ^ n1464 ;
  assign n15070 = n15069 ^ n13388 ^ n1781 ;
  assign n15071 = n7425 ^ n2348 ^ x100 ;
  assign n15072 = n15071 ^ n11767 ^ n775 ;
  assign n15073 = n15072 ^ n5619 ^ n4997 ;
  assign n15074 = ( n3316 & ~n7502 ) | ( n3316 & n15073 ) | ( ~n7502 & n15073 ) ;
  assign n15075 = n4224 | n6255 ;
  assign n15076 = n15075 ^ n2042 ^ 1'b0 ;
  assign n15077 = n15076 ^ n8006 ^ 1'b0 ;
  assign n15078 = n5592 | n15077 ;
  assign n15079 = n15078 ^ n3880 ^ n2033 ;
  assign n15082 = n7779 ^ n6642 ^ n1428 ;
  assign n15080 = ( n1617 & n7266 ) | ( n1617 & ~n9324 ) | ( n7266 & ~n9324 ) ;
  assign n15081 = n15080 ^ n3227 ^ n2292 ;
  assign n15083 = n15082 ^ n15081 ^ 1'b0 ;
  assign n15084 = n8694 ^ n4073 ^ n1184 ;
  assign n15085 = n9113 | n11716 ;
  assign n15086 = n11164 & ~n15085 ;
  assign n15087 = ( n12389 & ~n15084 ) | ( n12389 & n15086 ) | ( ~n15084 & n15086 ) ;
  assign n15088 = n11375 ^ n1794 ^ 1'b0 ;
  assign n15089 = n1955 & ~n15088 ;
  assign n15090 = n13125 ^ n5113 ^ n3642 ;
  assign n15091 = ( n2069 & ~n8907 ) | ( n2069 & n15090 ) | ( ~n8907 & n15090 ) ;
  assign n15092 = ( n8573 & n10270 ) | ( n8573 & n15091 ) | ( n10270 & n15091 ) ;
  assign n15093 = ( n3852 & n6090 ) | ( n3852 & n9829 ) | ( n6090 & n9829 ) ;
  assign n15094 = n1472 | n11379 ;
  assign n15095 = ( n3160 & ~n12924 ) | ( n3160 & n15094 ) | ( ~n12924 & n15094 ) ;
  assign n15107 = ( n2841 & n7694 ) | ( n2841 & ~n9753 ) | ( n7694 & ~n9753 ) ;
  assign n15108 = n15107 ^ n3509 ^ 1'b0 ;
  assign n15109 = n11513 & ~n15108 ;
  assign n15104 = ( n2177 & ~n7281 ) | ( n2177 & n10380 ) | ( ~n7281 & n10380 ) ;
  assign n15105 = n183 & ~n6424 ;
  assign n15106 = ~n15104 & n15105 ;
  assign n15098 = x43 & ~n4870 ;
  assign n15099 = n15098 ^ n356 ^ 1'b0 ;
  assign n15100 = n15099 ^ n8691 ^ n2971 ;
  assign n15096 = n7525 ^ n6930 ^ n5555 ;
  assign n15097 = n15096 ^ n4744 ^ 1'b0 ;
  assign n15101 = n15100 ^ n15097 ^ n6185 ;
  assign n15102 = n15101 ^ n11862 ^ n11711 ;
  assign n15103 = ( n3559 & n3976 ) | ( n3559 & ~n15102 ) | ( n3976 & ~n15102 ) ;
  assign n15110 = n15109 ^ n15106 ^ n15103 ;
  assign n15111 = n15110 ^ n2025 ^ x119 ;
  assign n15112 = n14611 ^ n3581 ^ 1'b0 ;
  assign n15113 = n6741 ^ n6277 ^ n6055 ;
  assign n15114 = n5946 | n15113 ;
  assign n15115 = n7036 & ~n15114 ;
  assign n15116 = n8503 & ~n13168 ;
  assign n15117 = ( n7993 & n15115 ) | ( n7993 & ~n15116 ) | ( n15115 & ~n15116 ) ;
  assign n15118 = n3607 ^ n2648 ^ 1'b0 ;
  assign n15119 = n296 & ~n15118 ;
  assign n15120 = n9839 ^ n6073 ^ x50 ;
  assign n15121 = n7344 ^ n4494 ^ n3142 ;
  assign n15122 = ( n13391 & n15120 ) | ( n13391 & n15121 ) | ( n15120 & n15121 ) ;
  assign n15123 = n10438 ^ n8932 ^ n2220 ;
  assign n15124 = n11965 ^ n10231 ^ n2633 ;
  assign n15125 = ( ~n2293 & n5533 ) | ( ~n2293 & n15124 ) | ( n5533 & n15124 ) ;
  assign n15126 = n15125 ^ n5600 ^ 1'b0 ;
  assign n15127 = n14609 ^ n11098 ^ n912 ;
  assign n15128 = n5451 ^ n4034 ^ n3569 ;
  assign n15129 = n15128 ^ n7329 ^ n4012 ;
  assign n15130 = ( n1903 & n10753 ) | ( n1903 & n11127 ) | ( n10753 & n11127 ) ;
  assign n15135 = n8129 ^ n1057 ^ 1'b0 ;
  assign n15136 = n12478 & n15135 ;
  assign n15132 = n2842 ^ n760 ^ n469 ;
  assign n15131 = n3374 & n4303 ;
  assign n15133 = n15132 ^ n15131 ^ 1'b0 ;
  assign n15134 = ( ~n7081 & n12932 ) | ( ~n7081 & n15133 ) | ( n12932 & n15133 ) ;
  assign n15137 = n15136 ^ n15134 ^ n231 ;
  assign n15138 = ( n7728 & n11800 ) | ( n7728 & n15137 ) | ( n11800 & n15137 ) ;
  assign n15139 = n14553 ^ n8479 ^ n6080 ;
  assign n15140 = n15139 ^ n8469 ^ n7938 ;
  assign n15141 = n15140 ^ n11712 ^ n4840 ;
  assign n15142 = ( ~n10191 & n11181 ) | ( ~n10191 & n15141 ) | ( n11181 & n15141 ) ;
  assign n15143 = ~n12187 & n12528 ;
  assign n15144 = n742 & n15143 ;
  assign n15145 = n15144 ^ n6325 ^ n5756 ;
  assign n15146 = ( n315 & ~n7186 ) | ( n315 & n10786 ) | ( ~n7186 & n10786 ) ;
  assign n15147 = n15146 ^ n9966 ^ n8882 ;
  assign n15148 = n5754 ^ n5386 ^ n2256 ;
  assign n15149 = n5062 ^ n1858 ^ n264 ;
  assign n15150 = ( n7561 & n15148 ) | ( n7561 & n15149 ) | ( n15148 & n15149 ) ;
  assign n15151 = ( n566 & n3656 ) | ( n566 & ~n7799 ) | ( n3656 & ~n7799 ) ;
  assign n15152 = ( n4769 & n9158 ) | ( n4769 & n13685 ) | ( n9158 & n13685 ) ;
  assign n15153 = ( ~n15150 & n15151 ) | ( ~n15150 & n15152 ) | ( n15151 & n15152 ) ;
  assign n15164 = n6895 ^ n2767 ^ n2236 ;
  assign n15165 = ( n6503 & n9552 ) | ( n6503 & ~n15164 ) | ( n9552 & ~n15164 ) ;
  assign n15154 = n14456 ^ n1669 ^ 1'b0 ;
  assign n15155 = ( n2847 & n6620 ) | ( n2847 & ~n13378 ) | ( n6620 & ~n13378 ) ;
  assign n15158 = n11813 ^ n4058 ^ 1'b0 ;
  assign n15156 = n7674 ^ n6562 ^ 1'b0 ;
  assign n15157 = n6800 & n15156 ;
  assign n15159 = n15158 ^ n15157 ^ n9636 ;
  assign n15160 = ( n11136 & ~n13946 ) | ( n11136 & n15159 ) | ( ~n13946 & n15159 ) ;
  assign n15161 = ( n15154 & ~n15155 ) | ( n15154 & n15160 ) | ( ~n15155 & n15160 ) ;
  assign n15162 = n15161 ^ n10900 ^ n761 ;
  assign n15163 = ( n4770 & n12963 ) | ( n4770 & ~n15162 ) | ( n12963 & ~n15162 ) ;
  assign n15166 = n15165 ^ n15163 ^ n11458 ;
  assign n15167 = ( ~n699 & n5425 ) | ( ~n699 & n8433 ) | ( n5425 & n8433 ) ;
  assign n15168 = n4884 ^ n2864 ^ n2372 ;
  assign n15169 = n15168 ^ n4174 ^ n2789 ;
  assign n15170 = n15169 ^ n11357 ^ n10157 ;
  assign n15171 = ( ~n8341 & n15167 ) | ( ~n8341 & n15170 ) | ( n15167 & n15170 ) ;
  assign n15172 = n7872 & n11422 ;
  assign n15173 = n8469 & n15172 ;
  assign n15174 = ( n570 & n1044 ) | ( n570 & n3776 ) | ( n1044 & n3776 ) ;
  assign n15175 = n15174 ^ n13649 ^ n7452 ;
  assign n15176 = n3896 | n15175 ;
  assign n15177 = n15176 ^ n3496 ^ 1'b0 ;
  assign n15178 = ( n2110 & ~n11249 ) | ( n2110 & n15177 ) | ( ~n11249 & n15177 ) ;
  assign n15179 = n15178 ^ n220 ^ 1'b0 ;
  assign n15180 = ~n6361 & n15179 ;
  assign n15181 = n1292 & n15180 ;
  assign n15182 = ( n1887 & n7697 ) | ( n1887 & ~n11785 ) | ( n7697 & ~n11785 ) ;
  assign n15183 = n8321 | n15182 ;
  assign n15184 = n2727 & ~n15183 ;
  assign n15185 = ( n2306 & n7773 ) | ( n2306 & ~n15184 ) | ( n7773 & ~n15184 ) ;
  assign n15186 = n10828 ^ n8455 ^ 1'b0 ;
  assign n15188 = n10328 ^ n9067 ^ n8695 ;
  assign n15187 = n13050 ^ n8495 ^ n7055 ;
  assign n15189 = n15188 ^ n15187 ^ 1'b0 ;
  assign n15190 = n8478 ^ n3313 ^ n2730 ;
  assign n15191 = n13054 ^ n2402 ^ 1'b0 ;
  assign n15192 = ( ~n2858 & n15190 ) | ( ~n2858 & n15191 ) | ( n15190 & n15191 ) ;
  assign n15193 = n13639 | n14768 ;
  assign n15194 = n15193 ^ n4803 ^ 1'b0 ;
  assign n15197 = ( n1045 & n2042 ) | ( n1045 & n3866 ) | ( n2042 & n3866 ) ;
  assign n15195 = n7264 ^ n1280 ^ n192 ;
  assign n15196 = n1866 & n15195 ;
  assign n15198 = n15197 ^ n15196 ^ 1'b0 ;
  assign n15199 = n9476 ^ n4465 ^ n3246 ;
  assign n15200 = ( n3330 & ~n8719 ) | ( n3330 & n15199 ) | ( ~n8719 & n15199 ) ;
  assign n15201 = n4234 ^ n4008 ^ n465 ;
  assign n15202 = ~n6151 & n15201 ;
  assign n15203 = n8128 ^ n4926 ^ 1'b0 ;
  assign n15204 = n10307 & ~n15203 ;
  assign n15205 = n14382 ^ n7241 ^ n6867 ;
  assign n15206 = n15205 ^ x13 ^ 1'b0 ;
  assign n15207 = ( ~n2876 & n14834 ) | ( ~n2876 & n15206 ) | ( n14834 & n15206 ) ;
  assign n15208 = n4599 ^ n4096 ^ 1'b0 ;
  assign n15209 = n15208 ^ n4641 ^ n3179 ;
  assign n15210 = n5593 ^ n2211 ^ 1'b0 ;
  assign n15211 = n9732 ^ n3953 ^ n3639 ;
  assign n15212 = n14490 ^ n1615 ^ n926 ;
  assign n15218 = n7979 ^ n2016 ^ 1'b0 ;
  assign n15219 = n15218 ^ n6194 ^ 1'b0 ;
  assign n15213 = ( n1940 & ~n2754 ) | ( n1940 & n10488 ) | ( ~n2754 & n10488 ) ;
  assign n15214 = n10404 ^ n1971 ^ n1386 ;
  assign n15215 = n15214 ^ n1729 ^ 1'b0 ;
  assign n15216 = n15213 | n15215 ;
  assign n15217 = n15216 ^ n8144 ^ n1539 ;
  assign n15220 = n15219 ^ n15217 ^ n11733 ;
  assign n15221 = n7873 ^ n1360 ^ 1'b0 ;
  assign n15222 = n15221 ^ n13464 ^ n8721 ;
  assign n15226 = n8412 & ~n13299 ;
  assign n15223 = ( n1842 & ~n2678 ) | ( n1842 & n4720 ) | ( ~n2678 & n4720 ) ;
  assign n15224 = ( ~n2877 & n7226 ) | ( ~n2877 & n8793 ) | ( n7226 & n8793 ) ;
  assign n15225 = n15223 & ~n15224 ;
  assign n15227 = n15226 ^ n15225 ^ n6412 ;
  assign n15228 = n5912 & ~n15107 ;
  assign n15229 = n2237 & ~n9861 ;
  assign n15230 = n15229 ^ n1490 ^ x112 ;
  assign n15231 = ( n4104 & ~n5033 ) | ( n4104 & n15230 ) | ( ~n5033 & n15230 ) ;
  assign n15232 = ( n9722 & n15228 ) | ( n9722 & ~n15231 ) | ( n15228 & ~n15231 ) ;
  assign n15233 = n3586 ^ n2988 ^ n799 ;
  assign n15234 = n4389 ^ n175 ^ 1'b0 ;
  assign n15235 = ( n14914 & n15233 ) | ( n14914 & n15234 ) | ( n15233 & n15234 ) ;
  assign n15236 = n15235 ^ n6824 ^ n4053 ;
  assign n15237 = ( n6099 & n6509 ) | ( n6099 & n7685 ) | ( n6509 & n7685 ) ;
  assign n15238 = n9861 | n14324 ;
  assign n15239 = n13028 ^ n4020 ^ 1'b0 ;
  assign n15240 = n7340 & n15239 ;
  assign n15241 = n15240 ^ n7904 ^ n653 ;
  assign n15242 = ( ~n3519 & n4392 ) | ( ~n3519 & n7957 ) | ( n4392 & n7957 ) ;
  assign n15243 = ( n4732 & n7258 ) | ( n4732 & ~n12372 ) | ( n7258 & ~n12372 ) ;
  assign n15244 = ( n10354 & n15242 ) | ( n10354 & ~n15243 ) | ( n15242 & ~n15243 ) ;
  assign n15245 = n5773 & n11441 ;
  assign n15246 = n15245 ^ n11834 ^ 1'b0 ;
  assign n15247 = ( ~n2774 & n3269 ) | ( ~n2774 & n5508 ) | ( n3269 & n5508 ) ;
  assign n15248 = n15247 ^ n440 ^ 1'b0 ;
  assign n15249 = n12083 & n15248 ;
  assign n15250 = ( n3640 & n4886 ) | ( n3640 & ~n9715 ) | ( n4886 & ~n9715 ) ;
  assign n15251 = n15250 ^ n12224 ^ n4373 ;
  assign n15252 = ( n2024 & n7315 ) | ( n2024 & ~n15251 ) | ( n7315 & ~n15251 ) ;
  assign n15253 = ( n4362 & n5943 ) | ( n4362 & n9911 ) | ( n5943 & n9911 ) ;
  assign n15254 = n15253 ^ n9051 ^ n4999 ;
  assign n15255 = n15254 ^ n11397 ^ n6499 ;
  assign n15257 = n9253 & n9414 ;
  assign n15258 = n15257 ^ n3580 ^ n2262 ;
  assign n15256 = n4676 & ~n6872 ;
  assign n15259 = n15258 ^ n15256 ^ 1'b0 ;
  assign n15269 = ( ~n1078 & n1728 ) | ( ~n1078 & n5526 ) | ( n1728 & n5526 ) ;
  assign n15265 = n4092 ^ n3138 ^ n2157 ;
  assign n15264 = ( n2132 & ~n2698 ) | ( n2132 & n3863 ) | ( ~n2698 & n3863 ) ;
  assign n15266 = n15265 ^ n15264 ^ n392 ;
  assign n15267 = n15266 ^ n2913 ^ 1'b0 ;
  assign n15268 = n7017 & n15267 ;
  assign n15260 = n2767 & n5627 ;
  assign n15261 = n11619 & n15260 ;
  assign n15262 = n15261 ^ n6413 ^ n2577 ;
  assign n15263 = ~n12048 & n15262 ;
  assign n15270 = n15269 ^ n15268 ^ n15263 ;
  assign n15271 = n7639 ^ n335 ^ 1'b0 ;
  assign n15272 = n753 & n15271 ;
  assign n15273 = n15272 ^ n2569 ^ n1979 ;
  assign n15276 = n2108 & ~n4756 ;
  assign n15277 = n15276 ^ n7351 ^ n379 ;
  assign n15278 = ( n2450 & n3030 ) | ( n2450 & n15277 ) | ( n3030 & n15277 ) ;
  assign n15274 = ( n6124 & ~n7515 ) | ( n6124 & n13400 ) | ( ~n7515 & n13400 ) ;
  assign n15275 = n15274 ^ n595 ^ 1'b0 ;
  assign n15279 = n15278 ^ n15275 ^ n2861 ;
  assign n15280 = ( ~n7566 & n8604 ) | ( ~n7566 & n12257 ) | ( n8604 & n12257 ) ;
  assign n15281 = n3172 ^ n2982 ^ n407 ;
  assign n15282 = n15281 ^ n7619 ^ n2681 ;
  assign n15283 = n8276 & ~n10925 ;
  assign n15284 = n6435 & n15283 ;
  assign n15285 = ~n5934 & n8158 ;
  assign n15286 = n15285 ^ n7201 ^ 1'b0 ;
  assign n15287 = n15286 ^ n3553 ^ n2871 ;
  assign n15288 = n8891 ^ n8027 ^ n4362 ;
  assign n15289 = ~n226 & n1862 ;
  assign n15290 = ( ~n1632 & n14087 ) | ( ~n1632 & n15289 ) | ( n14087 & n15289 ) ;
  assign n15293 = n4371 & ~n9707 ;
  assign n15294 = n15293 ^ n2235 ^ n1318 ;
  assign n15291 = n4471 & n5514 ;
  assign n15292 = n15291 ^ n13326 ^ 1'b0 ;
  assign n15295 = n15294 ^ n15292 ^ n5311 ;
  assign n15296 = ( n4154 & ~n15290 ) | ( n4154 & n15295 ) | ( ~n15290 & n15295 ) ;
  assign n15297 = n12683 ^ n5234 ^ n2039 ;
  assign n15299 = n2421 & n11651 ;
  assign n15298 = n11376 ^ n5113 ^ 1'b0 ;
  assign n15300 = n15299 ^ n15298 ^ n2559 ;
  assign n15301 = ( n2429 & n2484 ) | ( n2429 & n3251 ) | ( n2484 & n3251 ) ;
  assign n15302 = ( ~n3996 & n4153 ) | ( ~n3996 & n15301 ) | ( n4153 & n15301 ) ;
  assign n15303 = n15302 ^ n7478 ^ n4155 ;
  assign n15304 = n15303 ^ n10368 ^ n9744 ;
  assign n15305 = n5630 ^ n4205 ^ 1'b0 ;
  assign n15306 = n12760 & ~n15305 ;
  assign n15307 = n15306 ^ n3825 ^ 1'b0 ;
  assign n15308 = n13685 ^ n2750 ^ 1'b0 ;
  assign n15309 = ( n6745 & ~n8652 ) | ( n6745 & n12453 ) | ( ~n8652 & n12453 ) ;
  assign n15310 = n6211 ^ n4115 ^ n517 ;
  assign n15311 = n14691 | n15310 ;
  assign n15312 = n15311 ^ n13212 ^ n9616 ;
  assign n15313 = n15312 ^ n2873 ^ 1'b0 ;
  assign n15314 = ( ~n4080 & n11990 ) | ( ~n4080 & n15177 ) | ( n11990 & n15177 ) ;
  assign n15315 = ( n12449 & ~n14353 ) | ( n12449 & n15314 ) | ( ~n14353 & n15314 ) ;
  assign n15316 = n4127 ^ n3342 ^ n2398 ;
  assign n15317 = n15316 ^ n12781 ^ 1'b0 ;
  assign n15318 = n15317 ^ n2307 ^ 1'b0 ;
  assign n15319 = n6926 ^ n5579 ^ 1'b0 ;
  assign n15320 = n15319 ^ n3603 ^ n1079 ;
  assign n15321 = n15320 ^ n14729 ^ 1'b0 ;
  assign n15326 = n3039 ^ n379 ^ 1'b0 ;
  assign n15322 = n375 & ~n6173 ;
  assign n15323 = n11230 & ~n15322 ;
  assign n15324 = n15323 ^ n5710 ^ 1'b0 ;
  assign n15325 = n9809 & ~n15324 ;
  assign n15327 = n15326 ^ n15325 ^ 1'b0 ;
  assign n15328 = ( ~x97 & n8965 ) | ( ~x97 & n9660 ) | ( n8965 & n9660 ) ;
  assign n15329 = n7689 & ~n15328 ;
  assign n15330 = n3779 ^ n1664 ^ 1'b0 ;
  assign n15331 = n5982 & ~n15330 ;
  assign n15333 = n5983 ^ n1870 ^ 1'b0 ;
  assign n15334 = ~n7314 & n15333 ;
  assign n15332 = ( ~n3574 & n3855 ) | ( ~n3574 & n6679 ) | ( n3855 & n6679 ) ;
  assign n15335 = n15334 ^ n15332 ^ n11006 ;
  assign n15336 = n8719 ^ n3253 ^ 1'b0 ;
  assign n15340 = ( n822 & ~n1957 ) | ( n822 & n10108 ) | ( ~n1957 & n10108 ) ;
  assign n15341 = n10537 | n15340 ;
  assign n15337 = n9367 ^ n8329 ^ n229 ;
  assign n15338 = n6271 ^ n5266 ^ 1'b0 ;
  assign n15339 = n15337 & n15338 ;
  assign n15342 = n15341 ^ n15339 ^ 1'b0 ;
  assign n15343 = n2424 & n15214 ;
  assign n15344 = ( n6104 & n9476 ) | ( n6104 & ~n10150 ) | ( n9476 & ~n10150 ) ;
  assign n15345 = n13236 ^ n857 ^ 1'b0 ;
  assign n15346 = n11103 & n15345 ;
  assign n15347 = n1381 | n3727 ;
  assign n15348 = n2182 | n15347 ;
  assign n15349 = n672 | n3009 ;
  assign n15350 = n15349 ^ n8471 ^ 1'b0 ;
  assign n15351 = n12030 & n15350 ;
  assign n15352 = n15351 ^ n11304 ^ n4714 ;
  assign n15353 = ( ~n7467 & n15348 ) | ( ~n7467 & n15352 ) | ( n15348 & n15352 ) ;
  assign n15361 = n9664 ^ n3038 ^ n2973 ;
  assign n15354 = n6600 ^ n6214 ^ n1100 ;
  assign n15355 = n5670 ^ n4203 ^ n3862 ;
  assign n15356 = ( ~n4034 & n15354 ) | ( ~n4034 & n15355 ) | ( n15354 & n15355 ) ;
  assign n15357 = n8751 | n15356 ;
  assign n15358 = n15357 ^ n10189 ^ 1'b0 ;
  assign n15359 = n15358 ^ n12521 ^ 1'b0 ;
  assign n15360 = n3801 | n15359 ;
  assign n15362 = n15361 ^ n15360 ^ 1'b0 ;
  assign n15366 = n6824 ^ n3317 ^ n1906 ;
  assign n15363 = n4929 ^ n4732 ^ n1995 ;
  assign n15364 = n15363 ^ n7993 ^ n1271 ;
  assign n15365 = n15364 ^ n14236 ^ n6703 ;
  assign n15367 = n15366 ^ n15365 ^ n11928 ;
  assign n15368 = x72 & ~n461 ;
  assign n15369 = ~n4683 & n15368 ;
  assign n15370 = n15369 ^ n8439 ^ 1'b0 ;
  assign n15371 = ~n4121 & n15370 ;
  assign n15372 = ( ~n362 & n9445 ) | ( ~n362 & n15371 ) | ( n9445 & n15371 ) ;
  assign n15373 = n6315 | n11317 ;
  assign n15374 = n1709 | n15373 ;
  assign n15375 = n3888 ^ n2804 ^ n954 ;
  assign n15376 = n7930 & ~n12723 ;
  assign n15377 = ( n1188 & n10514 ) | ( n1188 & ~n11504 ) | ( n10514 & ~n11504 ) ;
  assign n15378 = ( n2643 & n4396 ) | ( n2643 & ~n15377 ) | ( n4396 & ~n15377 ) ;
  assign n15379 = ( n2239 & n4046 ) | ( n2239 & n4447 ) | ( n4046 & n4447 ) ;
  assign n15380 = n15379 ^ n5005 ^ n3278 ;
  assign n15381 = n15380 ^ n7804 ^ n374 ;
  assign n15382 = n5526 | n15381 ;
  assign n15384 = ~n1818 & n4163 ;
  assign n15385 = n15384 ^ n6615 ^ 1'b0 ;
  assign n15383 = n404 & ~n5052 ;
  assign n15386 = n15385 ^ n15383 ^ 1'b0 ;
  assign n15387 = n15386 ^ n5964 ^ n4554 ;
  assign n15388 = n2965 ^ n2310 ^ 1'b0 ;
  assign n15389 = n9020 & n15388 ;
  assign n15390 = n10419 ^ n6743 ^ n3779 ;
  assign n15391 = ( n4295 & n9449 ) | ( n4295 & ~n15390 ) | ( n9449 & ~n15390 ) ;
  assign n15392 = ( n5578 & ~n11701 ) | ( n5578 & n15391 ) | ( ~n11701 & n15391 ) ;
  assign n15393 = ( n8922 & n15389 ) | ( n8922 & n15392 ) | ( n15389 & n15392 ) ;
  assign n15394 = n15393 ^ n2733 ^ n1036 ;
  assign n15395 = n8883 ^ n7610 ^ n1291 ;
  assign n15396 = n9108 & n15395 ;
  assign n15397 = n15396 ^ n6403 ^ 1'b0 ;
  assign n15403 = n6550 ^ n3094 ^ n1247 ;
  assign n15400 = n9451 ^ n1342 ^ 1'b0 ;
  assign n15401 = n8518 & ~n15400 ;
  assign n15402 = n15401 ^ n233 ^ 1'b0 ;
  assign n15398 = n9044 ^ n4196 ^ n3485 ;
  assign n15399 = n8938 | n15398 ;
  assign n15404 = n15403 ^ n15402 ^ n15399 ;
  assign n15405 = ( n4156 & n4998 ) | ( n4156 & n6119 ) | ( n4998 & n6119 ) ;
  assign n15406 = n15405 ^ n4266 ^ n3229 ;
  assign n15407 = n15406 ^ n8672 ^ 1'b0 ;
  assign n15408 = n12992 ^ n5753 ^ n4199 ;
  assign n15409 = ( ~n11254 & n15407 ) | ( ~n11254 & n15408 ) | ( n15407 & n15408 ) ;
  assign n15410 = n15409 ^ n10325 ^ n6308 ;
  assign n15411 = n1863 & n2944 ;
  assign n15412 = ( ~n6651 & n9584 ) | ( ~n6651 & n10035 ) | ( n9584 & n10035 ) ;
  assign n15413 = n15412 ^ n14217 ^ n7756 ;
  assign n15415 = ~n4432 & n11829 ;
  assign n15414 = n11780 ^ n9110 ^ n7111 ;
  assign n15416 = n15415 ^ n15414 ^ n10385 ;
  assign n15417 = ( n2389 & n5295 ) | ( n2389 & ~n8006 ) | ( n5295 & ~n8006 ) ;
  assign n15418 = n4511 & n15417 ;
  assign n15419 = ~n9197 & n13918 ;
  assign n15420 = n9560 ^ n4717 ^ n1578 ;
  assign n15421 = n15420 ^ n4370 ^ n4273 ;
  assign n15422 = n3831 | n8508 ;
  assign n15423 = n7865 & ~n15422 ;
  assign n15424 = ( n11627 & ~n12859 ) | ( n11627 & n15423 ) | ( ~n12859 & n15423 ) ;
  assign n15425 = n5640 ^ n1874 ^ n582 ;
  assign n15426 = ( n2123 & n9378 ) | ( n2123 & ~n15425 ) | ( n9378 & ~n15425 ) ;
  assign n15427 = ( x24 & n1655 ) | ( x24 & ~n2557 ) | ( n1655 & ~n2557 ) ;
  assign n15428 = ( n2297 & n7071 ) | ( n2297 & n15427 ) | ( n7071 & n15427 ) ;
  assign n15429 = n5586 ^ n3867 ^ 1'b0 ;
  assign n15430 = n15429 ^ n4302 ^ 1'b0 ;
  assign n15431 = n15428 & ~n15430 ;
  assign n15432 = n14634 ^ n12505 ^ 1'b0 ;
  assign n15433 = n12121 & n13649 ;
  assign n15434 = ~n1227 & n2606 ;
  assign n15435 = n10683 & n15434 ;
  assign n15436 = n14414 ^ n5616 ^ n409 ;
  assign n15437 = ( n15433 & n15435 ) | ( n15433 & n15436 ) | ( n15435 & n15436 ) ;
  assign n15438 = n9122 ^ n4540 ^ n4376 ;
  assign n15439 = n4528 ^ n815 ^ 1'b0 ;
  assign n15440 = n1466 | n15439 ;
  assign n15441 = n15440 ^ n5974 ^ n1868 ;
  assign n15442 = ( ~n8504 & n11255 ) | ( ~n8504 & n15441 ) | ( n11255 & n15441 ) ;
  assign n15444 = n1712 | n5039 ;
  assign n15445 = ( ~n1108 & n8414 ) | ( ~n1108 & n15444 ) | ( n8414 & n15444 ) ;
  assign n15443 = n6356 ^ n2856 ^ 1'b0 ;
  assign n15446 = n15445 ^ n15443 ^ n4240 ;
  assign n15458 = ( n841 & n1089 ) | ( n841 & ~n12366 ) | ( n1089 & ~n12366 ) ;
  assign n15456 = n8785 ^ n8620 ^ 1'b0 ;
  assign n15457 = n2548 & n15456 ;
  assign n15459 = n15458 ^ n15457 ^ 1'b0 ;
  assign n15448 = n6530 ^ n5747 ^ n5194 ;
  assign n15447 = n10324 ^ n7581 ^ n553 ;
  assign n15449 = n15448 ^ n15447 ^ n10622 ;
  assign n15450 = n2065 & n6551 ;
  assign n15451 = n2038 & ~n2174 ;
  assign n15452 = ( n737 & n12126 ) | ( n737 & n15451 ) | ( n12126 & n15451 ) ;
  assign n15453 = n15450 & n15452 ;
  assign n15454 = ~n865 & n15453 ;
  assign n15455 = n15449 | n15454 ;
  assign n15460 = n15459 ^ n15455 ^ n6824 ;
  assign n15461 = n7400 ^ n6732 ^ n1499 ;
  assign n15462 = ~n2028 & n7894 ;
  assign n15463 = n15462 ^ n3750 ^ 1'b0 ;
  assign n15464 = ( n2358 & n12427 ) | ( n2358 & ~n15463 ) | ( n12427 & ~n15463 ) ;
  assign n15465 = n9183 ^ n3700 ^ n1482 ;
  assign n15466 = ( n6138 & n15464 ) | ( n6138 & n15465 ) | ( n15464 & n15465 ) ;
  assign n15469 = n4784 ^ n4479 ^ 1'b0 ;
  assign n15467 = ( n2555 & ~n5017 ) | ( n2555 & n8474 ) | ( ~n5017 & n8474 ) ;
  assign n15468 = ( n3396 & ~n5484 ) | ( n3396 & n15467 ) | ( ~n5484 & n15467 ) ;
  assign n15470 = n15469 ^ n15468 ^ n4063 ;
  assign n15471 = n7575 ^ n3967 ^ 1'b0 ;
  assign n15475 = ~n4836 & n10830 ;
  assign n15476 = n7984 & n15475 ;
  assign n15472 = n5107 & n9871 ;
  assign n15473 = n8568 ^ n3359 ^ 1'b0 ;
  assign n15474 = ( n7103 & n15472 ) | ( n7103 & ~n15473 ) | ( n15472 & ~n15473 ) ;
  assign n15477 = n15476 ^ n15474 ^ n8130 ;
  assign n15478 = ~n1828 & n11749 ;
  assign n15479 = n11157 ^ n2869 ^ 1'b0 ;
  assign n15480 = ( n7536 & ~n15478 ) | ( n7536 & n15479 ) | ( ~n15478 & n15479 ) ;
  assign n15487 = n8461 & n12377 ;
  assign n15488 = ( n1267 & n7908 ) | ( n1267 & ~n8429 ) | ( n7908 & ~n8429 ) ;
  assign n15489 = ~n15487 & n15488 ;
  assign n15485 = ( n3678 & n7837 ) | ( n3678 & n13415 ) | ( n7837 & n13415 ) ;
  assign n15486 = ( n11182 & n11927 ) | ( n11182 & n15485 ) | ( n11927 & n15485 ) ;
  assign n15483 = n4999 ^ n4637 ^ n4099 ;
  assign n15481 = n4920 ^ n4118 ^ n1147 ;
  assign n15482 = n1257 & ~n15481 ;
  assign n15484 = n15483 ^ n15482 ^ 1'b0 ;
  assign n15490 = n15489 ^ n15486 ^ n15484 ;
  assign n15491 = n14358 | n15123 ;
  assign n15492 = n15491 ^ x34 ^ 1'b0 ;
  assign n15493 = ~n3121 & n9612 ;
  assign n15494 = ( ~n1167 & n2402 ) | ( ~n1167 & n5192 ) | ( n2402 & n5192 ) ;
  assign n15495 = ( ~n6802 & n7403 ) | ( ~n6802 & n10733 ) | ( n7403 & n10733 ) ;
  assign n15496 = ( ~n1797 & n6590 ) | ( ~n1797 & n15380 ) | ( n6590 & n15380 ) ;
  assign n15497 = ( n12093 & n15495 ) | ( n12093 & ~n15496 ) | ( n15495 & ~n15496 ) ;
  assign n15498 = ( n155 & n5333 ) | ( n155 & n8996 ) | ( n5333 & n8996 ) ;
  assign n15499 = ~n12396 & n15498 ;
  assign n15500 = n15499 ^ n3425 ^ 1'b0 ;
  assign n15501 = n2585 | n12767 ;
  assign n15502 = n15501 ^ n14335 ^ 1'b0 ;
  assign n15503 = n15502 ^ n12869 ^ n4564 ;
  assign n15504 = n14965 & ~n15503 ;
  assign n15505 = n15504 ^ n5022 ^ 1'b0 ;
  assign n15510 = ~n9292 & n11396 ;
  assign n15511 = ~n5186 & n15510 ;
  assign n15509 = ~n1349 & n4175 ;
  assign n15512 = n15511 ^ n15509 ^ 1'b0 ;
  assign n15513 = n2926 & n8344 ;
  assign n15514 = ( ~x116 & n15512 ) | ( ~x116 & n15513 ) | ( n15512 & n15513 ) ;
  assign n15506 = n6708 & n11648 ;
  assign n15507 = n3318 & n15506 ;
  assign n15508 = ( n4542 & n5849 ) | ( n4542 & ~n15507 ) | ( n5849 & ~n15507 ) ;
  assign n15515 = n15514 ^ n15508 ^ n7501 ;
  assign n15516 = n7040 ^ n2934 ^ n1488 ;
  assign n15517 = ( n1200 & n3683 ) | ( n1200 & n4587 ) | ( n3683 & n4587 ) ;
  assign n15518 = n1356 | n8689 ;
  assign n15519 = n15517 & ~n15518 ;
  assign n15520 = ( n15063 & n15516 ) | ( n15063 & n15519 ) | ( n15516 & n15519 ) ;
  assign n15521 = n398 | n480 ;
  assign n15522 = ( n3308 & ~n4444 ) | ( n3308 & n15521 ) | ( ~n4444 & n15521 ) ;
  assign n15527 = n10160 ^ n5855 ^ n1469 ;
  assign n15523 = n5306 ^ n4962 ^ n2040 ;
  assign n15524 = n15523 ^ n3276 ^ n3258 ;
  assign n15525 = n5572 ^ n425 ^ 1'b0 ;
  assign n15526 = ( n2654 & n15524 ) | ( n2654 & n15525 ) | ( n15524 & n15525 ) ;
  assign n15528 = n15527 ^ n15526 ^ n3488 ;
  assign n15529 = n15528 ^ n14747 ^ n5479 ;
  assign n15530 = n15529 ^ n5020 ^ n3950 ;
  assign n15531 = n9975 ^ n8751 ^ x113 ;
  assign n15532 = ( n3047 & n3592 ) | ( n3047 & n8762 ) | ( n3592 & n8762 ) ;
  assign n15533 = n9662 ^ n2624 ^ n233 ;
  assign n15534 = n15533 ^ n6581 ^ 1'b0 ;
  assign n15535 = ~n6757 & n15534 ;
  assign n15536 = ( ~n6641 & n15532 ) | ( ~n6641 & n15535 ) | ( n15532 & n15535 ) ;
  assign n15537 = ( ~n7788 & n10217 ) | ( ~n7788 & n15536 ) | ( n10217 & n15536 ) ;
  assign n15538 = ~n3453 & n11510 ;
  assign n15539 = ( n15531 & ~n15537 ) | ( n15531 & n15538 ) | ( ~n15537 & n15538 ) ;
  assign n15540 = ( n3345 & n5729 ) | ( n3345 & ~n10711 ) | ( n5729 & ~n10711 ) ;
  assign n15541 = n5983 ^ n3505 ^ n2049 ;
  assign n15542 = n7370 ^ n7076 ^ 1'b0 ;
  assign n15543 = ( ~n1242 & n1984 ) | ( ~n1242 & n5708 ) | ( n1984 & n5708 ) ;
  assign n15544 = n15543 ^ n11809 ^ n8568 ;
  assign n15545 = n2879 ^ n1903 ^ n390 ;
  assign n15546 = n15545 ^ n11853 ^ 1'b0 ;
  assign n15547 = ~n3368 & n15546 ;
  assign n15548 = n2697 & n15547 ;
  assign n15549 = ( ~n1253 & n4154 ) | ( ~n1253 & n10143 ) | ( n4154 & n10143 ) ;
  assign n15550 = ~n14679 & n15549 ;
  assign n15551 = ~n10237 & n15550 ;
  assign n15552 = ( n2392 & n4895 ) | ( n2392 & ~n9983 ) | ( n4895 & ~n9983 ) ;
  assign n15553 = n13673 ^ n10908 ^ n8898 ;
  assign n15554 = n15553 ^ n13168 ^ n6356 ;
  assign n15555 = n13185 ^ n7253 ^ n6553 ;
  assign n15556 = ( ~n780 & n5528 ) | ( ~n780 & n7317 ) | ( n5528 & n7317 ) ;
  assign n15557 = n8534 & n13275 ;
  assign n15558 = ~n14163 & n15557 ;
  assign n15559 = n4466 ^ n3700 ^ n3385 ;
  assign n15562 = ( n3677 & n7206 ) | ( n3677 & n11554 ) | ( n7206 & n11554 ) ;
  assign n15560 = n450 ^ n186 ^ 1'b0 ;
  assign n15561 = n8827 & n15560 ;
  assign n15563 = n15562 ^ n15561 ^ 1'b0 ;
  assign n15564 = n15559 & ~n15563 ;
  assign n15565 = n10691 ^ n2695 ^ 1'b0 ;
  assign n15566 = n9438 | n15565 ;
  assign n15567 = n15566 ^ n5276 ^ n4264 ;
  assign n15568 = n8613 ^ n2583 ^ n1028 ;
  assign n15570 = n2051 | n8556 ;
  assign n15571 = n1314 & ~n15570 ;
  assign n15569 = n6677 ^ n6268 ^ 1'b0 ;
  assign n15572 = n15571 ^ n15569 ^ n5118 ;
  assign n15573 = ( n11404 & n15568 ) | ( n11404 & ~n15572 ) | ( n15568 & ~n15572 ) ;
  assign n15574 = n1674 | n3742 ;
  assign n15575 = ( ~n147 & n2624 ) | ( ~n147 & n2754 ) | ( n2624 & n2754 ) ;
  assign n15576 = ( n8199 & n8671 ) | ( n8199 & ~n15575 ) | ( n8671 & ~n15575 ) ;
  assign n15577 = ( ~n1632 & n15574 ) | ( ~n1632 & n15576 ) | ( n15574 & n15576 ) ;
  assign n15578 = n11232 ^ n6340 ^ x64 ;
  assign n15582 = n944 ^ n341 ^ 1'b0 ;
  assign n15579 = n1386 | n4131 ;
  assign n15580 = n15579 ^ n9092 ^ 1'b0 ;
  assign n15581 = ~n1230 & n15580 ;
  assign n15583 = n15582 ^ n15581 ^ n11438 ;
  assign n15584 = n15578 & ~n15583 ;
  assign n15585 = n15433 & n15584 ;
  assign n15586 = n15036 ^ n14326 ^ n4829 ;
  assign n15587 = n6197 ^ n4494 ^ x88 ;
  assign n15588 = ( n6071 & ~n13150 ) | ( n6071 & n15587 ) | ( ~n13150 & n15587 ) ;
  assign n15589 = n8364 ^ n5578 ^ n3610 ;
  assign n15590 = ( n3734 & n12114 ) | ( n3734 & ~n15589 ) | ( n12114 & ~n15589 ) ;
  assign n15591 = n15590 ^ n3012 ^ 1'b0 ;
  assign n15592 = ( n3498 & ~n5375 ) | ( n3498 & n10701 ) | ( ~n5375 & n10701 ) ;
  assign n15593 = n15592 ^ n11409 ^ n712 ;
  assign n15594 = n14760 & n15593 ;
  assign n15595 = ~n4879 & n15594 ;
  assign n15596 = ( ~n2452 & n2859 ) | ( ~n2452 & n12781 ) | ( n2859 & n12781 ) ;
  assign n15597 = ~n9198 & n13570 ;
  assign n15598 = n4858 & n15597 ;
  assign n15599 = n14743 ^ n13634 ^ n4905 ;
  assign n15600 = n15599 ^ n10046 ^ n8696 ;
  assign n15601 = ( n376 & n4038 ) | ( n376 & n15600 ) | ( n4038 & n15600 ) ;
  assign n15602 = n3526 & ~n11618 ;
  assign n15603 = n15602 ^ n548 ^ 1'b0 ;
  assign n15604 = n15603 ^ n15428 ^ n8211 ;
  assign n15605 = ( n4193 & n7364 ) | ( n4193 & ~n15604 ) | ( n7364 & ~n15604 ) ;
  assign n15606 = n12824 ^ n8217 ^ 1'b0 ;
  assign n15607 = ( n3579 & n13790 ) | ( n3579 & n15606 ) | ( n13790 & n15606 ) ;
  assign n15608 = ( ~n2699 & n7563 ) | ( ~n2699 & n12852 ) | ( n7563 & n12852 ) ;
  assign n15609 = n1965 & n3164 ;
  assign n15610 = n235 | n15609 ;
  assign n15611 = n15610 ^ n11855 ^ 1'b0 ;
  assign n15619 = ( n758 & ~n3335 ) | ( n758 & n6094 ) | ( ~n3335 & n6094 ) ;
  assign n15620 = n11627 | n15619 ;
  assign n15615 = n5579 ^ n2411 ^ n2356 ;
  assign n15616 = n15615 ^ n14187 ^ n10479 ;
  assign n15617 = n15616 ^ n8316 ^ n6930 ;
  assign n15613 = n12850 ^ n11677 ^ 1'b0 ;
  assign n15612 = ( n8699 & n9545 ) | ( n8699 & n9989 ) | ( n9545 & n9989 ) ;
  assign n15614 = n15613 ^ n15612 ^ n12305 ;
  assign n15618 = n15617 ^ n15614 ^ n5578 ;
  assign n15621 = n15620 ^ n15618 ^ n14938 ;
  assign n15622 = n10883 ^ n7582 ^ n6921 ;
  assign n15623 = ( n10740 & ~n13405 ) | ( n10740 & n15622 ) | ( ~n13405 & n15622 ) ;
  assign n15624 = ( ~n5185 & n7471 ) | ( ~n5185 & n14475 ) | ( n7471 & n14475 ) ;
  assign n15625 = n11152 | n11879 ;
  assign n15626 = n15625 ^ n7392 ^ 1'b0 ;
  assign n15627 = ~n4926 & n15626 ;
  assign n15628 = n11557 ^ n4384 ^ n575 ;
  assign n15629 = n1399 | n11200 ;
  assign n15630 = ( n2371 & ~n15340 ) | ( n2371 & n15629 ) | ( ~n15340 & n15629 ) ;
  assign n15631 = ~n4363 & n9885 ;
  assign n15632 = n10572 ^ n8140 ^ 1'b0 ;
  assign n15633 = ~n327 & n616 ;
  assign n15634 = n3584 & n15633 ;
  assign n15635 = n15634 ^ n5162 ^ n2938 ;
  assign n15636 = n6769 & n7586 ;
  assign n15637 = n15636 ^ n6423 ^ 1'b0 ;
  assign n15638 = ~n7251 & n15637 ;
  assign n15639 = n15638 ^ n5572 ^ 1'b0 ;
  assign n15640 = ( n3305 & n15635 ) | ( n3305 & ~n15639 ) | ( n15635 & ~n15639 ) ;
  assign n15641 = ( ~n3269 & n5293 ) | ( ~n3269 & n8319 ) | ( n5293 & n8319 ) ;
  assign n15642 = n4732 & n12068 ;
  assign n15643 = ~n8729 & n15642 ;
  assign n15644 = ( ~n1091 & n11016 ) | ( ~n1091 & n15643 ) | ( n11016 & n15643 ) ;
  assign n15645 = ( ~n12181 & n12434 ) | ( ~n12181 & n15644 ) | ( n12434 & n15644 ) ;
  assign n15646 = n13162 ^ n2458 ^ n1911 ;
  assign n15647 = n15646 ^ n9169 ^ 1'b0 ;
  assign n15648 = ( ~n1515 & n1946 ) | ( ~n1515 & n15647 ) | ( n1946 & n15647 ) ;
  assign n15649 = n15648 ^ n11891 ^ 1'b0 ;
  assign n15650 = n8341 & ~n15649 ;
  assign n15651 = n11573 ^ n6367 ^ n896 ;
  assign n15652 = n15651 ^ n11021 ^ n2297 ;
  assign n15653 = ( n10140 & n14097 ) | ( n10140 & n15652 ) | ( n14097 & n15652 ) ;
  assign n15654 = n7320 ^ n4259 ^ n2305 ;
  assign n15655 = ~n9652 & n11807 ;
  assign n15656 = n15655 ^ n4217 ^ 1'b0 ;
  assign n15657 = ( n12698 & n15654 ) | ( n12698 & n15656 ) | ( n15654 & n15656 ) ;
  assign n15658 = n15657 ^ n14721 ^ n1949 ;
  assign n15659 = n14814 ^ n9939 ^ n6896 ;
  assign n15660 = ( n1904 & ~n5753 ) | ( n1904 & n10143 ) | ( ~n5753 & n10143 ) ;
  assign n15661 = n15660 ^ n13857 ^ n13258 ;
  assign n15662 = ( n11952 & ~n15659 ) | ( n11952 & n15661 ) | ( ~n15659 & n15661 ) ;
  assign n15663 = n12553 ^ n12159 ^ 1'b0 ;
  assign n15666 = n1645 & ~n7842 ;
  assign n15667 = n15666 ^ n14125 ^ 1'b0 ;
  assign n15668 = n15667 ^ n13031 ^ 1'b0 ;
  assign n15664 = ( n7383 & ~n12151 ) | ( n7383 & n12355 ) | ( ~n12151 & n12355 ) ;
  assign n15665 = n15664 ^ n3025 ^ n1918 ;
  assign n15669 = n15668 ^ n15665 ^ n3165 ;
  assign n15670 = n13132 ^ n9777 ^ 1'b0 ;
  assign n15671 = n4733 | n15670 ;
  assign n15672 = n15671 ^ n7935 ^ 1'b0 ;
  assign n15675 = ( x99 & ~n946 ) | ( x99 & n1482 ) | ( ~n946 & n1482 ) ;
  assign n15674 = n2010 ^ n702 ^ 1'b0 ;
  assign n15673 = n4131 & ~n8529 ;
  assign n15676 = n15675 ^ n15674 ^ n15673 ;
  assign n15677 = n4879 & n5555 ;
  assign n15678 = ~n12946 & n15677 ;
  assign n15679 = n15678 ^ n10501 ^ n3656 ;
  assign n15680 = ( n2665 & n15676 ) | ( n2665 & n15679 ) | ( n15676 & n15679 ) ;
  assign n15681 = n12167 ^ n5731 ^ n1160 ;
  assign n15682 = ( n7760 & n9036 ) | ( n7760 & ~n15681 ) | ( n9036 & ~n15681 ) ;
  assign n15684 = ( n681 & n4146 ) | ( n681 & ~n14802 ) | ( n4146 & ~n14802 ) ;
  assign n15685 = n15684 ^ n6941 ^ n4450 ;
  assign n15683 = n15299 ^ n13165 ^ n9146 ;
  assign n15686 = n15685 ^ n15683 ^ n9429 ;
  assign n15687 = n13242 | n14637 ;
  assign n15688 = n15687 ^ n14560 ^ n4673 ;
  assign n15691 = ( n5722 & n9285 ) | ( n5722 & n13855 ) | ( n9285 & n13855 ) ;
  assign n15689 = ( ~n3776 & n5114 ) | ( ~n3776 & n14883 ) | ( n5114 & n14883 ) ;
  assign n15690 = ( ~n4817 & n14015 ) | ( ~n4817 & n15689 ) | ( n14015 & n15689 ) ;
  assign n15692 = n15691 ^ n15690 ^ n1723 ;
  assign n15693 = n12663 ^ n4432 ^ 1'b0 ;
  assign n15694 = ( n654 & n3291 ) | ( n654 & n11200 ) | ( n3291 & n11200 ) ;
  assign n15696 = n6895 ^ n5820 ^ n2010 ;
  assign n15695 = n15647 ^ n2077 ^ n1938 ;
  assign n15697 = n15696 ^ n15695 ^ n6350 ;
  assign n15698 = ( n2061 & n15694 ) | ( n2061 & n15697 ) | ( n15694 & n15697 ) ;
  assign n15699 = n7975 ^ n5246 ^ n2604 ;
  assign n15700 = n15699 ^ n14878 ^ n4769 ;
  assign n15701 = n7258 ^ n6807 ^ n5752 ;
  assign n15702 = n15701 ^ n5381 ^ n1503 ;
  assign n15703 = n15702 ^ n14509 ^ 1'b0 ;
  assign n15704 = n14155 | n14404 ;
  assign n15705 = ( n1395 & n15703 ) | ( n1395 & ~n15704 ) | ( n15703 & ~n15704 ) ;
  assign n15706 = n3023 ^ n1836 ^ n505 ;
  assign n15707 = n15706 ^ n9522 ^ n1295 ;
  assign n15708 = ( n2405 & n11545 ) | ( n2405 & ~n13650 ) | ( n11545 & ~n13650 ) ;
  assign n15709 = n12647 | n15708 ;
  assign n15710 = n15709 ^ n8763 ^ 1'b0 ;
  assign n15711 = n8781 | n15710 ;
  assign n15712 = n4216 & n4691 ;
  assign n15713 = n1258 & n15712 ;
  assign n15714 = ( ~n618 & n4020 ) | ( ~n618 & n4613 ) | ( n4020 & n4613 ) ;
  assign n15715 = ~n11505 & n15714 ;
  assign n15716 = n15715 ^ n4828 ^ 1'b0 ;
  assign n15717 = ( n253 & n2420 ) | ( n253 & n2918 ) | ( n2420 & n2918 ) ;
  assign n15718 = n7743 & ~n13731 ;
  assign n15719 = n15717 & n15718 ;
  assign n15721 = n174 & n2810 ;
  assign n15722 = n7195 ^ n2262 ^ n1165 ;
  assign n15723 = n11994 | n15722 ;
  assign n15724 = n15721 | n15723 ;
  assign n15720 = ~n4063 & n4911 ;
  assign n15725 = n15724 ^ n15720 ^ 1'b0 ;
  assign n15726 = ( ~n1479 & n6163 ) | ( ~n1479 & n11216 ) | ( n6163 & n11216 ) ;
  assign n15727 = n15726 ^ n5114 ^ n1084 ;
  assign n15728 = n15727 ^ n14803 ^ 1'b0 ;
  assign n15729 = n8629 & ~n15728 ;
  assign n15730 = n15090 & n15729 ;
  assign n15731 = n13015 ^ n3896 ^ n963 ;
  assign n15732 = n916 | n5026 ;
  assign n15733 = n13140 ^ n5479 ^ 1'b0 ;
  assign n15734 = ~n14654 & n15733 ;
  assign n15735 = n12631 ^ n8588 ^ n5251 ;
  assign n15736 = n1395 ^ n734 ^ 1'b0 ;
  assign n15737 = n6030 ^ n3935 ^ 1'b0 ;
  assign n15738 = n7639 & ~n15737 ;
  assign n15739 = n2938 ^ n2487 ^ n2449 ;
  assign n15740 = n1783 & ~n15739 ;
  assign n15741 = ~n15738 & n15740 ;
  assign n15742 = ( n15735 & n15736 ) | ( n15735 & ~n15741 ) | ( n15736 & ~n15741 ) ;
  assign n15743 = ( n2748 & n4835 ) | ( n2748 & n14081 ) | ( n4835 & n14081 ) ;
  assign n15744 = ~n2957 & n9380 ;
  assign n15745 = ~n11703 & n15744 ;
  assign n15746 = ( n237 & n2265 ) | ( n237 & n3653 ) | ( n2265 & n3653 ) ;
  assign n15747 = n15746 ^ n10333 ^ n3475 ;
  assign n15748 = n15747 ^ x61 ^ 1'b0 ;
  assign n15749 = n15748 ^ n10676 ^ n10584 ;
  assign n15750 = ( n2705 & n3382 ) | ( n2705 & n5546 ) | ( n3382 & n5546 ) ;
  assign n15751 = ( ~n2506 & n3696 ) | ( ~n2506 & n5606 ) | ( n3696 & n5606 ) ;
  assign n15752 = ( n9579 & ~n15750 ) | ( n9579 & n15751 ) | ( ~n15750 & n15751 ) ;
  assign n15753 = ( n1865 & n2755 ) | ( n1865 & ~n3991 ) | ( n2755 & ~n3991 ) ;
  assign n15754 = n3590 | n15533 ;
  assign n15755 = n15753 | n15754 ;
  assign n15756 = n12058 ^ n3149 ^ 1'b0 ;
  assign n15757 = ( n182 & ~n2915 ) | ( n182 & n15756 ) | ( ~n2915 & n15756 ) ;
  assign n15758 = n3724 | n5213 ;
  assign n15759 = n2004 | n15758 ;
  assign n15760 = ~n1295 & n15759 ;
  assign n15761 = ~n4920 & n15760 ;
  assign n15762 = ( ~n4941 & n8166 ) | ( ~n4941 & n15761 ) | ( n8166 & n15761 ) ;
  assign n15763 = ( n565 & n9627 ) | ( n565 & n15762 ) | ( n9627 & n15762 ) ;
  assign n15764 = ( n9335 & n12728 ) | ( n9335 & ~n12975 ) | ( n12728 & ~n12975 ) ;
  assign n15765 = n1657 & n6990 ;
  assign n15766 = n15765 ^ n12541 ^ 1'b0 ;
  assign n15767 = ~n15764 & n15766 ;
  assign n15768 = ( n1004 & ~n1109 ) | ( n1004 & n1476 ) | ( ~n1109 & n1476 ) ;
  assign n15769 = n2861 & ~n7909 ;
  assign n15770 = n15769 ^ n11557 ^ n3568 ;
  assign n15771 = n15770 ^ n4939 ^ n2495 ;
  assign n15772 = ( n186 & ~n7333 ) | ( n186 & n7482 ) | ( ~n7333 & n7482 ) ;
  assign n15773 = n15772 ^ n13135 ^ n5121 ;
  assign n15774 = n7228 ^ n4524 ^ n3631 ;
  assign n15775 = n15774 ^ n10027 ^ n9973 ;
  assign n15776 = n15775 ^ n4659 ^ n272 ;
  assign n15777 = ( n545 & n2495 ) | ( n545 & ~n15776 ) | ( n2495 & ~n15776 ) ;
  assign n15779 = ~n605 & n6707 ;
  assign n15780 = n15779 ^ n6981 ^ 1'b0 ;
  assign n15781 = n15780 ^ n1750 ^ 1'b0 ;
  assign n15778 = ( ~n8603 & n8854 ) | ( ~n8603 & n12993 ) | ( n8854 & n12993 ) ;
  assign n15782 = n15781 ^ n15778 ^ n9075 ;
  assign n15783 = n8961 ^ n4336 ^ 1'b0 ;
  assign n15784 = ~n4463 & n15783 ;
  assign n15785 = n13674 ^ n4548 ^ n1661 ;
  assign n15786 = ( n4037 & n9001 ) | ( n4037 & ~n15785 ) | ( n9001 & ~n15785 ) ;
  assign n15787 = ( ~n14711 & n15784 ) | ( ~n14711 & n15786 ) | ( n15784 & n15786 ) ;
  assign n15788 = n3615 ^ n2019 ^ 1'b0 ;
  assign n15789 = n14864 & ~n15788 ;
  assign n15790 = n3607 ^ n1821 ^ n1280 ;
  assign n15791 = n3206 & ~n15790 ;
  assign n15792 = n15791 ^ n2448 ^ 1'b0 ;
  assign n15793 = ( ~n5801 & n6910 ) | ( ~n5801 & n15792 ) | ( n6910 & n15792 ) ;
  assign n15794 = ( n2234 & ~n12562 ) | ( n2234 & n15793 ) | ( ~n12562 & n15793 ) ;
  assign n15795 = n2231 & ~n9335 ;
  assign n15796 = ~x46 & n15795 ;
  assign n15797 = ( ~n3827 & n11117 ) | ( ~n3827 & n15796 ) | ( n11117 & n15796 ) ;
  assign n15798 = ( n2990 & ~n13059 ) | ( n2990 & n15797 ) | ( ~n13059 & n15797 ) ;
  assign n15799 = ~n4480 & n4838 ;
  assign n15800 = ( n256 & n9636 ) | ( n256 & n12651 ) | ( n9636 & n12651 ) ;
  assign n15801 = ( n8092 & n15799 ) | ( n8092 & ~n15800 ) | ( n15799 & ~n15800 ) ;
  assign n15802 = ( n6177 & n8653 ) | ( n6177 & n15801 ) | ( n8653 & n15801 ) ;
  assign n15803 = n2400 & ~n4851 ;
  assign n15804 = ( ~n1032 & n6373 ) | ( ~n1032 & n15803 ) | ( n6373 & n15803 ) ;
  assign n15805 = ( ~n10046 & n13073 ) | ( ~n10046 & n15804 ) | ( n13073 & n15804 ) ;
  assign n15806 = ( n14973 & n15802 ) | ( n14973 & n15805 ) | ( n15802 & n15805 ) ;
  assign n15807 = n6660 | n7528 ;
  assign n15808 = n14270 | n15807 ;
  assign n15809 = n15808 ^ n11485 ^ 1'b0 ;
  assign n15810 = n15809 ^ n1316 ^ 1'b0 ;
  assign n15811 = ( ~n3013 & n5638 ) | ( ~n3013 & n13150 ) | ( n5638 & n13150 ) ;
  assign n15812 = n3327 & n5618 ;
  assign n15813 = n15812 ^ n4588 ^ 1'b0 ;
  assign n15814 = ( n270 & n6783 ) | ( n270 & n14743 ) | ( n6783 & n14743 ) ;
  assign n15815 = n12688 | n15354 ;
  assign n15816 = n8107 & ~n15815 ;
  assign n15817 = ( n15813 & n15814 ) | ( n15813 & n15816 ) | ( n15814 & n15816 ) ;
  assign n15818 = ( n2784 & ~n4241 ) | ( n2784 & n7541 ) | ( ~n4241 & n7541 ) ;
  assign n15819 = n9056 | n15818 ;
  assign n15820 = n15819 ^ n13756 ^ 1'b0 ;
  assign n15821 = n8074 ^ n1898 ^ n1467 ;
  assign n15822 = n356 & ~n15266 ;
  assign n15823 = n7827 & n8575 ;
  assign n15824 = ( n15821 & ~n15822 ) | ( n15821 & n15823 ) | ( ~n15822 & n15823 ) ;
  assign n15825 = ( n1167 & ~n3911 ) | ( n1167 & n12862 ) | ( ~n3911 & n12862 ) ;
  assign n15826 = ( n1337 & n9715 ) | ( n1337 & n14848 ) | ( n9715 & n14848 ) ;
  assign n15827 = n13294 ^ n8435 ^ 1'b0 ;
  assign n15828 = ( n15825 & ~n15826 ) | ( n15825 & n15827 ) | ( ~n15826 & n15827 ) ;
  assign n15829 = n15828 ^ n7986 ^ 1'b0 ;
  assign n15830 = n13930 ^ n7839 ^ n3733 ;
  assign n15833 = ( n1395 & n1629 ) | ( n1395 & ~n5960 ) | ( n1629 & ~n5960 ) ;
  assign n15834 = n15833 ^ n5320 ^ 1'b0 ;
  assign n15831 = n393 | n11853 ;
  assign n15832 = n10213 | n15831 ;
  assign n15835 = n15834 ^ n15832 ^ n6512 ;
  assign n15836 = ( n3882 & n13971 ) | ( n3882 & ~n15835 ) | ( n13971 & ~n15835 ) ;
  assign n15837 = n9340 ^ n6481 ^ 1'b0 ;
  assign n15838 = n186 & ~n15837 ;
  assign n15839 = n13009 ^ n8593 ^ n5064 ;
  assign n15840 = ( n5028 & n15838 ) | ( n5028 & n15839 ) | ( n15838 & n15839 ) ;
  assign n15841 = n15840 ^ n11749 ^ n11640 ;
  assign n15844 = ( n7020 & n11011 ) | ( n7020 & ~n12782 ) | ( n11011 & ~n12782 ) ;
  assign n15845 = n5650 & ~n15844 ;
  assign n15846 = ~x40 & n15845 ;
  assign n15847 = n15846 ^ n13802 ^ n2369 ;
  assign n15842 = ( n2441 & ~n3683 ) | ( n2441 & n8629 ) | ( ~n3683 & n8629 ) ;
  assign n15843 = n15842 ^ n15587 ^ n2137 ;
  assign n15848 = n15847 ^ n15843 ^ 1'b0 ;
  assign n15849 = n5239 & n8072 ;
  assign n15850 = ~n11902 & n15849 ;
  assign n15852 = n13042 ^ n3882 ^ n925 ;
  assign n15851 = n11425 ^ n5560 ^ n3066 ;
  assign n15853 = n15852 ^ n15851 ^ n865 ;
  assign n15854 = n15853 ^ n15592 ^ n4473 ;
  assign n15855 = ( n12000 & ~n15850 ) | ( n12000 & n15854 ) | ( ~n15850 & n15854 ) ;
  assign n15856 = n7003 ^ n2528 ^ 1'b0 ;
  assign n15857 = n7420 | n15856 ;
  assign n15858 = ( n2445 & n12932 ) | ( n2445 & n15178 ) | ( n12932 & n15178 ) ;
  assign n15859 = ( ~n8669 & n8716 ) | ( ~n8669 & n13306 ) | ( n8716 & n13306 ) ;
  assign n15860 = ( n592 & n3956 ) | ( n592 & ~n9303 ) | ( n3956 & ~n9303 ) ;
  assign n15861 = n15860 ^ n3171 ^ n3139 ;
  assign n15862 = n5748 & ~n15861 ;
  assign n15863 = n12344 & n15862 ;
  assign n15868 = ( n2313 & n7588 ) | ( n2313 & ~n11467 ) | ( n7588 & ~n11467 ) ;
  assign n15869 = n15868 ^ n4806 ^ n514 ;
  assign n15864 = n9349 ^ n3165 ^ 1'b0 ;
  assign n15865 = n3817 & n15864 ;
  assign n15866 = n15865 ^ x71 ^ 1'b0 ;
  assign n15867 = n15866 ^ n7476 ^ n5052 ;
  assign n15870 = n15869 ^ n15867 ^ n11447 ;
  assign n15871 = n13220 ^ n2958 ^ 1'b0 ;
  assign n15872 = n12249 ^ n7110 ^ n3950 ;
  assign n15873 = n1837 & ~n15872 ;
  assign n15874 = n15873 ^ n9652 ^ n3285 ;
  assign n15875 = ( n2086 & n2248 ) | ( n2086 & ~n15874 ) | ( n2248 & ~n15874 ) ;
  assign n15876 = ( n1174 & n4549 ) | ( n1174 & ~n8996 ) | ( n4549 & ~n8996 ) ;
  assign n15877 = n15876 ^ n12029 ^ 1'b0 ;
  assign n15879 = ( n516 & n6383 ) | ( n516 & n8261 ) | ( n6383 & n8261 ) ;
  assign n15880 = ( n902 & ~n3179 ) | ( n902 & n15879 ) | ( ~n3179 & n15879 ) ;
  assign n15878 = ( x38 & n4079 ) | ( x38 & ~n12484 ) | ( n4079 & ~n12484 ) ;
  assign n15881 = n15880 ^ n15878 ^ n6277 ;
  assign n15882 = n15881 ^ n10293 ^ n6416 ;
  assign n15883 = ( n359 & ~n3195 ) | ( n359 & n3959 ) | ( ~n3195 & n3959 ) ;
  assign n15884 = ( n10409 & n12572 ) | ( n10409 & n15498 ) | ( n12572 & n15498 ) ;
  assign n15885 = n5328 | n10107 ;
  assign n15886 = n15885 ^ n2108 ^ 1'b0 ;
  assign n15890 = n7557 | n7840 ;
  assign n15891 = ( n975 & ~n11563 ) | ( n975 & n15890 ) | ( ~n11563 & n15890 ) ;
  assign n15892 = ( n1019 & ~n15369 ) | ( n1019 & n15891 ) | ( ~n15369 & n15891 ) ;
  assign n15887 = n9599 | n12918 ;
  assign n15888 = ( n2190 & ~n9244 ) | ( n2190 & n15887 ) | ( ~n9244 & n15887 ) ;
  assign n15889 = n10355 & n15888 ;
  assign n15893 = n15892 ^ n15889 ^ 1'b0 ;
  assign n15894 = n8382 ^ n1805 ^ n1239 ;
  assign n15895 = n7735 ^ n6309 ^ n5464 ;
  assign n15896 = n15895 ^ n13855 ^ n1333 ;
  assign n15902 = n5721 ^ n775 ^ 1'b0 ;
  assign n15897 = n15132 ^ n5280 ^ n4169 ;
  assign n15898 = ( n1476 & n5248 ) | ( n1476 & n7284 ) | ( n5248 & n7284 ) ;
  assign n15899 = n15898 ^ n4915 ^ 1'b0 ;
  assign n15900 = n15897 | n15899 ;
  assign n15901 = n14285 & ~n15900 ;
  assign n15903 = n15902 ^ n15901 ^ 1'b0 ;
  assign n15904 = ~n14030 & n15903 ;
  assign n15905 = ( n3693 & n7646 ) | ( n3693 & n12579 ) | ( n7646 & n12579 ) ;
  assign n15906 = ( n3336 & n12512 ) | ( n3336 & ~n15905 ) | ( n12512 & ~n15905 ) ;
  assign n15907 = n4600 ^ n4482 ^ n2784 ;
  assign n15908 = n6713 ^ n2525 ^ n1007 ;
  assign n15909 = ( n5113 & ~n15793 ) | ( n5113 & n15908 ) | ( ~n15793 & n15908 ) ;
  assign n15910 = n5783 | n15517 ;
  assign n15911 = n4136 & ~n15910 ;
  assign n15912 = n15909 & ~n15911 ;
  assign n15913 = ( ~n8149 & n9322 ) | ( ~n8149 & n13279 ) | ( n9322 & n13279 ) ;
  assign n15915 = n12469 ^ n10322 ^ n592 ;
  assign n15914 = ( ~n503 & n5140 ) | ( ~n503 & n14640 ) | ( n5140 & n14640 ) ;
  assign n15916 = n15915 ^ n15914 ^ n892 ;
  assign n15917 = ( n11640 & ~n15913 ) | ( n11640 & n15916 ) | ( ~n15913 & n15916 ) ;
  assign n15918 = ( n5935 & n7124 ) | ( n5935 & n15133 ) | ( n7124 & n15133 ) ;
  assign n15919 = n13991 ^ n10621 ^ 1'b0 ;
  assign n15920 = n15918 | n15919 ;
  assign n15921 = ( n472 & n3623 ) | ( n472 & ~n6110 ) | ( n3623 & ~n6110 ) ;
  assign n15922 = n387 | n13702 ;
  assign n15923 = ( ~n3104 & n15921 ) | ( ~n3104 & n15922 ) | ( n15921 & n15922 ) ;
  assign n15924 = ( n796 & n1685 ) | ( n796 & n6948 ) | ( n1685 & n6948 ) ;
  assign n15925 = n15924 ^ n12993 ^ n1645 ;
  assign n15926 = ( n4664 & ~n7870 ) | ( n4664 & n15925 ) | ( ~n7870 & n15925 ) ;
  assign n15927 = n1472 | n11584 ;
  assign n15928 = n15927 ^ n9814 ^ 1'b0 ;
  assign n15929 = n15928 ^ n10385 ^ n2078 ;
  assign n15930 = n6753 ^ n4974 ^ n1201 ;
  assign n15931 = n15930 ^ n15523 ^ n13616 ;
  assign n15932 = ( n5000 & n11772 ) | ( n5000 & ~n15931 ) | ( n11772 & ~n15931 ) ;
  assign n15933 = n3142 & ~n15175 ;
  assign n15934 = n15932 & n15933 ;
  assign n15935 = ~n4348 & n15934 ;
  assign n15936 = ~n3045 & n3352 ;
  assign n15937 = n15936 ^ n9431 ^ 1'b0 ;
  assign n15938 = ~n3599 & n15937 ;
  assign n15939 = n15938 ^ n4392 ^ 1'b0 ;
  assign n15940 = n12333 & ~n15018 ;
  assign n15941 = n15940 ^ n3224 ^ 1'b0 ;
  assign n15942 = n1037 ^ n314 ^ 1'b0 ;
  assign n15943 = ( n2364 & ~n6233 ) | ( n2364 & n15942 ) | ( ~n6233 & n15942 ) ;
  assign n15944 = n15943 ^ n5840 ^ 1'b0 ;
  assign n15945 = n15941 & n15944 ;
  assign n15946 = n15945 ^ n13615 ^ n13464 ;
  assign n15947 = n7904 ^ n7266 ^ n2687 ;
  assign n15948 = n5608 ^ n2868 ^ n1973 ;
  assign n15949 = n15948 ^ n15704 ^ n13430 ;
  assign n15950 = n4844 & ~n15086 ;
  assign n15951 = n3862 & ~n9858 ;
  assign n15952 = n15951 ^ n9164 ^ 1'b0 ;
  assign n15953 = n1600 & n5216 ;
  assign n15954 = ( n5667 & n9826 ) | ( n5667 & n15953 ) | ( n9826 & n15953 ) ;
  assign n15955 = ( n4824 & n8096 ) | ( n4824 & ~n10274 ) | ( n8096 & ~n10274 ) ;
  assign n15958 = n8032 ^ n2525 ^ n1748 ;
  assign n15959 = n1511 | n15958 ;
  assign n15960 = n15959 ^ n6260 ^ 1'b0 ;
  assign n15956 = n2493 & ~n15634 ;
  assign n15957 = n15956 ^ n14886 ^ n6247 ;
  assign n15961 = n15960 ^ n15957 ^ n1894 ;
  assign n15962 = n13752 ^ n2333 ^ 1'b0 ;
  assign n15963 = n4249 ^ n2317 ^ n1792 ;
  assign n15964 = ( x35 & n5146 ) | ( x35 & n9628 ) | ( n5146 & n9628 ) ;
  assign n15965 = ( n3606 & n9854 ) | ( n3606 & n11246 ) | ( n9854 & n11246 ) ;
  assign n15966 = ( ~n7165 & n9322 ) | ( ~n7165 & n15965 ) | ( n9322 & n15965 ) ;
  assign n15967 = n558 & n3084 ;
  assign n15968 = n15967 ^ n1420 ^ 1'b0 ;
  assign n15969 = n15968 ^ n8164 ^ n7263 ;
  assign n15970 = n15969 ^ n12666 ^ n461 ;
  assign n15971 = ~n9416 & n12562 ;
  assign n15972 = n15971 ^ n10560 ^ 1'b0 ;
  assign n15979 = n10667 ^ n6034 ^ n5260 ;
  assign n15978 = ( n4504 & n11347 ) | ( n4504 & ~n14611 ) | ( n11347 & ~n14611 ) ;
  assign n15973 = n5599 ^ n2646 ^ n667 ;
  assign n15974 = n15973 ^ n8234 ^ n5743 ;
  assign n15975 = n2934 & n13313 ;
  assign n15976 = ~n15974 & n15975 ;
  assign n15977 = n8425 & ~n15976 ;
  assign n15980 = n15979 ^ n15978 ^ n15977 ;
  assign n15981 = n5948 ^ n3661 ^ x127 ;
  assign n15982 = n15981 ^ n2890 ^ n1635 ;
  assign n15983 = n8011 ^ n7034 ^ n1635 ;
  assign n15985 = n2732 | n14968 ;
  assign n15984 = ( ~n2083 & n12031 ) | ( ~n2083 & n13272 ) | ( n12031 & n13272 ) ;
  assign n15986 = n15985 ^ n15984 ^ 1'b0 ;
  assign n15987 = n8434 | n15986 ;
  assign n15988 = n11174 ^ n3036 ^ x5 ;
  assign n15989 = n15988 ^ n8307 ^ n2122 ;
  assign n15990 = n15989 ^ n7349 ^ n3926 ;
  assign n15991 = ( ~n5078 & n7051 ) | ( ~n5078 & n12694 ) | ( n7051 & n12694 ) ;
  assign n15992 = n15991 ^ n12145 ^ n3518 ;
  assign n15993 = n10793 ^ n10621 ^ n3432 ;
  assign n15994 = n15993 ^ n5748 ^ n1398 ;
  assign n15995 = n1958 & n9638 ;
  assign n15996 = ( ~n2389 & n9547 ) | ( ~n2389 & n12513 ) | ( n9547 & n12513 ) ;
  assign n15997 = ( n1272 & n15995 ) | ( n1272 & n15996 ) | ( n15995 & n15996 ) ;
  assign n15998 = ( n516 & n4848 ) | ( n516 & n15997 ) | ( n4848 & n15997 ) ;
  assign n15999 = n12228 & n15613 ;
  assign n16000 = ~n9650 & n15999 ;
  assign n16001 = n7319 | n15303 ;
  assign n16002 = n16001 ^ n15722 ^ 1'b0 ;
  assign n16003 = ( ~n3342 & n16000 ) | ( ~n3342 & n16002 ) | ( n16000 & n16002 ) ;
  assign n16004 = n14053 ^ n12633 ^ n8671 ;
  assign n16005 = ( n1166 & ~n10570 ) | ( n1166 & n15571 ) | ( ~n10570 & n15571 ) ;
  assign n16006 = n15000 ^ n13634 ^ n8707 ;
  assign n16007 = ~n12411 & n14640 ;
  assign n16008 = ~x101 & n16007 ;
  assign n16009 = n16008 ^ n3010 ^ n1044 ;
  assign n16010 = n5550 | n11292 ;
  assign n16011 = ( ~n448 & n2861 ) | ( ~n448 & n5435 ) | ( n2861 & n5435 ) ;
  assign n16012 = ( n3208 & ~n15036 ) | ( n3208 & n16011 ) | ( ~n15036 & n16011 ) ;
  assign n16013 = ( ~x18 & x21 ) | ( ~x18 & n5469 ) | ( x21 & n5469 ) ;
  assign n16014 = n298 | n16013 ;
  assign n16015 = n4627 & ~n16014 ;
  assign n16017 = n329 & n5003 ;
  assign n16018 = ( n287 & n5382 ) | ( n287 & ~n16017 ) | ( n5382 & ~n16017 ) ;
  assign n16016 = ( n4495 & n7305 ) | ( n4495 & ~n7343 ) | ( n7305 & ~n7343 ) ;
  assign n16019 = n16018 ^ n16016 ^ n15097 ;
  assign n16020 = ( n3389 & ~n16015 ) | ( n3389 & n16019 ) | ( ~n16015 & n16019 ) ;
  assign n16021 = ( ~n8753 & n16012 ) | ( ~n8753 & n16020 ) | ( n16012 & n16020 ) ;
  assign n16022 = n11087 ^ n9160 ^ x23 ;
  assign n16023 = n15609 ^ n4939 ^ 1'b0 ;
  assign n16024 = n16022 | n16023 ;
  assign n16025 = n5277 ^ n2871 ^ 1'b0 ;
  assign n16026 = ( n8260 & n12690 ) | ( n8260 & n13756 ) | ( n12690 & n13756 ) ;
  assign n16027 = n16026 ^ n475 ^ 1'b0 ;
  assign n16028 = ~n16025 & n16027 ;
  assign n16029 = n11330 ^ n10998 ^ n184 ;
  assign n16032 = n543 | n2312 ;
  assign n16033 = n16032 ^ n1150 ^ 1'b0 ;
  assign n16034 = n3760 ^ n2637 ^ 1'b0 ;
  assign n16035 = n16033 | n16034 ;
  assign n16030 = n4142 & ~n7230 ;
  assign n16031 = ( n2245 & n9897 ) | ( n2245 & n16030 ) | ( n9897 & n16030 ) ;
  assign n16036 = n16035 ^ n16031 ^ n13553 ;
  assign n16037 = n4664 ^ n4351 ^ 1'b0 ;
  assign n16038 = n6210 & n16037 ;
  assign n16039 = ( n7633 & ~n9232 ) | ( n7633 & n16038 ) | ( ~n9232 & n16038 ) ;
  assign n16040 = ( n3557 & n11376 ) | ( n3557 & ~n11467 ) | ( n11376 & ~n11467 ) ;
  assign n16041 = n16040 ^ n3846 ^ n1412 ;
  assign n16042 = n8495 ^ n939 ^ 1'b0 ;
  assign n16043 = ( n4171 & n4569 ) | ( n4171 & ~n5910 ) | ( n4569 & ~n5910 ) ;
  assign n16044 = n16043 ^ n8862 ^ n3867 ;
  assign n16045 = n16044 ^ n5605 ^ 1'b0 ;
  assign n16046 = ( n2630 & n5738 ) | ( n2630 & n5770 ) | ( n5738 & n5770 ) ;
  assign n16047 = ( n1879 & ~n5075 ) | ( n1879 & n16046 ) | ( ~n5075 & n16046 ) ;
  assign n16048 = ( n11544 & n15838 ) | ( n11544 & ~n16047 ) | ( n15838 & ~n16047 ) ;
  assign n16049 = ~n4496 & n13814 ;
  assign n16050 = n16049 ^ n11227 ^ 1'b0 ;
  assign n16051 = n14971 ^ n12905 ^ n9584 ;
  assign n16052 = n14234 ^ n4764 ^ 1'b0 ;
  assign n16053 = ( n4418 & n16051 ) | ( n4418 & ~n16052 ) | ( n16051 & ~n16052 ) ;
  assign n16054 = ( n3193 & n6645 ) | ( n3193 & n14464 ) | ( n6645 & n14464 ) ;
  assign n16055 = ( n4587 & ~n5381 ) | ( n4587 & n6499 ) | ( ~n5381 & n6499 ) ;
  assign n16056 = n7825 & n15354 ;
  assign n16057 = ( n3173 & n4494 ) | ( n3173 & n13088 ) | ( n4494 & n13088 ) ;
  assign n16058 = n16057 ^ n3227 ^ n2673 ;
  assign n16059 = n11375 & n13437 ;
  assign n16060 = n16059 ^ n1292 ^ 1'b0 ;
  assign n16061 = n16060 ^ n3323 ^ 1'b0 ;
  assign n16062 = n16058 & n16061 ;
  assign n16063 = n14450 ^ n2704 ^ 1'b0 ;
  assign n16064 = n6202 | n16063 ;
  assign n16065 = ( n12911 & n14673 ) | ( n12911 & ~n16064 ) | ( n14673 & ~n16064 ) ;
  assign n16066 = n1954 ^ n1836 ^ 1'b0 ;
  assign n16067 = n16066 ^ n6773 ^ n6182 ;
  assign n16068 = ( n7409 & n13354 ) | ( n7409 & n16067 ) | ( n13354 & n16067 ) ;
  assign n16069 = n13919 ^ n13258 ^ n7846 ;
  assign n16070 = n560 & ~n1042 ;
  assign n16071 = n16070 ^ n11603 ^ n4122 ;
  assign n16072 = n6957 ^ n6679 ^ n6360 ;
  assign n16073 = n2143 & ~n5407 ;
  assign n16074 = n16073 ^ n10524 ^ 1'b0 ;
  assign n16075 = n16074 ^ n5494 ^ n1433 ;
  assign n16076 = ( ~n2698 & n16072 ) | ( ~n2698 & n16075 ) | ( n16072 & n16075 ) ;
  assign n16077 = n912 & ~n4709 ;
  assign n16078 = ( n16071 & ~n16076 ) | ( n16071 & n16077 ) | ( ~n16076 & n16077 ) ;
  assign n16079 = n14023 ^ n8926 ^ n7614 ;
  assign n16080 = n16079 ^ n12196 ^ n4939 ;
  assign n16081 = ( ~n863 & n6731 ) | ( ~n863 & n14468 ) | ( n6731 & n14468 ) ;
  assign n16082 = n14109 ^ n6719 ^ n3391 ;
  assign n16083 = ( ~n4336 & n7465 ) | ( ~n4336 & n11138 ) | ( n7465 & n11138 ) ;
  assign n16084 = n8456 & n16083 ;
  assign n16085 = n16082 & n16084 ;
  assign n16086 = n14743 ^ n559 ^ 1'b0 ;
  assign n16087 = ( n12393 & n16085 ) | ( n12393 & n16086 ) | ( n16085 & n16086 ) ;
  assign n16088 = ( n5321 & n9210 ) | ( n5321 & ~n9695 ) | ( n9210 & ~n9695 ) ;
  assign n16093 = n14641 ^ n9828 ^ n5959 ;
  assign n16089 = n5637 ^ n2433 ^ 1'b0 ;
  assign n16090 = n9224 | n16089 ;
  assign n16091 = n16090 ^ n2898 ^ 1'b0 ;
  assign n16092 = ~n7235 & n16091 ;
  assign n16094 = n16093 ^ n16092 ^ n1688 ;
  assign n16095 = n3798 & n16094 ;
  assign n16096 = ~n13279 & n16095 ;
  assign n16098 = n10777 ^ n1917 ^ n498 ;
  assign n16099 = n16098 ^ n5701 ^ n2158 ;
  assign n16100 = ( n4363 & n8227 ) | ( n4363 & n11290 ) | ( n8227 & n11290 ) ;
  assign n16101 = ~n11056 & n16100 ;
  assign n16102 = ( n12557 & ~n16099 ) | ( n12557 & n16101 ) | ( ~n16099 & n16101 ) ;
  assign n16097 = n1913 & ~n7810 ;
  assign n16103 = n16102 ^ n16097 ^ 1'b0 ;
  assign n16104 = ( n2108 & ~n2163 ) | ( n2108 & n3255 ) | ( ~n2163 & n3255 ) ;
  assign n16105 = ( n1822 & n2302 ) | ( n1822 & ~n2671 ) | ( n2302 & ~n2671 ) ;
  assign n16106 = ( n13369 & ~n14160 ) | ( n13369 & n16105 ) | ( ~n14160 & n16105 ) ;
  assign n16107 = ( ~n396 & n14995 ) | ( ~n396 & n16106 ) | ( n14995 & n16106 ) ;
  assign n16108 = n16107 ^ n15427 ^ 1'b0 ;
  assign n16109 = n15572 | n16108 ;
  assign n16110 = ~n3656 & n9605 ;
  assign n16111 = ( ~n16104 & n16109 ) | ( ~n16104 & n16110 ) | ( n16109 & n16110 ) ;
  assign n16112 = n13049 ^ n8782 ^ x66 ;
  assign n16113 = n3531 ^ n1423 ^ 1'b0 ;
  assign n16114 = ( n1999 & n3147 ) | ( n1999 & n12223 ) | ( n3147 & n12223 ) ;
  assign n16115 = n4487 & n16114 ;
  assign n16116 = ( n13507 & ~n16113 ) | ( n13507 & n16115 ) | ( ~n16113 & n16115 ) ;
  assign n16117 = ~n2051 & n16116 ;
  assign n16121 = n13528 ^ n9308 ^ n2191 ;
  assign n16118 = ( ~n447 & n1045 ) | ( ~n447 & n5030 ) | ( n1045 & n5030 ) ;
  assign n16119 = n16118 ^ n1983 ^ n766 ;
  assign n16120 = n14060 | n16119 ;
  assign n16122 = n16121 ^ n16120 ^ n8918 ;
  assign n16123 = n3567 ^ x31 ^ 1'b0 ;
  assign n16124 = n2405 ^ n479 ^ 1'b0 ;
  assign n16125 = n16123 & ~n16124 ;
  assign n16126 = n1214 & ~n2566 ;
  assign n16127 = n16126 ^ n11368 ^ 1'b0 ;
  assign n16128 = n16127 ^ n4016 ^ 1'b0 ;
  assign n16129 = n14803 ^ n6403 ^ n1617 ;
  assign n16130 = n2769 & n16129 ;
  assign n16131 = ~n8572 & n14317 ;
  assign n16135 = n12651 ^ n3262 ^ n1264 ;
  assign n16132 = ( ~n972 & n1728 ) | ( ~n972 & n6104 ) | ( n1728 & n6104 ) ;
  assign n16133 = n16132 ^ n4108 ^ n2121 ;
  assign n16134 = ( x2 & n11166 ) | ( x2 & n16133 ) | ( n11166 & n16133 ) ;
  assign n16136 = n16135 ^ n16134 ^ n15549 ;
  assign n16137 = n3709 & n4471 ;
  assign n16138 = n9301 ^ n1499 ^ 1'b0 ;
  assign n16139 = ~n9656 & n16138 ;
  assign n16140 = n16139 ^ n12911 ^ 1'b0 ;
  assign n16142 = ( ~n3576 & n8513 ) | ( ~n3576 & n13318 ) | ( n8513 & n13318 ) ;
  assign n16141 = n5838 | n16123 ;
  assign n16143 = n16142 ^ n16141 ^ n346 ;
  assign n16144 = ( n3396 & n3744 ) | ( n3396 & n6067 ) | ( n3744 & n6067 ) ;
  assign n16145 = n10100 ^ n410 ^ 1'b0 ;
  assign n16146 = n16144 & n16145 ;
  assign n16147 = ( n2058 & ~n4838 ) | ( n2058 & n9885 ) | ( ~n4838 & n9885 ) ;
  assign n16148 = ( n857 & n5720 ) | ( n857 & ~n16147 ) | ( n5720 & ~n16147 ) ;
  assign n16149 = ( ~n219 & n16146 ) | ( ~n219 & n16148 ) | ( n16146 & n16148 ) ;
  assign n16150 = n7641 & n15887 ;
  assign n16151 = n16150 ^ n4435 ^ 1'b0 ;
  assign n16152 = n8688 | n16151 ;
  assign n16153 = ( n8699 & n9116 ) | ( n8699 & n16152 ) | ( n9116 & n16152 ) ;
  assign n16154 = ( ~x2 & n4782 ) | ( ~x2 & n5592 ) | ( n4782 & n5592 ) ;
  assign n16155 = ( x48 & n1574 ) | ( x48 & n5300 ) | ( n1574 & n5300 ) ;
  assign n16156 = ( n9248 & n16154 ) | ( n9248 & ~n16155 ) | ( n16154 & ~n16155 ) ;
  assign n16157 = ( ~n1830 & n15199 ) | ( ~n1830 & n16043 ) | ( n15199 & n16043 ) ;
  assign n16158 = n16157 ^ n14347 ^ n3204 ;
  assign n16159 = ~n2990 & n16158 ;
  assign n16160 = n16156 & n16159 ;
  assign n16161 = ( n488 & n8586 ) | ( n488 & ~n8649 ) | ( n8586 & ~n8649 ) ;
  assign n16173 = n2147 ^ n1716 ^ n436 ;
  assign n16162 = ~n3806 & n14370 ;
  assign n16163 = n16162 ^ n3657 ^ 1'b0 ;
  assign n16164 = n14704 ^ n5038 ^ n2337 ;
  assign n16165 = n16163 | n16164 ;
  assign n16166 = n16165 ^ n2720 ^ 1'b0 ;
  assign n16167 = n6772 ^ n4998 ^ n2122 ;
  assign n16168 = n15099 ^ n6450 ^ n1936 ;
  assign n16169 = n16168 ^ n9828 ^ n1369 ;
  assign n16170 = n16169 ^ n8964 ^ n4401 ;
  assign n16171 = ( n5370 & ~n16167 ) | ( n5370 & n16170 ) | ( ~n16167 & n16170 ) ;
  assign n16172 = ( n5487 & n16166 ) | ( n5487 & ~n16171 ) | ( n16166 & ~n16171 ) ;
  assign n16174 = n16173 ^ n16172 ^ n3540 ;
  assign n16175 = n16174 ^ n13051 ^ n2579 ;
  assign n16176 = n482 | n5546 ;
  assign n16177 = ( n1255 & n10314 ) | ( n1255 & n16176 ) | ( n10314 & n16176 ) ;
  assign n16178 = n5569 | n9750 ;
  assign n16179 = ( ~n2933 & n6695 ) | ( ~n2933 & n8628 ) | ( n6695 & n8628 ) ;
  assign n16180 = n13787 ^ n11054 ^ n6966 ;
  assign n16187 = n8028 ^ n1562 ^ n844 ;
  assign n16185 = n15218 ^ n6158 ^ n1892 ;
  assign n16183 = n1452 & ~n8573 ;
  assign n16184 = n3188 & n16183 ;
  assign n16186 = n16185 ^ n16184 ^ n4202 ;
  assign n16181 = n3292 | n12366 ;
  assign n16182 = n16181 ^ n14656 ^ 1'b0 ;
  assign n16188 = n16187 ^ n16186 ^ n16182 ;
  assign n16189 = ( n867 & n6044 ) | ( n867 & n10552 ) | ( n6044 & n10552 ) ;
  assign n16190 = n16189 ^ n11237 ^ n1742 ;
  assign n16191 = n5450 ^ n3088 ^ n3074 ;
  assign n16192 = n16191 ^ n6041 ^ n3460 ;
  assign n16195 = ( n2358 & n3659 ) | ( n2358 & n11189 ) | ( n3659 & n11189 ) ;
  assign n16196 = n16195 ^ n15178 ^ n14359 ;
  assign n16193 = n8595 ^ n1226 ^ 1'b0 ;
  assign n16194 = ( ~n8364 & n14381 ) | ( ~n8364 & n16193 ) | ( n14381 & n16193 ) ;
  assign n16197 = n16196 ^ n16194 ^ n6171 ;
  assign n16198 = ( n1717 & n16192 ) | ( n1717 & ~n16197 ) | ( n16192 & ~n16197 ) ;
  assign n16199 = ( n2879 & ~n11939 ) | ( n2879 & n14144 ) | ( ~n11939 & n14144 ) ;
  assign n16200 = ( ~n5131 & n14078 ) | ( ~n5131 & n16199 ) | ( n14078 & n16199 ) ;
  assign n16201 = n233 & ~n12227 ;
  assign n16202 = x80 | n8338 ;
  assign n16203 = n16202 ^ n14966 ^ n14950 ;
  assign n16204 = ~n8594 & n12383 ;
  assign n16205 = n16204 ^ n11774 ^ 1'b0 ;
  assign n16207 = n1125 & n11250 ;
  assign n16206 = n12249 ^ n8727 ^ n7827 ;
  assign n16208 = n16207 ^ n16206 ^ n8412 ;
  assign n16209 = ( ~n264 & n1800 ) | ( ~n264 & n3877 ) | ( n1800 & n3877 ) ;
  assign n16210 = n16209 ^ n10701 ^ n980 ;
  assign n16211 = n16210 ^ n13872 ^ n13106 ;
  assign n16212 = ( n1086 & ~n5106 ) | ( n1086 & n5653 ) | ( ~n5106 & n5653 ) ;
  assign n16213 = ( n1654 & n5026 ) | ( n1654 & ~n16212 ) | ( n5026 & ~n16212 ) ;
  assign n16214 = n16213 ^ n3107 ^ 1'b0 ;
  assign n16215 = ( n7604 & n7931 ) | ( n7604 & n9952 ) | ( n7931 & n9952 ) ;
  assign n16216 = ( n2905 & ~n16214 ) | ( n2905 & n16215 ) | ( ~n16214 & n16215 ) ;
  assign n16217 = ( n6214 & n9545 ) | ( n6214 & ~n16216 ) | ( n9545 & ~n16216 ) ;
  assign n16218 = n1496 & n2862 ;
  assign n16219 = ( n15674 & n16217 ) | ( n15674 & ~n16218 ) | ( n16217 & ~n16218 ) ;
  assign n16220 = ( n1679 & ~n9378 ) | ( n1679 & n13758 ) | ( ~n9378 & n13758 ) ;
  assign n16221 = n15427 ^ n13772 ^ n4590 ;
  assign n16222 = ~n579 & n5419 ;
  assign n16223 = n16222 ^ n1664 ^ 1'b0 ;
  assign n16224 = n5493 ^ n2050 ^ 1'b0 ;
  assign n16225 = ~n11609 & n16224 ;
  assign n16229 = ~n1699 & n3140 ;
  assign n16226 = ( n1655 & ~n5341 ) | ( n1655 & n7754 ) | ( ~n5341 & n7754 ) ;
  assign n16227 = ( ~n8682 & n12484 ) | ( ~n8682 & n16226 ) | ( n12484 & n16226 ) ;
  assign n16228 = n10935 & n16227 ;
  assign n16230 = n16229 ^ n16228 ^ 1'b0 ;
  assign n16231 = n2845 & n16230 ;
  assign n16232 = n5753 ^ n2486 ^ 1'b0 ;
  assign n16233 = ( n1109 & n8637 ) | ( n1109 & ~n16232 ) | ( n8637 & ~n16232 ) ;
  assign n16234 = n2932 & n12336 ;
  assign n16235 = ~n16233 & n16234 ;
  assign n16237 = n7600 ^ n153 ^ 1'b0 ;
  assign n16236 = ( n631 & ~n3493 ) | ( n631 & n15747 ) | ( ~n3493 & n15747 ) ;
  assign n16238 = n16237 ^ n16236 ^ n15000 ;
  assign n16239 = n1456 & ~n16238 ;
  assign n16240 = n16235 & n16239 ;
  assign n16241 = n10907 ^ n6202 ^ n3119 ;
  assign n16242 = n16241 ^ n13385 ^ n12430 ;
  assign n16243 = ( n577 & n7294 ) | ( n577 & n9280 ) | ( n7294 & n9280 ) ;
  assign n16244 = n16243 ^ n12784 ^ n11672 ;
  assign n16245 = n8956 | n12652 ;
  assign n16246 = n2953 & ~n16245 ;
  assign n16247 = n9436 & n13637 ;
  assign n16248 = n15532 & n16247 ;
  assign n16249 = n7468 ^ n3844 ^ n296 ;
  assign n16250 = n3757 & ~n16249 ;
  assign n16251 = ~n283 & n16250 ;
  assign n16252 = n16251 ^ n525 ^ 1'b0 ;
  assign n16253 = n16248 | n16252 ;
  assign n16254 = n10828 ^ n4035 ^ n3262 ;
  assign n16255 = n16254 ^ n14567 ^ n7074 ;
  assign n16256 = ( n9156 & ~n11893 ) | ( n9156 & n14896 ) | ( ~n11893 & n14896 ) ;
  assign n16257 = n16256 ^ n12071 ^ n4181 ;
  assign n16258 = n1296 | n5552 ;
  assign n16259 = x90 & ~n16258 ;
  assign n16260 = ( n527 & n2314 ) | ( n527 & ~n11584 ) | ( n2314 & ~n11584 ) ;
  assign n16261 = n5259 & n16260 ;
  assign n16262 = n16261 ^ n14261 ^ n13031 ;
  assign n16263 = ( ~n2419 & n3859 ) | ( ~n2419 & n4080 ) | ( n3859 & n4080 ) ;
  assign n16264 = n16263 ^ n8694 ^ n3870 ;
  assign n16267 = n7208 & n9054 ;
  assign n16265 = n7333 ^ n2545 ^ n1097 ;
  assign n16266 = n16265 ^ n4792 ^ n3091 ;
  assign n16268 = n16267 ^ n16266 ^ n11385 ;
  assign n16269 = n3419 & ~n7654 ;
  assign n16270 = n16269 ^ n669 ^ 1'b0 ;
  assign n16271 = n3710 | n16270 ;
  assign n16272 = ~n1678 & n16271 ;
  assign n16273 = ( n2130 & ~n5525 ) | ( n2130 & n6986 ) | ( ~n5525 & n6986 ) ;
  assign n16274 = n16273 ^ n8698 ^ 1'b0 ;
  assign n16275 = ( n2040 & ~n2361 ) | ( n2040 & n9806 ) | ( ~n2361 & n9806 ) ;
  assign n16276 = ( n10612 & n12689 ) | ( n10612 & ~n16275 ) | ( n12689 & ~n16275 ) ;
  assign n16277 = n15195 ^ n3639 ^ 1'b0 ;
  assign n16278 = n435 | n16277 ;
  assign n16279 = n8500 | n16278 ;
  assign n16280 = n5289 ^ n4055 ^ x34 ;
  assign n16286 = n8984 ^ n1503 ^ 1'b0 ;
  assign n16287 = n4791 | n16286 ;
  assign n16285 = n9391 ^ n7555 ^ n6433 ;
  assign n16288 = n16287 ^ n16285 ^ n7658 ;
  assign n16281 = ( n2456 & ~n3089 ) | ( n2456 & n7622 ) | ( ~n3089 & n7622 ) ;
  assign n16282 = ( n200 & n3621 ) | ( n200 & ~n5287 ) | ( n3621 & ~n5287 ) ;
  assign n16283 = ( n2554 & ~n9545 ) | ( n2554 & n16282 ) | ( ~n9545 & n16282 ) ;
  assign n16284 = ( n13247 & n16281 ) | ( n13247 & n16283 ) | ( n16281 & n16283 ) ;
  assign n16289 = n16288 ^ n16284 ^ n15879 ;
  assign n16290 = n16289 ^ n6487 ^ n478 ;
  assign n16291 = n16290 ^ n12222 ^ 1'b0 ;
  assign n16292 = n16280 & ~n16291 ;
  assign n16293 = ( n5272 & ~n11671 ) | ( n5272 & n15634 ) | ( ~n11671 & n15634 ) ;
  assign n16294 = n9303 ^ n4024 ^ 1'b0 ;
  assign n16295 = n747 & n16294 ;
  assign n16296 = ~n5625 & n16295 ;
  assign n16297 = n16293 & n16296 ;
  assign n16298 = ( n3015 & n3365 ) | ( n3015 & n16297 ) | ( n3365 & n16297 ) ;
  assign n16303 = n4252 ^ n1568 ^ 1'b0 ;
  assign n16299 = n9434 | n9542 ;
  assign n16300 = n1465 | n16299 ;
  assign n16301 = ~n176 & n16300 ;
  assign n16302 = n16301 ^ n14139 ^ 1'b0 ;
  assign n16304 = n16303 ^ n16302 ^ n7366 ;
  assign n16309 = ( n5421 & n5770 ) | ( n5421 & n12157 ) | ( n5770 & n12157 ) ;
  assign n16310 = n5404 & n16309 ;
  assign n16305 = n6358 ^ n1759 ^ 1'b0 ;
  assign n16306 = n14932 & ~n16305 ;
  assign n16307 = x111 & n16306 ;
  assign n16308 = n16307 ^ n3118 ^ 1'b0 ;
  assign n16311 = n16310 ^ n16308 ^ n8862 ;
  assign n16312 = n9773 & n13929 ;
  assign n16313 = n16312 ^ n959 ^ 1'b0 ;
  assign n16314 = n12325 | n16313 ;
  assign n16315 = n16314 ^ n2489 ^ 1'b0 ;
  assign n16316 = n15953 ^ n15221 ^ n4348 ;
  assign n16317 = n6773 | n16316 ;
  assign n16321 = n4836 ^ n2665 ^ n1056 ;
  assign n16322 = ( ~n8436 & n10226 ) | ( ~n8436 & n16321 ) | ( n10226 & n16321 ) ;
  assign n16318 = n11131 & ~n12780 ;
  assign n16319 = ~n3572 & n16318 ;
  assign n16320 = n8891 & n16319 ;
  assign n16323 = n16322 ^ n16320 ^ n12193 ;
  assign n16324 = ( ~n1063 & n9891 ) | ( ~n1063 & n10831 ) | ( n9891 & n10831 ) ;
  assign n16326 = n6972 ^ n1135 ^ 1'b0 ;
  assign n16327 = ~n209 & n16326 ;
  assign n16328 = n10251 ^ n9428 ^ n2609 ;
  assign n16329 = ( n12208 & ~n16327 ) | ( n12208 & n16328 ) | ( ~n16327 & n16328 ) ;
  assign n16325 = n12189 ^ n6548 ^ n1932 ;
  assign n16330 = n16329 ^ n16325 ^ n12114 ;
  assign n16331 = n16330 ^ n14609 ^ n11328 ;
  assign n16332 = ( n2478 & n2504 ) | ( n2478 & ~n8624 ) | ( n2504 & ~n8624 ) ;
  assign n16333 = ( n6571 & n10197 ) | ( n6571 & n16332 ) | ( n10197 & n16332 ) ;
  assign n16334 = n8006 ^ n5047 ^ n642 ;
  assign n16335 = n16334 ^ n14265 ^ n9093 ;
  assign n16336 = n306 & n9160 ;
  assign n16337 = n16335 & n16336 ;
  assign n16338 = n10722 ^ n6273 ^ 1'b0 ;
  assign n16339 = n3895 & ~n16338 ;
  assign n16340 = n9044 ^ n3262 ^ 1'b0 ;
  assign n16341 = n16340 ^ n9476 ^ n8068 ;
  assign n16342 = n13525 ^ n10659 ^ 1'b0 ;
  assign n16343 = n16341 & n16342 ;
  assign n16344 = n6026 ^ n5310 ^ 1'b0 ;
  assign n16345 = ( n2549 & n11297 ) | ( n2549 & ~n16344 ) | ( n11297 & ~n16344 ) ;
  assign n16347 = ( n2804 & n3339 ) | ( n2804 & n3574 ) | ( n3339 & n3574 ) ;
  assign n16348 = ( n3927 & n14669 ) | ( n3927 & ~n16347 ) | ( n14669 & ~n16347 ) ;
  assign n16346 = ( n6121 & n6716 ) | ( n6121 & ~n15265 ) | ( n6716 & ~n15265 ) ;
  assign n16349 = n16348 ^ n16346 ^ n13064 ;
  assign n16350 = ( n4917 & n15469 ) | ( n4917 & ~n16349 ) | ( n15469 & ~n16349 ) ;
  assign n16351 = ( n1952 & n15508 ) | ( n1952 & n16350 ) | ( n15508 & n16350 ) ;
  assign n16365 = ( n652 & ~n7590 ) | ( n652 & n9472 ) | ( ~n7590 & n9472 ) ;
  assign n16360 = ( n5661 & n7229 ) | ( n5661 & ~n7387 ) | ( n7229 & ~n7387 ) ;
  assign n16361 = n3060 ^ n441 ^ 1'b0 ;
  assign n16362 = n1659 & n16361 ;
  assign n16363 = n16360 & n16362 ;
  assign n16352 = n11898 ^ n11285 ^ n5747 ;
  assign n16353 = n3660 | n11557 ;
  assign n16354 = n16353 ^ n1757 ^ 1'b0 ;
  assign n16355 = n16354 ^ n4253 ^ n3712 ;
  assign n16356 = ( n2725 & n9300 ) | ( n2725 & n16355 ) | ( n9300 & n16355 ) ;
  assign n16357 = ( n4423 & ~n9712 ) | ( n4423 & n16356 ) | ( ~n9712 & n16356 ) ;
  assign n16358 = ( ~n2004 & n16352 ) | ( ~n2004 & n16357 ) | ( n16352 & n16357 ) ;
  assign n16359 = n16358 ^ n14095 ^ n1745 ;
  assign n16364 = n16363 ^ n16359 ^ n13833 ;
  assign n16366 = n16365 ^ n16364 ^ n2291 ;
  assign n16367 = n6344 ^ n3847 ^ n141 ;
  assign n16368 = n7399 ^ n3689 ^ 1'b0 ;
  assign n16369 = n16367 | n16368 ;
  assign n16370 = n16369 ^ n3600 ^ n331 ;
  assign n16371 = n3742 & n10543 ;
  assign n16372 = n16371 ^ n12040 ^ 1'b0 ;
  assign n16373 = ~n7950 & n14024 ;
  assign n16374 = n16373 ^ n2419 ^ 1'b0 ;
  assign n16375 = n4096 | n15993 ;
  assign n16376 = n16374 & ~n16375 ;
  assign n16378 = n6697 & n9869 ;
  assign n16377 = ( n2504 & n6942 ) | ( n2504 & n12491 ) | ( n6942 & n12491 ) ;
  assign n16379 = n16378 ^ n16377 ^ n7891 ;
  assign n16382 = ( n5280 & ~n6653 ) | ( n5280 & n10922 ) | ( ~n6653 & n10922 ) ;
  assign n16381 = n5552 | n5896 ;
  assign n16383 = n16382 ^ n16381 ^ 1'b0 ;
  assign n16380 = n7003 ^ n1350 ^ 1'b0 ;
  assign n16384 = n16383 ^ n16380 ^ 1'b0 ;
  assign n16385 = ( n4711 & ~n8303 ) | ( n4711 & n16384 ) | ( ~n8303 & n16384 ) ;
  assign n16391 = n6601 ^ n3859 ^ n360 ;
  assign n16392 = n258 & ~n2082 ;
  assign n16393 = n16392 ^ n11891 ^ 1'b0 ;
  assign n16394 = ( ~n5193 & n16391 ) | ( ~n5193 & n16393 ) | ( n16391 & n16393 ) ;
  assign n16395 = n3762 | n16394 ;
  assign n16387 = n14559 ^ n11813 ^ n1560 ;
  assign n16386 = ( n477 & n931 ) | ( n477 & n12928 ) | ( n931 & n12928 ) ;
  assign n16388 = n16387 ^ n16386 ^ n705 ;
  assign n16389 = ~n705 & n3088 ;
  assign n16390 = ( ~n11555 & n16388 ) | ( ~n11555 & n16389 ) | ( n16388 & n16389 ) ;
  assign n16396 = n16395 ^ n16390 ^ n163 ;
  assign n16397 = ( x100 & ~n3180 ) | ( x100 & n7481 ) | ( ~n3180 & n7481 ) ;
  assign n16398 = n7839 ^ n4479 ^ n2212 ;
  assign n16399 = n2488 | n16398 ;
  assign n16400 = n16397 | n16399 ;
  assign n16401 = ( n4624 & n10101 ) | ( n4624 & n16400 ) | ( n10101 & n16400 ) ;
  assign n16402 = n12847 ^ n9443 ^ 1'b0 ;
  assign n16403 = n9127 & ~n16402 ;
  assign n16404 = ( n3470 & ~n11459 ) | ( n3470 & n12794 ) | ( ~n11459 & n12794 ) ;
  assign n16405 = ( n1685 & n15965 ) | ( n1685 & n16404 ) | ( n15965 & n16404 ) ;
  assign n16406 = n16405 ^ n15024 ^ n2982 ;
  assign n16407 = n12265 ^ n8699 ^ n5662 ;
  assign n16408 = n10182 ^ n5211 ^ n2068 ;
  assign n16409 = n4527 & n16408 ;
  assign n16410 = ~n8668 & n16409 ;
  assign n16411 = n7567 ^ n4555 ^ n565 ;
  assign n16412 = ( n15290 & n16410 ) | ( n15290 & ~n16411 ) | ( n16410 & ~n16411 ) ;
  assign n16413 = n14222 ^ n11704 ^ n9957 ;
  assign n16414 = n10819 ^ n3927 ^ n3266 ;
  assign n16415 = n1761 | n16414 ;
  assign n16416 = n16415 ^ n6571 ^ n5879 ;
  assign n16417 = n2446 & ~n12351 ;
  assign n16418 = n16416 & n16417 ;
  assign n16419 = n13152 ^ n3175 ^ n2178 ;
  assign n16420 = ( n5702 & ~n8986 ) | ( n5702 & n16419 ) | ( ~n8986 & n16419 ) ;
  assign n16421 = n567 & ~n16420 ;
  assign n16422 = n468 | n13326 ;
  assign n16423 = n5584 & ~n11855 ;
  assign n16424 = n16423 ^ n6241 ^ 1'b0 ;
  assign n16425 = n11052 ^ n6005 ^ n3820 ;
  assign n16426 = n16425 ^ n3243 ^ 1'b0 ;
  assign n16427 = n713 & ~n16426 ;
  assign n16428 = ( n2292 & n16424 ) | ( n2292 & ~n16427 ) | ( n16424 & ~n16427 ) ;
  assign n16429 = ( n3196 & n8017 ) | ( n3196 & n16428 ) | ( n8017 & n16428 ) ;
  assign n16430 = n16422 & ~n16429 ;
  assign n16431 = n16167 ^ n9506 ^ n5931 ;
  assign n16432 = ~n3987 & n8639 ;
  assign n16433 = ~n16431 & n16432 ;
  assign n16436 = ( n4320 & n6779 ) | ( n4320 & n13365 ) | ( n6779 & n13365 ) ;
  assign n16434 = ( ~n1607 & n7403 ) | ( ~n1607 & n9064 ) | ( n7403 & n9064 ) ;
  assign n16435 = n16434 ^ n4985 ^ n4104 ;
  assign n16437 = n16436 ^ n16435 ^ 1'b0 ;
  assign n16438 = n13917 ^ n3499 ^ n3193 ;
  assign n16439 = ( n2316 & n4243 ) | ( n2316 & ~n10054 ) | ( n4243 & ~n10054 ) ;
  assign n16446 = n6260 ^ n4560 ^ n3995 ;
  assign n16440 = n14249 ^ n13074 ^ 1'b0 ;
  assign n16441 = n8562 | n16440 ;
  assign n16442 = n970 | n4598 ;
  assign n16443 = n16442 ^ n7731 ^ n6721 ;
  assign n16444 = n13437 & n16443 ;
  assign n16445 = n16441 & n16444 ;
  assign n16447 = n16446 ^ n16445 ^ 1'b0 ;
  assign n16448 = ( n2842 & n16439 ) | ( n2842 & n16447 ) | ( n16439 & n16447 ) ;
  assign n16449 = n13552 ^ n9302 ^ n4351 ;
  assign n16450 = n5664 & n14387 ;
  assign n16451 = n16450 ^ n11973 ^ 1'b0 ;
  assign n16452 = n16451 ^ n8536 ^ n8510 ;
  assign n16453 = ( ~n13898 & n16449 ) | ( ~n13898 & n16452 ) | ( n16449 & n16452 ) ;
  assign n16454 = n6113 | n6202 ;
  assign n16455 = n9269 & ~n16454 ;
  assign n16456 = n3987 | n16455 ;
  assign n16457 = n6953 & ~n16456 ;
  assign n16458 = n3557 & n12012 ;
  assign n16459 = ~n7741 & n16458 ;
  assign n16460 = n16459 ^ n10416 ^ n319 ;
  assign n16461 = n16460 ^ n11516 ^ n7023 ;
  assign n16462 = n8063 ^ n3843 ^ n3230 ;
  assign n16463 = ( ~n4974 & n12913 ) | ( ~n4974 & n16462 ) | ( n12913 & n16462 ) ;
  assign n16464 = n16463 ^ n3883 ^ 1'b0 ;
  assign n16465 = ~n16461 & n16464 ;
  assign n16466 = ( ~n1675 & n11125 ) | ( ~n1675 & n16442 ) | ( n11125 & n16442 ) ;
  assign n16467 = n16466 ^ n8061 ^ n6482 ;
  assign n16468 = ( n1822 & n6107 ) | ( n1822 & ~n16467 ) | ( n6107 & ~n16467 ) ;
  assign n16469 = ( ~n5735 & n10711 ) | ( ~n5735 & n14645 ) | ( n10711 & n14645 ) ;
  assign n16479 = ( n2674 & n6413 ) | ( n2674 & ~n6802 ) | ( n6413 & ~n6802 ) ;
  assign n16478 = n8974 ^ n4697 ^ n652 ;
  assign n16470 = n3045 ^ n2540 ^ n2186 ;
  assign n16471 = n2391 & ~n3866 ;
  assign n16472 = ~n1084 & n15907 ;
  assign n16473 = n11814 & n16472 ;
  assign n16474 = n16471 | n16473 ;
  assign n16475 = n16470 & ~n16474 ;
  assign n16476 = n16475 ^ n6244 ^ n775 ;
  assign n16477 = n16476 ^ n14971 ^ n4752 ;
  assign n16480 = n16479 ^ n16478 ^ n16477 ;
  assign n16481 = n11140 ^ n746 ^ 1'b0 ;
  assign n16482 = n16481 ^ n10913 ^ 1'b0 ;
  assign n16483 = n16482 ^ n4838 ^ n3576 ;
  assign n16484 = n16483 ^ n11702 ^ n4891 ;
  assign n16485 = n2230 ^ n1833 ^ n1665 ;
  assign n16486 = ( ~n1822 & n5260 ) | ( ~n1822 & n16485 ) | ( n5260 & n16485 ) ;
  assign n16487 = ( n6793 & n9469 ) | ( n6793 & ~n16486 ) | ( n9469 & ~n16486 ) ;
  assign n16488 = n6200 ^ n3000 ^ n2639 ;
  assign n16489 = n15768 ^ n8525 ^ 1'b0 ;
  assign n16490 = n5458 & n13002 ;
  assign n16491 = n5022 ^ n4701 ^ 1'b0 ;
  assign n16492 = ~n11650 & n15354 ;
  assign n16493 = n16492 ^ n3951 ^ 1'b0 ;
  assign n16494 = n6465 | n16493 ;
  assign n16495 = ( n2649 & ~n3520 ) | ( n2649 & n4235 ) | ( ~n3520 & n4235 ) ;
  assign n16496 = n16495 ^ n15268 ^ n7710 ;
  assign n16497 = ( ~n5603 & n11826 ) | ( ~n5603 & n12478 ) | ( n11826 & n12478 ) ;
  assign n16498 = n2068 & n16497 ;
  assign n16499 = ( n153 & n3186 ) | ( n153 & ~n7532 ) | ( n3186 & ~n7532 ) ;
  assign n16500 = ~n4804 & n16499 ;
  assign n16501 = n16500 ^ n5181 ^ 1'b0 ;
  assign n16502 = n14459 & n16501 ;
  assign n16503 = n16502 ^ n4032 ^ n2130 ;
  assign n16504 = n8637 ^ n1462 ^ x29 ;
  assign n16505 = n8418 ^ n5365 ^ 1'b0 ;
  assign n16506 = n1386 | n16505 ;
  assign n16507 = ( n1134 & n6272 ) | ( n1134 & n14477 ) | ( n6272 & n14477 ) ;
  assign n16508 = ( n9010 & ~n16506 ) | ( n9010 & n16507 ) | ( ~n16506 & n16507 ) ;
  assign n16509 = n16508 ^ n1186 ^ 1'b0 ;
  assign n16510 = ~n2549 & n16509 ;
  assign n16511 = n14677 ^ n5655 ^ n2042 ;
  assign n16512 = n1688 | n5892 ;
  assign n16513 = n16512 ^ n13536 ^ 1'b0 ;
  assign n16514 = n16513 ^ n3022 ^ 1'b0 ;
  assign n16515 = ~n16511 & n16514 ;
  assign n16516 = n9417 ^ n5246 ^ n489 ;
  assign n16517 = n16516 ^ n5216 ^ n520 ;
  assign n16518 = ( n892 & n9564 ) | ( n892 & ~n16517 ) | ( n9564 & ~n16517 ) ;
  assign n16519 = n16518 ^ n12742 ^ n2086 ;
  assign n16520 = n4899 & ~n16031 ;
  assign n16521 = ~n4995 & n16520 ;
  assign n16522 = ( n1427 & n12185 ) | ( n1427 & n16521 ) | ( n12185 & n16521 ) ;
  assign n16523 = n5625 ^ n3200 ^ n1104 ;
  assign n16524 = n4148 & ~n6469 ;
  assign n16525 = n16524 ^ n2421 ^ 1'b0 ;
  assign n16526 = ~n5038 & n7195 ;
  assign n16527 = n16525 & n16526 ;
  assign n16528 = ( n4247 & n11404 ) | ( n4247 & ~n16527 ) | ( n11404 & ~n16527 ) ;
  assign n16529 = n12500 ^ n5380 ^ 1'b0 ;
  assign n16532 = n11460 ^ n9119 ^ n8756 ;
  assign n16530 = n8041 ^ n6560 ^ n3454 ;
  assign n16531 = ( n3695 & n10878 ) | ( n3695 & n16530 ) | ( n10878 & n16530 ) ;
  assign n16533 = n16532 ^ n16531 ^ n10472 ;
  assign n16534 = ( n633 & ~n1005 ) | ( n633 & n1300 ) | ( ~n1005 & n1300 ) ;
  assign n16535 = ( n1567 & n4868 ) | ( n1567 & n16534 ) | ( n4868 & n16534 ) ;
  assign n16536 = n1027 | n6679 ;
  assign n16537 = ( n3566 & ~n11069 ) | ( n3566 & n16536 ) | ( ~n11069 & n16536 ) ;
  assign n16538 = ( n3678 & n11909 ) | ( n3678 & ~n16537 ) | ( n11909 & ~n16537 ) ;
  assign n16539 = ( n14608 & ~n16535 ) | ( n14608 & n16538 ) | ( ~n16535 & n16538 ) ;
  assign n16540 = n14560 ^ n2348 ^ n2237 ;
  assign n16541 = n16540 ^ n5592 ^ 1'b0 ;
  assign n16542 = ~n4954 & n16541 ;
  assign n16543 = n16542 ^ n13946 ^ 1'b0 ;
  assign n16544 = n12657 ^ n6930 ^ n6509 ;
  assign n16545 = n16544 ^ n7280 ^ 1'b0 ;
  assign n16546 = n14552 & ~n16545 ;
  assign n16547 = n12491 ^ n11700 ^ n7397 ;
  assign n16553 = n3671 ^ n654 ^ n454 ;
  assign n16554 = n16553 ^ n6262 ^ n941 ;
  assign n16555 = n16554 ^ n14644 ^ n3547 ;
  assign n16548 = n3068 & ~n11717 ;
  assign n16549 = n4501 | n16548 ;
  assign n16550 = n16549 ^ n234 ^ 1'b0 ;
  assign n16551 = ( ~n4936 & n5989 ) | ( ~n4936 & n16550 ) | ( n5989 & n16550 ) ;
  assign n16552 = ( n244 & n11678 ) | ( n244 & n16551 ) | ( n11678 & n16551 ) ;
  assign n16556 = n16555 ^ n16552 ^ n7826 ;
  assign n16557 = n3367 & n6429 ;
  assign n16558 = n16557 ^ n3403 ^ 1'b0 ;
  assign n16559 = n3255 & n14504 ;
  assign n16560 = ( ~n2701 & n2734 ) | ( ~n2701 & n16559 ) | ( n2734 & n16559 ) ;
  assign n16561 = ~n7270 & n16560 ;
  assign n16562 = n16558 & n16561 ;
  assign n16567 = n1949 & ~n13116 ;
  assign n16563 = n8838 ^ n8563 ^ n2016 ;
  assign n16564 = n8294 ^ n3278 ^ 1'b0 ;
  assign n16565 = n349 & n16564 ;
  assign n16566 = ( ~n3251 & n16563 ) | ( ~n3251 & n16565 ) | ( n16563 & n16565 ) ;
  assign n16568 = n16567 ^ n16566 ^ n470 ;
  assign n16569 = ~n4214 & n6052 ;
  assign n16570 = n16569 ^ n9125 ^ 1'b0 ;
  assign n16571 = ~n12912 & n16570 ;
  assign n16572 = n16571 ^ n6590 ^ 1'b0 ;
  assign n16573 = n11898 ^ n1610 ^ n573 ;
  assign n16574 = ~n5484 & n16573 ;
  assign n16575 = ( n2991 & ~n5340 ) | ( n2991 & n15974 ) | ( ~n5340 & n15974 ) ;
  assign n16576 = n16575 ^ n8011 ^ 1'b0 ;
  assign n16577 = n16574 & n16576 ;
  assign n16578 = n4817 ^ n2237 ^ 1'b0 ;
  assign n16579 = n16578 ^ n15913 ^ n13743 ;
  assign n16589 = n5441 & n11420 ;
  assign n16580 = n16226 ^ n3086 ^ x4 ;
  assign n16581 = ( n5733 & n12647 ) | ( n5733 & n16580 ) | ( n12647 & n16580 ) ;
  assign n16582 = n13380 | n16581 ;
  assign n16583 = n11565 & ~n16582 ;
  assign n16584 = n1982 & ~n16553 ;
  assign n16585 = ( ~n3174 & n3912 ) | ( ~n3174 & n13695 ) | ( n3912 & n13695 ) ;
  assign n16586 = n5608 ^ n4068 ^ 1'b0 ;
  assign n16587 = ( n16584 & ~n16585 ) | ( n16584 & n16586 ) | ( ~n16585 & n16586 ) ;
  assign n16588 = ( n9479 & n16583 ) | ( n9479 & n16587 ) | ( n16583 & n16587 ) ;
  assign n16590 = n16589 ^ n16588 ^ 1'b0 ;
  assign n16592 = ( n7058 & n9207 ) | ( n7058 & n10606 ) | ( n9207 & n10606 ) ;
  assign n16593 = ( n1418 & n12887 ) | ( n1418 & ~n16592 ) | ( n12887 & ~n16592 ) ;
  assign n16591 = n766 & ~n13708 ;
  assign n16594 = n16593 ^ n16591 ^ 1'b0 ;
  assign n16599 = ( ~n395 & n8944 ) | ( ~n395 & n10210 ) | ( n8944 & n10210 ) ;
  assign n16595 = n5072 ^ n3618 ^ n3561 ;
  assign n16596 = ~n2726 & n15890 ;
  assign n16597 = n12384 & n16596 ;
  assign n16598 = n16595 & ~n16597 ;
  assign n16600 = n16599 ^ n16598 ^ n11589 ;
  assign n16601 = n10280 ^ n6442 ^ n3865 ;
  assign n16602 = n8339 ^ n1860 ^ 1'b0 ;
  assign n16603 = n2598 | n16602 ;
  assign n16604 = ( ~n1451 & n16601 ) | ( ~n1451 & n16603 ) | ( n16601 & n16603 ) ;
  assign n16605 = n1495 & ~n1912 ;
  assign n16606 = n16605 ^ n171 ^ 1'b0 ;
  assign n16607 = ( n3105 & n4176 ) | ( n3105 & ~n16606 ) | ( n4176 & ~n16606 ) ;
  assign n16608 = n16607 ^ n4793 ^ n235 ;
  assign n16609 = ( n551 & n7496 ) | ( n551 & n16608 ) | ( n7496 & n16608 ) ;
  assign n16610 = n16609 ^ n14665 ^ n2859 ;
  assign n16611 = n16610 ^ n14288 ^ 1'b0 ;
  assign n16612 = n3878 & n16611 ;
  assign n16613 = n857 & n4866 ;
  assign n16614 = ( ~n5658 & n7182 ) | ( ~n5658 & n16613 ) | ( n7182 & n16613 ) ;
  assign n16615 = n16614 ^ n11612 ^ n1642 ;
  assign n16616 = ( n10638 & n11259 ) | ( n10638 & ~n12133 ) | ( n11259 & ~n12133 ) ;
  assign n16617 = n7784 ^ n4519 ^ 1'b0 ;
  assign n16618 = n16617 ^ n8962 ^ n8956 ;
  assign n16619 = ( n7951 & n12499 ) | ( n7951 & ~n16618 ) | ( n12499 & ~n16618 ) ;
  assign n16620 = ( n1794 & n2496 ) | ( n1794 & n8251 ) | ( n2496 & n8251 ) ;
  assign n16621 = ( n14525 & ~n16619 ) | ( n14525 & n16620 ) | ( ~n16619 & n16620 ) ;
  assign n16622 = n4993 ^ n3822 ^ n344 ;
  assign n16623 = n689 & ~n2028 ;
  assign n16624 = ~n14518 & n16623 ;
  assign n16625 = n15617 ^ n11811 ^ n253 ;
  assign n16628 = ( n2555 & ~n7847 ) | ( n2555 & n16025 ) | ( ~n7847 & n16025 ) ;
  assign n16626 = ( n3173 & ~n9637 ) | ( n3173 & n12729 ) | ( ~n9637 & n12729 ) ;
  assign n16627 = n7003 & n16626 ;
  assign n16629 = n16628 ^ n16627 ^ n2237 ;
  assign n16630 = n16584 ^ n12653 ^ 1'b0 ;
  assign n16631 = n11912 | n16630 ;
  assign n16632 = ( n2041 & n16534 ) | ( n2041 & ~n16631 ) | ( n16534 & ~n16631 ) ;
  assign n16633 = n16632 ^ n8904 ^ n2797 ;
  assign n16634 = ( x28 & n2670 ) | ( x28 & ~n7274 ) | ( n2670 & ~n7274 ) ;
  assign n16635 = n4251 ^ n2990 ^ 1'b0 ;
  assign n16636 = n16635 ^ n12158 ^ n6079 ;
  assign n16637 = ( n1416 & ~n16634 ) | ( n1416 & n16636 ) | ( ~n16634 & n16636 ) ;
  assign n16638 = ( n4529 & ~n5125 ) | ( n4529 & n9345 ) | ( ~n5125 & n9345 ) ;
  assign n16639 = ( n8909 & ~n12554 ) | ( n8909 & n16638 ) | ( ~n12554 & n16638 ) ;
  assign n16640 = ( n3731 & n6514 ) | ( n3731 & n9686 ) | ( n6514 & n9686 ) ;
  assign n16641 = ( n13220 & n15681 ) | ( n13220 & ~n16640 ) | ( n15681 & ~n16640 ) ;
  assign n16642 = ( n5473 & n7477 ) | ( n5473 & ~n7728 ) | ( n7477 & ~n7728 ) ;
  assign n16643 = n13531 | n16642 ;
  assign n16644 = n12158 ^ n8380 ^ 1'b0 ;
  assign n16645 = n16644 ^ n11217 ^ n754 ;
  assign n16646 = n5358 | n16645 ;
  assign n16649 = n9568 ^ n6742 ^ n4804 ;
  assign n16647 = n2716 | n3213 ;
  assign n16648 = ( n12633 & n12979 ) | ( n12633 & ~n16647 ) | ( n12979 & ~n16647 ) ;
  assign n16650 = n16649 ^ n16648 ^ 1'b0 ;
  assign n16651 = n12423 ^ n4133 ^ n3077 ;
  assign n16652 = ( ~n6914 & n7174 ) | ( ~n6914 & n16113 ) | ( n7174 & n16113 ) ;
  assign n16653 = n16651 & n16652 ;
  assign n16655 = n3243 & n3289 ;
  assign n16656 = n2335 & n16655 ;
  assign n16657 = n16656 ^ n10536 ^ n8330 ;
  assign n16654 = n6520 ^ n3586 ^ n1534 ;
  assign n16658 = n16657 ^ n16654 ^ 1'b0 ;
  assign n16659 = n1568 | n2036 ;
  assign n16660 = n16659 ^ n8730 ^ 1'b0 ;
  assign n16661 = n155 & n582 ;
  assign n16662 = n16660 & n16661 ;
  assign n16665 = n9841 & ~n16209 ;
  assign n16666 = n16665 ^ n11436 ^ 1'b0 ;
  assign n16663 = ( n1847 & ~n3518 ) | ( n1847 & n5641 ) | ( ~n3518 & n5641 ) ;
  assign n16664 = ( n8136 & n9854 ) | ( n8136 & n16663 ) | ( n9854 & n16663 ) ;
  assign n16667 = n16666 ^ n16664 ^ n3046 ;
  assign n16668 = ~n1688 & n4640 ;
  assign n16669 = n14152 ^ n2708 ^ 1'b0 ;
  assign n16670 = ~n7020 & n7817 ;
  assign n16671 = ~n16669 & n16670 ;
  assign n16672 = ( n13634 & ~n16363 ) | ( n13634 & n16671 ) | ( ~n16363 & n16671 ) ;
  assign n16673 = ( n6812 & n16668 ) | ( n6812 & n16672 ) | ( n16668 & n16672 ) ;
  assign n16676 = n11848 ^ n10579 ^ n3493 ;
  assign n16674 = ~n3931 & n7086 ;
  assign n16675 = n16674 ^ n8360 ^ 1'b0 ;
  assign n16677 = n16676 ^ n16675 ^ 1'b0 ;
  assign n16678 = ( n2602 & n7555 ) | ( n2602 & n9783 ) | ( n7555 & n9783 ) ;
  assign n16679 = n1664 & n8922 ;
  assign n16680 = ( n1076 & ~n8817 ) | ( n1076 & n16679 ) | ( ~n8817 & n16679 ) ;
  assign n16681 = ( n2758 & n10841 ) | ( n2758 & ~n16680 ) | ( n10841 & ~n16680 ) ;
  assign n16685 = n8106 ^ n6085 ^ n4951 ;
  assign n16686 = n16685 ^ n16066 ^ 1'b0 ;
  assign n16682 = n15029 ^ n13463 ^ n11410 ;
  assign n16683 = n16682 ^ n10865 ^ 1'b0 ;
  assign n16684 = n10610 & ~n16683 ;
  assign n16687 = n16686 ^ n16684 ^ n8006 ;
  assign n16688 = n4496 ^ n3236 ^ n881 ;
  assign n16689 = n2218 & ~n11654 ;
  assign n16690 = ~n16688 & n16689 ;
  assign n16693 = n4566 & n9854 ;
  assign n16694 = n16693 ^ n1244 ^ 1'b0 ;
  assign n16691 = ( n9160 & n11377 ) | ( n9160 & ~n14645 ) | ( n11377 & ~n14645 ) ;
  assign n16692 = ~n11454 & n16691 ;
  assign n16695 = n16694 ^ n16692 ^ 1'b0 ;
  assign n16696 = n5830 ^ n1542 ^ 1'b0 ;
  assign n16697 = ~n14359 & n16696 ;
  assign n16698 = n16697 ^ n15121 ^ n7889 ;
  assign n16699 = ( n6755 & n14262 ) | ( n6755 & ~n16290 ) | ( n14262 & ~n16290 ) ;
  assign n16700 = n7869 ^ n6148 ^ n1589 ;
  assign n16702 = ( n4707 & ~n5678 ) | ( n4707 & n8056 ) | ( ~n5678 & n8056 ) ;
  assign n16701 = ( n1813 & ~n6487 ) | ( n1813 & n7896 ) | ( ~n6487 & n7896 ) ;
  assign n16703 = n16702 ^ n16701 ^ n16684 ;
  assign n16704 = n7004 & n10385 ;
  assign n16705 = ( n6855 & n10390 ) | ( n6855 & n16704 ) | ( n10390 & n16704 ) ;
  assign n16706 = n14615 ^ n8599 ^ 1'b0 ;
  assign n16707 = n506 & ~n16706 ;
  assign n16714 = ~n2414 & n4781 ;
  assign n16715 = n8071 & n16714 ;
  assign n16708 = n2036 & ~n3519 ;
  assign n16711 = n14401 ^ n9298 ^ x86 ;
  assign n16709 = ( n5500 & ~n7022 ) | ( n5500 & n8949 ) | ( ~n7022 & n8949 ) ;
  assign n16710 = ~n12850 & n16709 ;
  assign n16712 = n16711 ^ n16710 ^ 1'b0 ;
  assign n16713 = n16708 | n16712 ;
  assign n16716 = n16715 ^ n16713 ^ n13294 ;
  assign n16717 = ( n1539 & n9863 ) | ( n1539 & n15355 ) | ( n9863 & n15355 ) ;
  assign n16718 = n16717 ^ n15909 ^ 1'b0 ;
  assign n16719 = n16619 ^ n5568 ^ x66 ;
  assign n16720 = ~n6852 & n16719 ;
  assign n16721 = n5246 ^ n4139 ^ n1576 ;
  assign n16722 = n2890 | n16721 ;
  assign n16723 = n10643 | n16722 ;
  assign n16724 = n16723 ^ n14712 ^ n10710 ;
  assign n16725 = n16724 ^ n9060 ^ 1'b0 ;
  assign n16726 = n3688 ^ n2864 ^ n2686 ;
  assign n16727 = ~n1448 & n16726 ;
  assign n16728 = n13196 & n16727 ;
  assign n16729 = ( x109 & n4810 ) | ( x109 & n9341 ) | ( n4810 & n9341 ) ;
  assign n16730 = ~n412 & n16729 ;
  assign n16731 = n6915 | n16730 ;
  assign n16732 = n6887 ^ n4535 ^ 1'b0 ;
  assign n16733 = n13562 ^ n11754 ^ n10863 ;
  assign n16734 = ( n16574 & ~n16732 ) | ( n16574 & n16733 ) | ( ~n16732 & n16733 ) ;
  assign n16735 = ( n3588 & ~n10948 ) | ( n3588 & n11810 ) | ( ~n10948 & n11810 ) ;
  assign n16736 = ~n2636 & n10635 ;
  assign n16737 = n16736 ^ n3092 ^ 1'b0 ;
  assign n16738 = n10299 & n10977 ;
  assign n16739 = n16737 & n16738 ;
  assign n16740 = n16739 ^ n2236 ^ n1299 ;
  assign n16742 = ( n933 & ~n3228 ) | ( n933 & n3734 ) | ( ~n3228 & n3734 ) ;
  assign n16741 = ~n8199 & n9408 ;
  assign n16743 = n16742 ^ n16741 ^ 1'b0 ;
  assign n16744 = n11722 | n16743 ;
  assign n16745 = ~n1946 & n5850 ;
  assign n16746 = n16745 ^ n4263 ^ n3846 ;
  assign n16747 = n7238 | n16746 ;
  assign n16748 = n7083 | n13252 ;
  assign n16749 = ( x49 & n16747 ) | ( x49 & ~n16748 ) | ( n16747 & ~n16748 ) ;
  assign n16750 = n16749 ^ n8168 ^ n3224 ;
  assign n16751 = ~n9451 & n9664 ;
  assign n16752 = n1054 & ~n16751 ;
  assign n16753 = n16752 ^ n15691 ^ 1'b0 ;
  assign n16754 = ( ~n6874 & n9931 ) | ( ~n6874 & n16306 ) | ( n9931 & n16306 ) ;
  assign n16755 = ( ~n7437 & n12005 ) | ( ~n7437 & n16754 ) | ( n12005 & n16754 ) ;
  assign n16756 = n11397 ^ n10162 ^ n516 ;
  assign n16757 = n15814 ^ n5268 ^ n2464 ;
  assign n16758 = ( n3136 & n4333 ) | ( n3136 & ~n6654 ) | ( n4333 & ~n6654 ) ;
  assign n16759 = n16758 ^ n10000 ^ n9564 ;
  assign n16760 = ( n374 & n1750 ) | ( n374 & ~n2478 ) | ( n1750 & ~n2478 ) ;
  assign n16761 = n16760 ^ n14559 ^ n9506 ;
  assign n16762 = n16610 ^ n6116 ^ 1'b0 ;
  assign n16763 = n1362 & ~n16762 ;
  assign n16764 = n16763 ^ n4674 ^ 1'b0 ;
  assign n16765 = ( n1477 & n2920 ) | ( n1477 & ~n7254 ) | ( n2920 & ~n7254 ) ;
  assign n16766 = n4294 | n16765 ;
  assign n16767 = n7950 & ~n16766 ;
  assign n16768 = n16767 ^ n3384 ^ n723 ;
  assign n16769 = n14858 & ~n16768 ;
  assign n16771 = ( ~n5153 & n6886 ) | ( ~n5153 & n8338 ) | ( n6886 & n8338 ) ;
  assign n16770 = x55 & ~n2579 ;
  assign n16772 = n16771 ^ n16770 ^ 1'b0 ;
  assign n16773 = n16772 ^ n13620 ^ n3688 ;
  assign n16774 = n4186 | n4969 ;
  assign n16779 = n11595 ^ n9665 ^ 1'b0 ;
  assign n16780 = n1086 & ~n16779 ;
  assign n16778 = ( n2348 & n3365 ) | ( n2348 & n8016 ) | ( n3365 & n8016 ) ;
  assign n16775 = n2629 ^ n746 ^ 1'b0 ;
  assign n16776 = n9514 | n16775 ;
  assign n16777 = n4782 | n16776 ;
  assign n16781 = n16780 ^ n16778 ^ n16777 ;
  assign n16785 = n4129 & n7826 ;
  assign n16786 = ~n4187 & n16785 ;
  assign n16782 = ( n818 & n3695 ) | ( n818 & ~n10481 ) | ( n3695 & ~n10481 ) ;
  assign n16783 = n16782 ^ n4423 ^ 1'b0 ;
  assign n16784 = ~n13481 & n16783 ;
  assign n16787 = n16786 ^ n16784 ^ n6662 ;
  assign n16788 = n10883 & ~n16787 ;
  assign n16789 = n13750 & n16788 ;
  assign n16790 = n6216 ^ n5295 ^ n2186 ;
  assign n16791 = n2725 | n16790 ;
  assign n16792 = n16791 ^ n8890 ^ n5111 ;
  assign n16793 = n9474 & n15352 ;
  assign n16794 = ~n16792 & n16793 ;
  assign n16795 = ~n6508 & n9372 ;
  assign n16796 = ~n11612 & n16795 ;
  assign n16797 = n16796 ^ n16167 ^ 1'b0 ;
  assign n16806 = ( ~n4868 & n10649 ) | ( ~n4868 & n11650 ) | ( n10649 & n11650 ) ;
  assign n16807 = n15173 ^ n8684 ^ 1'b0 ;
  assign n16808 = n16806 | n16807 ;
  assign n16800 = n5227 & n10489 ;
  assign n16801 = n3877 & n16800 ;
  assign n16802 = n2305 | n3787 ;
  assign n16803 = n16801 & ~n16802 ;
  assign n16798 = n265 | n850 ;
  assign n16799 = n16798 ^ n10929 ^ n10742 ;
  assign n16804 = n16803 ^ n16799 ^ n7896 ;
  assign n16805 = n3769 & ~n16804 ;
  assign n16809 = n16808 ^ n16805 ^ 1'b0 ;
  assign n16810 = ( ~n1762 & n7483 ) | ( ~n1762 & n9191 ) | ( n7483 & n9191 ) ;
  assign n16811 = n1735 & ~n16810 ;
  assign n16812 = n16811 ^ n9285 ^ 1'b0 ;
  assign n16813 = ( n7407 & n7918 ) | ( n7407 & n8495 ) | ( n7918 & n8495 ) ;
  assign n16814 = ( n3983 & n13847 ) | ( n3983 & ~n16813 ) | ( n13847 & ~n16813 ) ;
  assign n16815 = n16814 ^ n9912 ^ n6693 ;
  assign n16816 = n11661 ^ n2489 ^ n216 ;
  assign n16817 = n2372 | n4806 ;
  assign n16818 = n16817 ^ n12307 ^ n5603 ;
  assign n16819 = n16818 ^ n9972 ^ 1'b0 ;
  assign n16820 = n13558 & ~n16819 ;
  assign n16821 = n9286 & ~n13061 ;
  assign n16822 = n16821 ^ n11873 ^ 1'b0 ;
  assign n16823 = ( n1496 & n16820 ) | ( n1496 & n16822 ) | ( n16820 & n16822 ) ;
  assign n16824 = n16823 ^ n12549 ^ n11682 ;
  assign n16825 = ~n16816 & n16824 ;
  assign n16826 = ( n6241 & ~n6378 ) | ( n6241 & n6926 ) | ( ~n6378 & n6926 ) ;
  assign n16827 = ( n641 & n2004 ) | ( n641 & ~n2539 ) | ( n2004 & ~n2539 ) ;
  assign n16828 = n16827 ^ n472 ^ 1'b0 ;
  assign n16829 = n16826 | n16828 ;
  assign n16831 = ( ~n2201 & n5843 ) | ( ~n2201 & n6262 ) | ( n5843 & n6262 ) ;
  assign n16830 = n14517 ^ n4136 ^ n336 ;
  assign n16832 = n16831 ^ n16830 ^ n6781 ;
  assign n16835 = n758 & n4767 ;
  assign n16836 = n16835 ^ n12114 ^ n10002 ;
  assign n16833 = n10574 ^ n5854 ^ n4861 ;
  assign n16834 = x54 & n16833 ;
  assign n16837 = n16836 ^ n16834 ^ 1'b0 ;
  assign n16838 = ( n3286 & ~n6804 ) | ( n3286 & n15579 ) | ( ~n6804 & n15579 ) ;
  assign n16839 = n14120 ^ n12911 ^ n8782 ;
  assign n16840 = ( n2094 & ~n16838 ) | ( n2094 & n16839 ) | ( ~n16838 & n16839 ) ;
  assign n16841 = n3633 & n7887 ;
  assign n16842 = n11709 ^ n7176 ^ n761 ;
  assign n16843 = ( n295 & n16841 ) | ( n295 & ~n16842 ) | ( n16841 & ~n16842 ) ;
  assign n16844 = n1606 | n16843 ;
  assign n16845 = n16840 | n16844 ;
  assign n16846 = ( n2178 & ~n4225 ) | ( n2178 & n11369 ) | ( ~n4225 & n11369 ) ;
  assign n16847 = n11767 ^ n992 ^ 1'b0 ;
  assign n16848 = n16847 ^ n3803 ^ n1499 ;
  assign n16849 = ( n4291 & n7939 ) | ( n4291 & n10748 ) | ( n7939 & n10748 ) ;
  assign n16850 = n16849 ^ n16536 ^ n8148 ;
  assign n16851 = x43 & n4998 ;
  assign n16853 = n15381 ^ n8618 ^ n4759 ;
  assign n16852 = ( n6649 & ~n7968 ) | ( n6649 & n10291 ) | ( ~n7968 & n10291 ) ;
  assign n16854 = n16853 ^ n16852 ^ n4779 ;
  assign n16855 = ~n7230 & n13978 ;
  assign n16856 = n16855 ^ n3486 ^ 1'b0 ;
  assign n16857 = n10681 ^ n291 ^ 1'b0 ;
  assign n16858 = ( ~n5415 & n6172 ) | ( ~n5415 & n16857 ) | ( n6172 & n16857 ) ;
  assign n16859 = ( n1612 & n13011 ) | ( n1612 & ~n16858 ) | ( n13011 & ~n16858 ) ;
  assign n16860 = n16859 ^ n2091 ^ 1'b0 ;
  assign n16861 = ( n15233 & ~n16481 ) | ( n15233 & n16860 ) | ( ~n16481 & n16860 ) ;
  assign n16862 = n9153 ^ n2903 ^ n1847 ;
  assign n16863 = n16862 ^ n9468 ^ n668 ;
  assign n16864 = ( ~n8348 & n14417 ) | ( ~n8348 & n16863 ) | ( n14417 & n16863 ) ;
  assign n16865 = n9833 ^ n9348 ^ 1'b0 ;
  assign n16866 = n1333 & n16865 ;
  assign n16867 = n9465 ^ n3580 ^ 1'b0 ;
  assign n16868 = x79 & n16867 ;
  assign n16869 = ( n5909 & n15591 ) | ( n5909 & n16868 ) | ( n15591 & n16868 ) ;
  assign n16870 = n4372 ^ n3968 ^ n2468 ;
  assign n16871 = n16870 ^ n732 ^ 1'b0 ;
  assign n16872 = n10938 | n16871 ;
  assign n16873 = n237 & ~n4270 ;
  assign n16874 = n16873 ^ n7833 ^ 1'b0 ;
  assign n16875 = n16092 ^ n2367 ^ n1093 ;
  assign n16876 = ( n16872 & n16874 ) | ( n16872 & ~n16875 ) | ( n16874 & ~n16875 ) ;
  assign n16877 = ( ~n4714 & n12897 ) | ( ~n4714 & n16876 ) | ( n12897 & n16876 ) ;
  assign n16878 = n9159 ^ n5930 ^ n2948 ;
  assign n16879 = n4562 ^ n3249 ^ n2631 ;
  assign n16880 = ( n2043 & n12959 ) | ( n2043 & ~n14877 ) | ( n12959 & ~n14877 ) ;
  assign n16881 = n5250 ^ n2475 ^ n2379 ;
  assign n16882 = ( n7963 & n9347 ) | ( n7963 & ~n16881 ) | ( n9347 & ~n16881 ) ;
  assign n16885 = n11949 ^ n10589 ^ n4200 ;
  assign n16886 = ( ~n8438 & n13131 ) | ( ~n8438 & n16885 ) | ( n13131 & n16885 ) ;
  assign n16883 = n16382 ^ n5879 ^ n936 ;
  assign n16884 = n13615 & n16883 ;
  assign n16887 = n16886 ^ n16884 ^ 1'b0 ;
  assign n16888 = n4137 | n13734 ;
  assign n16889 = ( n6044 & n8174 ) | ( n6044 & ~n12509 ) | ( n8174 & ~n12509 ) ;
  assign n16890 = ( n14795 & n16888 ) | ( n14795 & ~n16889 ) | ( n16888 & ~n16889 ) ;
  assign n16891 = n16098 ^ n3268 ^ n2281 ;
  assign n16892 = ( n3927 & n4964 ) | ( n3927 & n10572 ) | ( n4964 & n10572 ) ;
  assign n16893 = n14498 ^ n14317 ^ n1865 ;
  assign n16894 = ( ~n1531 & n16892 ) | ( ~n1531 & n16893 ) | ( n16892 & n16893 ) ;
  assign n16895 = n8351 ^ n2117 ^ n1350 ;
  assign n16896 = ( n4678 & ~n8035 ) | ( n4678 & n13634 ) | ( ~n8035 & n13634 ) ;
  assign n16897 = n16896 ^ n9131 ^ n195 ;
  assign n16898 = n16897 ^ n5879 ^ n2214 ;
  assign n16899 = n11704 ^ n10694 ^ n2555 ;
  assign n16900 = ( n305 & n4743 ) | ( n305 & n8435 ) | ( n4743 & n8435 ) ;
  assign n16901 = ( ~n16898 & n16899 ) | ( ~n16898 & n16900 ) | ( n16899 & n16900 ) ;
  assign n16902 = ~n5464 & n8603 ;
  assign n16903 = n16902 ^ n4400 ^ 1'b0 ;
  assign n16904 = n9402 & n16903 ;
  assign n16905 = n16904 ^ n12076 ^ 1'b0 ;
  assign n16906 = ( ~n3680 & n9131 ) | ( ~n3680 & n15860 ) | ( n9131 & n15860 ) ;
  assign n16907 = ( n9951 & n11769 ) | ( n9951 & n16906 ) | ( n11769 & n16906 ) ;
  assign n16908 = ( n5295 & ~n15443 ) | ( n5295 & n16640 ) | ( ~n15443 & n16640 ) ;
  assign n16915 = n5351 & n10616 ;
  assign n16916 = n16915 ^ n3619 ^ 1'b0 ;
  assign n16917 = ( n8113 & n9627 ) | ( n8113 & n16916 ) | ( n9627 & n16916 ) ;
  assign n16912 = n13394 ^ n8649 ^ n3521 ;
  assign n16909 = n9202 ^ n5937 ^ n5329 ;
  assign n16910 = n4414 & ~n16909 ;
  assign n16911 = n12592 & n16910 ;
  assign n16913 = n16912 ^ n16911 ^ n2595 ;
  assign n16914 = n7736 & n16913 ;
  assign n16918 = n16917 ^ n16914 ^ 1'b0 ;
  assign n16919 = n4673 | n5411 ;
  assign n16920 = n3191 | n16919 ;
  assign n16921 = ( n2506 & ~n6508 ) | ( n2506 & n8161 ) | ( ~n6508 & n8161 ) ;
  assign n16922 = n16921 ^ n12740 ^ n1830 ;
  assign n16923 = n12316 | n12434 ;
  assign n16924 = n16923 ^ n9117 ^ 1'b0 ;
  assign n16925 = ( n9662 & n15295 ) | ( n9662 & n16924 ) | ( n15295 & n16924 ) ;
  assign n16928 = n9998 ^ n1776 ^ n1205 ;
  assign n16926 = ( ~n2346 & n3231 ) | ( ~n2346 & n6409 ) | ( n3231 & n6409 ) ;
  assign n16927 = ( ~n1174 & n8534 ) | ( ~n1174 & n16926 ) | ( n8534 & n16926 ) ;
  assign n16929 = n16928 ^ n16927 ^ n6966 ;
  assign n16930 = n4646 ^ n2774 ^ 1'b0 ;
  assign n16931 = x118 & ~n16930 ;
  assign n16932 = n13390 & n16931 ;
  assign n16933 = n8431 | n13731 ;
  assign n16934 = n1760 & ~n16193 ;
  assign n16938 = n7281 ^ n1324 ^ n730 ;
  assign n16936 = n7939 ^ n900 ^ 1'b0 ;
  assign n16937 = n5789 | n16936 ;
  assign n16939 = n16938 ^ n16937 ^ n10421 ;
  assign n16935 = n3842 & n7631 ;
  assign n16940 = n16939 ^ n16935 ^ 1'b0 ;
  assign n16941 = n9666 ^ n4496 ^ n2790 ;
  assign n16942 = n1580 & ~n16941 ;
  assign n16943 = ~n1218 & n7967 ;
  assign n16944 = n16943 ^ n748 ^ 1'b0 ;
  assign n16945 = n16944 ^ n16504 ^ 1'b0 ;
  assign n16946 = ~n16942 & n16945 ;
  assign n16947 = n8973 | n14082 ;
  assign n16948 = n10712 & ~n16947 ;
  assign n16949 = n16948 ^ n4648 ^ 1'b0 ;
  assign n16950 = n16949 ^ x63 ^ 1'b0 ;
  assign n16954 = n4559 ^ n3607 ^ n2568 ;
  assign n16955 = n16954 ^ n5120 ^ 1'b0 ;
  assign n16956 = ~n15775 & n16955 ;
  assign n16951 = n5289 ^ n4673 ^ 1'b0 ;
  assign n16952 = n16951 ^ n3225 ^ 1'b0 ;
  assign n16953 = ( n11538 & n14532 ) | ( n11538 & n16952 ) | ( n14532 & n16952 ) ;
  assign n16957 = n16956 ^ n16953 ^ n3656 ;
  assign n16958 = n3927 ^ n944 ^ n326 ;
  assign n16959 = n16958 ^ n4127 ^ n1464 ;
  assign n16960 = n16959 ^ n10189 ^ n9159 ;
  assign n16962 = n3976 & n6652 ;
  assign n16963 = n16962 ^ n6701 ^ 1'b0 ;
  assign n16961 = ( ~n4088 & n7863 ) | ( ~n4088 & n14819 ) | ( n7863 & n14819 ) ;
  assign n16964 = n16963 ^ n16961 ^ n4950 ;
  assign n16966 = n5022 & ~n16154 ;
  assign n16967 = n266 & n16966 ;
  assign n16965 = n469 | n15850 ;
  assign n16968 = n16967 ^ n16965 ^ 1'b0 ;
  assign n16969 = n1342 & ~n15683 ;
  assign n16970 = n16969 ^ n6793 ^ 1'b0 ;
  assign n16971 = n10255 & ~n16970 ;
  assign n16972 = n16971 ^ n12608 ^ 1'b0 ;
  assign n16973 = n15753 ^ n7202 ^ n782 ;
  assign n16974 = ( n4581 & n15685 ) | ( n4581 & n16438 ) | ( n15685 & n16438 ) ;
  assign n16975 = n12274 ^ n7529 ^ 1'b0 ;
  assign n16976 = n1437 & n15988 ;
  assign n16977 = ~n16975 & n16976 ;
  assign n16978 = n16977 ^ n8965 ^ n5126 ;
  assign n16979 = ( n1790 & ~n5323 ) | ( n1790 & n9913 ) | ( ~n5323 & n9913 ) ;
  assign n16980 = n14931 ^ n6364 ^ n2411 ;
  assign n16981 = ( ~n7806 & n16979 ) | ( ~n7806 & n16980 ) | ( n16979 & n16980 ) ;
  assign n16982 = ( n686 & ~n1352 ) | ( n686 & n6137 ) | ( ~n1352 & n6137 ) ;
  assign n16983 = ~n2255 & n2577 ;
  assign n16984 = ( n10264 & n16982 ) | ( n10264 & ~n16983 ) | ( n16982 & ~n16983 ) ;
  assign n16985 = ~n7942 & n12103 ;
  assign n16986 = n16985 ^ n3994 ^ 1'b0 ;
  assign n16987 = n14244 ^ n3787 ^ n2922 ;
  assign n16988 = ( ~n5259 & n8495 ) | ( ~n5259 & n14094 ) | ( n8495 & n14094 ) ;
  assign n16989 = ( n15099 & ~n16987 ) | ( n15099 & n16988 ) | ( ~n16987 & n16988 ) ;
  assign n16990 = n14033 ^ n8737 ^ 1'b0 ;
  assign n16991 = n4991 & ~n16990 ;
  assign n16992 = n16991 ^ n11995 ^ n1918 ;
  assign n16993 = n6221 ^ n4617 ^ 1'b0 ;
  assign n16994 = n16993 ^ n14055 ^ n11826 ;
  assign n16995 = n16994 ^ n14261 ^ n237 ;
  assign n16996 = n7041 & n16995 ;
  assign n16997 = n5223 ^ n238 ^ 1'b0 ;
  assign n16998 = n4480 & n16997 ;
  assign n16999 = n810 & ~n2103 ;
  assign n17000 = ~n16998 & n16999 ;
  assign n17001 = n17000 ^ n6696 ^ 1'b0 ;
  assign n17002 = n13138 ^ n5988 ^ n5459 ;
  assign n17003 = n17002 ^ n2157 ^ 1'b0 ;
  assign n17004 = ( ~n1578 & n4032 ) | ( ~n1578 & n9345 ) | ( n4032 & n9345 ) ;
  assign n17007 = ( n4508 & n7513 ) | ( n4508 & n8330 ) | ( n7513 & n8330 ) ;
  assign n17005 = n14795 ^ n5572 ^ n354 ;
  assign n17006 = n17005 ^ n12342 ^ n9743 ;
  assign n17008 = n17007 ^ n17006 ^ n12385 ;
  assign n17009 = ~n3762 & n6796 ;
  assign n17010 = n15694 ^ n11715 ^ n8993 ;
  assign n17011 = n4557 | n13383 ;
  assign n17012 = n17011 ^ n12633 ^ 1'b0 ;
  assign n17013 = n17012 ^ n12125 ^ 1'b0 ;
  assign n17014 = n17010 | n17013 ;
  assign n17017 = ( n441 & n3218 ) | ( n441 & n4370 ) | ( n3218 & n4370 ) ;
  assign n17015 = n11114 ^ n7303 ^ 1'b0 ;
  assign n17016 = ( n5851 & n12391 ) | ( n5851 & ~n17015 ) | ( n12391 & ~n17015 ) ;
  assign n17018 = n17017 ^ n17016 ^ n7692 ;
  assign n17019 = n11686 ^ n9839 ^ n5114 ;
  assign n17020 = n1504 & n11032 ;
  assign n17021 = n17020 ^ n13123 ^ n9335 ;
  assign n17027 = n1213 & ~n4835 ;
  assign n17028 = ( n3583 & ~n12599 ) | ( n3583 & n17027 ) | ( ~n12599 & n17027 ) ;
  assign n17022 = n9073 ^ n4299 ^ n1865 ;
  assign n17023 = n13734 | n17022 ;
  assign n17024 = n17023 ^ n2988 ^ 1'b0 ;
  assign n17025 = n17024 ^ n1940 ^ 1'b0 ;
  assign n17026 = n2971 & n17025 ;
  assign n17029 = n17028 ^ n17026 ^ n9322 ;
  assign n17030 = n17029 ^ n4216 ^ n1089 ;
  assign n17031 = x124 & ~n4430 ;
  assign n17032 = n17031 ^ n5047 ^ n3044 ;
  assign n17033 = n17032 ^ n985 ^ 1'b0 ;
  assign n17034 = n8355 ^ n8227 ^ 1'b0 ;
  assign n17035 = n17034 ^ n9290 ^ n6598 ;
  assign n17036 = n9110 | n11769 ;
  assign n17037 = n12473 | n17036 ;
  assign n17039 = ( n983 & n8651 ) | ( n983 & ~n16066 ) | ( n8651 & ~n16066 ) ;
  assign n17038 = n6667 & n12277 ;
  assign n17040 = n17039 ^ n17038 ^ 1'b0 ;
  assign n17041 = n13266 ^ n3466 ^ 1'b0 ;
  assign n17042 = ( n5494 & ~n11508 ) | ( n5494 & n17041 ) | ( ~n11508 & n17041 ) ;
  assign n17043 = n17042 ^ n16648 ^ n7817 ;
  assign n17044 = n15943 ^ n1625 ^ 1'b0 ;
  assign n17045 = n13929 & n17044 ;
  assign n17047 = ( n3710 & n4689 ) | ( n3710 & n7469 ) | ( n4689 & n7469 ) ;
  assign n17046 = n11370 ^ n6798 ^ n4689 ;
  assign n17048 = n17047 ^ n17046 ^ 1'b0 ;
  assign n17050 = n4083 & n11856 ;
  assign n17051 = n17050 ^ n7173 ^ n4407 ;
  assign n17049 = n10404 ^ n4569 ^ n1642 ;
  assign n17052 = n17051 ^ n17049 ^ 1'b0 ;
  assign n17053 = n17048 & ~n17052 ;
  assign n17054 = n8750 ^ n7810 ^ n6275 ;
  assign n17055 = n17054 ^ n14349 ^ n8120 ;
  assign n17056 = ( n8870 & ~n11122 ) | ( n8870 & n15844 ) | ( ~n11122 & n15844 ) ;
  assign n17059 = n12112 ^ n2668 ^ 1'b0 ;
  assign n17060 = ~n3839 & n17059 ;
  assign n17061 = n17060 ^ n9298 ^ 1'b0 ;
  assign n17058 = ( n2434 & ~n2737 ) | ( n2434 & n14890 ) | ( ~n2737 & n14890 ) ;
  assign n17057 = n13537 ^ n8039 ^ n6553 ;
  assign n17062 = n17061 ^ n17058 ^ n17057 ;
  assign n17063 = ( ~x45 & n2673 ) | ( ~x45 & n4445 ) | ( n2673 & n4445 ) ;
  assign n17064 = n15120 & ~n17063 ;
  assign n17065 = n8287 ^ n2734 ^ 1'b0 ;
  assign n17066 = n17065 ^ n8662 ^ n1656 ;
  assign n17067 = n16553 ^ n2448 ^ 1'b0 ;
  assign n17068 = n2175 & ~n2766 ;
  assign n17069 = n17068 ^ n5299 ^ 1'b0 ;
  assign n17070 = ( n2304 & n2792 ) | ( n2304 & ~n7408 ) | ( n2792 & ~n7408 ) ;
  assign n17071 = ( x72 & n2740 ) | ( x72 & n17070 ) | ( n2740 & n17070 ) ;
  assign n17072 = ( n2461 & n8006 ) | ( n2461 & ~n17071 ) | ( n8006 & ~n17071 ) ;
  assign n17073 = ( ~n11975 & n17069 ) | ( ~n11975 & n17072 ) | ( n17069 & n17072 ) ;
  assign n17074 = ( n2729 & ~n10182 ) | ( n2729 & n11372 ) | ( ~n10182 & n11372 ) ;
  assign n17075 = ~n15410 & n17074 ;
  assign n17076 = ~n3263 & n17075 ;
  assign n17077 = ( n1194 & ~n2481 ) | ( n1194 & n4831 ) | ( ~n2481 & n4831 ) ;
  assign n17078 = n17077 ^ n1035 ^ 1'b0 ;
  assign n17079 = n17078 ^ n15412 ^ n10788 ;
  assign n17080 = n4183 ^ n4162 ^ n2258 ;
  assign n17081 = n2800 ^ n1181 ^ n323 ;
  assign n17082 = ( x5 & n12453 ) | ( x5 & n17081 ) | ( n12453 & n17081 ) ;
  assign n17083 = ( ~n5859 & n17080 ) | ( ~n5859 & n17082 ) | ( n17080 & n17082 ) ;
  assign n17084 = ~n5677 & n16133 ;
  assign n17085 = x23 & n8303 ;
  assign n17086 = ( n1944 & ~n7375 ) | ( n1944 & n17085 ) | ( ~n7375 & n17085 ) ;
  assign n17087 = ( n2314 & ~n17084 ) | ( n2314 & n17086 ) | ( ~n17084 & n17086 ) ;
  assign n17088 = ( n5843 & n9876 ) | ( n5843 & n14617 ) | ( n9876 & n14617 ) ;
  assign n17089 = n7351 ^ n6989 ^ n4514 ;
  assign n17090 = n753 ^ n646 ^ 1'b0 ;
  assign n17091 = ( n1607 & n13822 ) | ( n1607 & ~n17090 ) | ( n13822 & ~n17090 ) ;
  assign n17092 = n17091 ^ n7503 ^ n2285 ;
  assign n17093 = n3134 | n3310 ;
  assign n17094 = n17093 ^ n1658 ^ 1'b0 ;
  assign n17095 = ( n719 & n6158 ) | ( n719 & n8158 ) | ( n6158 & n8158 ) ;
  assign n17096 = n8354 & ~n9457 ;
  assign n17097 = ( n17094 & n17095 ) | ( n17094 & n17096 ) | ( n17095 & n17096 ) ;
  assign n17098 = n2511 | n2662 ;
  assign n17099 = n15821 & ~n17098 ;
  assign n17100 = n17099 ^ n8836 ^ n6158 ;
  assign n17101 = n6598 & n12860 ;
  assign n17102 = n17100 & n17101 ;
  assign n17103 = ( n1896 & n11382 ) | ( n1896 & ~n12980 ) | ( n11382 & ~n12980 ) ;
  assign n17104 = n15406 ^ n10334 ^ 1'b0 ;
  assign n17105 = ( n2948 & ~n7070 ) | ( n2948 & n8634 ) | ( ~n7070 & n8634 ) ;
  assign n17106 = ( n970 & n10481 ) | ( n970 & n17105 ) | ( n10481 & n17105 ) ;
  assign n17107 = ( n1114 & n15084 ) | ( n1114 & ~n15322 ) | ( n15084 & ~n15322 ) ;
  assign n17108 = n15242 ^ n5818 ^ 1'b0 ;
  assign n17109 = n17108 ^ n7327 ^ 1'b0 ;
  assign n17110 = n17107 | n17109 ;
  assign n17111 = n17110 ^ n16107 ^ n4205 ;
  assign n17112 = n10069 ^ n3754 ^ 1'b0 ;
  assign n17113 = n16365 | n17112 ;
  assign n17114 = n6368 ^ n4940 ^ n1950 ;
  assign n17115 = n17114 ^ n13252 ^ n5550 ;
  assign n17116 = n4452 & n17115 ;
  assign n17117 = n17116 ^ n16681 ^ 1'b0 ;
  assign n17118 = n15331 ^ n4261 ^ n1908 ;
  assign n17119 = n17118 ^ n8866 ^ n1182 ;
  assign n17120 = ~n961 & n7343 ;
  assign n17121 = n17120 ^ n11568 ^ n4804 ;
  assign n17122 = ( ~n153 & n732 ) | ( ~n153 & n17121 ) | ( n732 & n17121 ) ;
  assign n17123 = ( n3186 & n8871 ) | ( n3186 & ~n17122 ) | ( n8871 & ~n17122 ) ;
  assign n17124 = ( n1300 & n10738 ) | ( n1300 & ~n17123 ) | ( n10738 & ~n17123 ) ;
  assign n17125 = n16411 ^ n13217 ^ n3305 ;
  assign n17127 = n15908 ^ n6203 ^ n1518 ;
  assign n17128 = n1475 & ~n9351 ;
  assign n17129 = ~n17127 & n17128 ;
  assign n17126 = ( n2588 & ~n10266 ) | ( n2588 & n15019 ) | ( ~n10266 & n15019 ) ;
  assign n17130 = n17129 ^ n17126 ^ n5982 ;
  assign n17131 = n16685 ^ n15100 ^ n3307 ;
  assign n17132 = n9341 ^ n7973 ^ n5127 ;
  assign n17133 = ( n7411 & n14300 ) | ( n7411 & ~n17132 ) | ( n14300 & ~n17132 ) ;
  assign n17134 = ( n3081 & n17131 ) | ( n3081 & ~n17133 ) | ( n17131 & ~n17133 ) ;
  assign n17135 = ( n8225 & n17130 ) | ( n8225 & n17134 ) | ( n17130 & n17134 ) ;
  assign n17143 = ( n970 & ~n1962 ) | ( n970 & n6510 ) | ( ~n1962 & n6510 ) ;
  assign n17144 = n6827 & n10489 ;
  assign n17145 = ( n3555 & n17143 ) | ( n3555 & ~n17144 ) | ( n17143 & ~n17144 ) ;
  assign n17139 = ( n2172 & ~n5024 ) | ( n2172 & n6553 ) | ( ~n5024 & n6553 ) ;
  assign n17140 = n17139 ^ n8469 ^ n5209 ;
  assign n17136 = n15174 ^ n8092 ^ n640 ;
  assign n17137 = ( ~n2307 & n8004 ) | ( ~n2307 & n17136 ) | ( n8004 & n17136 ) ;
  assign n17138 = n17137 ^ n3516 ^ n1669 ;
  assign n17141 = n17140 ^ n17138 ^ n4486 ;
  assign n17142 = n17141 ^ n15026 ^ n6018 ;
  assign n17146 = n17145 ^ n17142 ^ n7963 ;
  assign n17149 = ( n1806 & ~n2670 ) | ( n1806 & n9712 ) | ( ~n2670 & n9712 ) ;
  assign n17147 = ~n1187 & n1664 ;
  assign n17148 = n1329 | n17147 ;
  assign n17150 = n17149 ^ n17148 ^ 1'b0 ;
  assign n17151 = n17150 ^ n8176 ^ 1'b0 ;
  assign n17152 = n4544 & n14743 ;
  assign n17153 = n15175 & n17152 ;
  assign n17154 = n3646 & ~n17153 ;
  assign n17155 = n17154 ^ n14871 ^ n6580 ;
  assign n17156 = n3885 ^ n2698 ^ n2028 ;
  assign n17157 = ( ~n1642 & n2974 ) | ( ~n1642 & n12864 ) | ( n2974 & n12864 ) ;
  assign n17158 = n17156 & ~n17157 ;
  assign n17159 = n9412 | n17158 ;
  assign n17160 = n17159 ^ n8591 ^ 1'b0 ;
  assign n17161 = ( ~n7981 & n8111 ) | ( ~n7981 & n14047 ) | ( n8111 & n14047 ) ;
  assign n17162 = ( n2237 & n13326 ) | ( n2237 & ~n15097 ) | ( n13326 & ~n15097 ) ;
  assign n17163 = ( n4369 & ~n10314 ) | ( n4369 & n17162 ) | ( ~n10314 & n17162 ) ;
  assign n17164 = n4351 & ~n14882 ;
  assign n17165 = ~n16040 & n17164 ;
  assign n17166 = n1413 & n16814 ;
  assign n17167 = n17166 ^ n3651 ^ 1'b0 ;
  assign n17168 = n12908 | n17167 ;
  assign n17169 = n17165 & ~n17168 ;
  assign n17170 = ( n10858 & n17163 ) | ( n10858 & ~n17169 ) | ( n17163 & ~n17169 ) ;
  assign n17171 = n1435 | n9283 ;
  assign n17172 = n450 | n17171 ;
  assign n17177 = ( n2179 & n3858 ) | ( n2179 & ~n4730 ) | ( n3858 & ~n4730 ) ;
  assign n17173 = ( n254 & n8175 ) | ( n254 & ~n14890 ) | ( n8175 & ~n14890 ) ;
  assign n17174 = n17173 ^ n11892 ^ n2164 ;
  assign n17175 = n5101 & ~n17174 ;
  assign n17176 = n17175 ^ n13708 ^ 1'b0 ;
  assign n17178 = n17177 ^ n17176 ^ 1'b0 ;
  assign n17179 = n10479 | n17178 ;
  assign n17180 = n2039 ^ n1135 ^ 1'b0 ;
  assign n17181 = n1058 & ~n17180 ;
  assign n17182 = n17181 ^ n4541 ^ 1'b0 ;
  assign n17183 = ( n130 & ~n454 ) | ( n130 & n17182 ) | ( ~n454 & n17182 ) ;
  assign n17184 = n14745 ^ n8655 ^ 1'b0 ;
  assign n17185 = ( n4384 & n14940 ) | ( n4384 & n17184 ) | ( n14940 & n17184 ) ;
  assign n17186 = n3094 & n5638 ;
  assign n17187 = n17186 ^ n5774 ^ 1'b0 ;
  assign n17188 = n17187 ^ n11189 ^ n3769 ;
  assign n17190 = n4134 | n8722 ;
  assign n17191 = n2530 & ~n17190 ;
  assign n17189 = n2595 & ~n9331 ;
  assign n17192 = n17191 ^ n17189 ^ 1'b0 ;
  assign n17193 = n11601 ^ n9057 ^ n5319 ;
  assign n17194 = n17193 ^ n8449 ^ 1'b0 ;
  assign n17195 = n15569 ^ n14324 ^ 1'b0 ;
  assign n17196 = ( n5246 & n17194 ) | ( n5246 & n17195 ) | ( n17194 & n17195 ) ;
  assign n17197 = n511 & n15825 ;
  assign n17198 = x126 & n3190 ;
  assign n17199 = n17198 ^ n4677 ^ 1'b0 ;
  assign n17200 = n17199 ^ n7418 ^ n2989 ;
  assign n17201 = n17200 ^ n2137 ^ 1'b0 ;
  assign n17202 = n17197 & n17201 ;
  assign n17203 = n17202 ^ n10256 ^ n8069 ;
  assign n17204 = ( ~n683 & n3382 ) | ( ~n683 & n6443 ) | ( n3382 & n6443 ) ;
  assign n17205 = n17204 ^ n3854 ^ n1024 ;
  assign n17215 = n2279 & ~n10982 ;
  assign n17216 = n17215 ^ n7826 ^ 1'b0 ;
  assign n17214 = x24 & n3748 ;
  assign n17217 = n17216 ^ n17214 ^ 1'b0 ;
  assign n17218 = ( n2326 & n3035 ) | ( n2326 & n17217 ) | ( n3035 & n17217 ) ;
  assign n17219 = n12060 ^ n3911 ^ n1791 ;
  assign n17220 = ( n10847 & n17218 ) | ( n10847 & n17219 ) | ( n17218 & n17219 ) ;
  assign n17221 = n5215 & ~n8521 ;
  assign n17222 = ~n17220 & n17221 ;
  assign n17206 = n3088 ^ n1822 ^ 1'b0 ;
  assign n17207 = ~n244 & n17206 ;
  assign n17208 = n17207 ^ n5098 ^ n1896 ;
  assign n17209 = n17208 ^ n4624 ^ n3553 ;
  assign n17210 = n17209 ^ n6076 ^ 1'b0 ;
  assign n17211 = n16098 & ~n17210 ;
  assign n17212 = ( n2708 & n3531 ) | ( n2708 & n7308 ) | ( n3531 & n7308 ) ;
  assign n17213 = ( ~n8089 & n17211 ) | ( ~n8089 & n17212 ) | ( n17211 & n17212 ) ;
  assign n17223 = n17222 ^ n17213 ^ n885 ;
  assign n17224 = ( n343 & n6813 ) | ( n343 & n10394 ) | ( n6813 & n10394 ) ;
  assign n17225 = ( n14178 & n16094 ) | ( n14178 & n17224 ) | ( n16094 & n17224 ) ;
  assign n17226 = n16135 ^ n11465 ^ 1'b0 ;
  assign n17227 = n6356 | n17226 ;
  assign n17228 = n17227 ^ n13271 ^ 1'b0 ;
  assign n17233 = ( n1825 & ~n3987 ) | ( n1825 & n6033 ) | ( ~n3987 & n6033 ) ;
  assign n17234 = ( n1942 & ~n4304 ) | ( n1942 & n8573 ) | ( ~n4304 & n8573 ) ;
  assign n17235 = x69 & ~n8429 ;
  assign n17236 = ( n4042 & n17234 ) | ( n4042 & n17235 ) | ( n17234 & n17235 ) ;
  assign n17237 = ( ~n820 & n17233 ) | ( ~n820 & n17236 ) | ( n17233 & n17236 ) ;
  assign n17238 = ( n5429 & ~n14108 ) | ( n5429 & n17237 ) | ( ~n14108 & n17237 ) ;
  assign n17229 = ( n1688 & ~n6983 ) | ( n1688 & n14093 ) | ( ~n6983 & n14093 ) ;
  assign n17230 = ( n1525 & ~n3784 ) | ( n1525 & n14429 ) | ( ~n3784 & n14429 ) ;
  assign n17231 = n17230 ^ n13931 ^ n11380 ;
  assign n17232 = ( n9051 & ~n17229 ) | ( n9051 & n17231 ) | ( ~n17229 & n17231 ) ;
  assign n17239 = n17238 ^ n17232 ^ n573 ;
  assign n17240 = n14092 ^ n8157 ^ n8069 ;
  assign n17241 = ( n2297 & n9547 ) | ( n2297 & n17240 ) | ( n9547 & n17240 ) ;
  assign n17246 = ( ~n859 & n8056 ) | ( ~n859 & n13700 ) | ( n8056 & n13700 ) ;
  assign n17245 = n12233 & ~n17022 ;
  assign n17242 = n3810 ^ n924 ^ 1'b0 ;
  assign n17243 = n17242 ^ n5571 ^ n4196 ;
  assign n17244 = n17243 ^ n11845 ^ n7864 ;
  assign n17247 = n17246 ^ n17245 ^ n17244 ;
  assign n17248 = n3750 ^ n1983 ^ 1'b0 ;
  assign n17249 = ( n1647 & ~n2800 ) | ( n1647 & n6203 ) | ( ~n2800 & n6203 ) ;
  assign n17250 = n17249 ^ n16085 ^ n10552 ;
  assign n17251 = n17248 | n17250 ;
  assign n17252 = ( n10876 & n14645 ) | ( n10876 & n16636 ) | ( n14645 & n16636 ) ;
  assign n17253 = n17252 ^ n14599 ^ n10233 ;
  assign n17254 = ~n2883 & n14087 ;
  assign n17255 = n11808 & n17254 ;
  assign n17256 = ( n5171 & n12727 ) | ( n5171 & ~n14920 ) | ( n12727 & ~n14920 ) ;
  assign n17257 = ( n10062 & ~n13555 ) | ( n10062 & n17256 ) | ( ~n13555 & n17256 ) ;
  assign n17258 = n16209 ^ n8847 ^ n8726 ;
  assign n17259 = ( n536 & ~n4036 ) | ( n536 & n16573 ) | ( ~n4036 & n16573 ) ;
  assign n17260 = ( n5451 & n7372 ) | ( n5451 & ~n17259 ) | ( n7372 & ~n17259 ) ;
  assign n17261 = ( n1306 & n3689 ) | ( n1306 & n17260 ) | ( n3689 & n17260 ) ;
  assign n17262 = n14487 ^ n3101 ^ 1'b0 ;
  assign n17263 = ( n2040 & ~n2478 ) | ( n2040 & n3754 ) | ( ~n2478 & n3754 ) ;
  assign n17264 = n8339 ^ n4881 ^ n3087 ;
  assign n17265 = ( n2238 & n17263 ) | ( n2238 & n17264 ) | ( n17263 & n17264 ) ;
  assign n17266 = ( n17261 & n17262 ) | ( n17261 & ~n17265 ) | ( n17262 & ~n17265 ) ;
  assign n17267 = ( n2255 & n8326 ) | ( n2255 & ~n15072 ) | ( n8326 & ~n15072 ) ;
  assign n17268 = n17267 ^ n6658 ^ n1701 ;
  assign n17269 = ( ~n10217 & n11322 ) | ( ~n10217 & n16697 ) | ( n11322 & n16697 ) ;
  assign n17272 = n9767 ^ n3049 ^ 1'b0 ;
  assign n17273 = n1411 & n17272 ;
  assign n17270 = n8020 & n9929 ;
  assign n17271 = n17270 ^ n7851 ^ 1'b0 ;
  assign n17274 = n17273 ^ n17271 ^ n13801 ;
  assign n17275 = ( n8737 & n9202 ) | ( n8737 & ~n10907 ) | ( n9202 & ~n10907 ) ;
  assign n17276 = ~n1446 & n17275 ;
  assign n17277 = n8986 ^ n5211 ^ x21 ;
  assign n17278 = n17277 ^ n12609 ^ n12480 ;
  assign n17279 = n7085 & ~n17278 ;
  assign n17280 = ~n15965 & n17279 ;
  assign n17281 = n16094 ^ n13550 ^ n10505 ;
  assign n17282 = ( ~n6499 & n7901 ) | ( ~n6499 & n17281 ) | ( n7901 & n17281 ) ;
  assign n17283 = n9336 ^ n6514 ^ 1'b0 ;
  assign n17284 = ( n3782 & n9824 ) | ( n3782 & n9850 ) | ( n9824 & n9850 ) ;
  assign n17285 = n17284 ^ n16789 ^ n9777 ;
  assign n17286 = n15768 ^ n14487 ^ 1'b0 ;
  assign n17287 = ~n4685 & n17286 ;
  assign n17288 = n6745 & n17287 ;
  assign n17289 = ( n4730 & ~n10309 ) | ( n4730 & n17288 ) | ( ~n10309 & n17288 ) ;
  assign n17290 = n9159 ^ n6008 ^ 1'b0 ;
  assign n17291 = n7518 ^ n6977 ^ 1'b0 ;
  assign n17292 = n9375 & ~n17291 ;
  assign n17293 = n17292 ^ n11426 ^ 1'b0 ;
  assign n17298 = n14860 ^ n7792 ^ n4899 ;
  assign n17294 = n3359 ^ n2092 ^ 1'b0 ;
  assign n17295 = ~n5092 & n17294 ;
  assign n17296 = ~n14416 & n17295 ;
  assign n17297 = n6573 & n17296 ;
  assign n17299 = n17298 ^ n17297 ^ n1755 ;
  assign n17300 = n8418 ^ n7091 ^ n2572 ;
  assign n17301 = n17300 ^ n3748 ^ 1'b0 ;
  assign n17302 = ( ~n1707 & n5648 ) | ( ~n1707 & n17301 ) | ( n5648 & n17301 ) ;
  assign n17303 = n17302 ^ n1470 ^ 1'b0 ;
  assign n17304 = ( ~n11398 & n13355 ) | ( ~n11398 & n17303 ) | ( n13355 & n17303 ) ;
  assign n17305 = ( n5808 & n9187 ) | ( n5808 & n12630 ) | ( n9187 & n12630 ) ;
  assign n17306 = ( n13544 & ~n14244 ) | ( n13544 & n17305 ) | ( ~n14244 & n17305 ) ;
  assign n17307 = n17306 ^ n17010 ^ 1'b0 ;
  assign n17311 = n6606 & ~n11549 ;
  assign n17308 = n3283 & ~n12752 ;
  assign n17309 = ( n182 & n2074 ) | ( n182 & n17308 ) | ( n2074 & n17308 ) ;
  assign n17310 = ( n7263 & n9903 ) | ( n7263 & ~n17309 ) | ( n9903 & ~n17309 ) ;
  assign n17312 = n17311 ^ n17310 ^ n4277 ;
  assign n17313 = ( n5063 & n15348 ) | ( n5063 & n17312 ) | ( n15348 & n17312 ) ;
  assign n17314 = n2352 | n17313 ;
  assign n17315 = n16090 & ~n17314 ;
  assign n17316 = ~n3066 & n6406 ;
  assign n17317 = n17316 ^ n12206 ^ 1'b0 ;
  assign n17318 = n3652 | n17317 ;
  assign n17319 = n4222 & ~n17318 ;
  assign n17320 = ~x123 & n17319 ;
  assign n17321 = n6113 ^ n6102 ^ n4494 ;
  assign n17322 = ( n2163 & n6029 ) | ( n2163 & n17321 ) | ( n6029 & n17321 ) ;
  assign n17323 = n6616 & ~n17322 ;
  assign n17324 = ( n9413 & n10612 ) | ( n9413 & n17323 ) | ( n10612 & n17323 ) ;
  assign n17325 = n516 & ~n5088 ;
  assign n17326 = ( ~n6447 & n7805 ) | ( ~n6447 & n14364 ) | ( n7805 & n14364 ) ;
  assign n17327 = ( ~n2270 & n17325 ) | ( ~n2270 & n17326 ) | ( n17325 & n17326 ) ;
  assign n17329 = n5446 ^ n2199 ^ n1745 ;
  assign n17330 = n17329 ^ n6360 ^ n936 ;
  assign n17328 = n11707 ^ n5803 ^ n5183 ;
  assign n17331 = n17330 ^ n17328 ^ n1007 ;
  assign n17332 = n3704 & ~n4581 ;
  assign n17333 = ( n1876 & n2076 ) | ( n1876 & ~n13242 ) | ( n2076 & ~n13242 ) ;
  assign n17334 = ( ~n5700 & n17332 ) | ( ~n5700 & n17333 ) | ( n17332 & n17333 ) ;
  assign n17335 = ( ~n1965 & n14634 ) | ( ~n1965 & n17334 ) | ( n14634 & n17334 ) ;
  assign n17336 = n12389 ^ n2008 ^ x97 ;
  assign n17337 = ( n7324 & n12493 ) | ( n7324 & ~n17336 ) | ( n12493 & ~n17336 ) ;
  assign n17338 = n17337 ^ n2603 ^ 1'b0 ;
  assign n17339 = n8597 | n17338 ;
  assign n17340 = ( n9227 & ~n9286 ) | ( n9227 & n16958 ) | ( ~n9286 & n16958 ) ;
  assign n17341 = n1171 ^ n252 ^ 1'b0 ;
  assign n17342 = ( n5876 & n7349 ) | ( n5876 & ~n17341 ) | ( n7349 & ~n17341 ) ;
  assign n17343 = n2854 & n14085 ;
  assign n17344 = ( n752 & n7248 ) | ( n752 & n11467 ) | ( n7248 & n11467 ) ;
  assign n17345 = n8825 & n11778 ;
  assign n17346 = ~n10562 & n17345 ;
  assign n17347 = n15511 ^ n12464 ^ 1'b0 ;
  assign n17348 = n15009 | n17347 ;
  assign n17355 = n15013 ^ n3200 ^ n2439 ;
  assign n17354 = n15281 ^ n8383 ^ n4249 ;
  assign n17349 = ~n4795 & n5221 ;
  assign n17350 = n10564 & n17349 ;
  assign n17351 = n6374 ^ n5566 ^ 1'b0 ;
  assign n17352 = ~n17350 & n17351 ;
  assign n17353 = n17352 ^ n8743 ^ 1'b0 ;
  assign n17356 = n17355 ^ n17354 ^ n17353 ;
  assign n17357 = ( x49 & n437 ) | ( x49 & ~n5342 ) | ( n437 & ~n5342 ) ;
  assign n17358 = ( n1424 & n1726 ) | ( n1424 & n17357 ) | ( n1726 & n17357 ) ;
  assign n17359 = n8896 ^ n7325 ^ n6762 ;
  assign n17360 = n7292 & ~n17359 ;
  assign n17362 = ( n1457 & ~n2990 ) | ( n1457 & n11844 ) | ( ~n2990 & n11844 ) ;
  assign n17363 = n5866 & n17362 ;
  assign n17361 = n14337 ^ n11132 ^ n5382 ;
  assign n17364 = n17363 ^ n17361 ^ n4011 ;
  assign n17365 = n17364 ^ n13028 ^ 1'b0 ;
  assign n17366 = n4663 | n8703 ;
  assign n17367 = n17366 ^ n14114 ^ 1'b0 ;
  assign n17368 = n17365 | n17367 ;
  assign n17369 = n17368 ^ n7379 ^ n6299 ;
  assign n17370 = n15761 ^ n15687 ^ n12384 ;
  assign n17372 = ( n924 & n6848 ) | ( n924 & ~n8839 ) | ( n6848 & ~n8839 ) ;
  assign n17371 = n12238 ^ n7283 ^ n2074 ;
  assign n17373 = n17372 ^ n17371 ^ n4729 ;
  assign n17378 = n10952 ^ n7987 ^ n4641 ;
  assign n17374 = n12240 ^ n5316 ^ n2532 ;
  assign n17375 = n14539 ^ n7289 ^ 1'b0 ;
  assign n17376 = ~n17374 & n17375 ;
  assign n17377 = n11145 & n17376 ;
  assign n17379 = n17378 ^ n17377 ^ 1'b0 ;
  assign n17380 = ( n3473 & n17373 ) | ( n3473 & n17379 ) | ( n17373 & n17379 ) ;
  assign n17381 = ( n1331 & n2348 ) | ( n1331 & n17303 ) | ( n2348 & n17303 ) ;
  assign n17382 = n676 | n9735 ;
  assign n17383 = n17382 ^ n15448 ^ n6931 ;
  assign n17384 = ( n5517 & n9351 ) | ( n5517 & ~n17383 ) | ( n9351 & ~n17383 ) ;
  assign n17385 = n14541 ^ n12297 ^ n12293 ;
  assign n17391 = n6020 ^ n2540 ^ 1'b0 ;
  assign n17392 = n1848 & ~n7772 ;
  assign n17393 = n17391 & n17392 ;
  assign n17389 = n3363 & ~n6992 ;
  assign n17390 = n17389 ^ n9756 ^ 1'b0 ;
  assign n17386 = x52 & ~n9153 ;
  assign n17387 = n8815 & ~n14755 ;
  assign n17388 = ~n17386 & n17387 ;
  assign n17394 = n17393 ^ n17390 ^ n17388 ;
  assign n17396 = ~n1932 & n3409 ;
  assign n17397 = n6076 ^ n2621 ^ 1'b0 ;
  assign n17398 = n17396 & n17397 ;
  assign n17395 = n3801 & ~n9082 ;
  assign n17399 = n17398 ^ n17395 ^ n3649 ;
  assign n17400 = ~n1318 & n10877 ;
  assign n17401 = n17400 ^ n631 ^ 1'b0 ;
  assign n17402 = n17401 ^ n3287 ^ n452 ;
  assign n17403 = ( n1064 & n2539 ) | ( n1064 & n8237 ) | ( n2539 & n8237 ) ;
  assign n17404 = ( ~n14978 & n15355 ) | ( ~n14978 & n17403 ) | ( n15355 & n17403 ) ;
  assign n17405 = n9501 & n17404 ;
  assign n17409 = ( ~n4541 & n7233 ) | ( ~n4541 & n9792 ) | ( n7233 & n9792 ) ;
  assign n17410 = n13084 ^ n7481 ^ n4251 ;
  assign n17411 = n11019 ^ n6228 ^ n4959 ;
  assign n17412 = n17411 ^ n12843 ^ n3318 ;
  assign n17413 = ( n17409 & ~n17410 ) | ( n17409 & n17412 ) | ( ~n17410 & n17412 ) ;
  assign n17408 = n9053 ^ n4619 ^ n1298 ;
  assign n17406 = n10507 | n14810 ;
  assign n17407 = n17406 ^ n3838 ^ n2936 ;
  assign n17414 = n17413 ^ n17408 ^ n17407 ;
  assign n17415 = n14460 | n17414 ;
  assign n17416 = n17405 & ~n17415 ;
  assign n17419 = n8113 ^ n1319 ^ n333 ;
  assign n17417 = n2432 | n12534 ;
  assign n17418 = ( ~n538 & n686 ) | ( ~n538 & n17417 ) | ( n686 & n17417 ) ;
  assign n17420 = n17419 ^ n17418 ^ n13976 ;
  assign n17421 = ( ~n5686 & n17416 ) | ( ~n5686 & n17420 ) | ( n17416 & n17420 ) ;
  assign n17422 = x13 & ~n5389 ;
  assign n17423 = ~n5250 & n17422 ;
  assign n17424 = n2131 & ~n17423 ;
  assign n17425 = n17424 ^ n4945 ^ 1'b0 ;
  assign n17426 = n6391 ^ n2882 ^ 1'b0 ;
  assign n17427 = ( n2524 & n4160 ) | ( n2524 & n8012 ) | ( n4160 & n8012 ) ;
  assign n17428 = n17427 ^ n7479 ^ n3928 ;
  assign n17429 = n17428 ^ n4079 ^ n3670 ;
  assign n17435 = ( n496 & ~n12048 ) | ( n496 & n16070 ) | ( ~n12048 & n16070 ) ;
  assign n17433 = n2248 | n7053 ;
  assign n17434 = n17433 ^ n15417 ^ n11458 ;
  assign n17431 = ( x28 & ~n6493 ) | ( x28 & n6603 ) | ( ~n6493 & n6603 ) ;
  assign n17430 = n5440 ^ n3972 ^ n1057 ;
  assign n17432 = n17431 ^ n17430 ^ n16011 ;
  assign n17436 = n17435 ^ n17434 ^ n17432 ;
  assign n17437 = n7794 ^ n5317 ^ 1'b0 ;
  assign n17438 = ~n5490 & n17437 ;
  assign n17439 = n9152 & n17438 ;
  assign n17440 = ~n15247 & n17439 ;
  assign n17441 = ~n6303 & n9590 ;
  assign n17442 = ~n10052 & n12011 ;
  assign n17443 = n17442 ^ n9348 ^ n562 ;
  assign n17444 = n1868 & ~n17443 ;
  assign n17445 = n17444 ^ n3842 ^ n2861 ;
  assign n17448 = ( n4040 & n8651 ) | ( n4040 & ~n12085 ) | ( n8651 & ~n12085 ) ;
  assign n17447 = ( n2694 & n3346 ) | ( n2694 & n5476 ) | ( n3346 & n5476 ) ;
  assign n17446 = n17126 ^ n14977 ^ n2984 ;
  assign n17449 = n17448 ^ n17447 ^ n17446 ;
  assign n17452 = n9672 ^ n7387 ^ 1'b0 ;
  assign n17450 = n7381 ^ n6667 ^ n4941 ;
  assign n17451 = n17450 ^ n10397 ^ n2356 ;
  assign n17453 = n17452 ^ n17451 ^ n10167 ;
  assign n17454 = n6867 & n15199 ;
  assign n17455 = n17454 ^ n1988 ^ 1'b0 ;
  assign n17456 = ( n8255 & ~n12217 ) | ( n8255 & n17455 ) | ( ~n12217 & n17455 ) ;
  assign n17457 = n11701 ^ n7007 ^ 1'b0 ;
  assign n17458 = n4560 & n17457 ;
  assign n17463 = n2251 ^ n1316 ^ n885 ;
  assign n17459 = n4017 ^ n2429 ^ 1'b0 ;
  assign n17460 = n12663 | n17459 ;
  assign n17461 = n17460 ^ n4083 ^ 1'b0 ;
  assign n17462 = n680 & ~n17461 ;
  assign n17464 = n17463 ^ n17462 ^ 1'b0 ;
  assign n17465 = n17129 ^ n2659 ^ 1'b0 ;
  assign n17466 = ( ~n13890 & n14779 ) | ( ~n13890 & n17465 ) | ( n14779 & n17465 ) ;
  assign n17467 = n5691 ^ n2575 ^ 1'b0 ;
  assign n17468 = ( x61 & n1134 ) | ( x61 & n1761 ) | ( n1134 & n1761 ) ;
  assign n17469 = n17468 ^ n2853 ^ n1125 ;
  assign n17470 = n17469 ^ n15835 ^ n1102 ;
  assign n17471 = ( n2874 & n17467 ) | ( n2874 & ~n17470 ) | ( n17467 & ~n17470 ) ;
  assign n17472 = ( n2866 & ~n5052 ) | ( n2866 & n17471 ) | ( ~n5052 & n17471 ) ;
  assign n17473 = n5417 ^ n3992 ^ n3918 ;
  assign n17474 = ( ~n2495 & n5146 ) | ( ~n2495 & n14229 ) | ( n5146 & n14229 ) ;
  assign n17475 = ( n15809 & ~n17473 ) | ( n15809 & n17474 ) | ( ~n17473 & n17474 ) ;
  assign n17476 = n14981 ^ n11370 ^ n7644 ;
  assign n17477 = n11984 ^ n10073 ^ 1'b0 ;
  assign n17478 = ( n7692 & n8031 ) | ( n7692 & ~n12892 ) | ( n8031 & ~n12892 ) ;
  assign n17480 = n13890 ^ n11337 ^ n10265 ;
  assign n17479 = ( ~n1409 & n4910 ) | ( ~n1409 & n7937 ) | ( n4910 & n7937 ) ;
  assign n17481 = n17480 ^ n17479 ^ n801 ;
  assign n17482 = ( n149 & n17478 ) | ( n149 & ~n17481 ) | ( n17478 & ~n17481 ) ;
  assign n17483 = ( n275 & n5416 ) | ( n275 & ~n9817 ) | ( n5416 & ~n9817 ) ;
  assign n17484 = n17483 ^ n13825 ^ x77 ;
  assign n17489 = ( n10104 & n10629 ) | ( n10104 & ~n17143 ) | ( n10629 & ~n17143 ) ;
  assign n17485 = n12983 ^ n8861 ^ 1'b0 ;
  assign n17486 = n15768 | n17485 ;
  assign n17487 = n3021 ^ n1229 ^ 1'b0 ;
  assign n17488 = ~n17486 & n17487 ;
  assign n17490 = n17489 ^ n17488 ^ n14603 ;
  assign n17491 = n8296 ^ n4838 ^ n3856 ;
  assign n17492 = n17491 ^ n12598 ^ 1'b0 ;
  assign n17493 = n17492 ^ n8962 ^ n5843 ;
  assign n17496 = ~n1568 & n7191 ;
  assign n17494 = n5293 ^ n3034 ^ 1'b0 ;
  assign n17495 = ~n1611 & n17494 ;
  assign n17497 = n17496 ^ n17495 ^ n6330 ;
  assign n17499 = n9520 ^ n7840 ^ n1465 ;
  assign n17500 = n17499 ^ n12976 ^ n5408 ;
  assign n17498 = ( ~n1969 & n11543 ) | ( ~n1969 & n16044 ) | ( n11543 & n16044 ) ;
  assign n17501 = n17500 ^ n17498 ^ n10420 ;
  assign n17502 = n2586 & n8420 ;
  assign n17503 = n13892 ^ n10409 ^ 1'b0 ;
  assign n17504 = n2609 & n17503 ;
  assign n17505 = ( n164 & n2303 ) | ( n164 & n3105 ) | ( n2303 & n3105 ) ;
  assign n17506 = ~n14277 & n17505 ;
  assign n17507 = ( n10730 & n17504 ) | ( n10730 & ~n17506 ) | ( n17504 & ~n17506 ) ;
  assign n17508 = n11902 & n12023 ;
  assign n17509 = ( n246 & n5528 ) | ( n246 & n17508 ) | ( n5528 & n17508 ) ;
  assign n17510 = n17509 ^ n12401 ^ n7266 ;
  assign n17511 = n10646 ^ n8862 ^ n1956 ;
  assign n17512 = n8349 | n17511 ;
  assign n17513 = n4614 | n17512 ;
  assign n17514 = ( n4900 & n15175 ) | ( n4900 & n17513 ) | ( n15175 & n17513 ) ;
  assign n17515 = n12293 ^ n7699 ^ n1574 ;
  assign n17516 = n17515 ^ n16859 ^ n8031 ;
  assign n17517 = n9502 ^ n8349 ^ 1'b0 ;
  assign n17518 = n12239 | n17517 ;
  assign n17519 = ( n7269 & n9251 ) | ( n7269 & ~n15247 ) | ( n9251 & ~n15247 ) ;
  assign n17520 = n4342 | n6177 ;
  assign n17521 = n17519 | n17520 ;
  assign n17522 = n15954 ^ n14970 ^ n12600 ;
  assign n17523 = n14530 ^ n7458 ^ 1'b0 ;
  assign n17530 = ( n9935 & ~n15320 ) | ( n9935 & n15487 ) | ( ~n15320 & n15487 ) ;
  assign n17524 = n8673 ^ n3705 ^ n549 ;
  assign n17525 = ~n9325 & n17524 ;
  assign n17526 = n17525 ^ n1660 ^ 1'b0 ;
  assign n17527 = n17526 ^ n4369 ^ n1123 ;
  assign n17528 = ( n7125 & ~n9050 ) | ( n7125 & n14878 ) | ( ~n9050 & n14878 ) ;
  assign n17529 = ~n17527 & n17528 ;
  assign n17531 = n17530 ^ n17529 ^ 1'b0 ;
  assign n17532 = n7303 ^ n5631 ^ n4362 ;
  assign n17533 = n3011 & ~n16217 ;
  assign n17534 = n17532 & n17533 ;
  assign n17535 = n13632 & ~n17534 ;
  assign n17536 = n17535 ^ n15028 ^ 1'b0 ;
  assign n17537 = n7164 ^ n5595 ^ n3327 ;
  assign n17538 = n17537 ^ n6407 ^ n729 ;
  assign n17539 = n8637 & ~n9061 ;
  assign n17540 = n17539 ^ n13218 ^ 1'b0 ;
  assign n17541 = n7063 & n17540 ;
  assign n17542 = ~n2650 & n17541 ;
  assign n17543 = n16168 ^ n10182 ^ n6421 ;
  assign n17544 = n6806 ^ n5185 ^ 1'b0 ;
  assign n17545 = n4588 & ~n17544 ;
  assign n17546 = ( n4975 & n9258 ) | ( n4975 & ~n16325 ) | ( n9258 & ~n16325 ) ;
  assign n17547 = n17546 ^ n13184 ^ n1126 ;
  assign n17549 = ( ~n11597 & n11872 ) | ( ~n11597 & n14182 ) | ( n11872 & n14182 ) ;
  assign n17548 = n6611 | n12910 ;
  assign n17550 = n17549 ^ n17548 ^ 1'b0 ;
  assign n17551 = n14089 ^ n4544 ^ n1699 ;
  assign n17552 = n17551 ^ n15398 ^ n8085 ;
  assign n17553 = ( n157 & n513 ) | ( n157 & n1520 ) | ( n513 & n1520 ) ;
  assign n17554 = n11333 & ~n17553 ;
  assign n17555 = ( n7980 & ~n11716 ) | ( n7980 & n17554 ) | ( ~n11716 & n17554 ) ;
  assign n17556 = n8273 ^ n7307 ^ n3171 ;
  assign n17557 = n13303 & ~n17556 ;
  assign n17558 = n17557 ^ n11543 ^ n8416 ;
  assign n17559 = ( ~n1193 & n8319 ) | ( ~n1193 & n17558 ) | ( n8319 & n17558 ) ;
  assign n17560 = ( x126 & n6923 ) | ( x126 & n14466 ) | ( n6923 & n14466 ) ;
  assign n17561 = n11834 & n17560 ;
  assign n17562 = ~n3967 & n17561 ;
  assign n17563 = n8560 & ~n11435 ;
  assign n17564 = n17563 ^ n16015 ^ 1'b0 ;
  assign n17565 = ( n5379 & n8194 ) | ( n5379 & ~n10190 ) | ( n8194 & ~n10190 ) ;
  assign n17566 = n11195 ^ n7742 ^ n5045 ;
  assign n17567 = ( n4125 & n4190 ) | ( n4125 & n5884 ) | ( n4190 & n5884 ) ;
  assign n17568 = n4717 ^ n2444 ^ 1'b0 ;
  assign n17569 = ( ~n4971 & n9458 ) | ( ~n4971 & n9707 ) | ( n9458 & n9707 ) ;
  assign n17570 = ( n4601 & n5047 ) | ( n4601 & ~n17569 ) | ( n5047 & ~n17569 ) ;
  assign n17571 = n17566 | n17570 ;
  assign n17572 = n14547 ^ n8456 ^ n6736 ;
  assign n17573 = ( n14436 & n15305 ) | ( n14436 & n17572 ) | ( n15305 & n17572 ) ;
  assign n17574 = ( n2733 & n3207 ) | ( n2733 & n3895 ) | ( n3207 & n3895 ) ;
  assign n17575 = ( ~n1860 & n3307 ) | ( ~n1860 & n17574 ) | ( n3307 & n17574 ) ;
  assign n17576 = n2549 ^ n2524 ^ n1008 ;
  assign n17577 = n17576 ^ n10948 ^ n7039 ;
  assign n17578 = n11909 & ~n17577 ;
  assign n17582 = ( ~n2000 & n4650 ) | ( ~n2000 & n10142 ) | ( n4650 & n10142 ) ;
  assign n17579 = n1020 & ~n2234 ;
  assign n17580 = n1027 & n17579 ;
  assign n17581 = n17580 ^ n11654 ^ n856 ;
  assign n17583 = n17582 ^ n17581 ^ n14530 ;
  assign n17584 = ( n1319 & ~n5437 ) | ( n1319 & n6438 ) | ( ~n5437 & n6438 ) ;
  assign n17585 = ~n4992 & n6986 ;
  assign n17588 = n4918 & n5622 ;
  assign n17589 = n17588 ^ n4476 ^ 1'b0 ;
  assign n17586 = ( ~n831 & n3152 ) | ( ~n831 & n12059 ) | ( n3152 & n12059 ) ;
  assign n17587 = n10675 & n17586 ;
  assign n17590 = n17589 ^ n17587 ^ 1'b0 ;
  assign n17591 = n13045 ^ n7887 ^ n4672 ;
  assign n17592 = ( n383 & ~n1035 ) | ( n383 & n1123 ) | ( ~n1035 & n1123 ) ;
  assign n17593 = n3363 & n17592 ;
  assign n17594 = n1776 & n17593 ;
  assign n17595 = n17594 ^ n3784 ^ 1'b0 ;
  assign n17596 = n17591 & ~n17595 ;
  assign n17597 = n7589 ^ n3975 ^ n708 ;
  assign n17598 = ( n6482 & n11101 ) | ( n6482 & ~n13027 ) | ( n11101 & ~n13027 ) ;
  assign n17599 = n6761 | n6957 ;
  assign n17600 = n17599 ^ n1364 ^ 1'b0 ;
  assign n17601 = n17600 ^ n15976 ^ n6715 ;
  assign n17602 = n17598 | n17601 ;
  assign n17603 = n16290 ^ n5844 ^ 1'b0 ;
  assign n17604 = n1812 | n17603 ;
  assign n17605 = n17604 ^ n2738 ^ 1'b0 ;
  assign n17606 = n17605 ^ n6598 ^ 1'b0 ;
  assign n17607 = ( n1909 & n6415 ) | ( n1909 & ~n17002 ) | ( n6415 & ~n17002 ) ;
  assign n17608 = n951 & n11778 ;
  assign n17609 = ~n13278 & n17608 ;
  assign n17610 = n17609 ^ n15908 ^ n11619 ;
  assign n17613 = n16584 ^ n14368 ^ n14093 ;
  assign n17611 = ( ~n7276 & n11872 ) | ( ~n7276 & n13405 ) | ( n11872 & n13405 ) ;
  assign n17612 = n17611 ^ n5329 ^ 1'b0 ;
  assign n17614 = n17613 ^ n17612 ^ n1940 ;
  assign n17615 = n1576 & n2876 ;
  assign n17616 = n17615 ^ n8703 ^ 1'b0 ;
  assign n17617 = n17616 ^ n2945 ^ n2918 ;
  assign n17618 = n5804 & ~n15406 ;
  assign n17619 = n17618 ^ n14023 ^ 1'b0 ;
  assign n17620 = n11064 ^ n4928 ^ 1'b0 ;
  assign n17621 = n15675 ^ n3166 ^ n1225 ;
  assign n17622 = n17621 ^ n7657 ^ n2888 ;
  assign n17623 = ( n8312 & ~n12695 ) | ( n8312 & n17622 ) | ( ~n12695 & n17622 ) ;
  assign n17624 = ( n8063 & n9391 ) | ( n8063 & n13293 ) | ( n9391 & n13293 ) ;
  assign n17625 = n17417 ^ n16776 ^ n2482 ;
  assign n17626 = n11665 ^ n9948 ^ 1'b0 ;
  assign n17627 = n8152 | n17626 ;
  assign n17628 = ( ~n2662 & n6546 ) | ( ~n2662 & n17376 ) | ( n6546 & n17376 ) ;
  assign n17629 = ( n9568 & n15197 ) | ( n9568 & n17628 ) | ( n15197 & n17628 ) ;
  assign n17632 = n9127 & n17401 ;
  assign n17630 = n11422 ^ n7125 ^ n2272 ;
  assign n17631 = n17630 ^ n13041 ^ n12559 ;
  assign n17633 = n17632 ^ n17631 ^ n9908 ;
  assign n17634 = ~n5196 & n12002 ;
  assign n17635 = ( n6290 & n7919 ) | ( n6290 & ~n17634 ) | ( n7919 & ~n17634 ) ;
  assign n17636 = n17635 ^ n16619 ^ n4382 ;
  assign n17637 = n17636 ^ n8932 ^ n8398 ;
  assign n17638 = n10099 ^ n9183 ^ n714 ;
  assign n17639 = n3574 & n13176 ;
  assign n17640 = n8006 & n17639 ;
  assign n17641 = n7684 ^ n5422 ^ 1'b0 ;
  assign n17642 = n17640 | n17641 ;
  assign n17643 = n17642 ^ n13713 ^ n5858 ;
  assign n17644 = n10511 ^ n4664 ^ n1479 ;
  assign n17645 = n3365 ^ n3128 ^ 1'b0 ;
  assign n17646 = ~n2233 & n17645 ;
  assign n17647 = n12843 ^ n2613 ^ 1'b0 ;
  assign n17648 = n17646 & ~n17647 ;
  assign n17649 = ( ~n7432 & n17644 ) | ( ~n7432 & n17648 ) | ( n17644 & n17648 ) ;
  assign n17651 = n626 & ~n8016 ;
  assign n17650 = n4190 & n12070 ;
  assign n17652 = n17651 ^ n17650 ^ 1'b0 ;
  assign n17653 = ( n4772 & n7406 ) | ( n4772 & n10559 ) | ( n7406 & n10559 ) ;
  assign n17654 = n8374 & n17653 ;
  assign n17655 = ~n8534 & n17654 ;
  assign n17656 = ( ~n372 & n17652 ) | ( ~n372 & n17655 ) | ( n17652 & n17655 ) ;
  assign n17657 = n1772 | n3286 ;
  assign n17658 = ( n1816 & n6378 ) | ( n1816 & n17657 ) | ( n6378 & n17657 ) ;
  assign n17659 = ~n380 & n2786 ;
  assign n17660 = n17659 ^ n157 ^ 1'b0 ;
  assign n17661 = ( ~n3911 & n4388 ) | ( ~n3911 & n17660 ) | ( n4388 & n17660 ) ;
  assign n17662 = n17661 ^ n2651 ^ n1899 ;
  assign n17663 = n17662 ^ n1421 ^ 1'b0 ;
  assign n17664 = n14925 & n17663 ;
  assign n17665 = ( ~n577 & n7454 ) | ( ~n577 & n14992 ) | ( n7454 & n14992 ) ;
  assign n17666 = n12049 ^ n5978 ^ 1'b0 ;
  assign n17667 = n12382 ^ n2771 ^ 1'b0 ;
  assign n17668 = n9316 & n17667 ;
  assign n17669 = n11858 ^ n239 ^ 1'b0 ;
  assign n17670 = ( n12944 & n17668 ) | ( n12944 & ~n17669 ) | ( n17668 & ~n17669 ) ;
  assign n17671 = ~n10904 & n17670 ;
  assign n17672 = n7849 & ~n17177 ;
  assign n17673 = n17672 ^ n7577 ^ 1'b0 ;
  assign n17677 = ( n2292 & n4505 ) | ( n2292 & ~n6292 ) | ( n4505 & ~n6292 ) ;
  assign n17678 = n17677 ^ n7457 ^ n6742 ;
  assign n17674 = n16495 ^ n8558 ^ n4569 ;
  assign n17675 = n9229 ^ n7142 ^ n5063 ;
  assign n17676 = n17674 | n17675 ;
  assign n17679 = n17678 ^ n17676 ^ 1'b0 ;
  assign n17680 = n5151 | n10659 ;
  assign n17681 = n17680 ^ n11801 ^ 1'b0 ;
  assign n17682 = n17149 ^ n4281 ^ n2733 ;
  assign n17683 = n17681 & n17682 ;
  assign n17684 = n17683 ^ n2341 ^ 1'b0 ;
  assign n17685 = ~n759 & n9826 ;
  assign n17686 = ( n3378 & n7731 ) | ( n3378 & ~n12224 ) | ( n7731 & ~n12224 ) ;
  assign n17687 = n4850 ^ n3423 ^ n2273 ;
  assign n17688 = x56 & ~n14393 ;
  assign n17689 = n17687 & n17688 ;
  assign n17690 = n15891 ^ n10640 ^ n8926 ;
  assign n17691 = n17690 ^ n14230 ^ n4996 ;
  assign n17692 = n16157 ^ n14501 ^ n10613 ;
  assign n17693 = n6865 & n14904 ;
  assign n17694 = n17693 ^ n9739 ^ n6516 ;
  assign n17695 = n12980 ^ n9482 ^ n4850 ;
  assign n17696 = ( n868 & n8357 ) | ( n868 & ~n17695 ) | ( n8357 & ~n17695 ) ;
  assign n17697 = ( n3720 & n3983 ) | ( n3720 & ~n17696 ) | ( n3983 & ~n17696 ) ;
  assign n17698 = n5824 ^ n144 ^ 1'b0 ;
  assign n17699 = ~n4429 & n17698 ;
  assign n17700 = n17664 ^ n13172 ^ 1'b0 ;
  assign n17701 = n17699 & ~n17700 ;
  assign n17702 = ( x119 & n3956 ) | ( x119 & ~n11232 ) | ( n3956 & ~n11232 ) ;
  assign n17703 = n8157 ^ n4646 ^ n470 ;
  assign n17704 = n17703 ^ n1367 ^ 1'b0 ;
  assign n17705 = ( n5058 & ~n17702 ) | ( n5058 & n17704 ) | ( ~n17702 & n17704 ) ;
  assign n17706 = n17705 ^ n10285 ^ 1'b0 ;
  assign n17707 = n9811 & ~n17706 ;
  assign n17709 = n14209 ^ n2098 ^ 1'b0 ;
  assign n17708 = ( n2398 & n3365 ) | ( n2398 & n6886 ) | ( n3365 & n6886 ) ;
  assign n17710 = n17709 ^ n17708 ^ n6312 ;
  assign n17711 = n10485 ^ n8775 ^ n5072 ;
  assign n17712 = n5946 | n11584 ;
  assign n17713 = n17712 ^ n4299 ^ 1'b0 ;
  assign n17714 = n3253 | n17713 ;
  assign n17715 = n17711 | n17714 ;
  assign n17716 = ( n3042 & ~n16436 ) | ( n3042 & n17715 ) | ( ~n16436 & n17715 ) ;
  assign n17717 = n17710 | n17716 ;
  assign n17718 = n6226 ^ n2103 ^ n1291 ;
  assign n17719 = ( n11194 & ~n13443 ) | ( n11194 & n16367 ) | ( ~n13443 & n16367 ) ;
  assign n17720 = ( n4557 & n6180 ) | ( n4557 & n17719 ) | ( n6180 & n17719 ) ;
  assign n17721 = n4388 & ~n7651 ;
  assign n17722 = n17720 & n17721 ;
  assign n17723 = n13781 ^ n12408 ^ n1549 ;
  assign n17724 = n9667 ^ n5020 ^ n4724 ;
  assign n17725 = ( ~n11199 & n12902 ) | ( ~n11199 & n17724 ) | ( n12902 & n17724 ) ;
  assign n17726 = ( n17722 & ~n17723 ) | ( n17722 & n17725 ) | ( ~n17723 & n17725 ) ;
  assign n17727 = n885 & n4982 ;
  assign n17730 = ~n11373 & n15386 ;
  assign n17731 = n9509 ^ n2665 ^ n2581 ;
  assign n17732 = n2346 & ~n17731 ;
  assign n17733 = n17730 & n17732 ;
  assign n17728 = ( x25 & ~n1903 ) | ( x25 & n8818 ) | ( ~n1903 & n8818 ) ;
  assign n17729 = ~n9732 & n17728 ;
  assign n17734 = n17733 ^ n17729 ^ n946 ;
  assign n17735 = x114 & n8786 ;
  assign n17736 = n17735 ^ n3699 ^ 1'b0 ;
  assign n17737 = n17736 ^ n15985 ^ n11743 ;
  assign n17738 = ( n3042 & ~n5676 ) | ( n3042 & n6220 ) | ( ~n5676 & n6220 ) ;
  assign n17739 = n17738 ^ n11158 ^ n1591 ;
  assign n17740 = ( n1098 & n2085 ) | ( n1098 & n3392 ) | ( n2085 & n3392 ) ;
  assign n17741 = ~n4390 & n17740 ;
  assign n17742 = ~n9333 & n17741 ;
  assign n17743 = n17742 ^ n5359 ^ n1025 ;
  assign n17744 = n17743 ^ n13340 ^ n7796 ;
  assign n17745 = ( n1153 & n2957 ) | ( n1153 & ~n17744 ) | ( n2957 & ~n17744 ) ;
  assign n17746 = ( n2307 & ~n17739 ) | ( n2307 & n17745 ) | ( ~n17739 & n17745 ) ;
  assign n17747 = ( n1664 & n4640 ) | ( n1664 & ~n8684 ) | ( n4640 & ~n8684 ) ;
  assign n17748 = ( n671 & ~n1582 ) | ( n671 & n17747 ) | ( ~n1582 & n17747 ) ;
  assign n17749 = ( n6211 & ~n7004 ) | ( n6211 & n7718 ) | ( ~n7004 & n7718 ) ;
  assign n17750 = ( n7964 & ~n17748 ) | ( n7964 & n17749 ) | ( ~n17748 & n17749 ) ;
  assign n17752 = ( n1645 & n4756 ) | ( n1645 & n8172 ) | ( n4756 & n8172 ) ;
  assign n17751 = n3915 & ~n6340 ;
  assign n17753 = n17752 ^ n17751 ^ n7613 ;
  assign n17754 = ( ~n3910 & n6626 ) | ( ~n3910 & n17753 ) | ( n6626 & n17753 ) ;
  assign n17756 = ( n1719 & n3737 ) | ( n1719 & n5415 ) | ( n3737 & n5415 ) ;
  assign n17757 = ( n339 & n5520 ) | ( n339 & ~n17756 ) | ( n5520 & ~n17756 ) ;
  assign n17758 = n17757 ^ n10765 ^ n8022 ;
  assign n17755 = n2146 & ~n8644 ;
  assign n17759 = n17758 ^ n17755 ^ n8533 ;
  assign n17760 = ( ~n2792 & n5484 ) | ( ~n2792 & n17759 ) | ( n5484 & n17759 ) ;
  assign n17763 = n15907 ^ n10589 ^ 1'b0 ;
  assign n17764 = ~n4124 & n17763 ;
  assign n17761 = n15354 ^ n7911 ^ 1'b0 ;
  assign n17762 = ~n333 & n17761 ;
  assign n17765 = n17764 ^ n17762 ^ n10182 ;
  assign n17766 = ( n9672 & n10731 ) | ( n9672 & ~n17765 ) | ( n10731 & ~n17765 ) ;
  assign n17767 = n820 & n17766 ;
  assign n17768 = n12672 ^ n4987 ^ n1800 ;
  assign n17769 = n5109 | n10343 ;
  assign n17770 = n11469 & ~n17769 ;
  assign n17771 = n16012 ^ n13173 ^ n558 ;
  assign n17772 = ( n3705 & ~n7255 ) | ( n3705 & n13966 ) | ( ~n7255 & n13966 ) ;
  assign n17773 = ( ~n4804 & n17771 ) | ( ~n4804 & n17772 ) | ( n17771 & n17772 ) ;
  assign n17775 = n3846 | n12502 ;
  assign n17774 = n2665 & ~n13072 ;
  assign n17776 = n17775 ^ n17774 ^ n310 ;
  assign n17777 = n6365 ^ n2615 ^ 1'b0 ;
  assign n17778 = ~n12334 & n17777 ;
  assign n17779 = n17778 ^ n10554 ^ n1159 ;
  assign n17780 = n17779 ^ n11199 ^ n8053 ;
  assign n17781 = ( n2808 & n8254 ) | ( n2808 & ~n17780 ) | ( n8254 & ~n17780 ) ;
  assign n17782 = ( n3700 & ~n10534 ) | ( n3700 & n17781 ) | ( ~n10534 & n17781 ) ;
  assign n17783 = ( n4985 & n14379 ) | ( n4985 & ~n17782 ) | ( n14379 & ~n17782 ) ;
  assign n17784 = n4764 | n6721 ;
  assign n17785 = n14107 | n17784 ;
  assign n17786 = n4406 ^ n3088 ^ n214 ;
  assign n17787 = ( n8568 & n17785 ) | ( n8568 & ~n17786 ) | ( n17785 & ~n17786 ) ;
  assign n17792 = ~n2397 & n9792 ;
  assign n17788 = n7404 | n9958 ;
  assign n17789 = ( n5377 & n10708 ) | ( n5377 & ~n17788 ) | ( n10708 & ~n17788 ) ;
  assign n17790 = n17789 ^ n15474 ^ n3109 ;
  assign n17791 = n17790 ^ n7121 ^ n4183 ;
  assign n17793 = n17792 ^ n17791 ^ n6092 ;
  assign n17794 = ( ~n1324 & n8994 ) | ( ~n1324 & n17793 ) | ( n8994 & n17793 ) ;
  assign n17795 = n6071 ^ n4451 ^ 1'b0 ;
  assign n17796 = n9524 & ~n17795 ;
  assign n17797 = n1361 ^ n1042 ^ 1'b0 ;
  assign n17798 = n3986 | n17797 ;
  assign n17799 = n7041 ^ n5724 ^ n1820 ;
  assign n17800 = n10161 ^ n7350 ^ n4641 ;
  assign n17801 = n5200 ^ n2757 ^ 1'b0 ;
  assign n17802 = n4947 & n17801 ;
  assign n17803 = ( n17799 & n17800 ) | ( n17799 & n17802 ) | ( n17800 & n17802 ) ;
  assign n17804 = ( n7059 & n8169 ) | ( n7059 & n8349 ) | ( n8169 & n8349 ) ;
  assign n17805 = ( n4039 & n7364 ) | ( n4039 & ~n9426 ) | ( n7364 & ~n9426 ) ;
  assign n17806 = ( ~n896 & n6106 ) | ( ~n896 & n17805 ) | ( n6106 & n17805 ) ;
  assign n17807 = n17804 & n17806 ;
  assign n17808 = n17807 ^ n17577 ^ 1'b0 ;
  assign n17813 = n3525 & n13917 ;
  assign n17814 = n17813 ^ n9708 ^ 1'b0 ;
  assign n17809 = n11425 ^ n1021 ^ 1'b0 ;
  assign n17810 = ( n337 & ~n4114 ) | ( n337 & n17809 ) | ( ~n4114 & n17809 ) ;
  assign n17811 = n1537 & ~n17810 ;
  assign n17812 = n4673 & n17811 ;
  assign n17815 = n17814 ^ n17812 ^ n270 ;
  assign n17816 = n7507 ^ n5871 ^ n3735 ;
  assign n17817 = n14401 | n17816 ;
  assign n17818 = n2073 | n17817 ;
  assign n17819 = ( n1849 & n9221 ) | ( n1849 & n15481 ) | ( n9221 & n15481 ) ;
  assign n17820 = n12265 ^ n8474 ^ n3820 ;
  assign n17821 = n17820 ^ n5903 ^ x76 ;
  assign n17822 = n17821 ^ n12869 ^ n6689 ;
  assign n17823 = ( n17818 & ~n17819 ) | ( n17818 & n17822 ) | ( ~n17819 & n17822 ) ;
  assign n17824 = ~n2115 & n6636 ;
  assign n17825 = ~n150 & n17824 ;
  assign n17826 = n17825 ^ n11165 ^ n5192 ;
  assign n17827 = ( ~n6861 & n11779 ) | ( ~n6861 & n13875 ) | ( n11779 & n13875 ) ;
  assign n17828 = ( n198 & ~n6077 ) | ( n198 & n17827 ) | ( ~n6077 & n17827 ) ;
  assign n17829 = n14716 & n17828 ;
  assign n17830 = ~n1269 & n4213 ;
  assign n17831 = n17830 ^ n9007 ^ 1'b0 ;
  assign n17832 = ( n3488 & n16265 ) | ( n3488 & n17831 ) | ( n16265 & n17831 ) ;
  assign n17833 = n17264 ^ n13152 ^ 1'b0 ;
  assign n17834 = ~n17832 & n17833 ;
  assign n17835 = n17834 ^ n459 ^ 1'b0 ;
  assign n17836 = ~n1501 & n17835 ;
  assign n17837 = n6755 ^ n1643 ^ n567 ;
  assign n17838 = n17837 ^ n16746 ^ 1'b0 ;
  assign n17839 = n2932 & ~n17838 ;
  assign n17840 = n7972 ^ n3867 ^ x46 ;
  assign n17841 = n17840 ^ n6106 ^ n2692 ;
  assign n17842 = n8763 ^ n7273 ^ 1'b0 ;
  assign n17843 = ( n9674 & ~n11765 ) | ( n9674 & n15293 ) | ( ~n11765 & n15293 ) ;
  assign n17852 = n7585 ^ n5763 ^ n2096 ;
  assign n17853 = ( n1124 & ~n10488 ) | ( n1124 & n17852 ) | ( ~n10488 & n17852 ) ;
  assign n17854 = ( n4487 & n8810 ) | ( n4487 & ~n17853 ) | ( n8810 & ~n17853 ) ;
  assign n17855 = ~n3703 & n17854 ;
  assign n17849 = x83 & n5667 ;
  assign n17850 = n17849 ^ n3545 ^ 1'b0 ;
  assign n17851 = n17850 ^ n7151 ^ n1847 ;
  assign n17844 = ( n143 & ~n756 ) | ( n143 & n11772 ) | ( ~n756 & n11772 ) ;
  assign n17845 = ~n735 & n17844 ;
  assign n17846 = n6148 ^ n4011 ^ n2431 ;
  assign n17847 = n17846 ^ n7847 ^ n7380 ;
  assign n17848 = ( n3092 & n17845 ) | ( n3092 & n17847 ) | ( n17845 & n17847 ) ;
  assign n17856 = n17855 ^ n17851 ^ n17848 ;
  assign n17857 = ( n486 & n8479 ) | ( n486 & ~n16431 ) | ( n8479 & ~n16431 ) ;
  assign n17858 = n13296 | n17857 ;
  assign n17859 = n17858 ^ n3699 ^ 1'b0 ;
  assign n17860 = ( n4434 & ~n9229 ) | ( n4434 & n13108 ) | ( ~n9229 & n13108 ) ;
  assign n17861 = n8484 ^ n4536 ^ n2897 ;
  assign n17862 = ( n2908 & n5273 ) | ( n2908 & ~n13652 ) | ( n5273 & ~n13652 ) ;
  assign n17863 = ( n6425 & n7196 ) | ( n6425 & ~n17862 ) | ( n7196 & ~n17862 ) ;
  assign n17864 = ( ~n4623 & n9544 ) | ( ~n4623 & n12654 ) | ( n9544 & n12654 ) ;
  assign n17865 = n17864 ^ n15072 ^ n13462 ;
  assign n17866 = ~n2573 & n17865 ;
  assign n17867 = n3264 & ~n5356 ;
  assign n17868 = n17867 ^ n1689 ^ 1'b0 ;
  assign n17869 = ( n8268 & ~n12017 ) | ( n8268 & n16993 ) | ( ~n12017 & n16993 ) ;
  assign n17870 = ( n8350 & n15514 ) | ( n8350 & n17869 ) | ( n15514 & n17869 ) ;
  assign n17871 = n17516 ^ n6511 ^ 1'b0 ;
  assign n17872 = ( n1109 & n6029 ) | ( n1109 & ~n15825 ) | ( n6029 & ~n15825 ) ;
  assign n17873 = ( n3462 & ~n4166 ) | ( n3462 & n17872 ) | ( ~n4166 & n17872 ) ;
  assign n17874 = ~n8078 & n14103 ;
  assign n17880 = n11322 ^ n11083 ^ n8491 ;
  assign n17875 = n5312 & ~n5995 ;
  assign n17876 = n17875 ^ n5134 ^ 1'b0 ;
  assign n17877 = ~n2696 & n17876 ;
  assign n17878 = ~n1659 & n17877 ;
  assign n17879 = ( ~n162 & n8124 ) | ( ~n162 & n17878 ) | ( n8124 & n17878 ) ;
  assign n17881 = n17880 ^ n17879 ^ n3817 ;
  assign n17882 = n11871 ^ n9104 ^ n3600 ;
  assign n17891 = n7727 ^ n3924 ^ n3604 ;
  assign n17888 = n5425 | n11459 ;
  assign n17889 = ( n12393 & n12488 ) | ( n12393 & n17888 ) | ( n12488 & n17888 ) ;
  assign n17890 = ~n3518 & n17889 ;
  assign n17892 = n17891 ^ n17890 ^ n16139 ;
  assign n17883 = ( n2147 & n3355 ) | ( n2147 & n3771 ) | ( n3355 & n3771 ) ;
  assign n17884 = n17883 ^ n1335 ^ 1'b0 ;
  assign n17885 = n17884 ^ n14382 ^ n6429 ;
  assign n17886 = ( ~n1081 & n17513 ) | ( ~n1081 & n17885 ) | ( n17513 & n17885 ) ;
  assign n17887 = n8773 | n17886 ;
  assign n17893 = n17892 ^ n17887 ^ 1'b0 ;
  assign n17894 = n15301 ^ n8679 ^ 1'b0 ;
  assign n17895 = n13491 | n17894 ;
  assign n17896 = ~n2832 & n5044 ;
  assign n17897 = n14865 & n17896 ;
  assign n17898 = ~n3562 & n17897 ;
  assign n17899 = ( n3861 & ~n8321 ) | ( n3861 & n17898 ) | ( ~n8321 & n17898 ) ;
  assign n17900 = n2391 & n8176 ;
  assign n17901 = n17900 ^ n16501 ^ 1'b0 ;
  assign n17902 = n17899 & ~n17901 ;
  assign n17903 = n9631 ^ n4857 ^ n1087 ;
  assign n17904 = n8223 ^ n4038 ^ 1'b0 ;
  assign n17905 = ( n4364 & ~n16824 ) | ( n4364 & n17904 ) | ( ~n16824 & n17904 ) ;
  assign n17906 = n7864 ^ n4361 ^ 1'b0 ;
  assign n17907 = n10606 & n17906 ;
  assign n17908 = n10803 ^ n1788 ^ 1'b0 ;
  assign n17909 = n6015 | n17908 ;
  assign n17910 = ( n8834 & n15054 ) | ( n8834 & n17909 ) | ( n15054 & n17909 ) ;
  assign n17911 = ( ~n3277 & n9421 ) | ( ~n3277 & n11799 ) | ( n9421 & n11799 ) ;
  assign n17912 = n17911 ^ n9046 ^ n629 ;
  assign n17913 = ( ~x124 & n5868 ) | ( ~x124 & n11885 ) | ( n5868 & n11885 ) ;
  assign n17914 = n5073 ^ n3578 ^ n2982 ;
  assign n17915 = ( n3985 & ~n5837 ) | ( n3985 & n15638 ) | ( ~n5837 & n15638 ) ;
  assign n17916 = n17914 & n17915 ;
  assign n17917 = ~n8996 & n17916 ;
  assign n17918 = ( n707 & n17913 ) | ( n707 & n17917 ) | ( n17913 & n17917 ) ;
  assign n17919 = ( ~n12149 & n17912 ) | ( ~n12149 & n17918 ) | ( n17912 & n17918 ) ;
  assign n17923 = n13740 ^ n11432 ^ n8821 ;
  assign n17922 = ( n1282 & n1804 ) | ( n1282 & ~n8996 ) | ( n1804 & ~n8996 ) ;
  assign n17924 = n17923 ^ n17922 ^ n11279 ;
  assign n17920 = n12468 ^ n7198 ^ n7145 ;
  assign n17921 = n17920 ^ n14367 ^ n4763 ;
  assign n17925 = n17924 ^ n17921 ^ n13473 ;
  assign n17926 = n8685 ^ n7848 ^ n5865 ;
  assign n17928 = n9759 ^ n8065 ^ n2085 ;
  assign n17927 = n1760 & n2593 ;
  assign n17929 = n17928 ^ n17927 ^ n16359 ;
  assign n17930 = ( ~n3597 & n5622 ) | ( ~n3597 & n6544 ) | ( n5622 & n6544 ) ;
  assign n17931 = n17930 ^ n14045 ^ n10039 ;
  assign n17932 = n16830 ^ n9526 ^ n4302 ;
  assign n17933 = n6874 ^ n255 ^ 1'b0 ;
  assign n17934 = n16022 & n17933 ;
  assign n17935 = n17934 ^ n17309 ^ n12305 ;
  assign n17936 = n2477 ^ n920 ^ 1'b0 ;
  assign n17937 = ~n4585 & n17936 ;
  assign n17938 = n17937 ^ n5525 ^ 1'b0 ;
  assign n17939 = ( n3854 & n15748 ) | ( n3854 & ~n17938 ) | ( n15748 & ~n17938 ) ;
  assign n17940 = n11985 ^ n7903 ^ n2720 ;
  assign n17941 = n11212 ^ n2812 ^ n1776 ;
  assign n17942 = ( n3378 & ~n11439 ) | ( n3378 & n17941 ) | ( ~n11439 & n17941 ) ;
  assign n17945 = n14015 ^ n7397 ^ n5301 ;
  assign n17943 = ( n3093 & n4069 ) | ( n3093 & ~n9266 ) | ( n4069 & ~n9266 ) ;
  assign n17944 = ( ~n8822 & n9556 ) | ( ~n8822 & n17943 ) | ( n9556 & n17943 ) ;
  assign n17946 = n17945 ^ n17944 ^ n3859 ;
  assign n17947 = n16295 ^ n10762 ^ n8134 ;
  assign n17948 = n13205 ^ n2050 ^ 1'b0 ;
  assign n17949 = n17947 | n17948 ;
  assign n17950 = ( n4434 & n5068 ) | ( n4434 & ~n12357 ) | ( n5068 & ~n12357 ) ;
  assign n17951 = n9846 ^ n2804 ^ 1'b0 ;
  assign n17952 = n17950 & ~n17951 ;
  assign n17953 = ( ~n2723 & n3267 ) | ( ~n2723 & n7154 ) | ( n3267 & n7154 ) ;
  assign n17954 = n6185 & n17953 ;
  assign n17955 = n17954 ^ n6370 ^ 1'b0 ;
  assign n17956 = n1494 ^ n1242 ^ 1'b0 ;
  assign n17957 = n10269 & ~n17956 ;
  assign n17958 = ~n4433 & n17957 ;
  assign n17959 = ( n10714 & n17955 ) | ( n10714 & ~n17958 ) | ( n17955 & ~n17958 ) ;
  assign n17960 = ( n3515 & n11547 ) | ( n3515 & ~n12878 ) | ( n11547 & ~n12878 ) ;
  assign n17961 = n17792 ^ n10861 ^ n5662 ;
  assign n17962 = ( n8799 & ~n17960 ) | ( n8799 & n17961 ) | ( ~n17960 & n17961 ) ;
  assign n17963 = n17805 ^ n12878 ^ n3096 ;
  assign n17964 = n16154 | n17963 ;
  assign n17965 = ( n2881 & n3835 ) | ( n2881 & n5997 ) | ( n3835 & n5997 ) ;
  assign n17966 = n17965 ^ n4892 ^ n1677 ;
  assign n17967 = n8235 & ~n10778 ;
  assign n17968 = n17966 & n17967 ;
  assign n17969 = n13247 ^ n3986 ^ n2837 ;
  assign n17970 = n17969 ^ n339 ^ 1'b0 ;
  assign n17971 = ( n6432 & ~n14271 ) | ( n6432 & n16953 ) | ( ~n14271 & n16953 ) ;
  assign n17972 = n14881 ^ n13763 ^ 1'b0 ;
  assign n17973 = ( ~n2988 & n5361 ) | ( ~n2988 & n8253 ) | ( n5361 & n8253 ) ;
  assign n17974 = n17973 ^ n6186 ^ n2106 ;
  assign n17975 = n10925 ^ n3620 ^ 1'b0 ;
  assign n17976 = n16104 ^ n1674 ^ 1'b0 ;
  assign n17977 = ( n3128 & n15028 ) | ( n3128 & ~n17976 ) | ( n15028 & ~n17976 ) ;
  assign n17978 = ~n5568 & n6908 ;
  assign n17979 = n17978 ^ n14254 ^ 1'b0 ;
  assign n17982 = n12672 ^ n10701 ^ n424 ;
  assign n17980 = n9865 ^ n818 ^ 1'b0 ;
  assign n17981 = n8054 | n17980 ;
  assign n17983 = n17982 ^ n17981 ^ n12856 ;
  assign n17984 = ( n809 & ~n1767 ) | ( n809 & n14659 ) | ( ~n1767 & n14659 ) ;
  assign n17985 = n17984 ^ n7773 ^ n673 ;
  assign n17986 = ( n2868 & n9757 ) | ( n2868 & n10698 ) | ( n9757 & n10698 ) ;
  assign n17987 = ( n6636 & n10512 ) | ( n6636 & n17986 ) | ( n10512 & n17986 ) ;
  assign n17988 = n10406 ^ n5117 ^ 1'b0 ;
  assign n17989 = ~n8570 & n17988 ;
  assign n17990 = ( ~n903 & n4603 ) | ( ~n903 & n17989 ) | ( n4603 & n17989 ) ;
  assign n17991 = n8679 ^ n5392 ^ n3910 ;
  assign n17993 = n8350 ^ n4864 ^ n2374 ;
  assign n17992 = n1748 ^ n1527 ^ 1'b0 ;
  assign n17994 = n17993 ^ n17992 ^ 1'b0 ;
  assign n17995 = ~n17991 & n17994 ;
  assign n17996 = n17995 ^ n8870 ^ n814 ;
  assign n17997 = ( n9772 & n13205 ) | ( n9772 & ~n15654 ) | ( n13205 & ~n15654 ) ;
  assign n17998 = n17211 ^ n9560 ^ n3580 ;
  assign n17999 = n17998 ^ n14925 ^ n3633 ;
  assign n18000 = ( n1437 & n17261 ) | ( n1437 & n17999 ) | ( n17261 & n17999 ) ;
  assign n18001 = ( n3932 & n5005 ) | ( n3932 & ~n12212 ) | ( n5005 & ~n12212 ) ;
  assign n18002 = ( n734 & ~n1536 ) | ( n734 & n18001 ) | ( ~n1536 & n18001 ) ;
  assign n18003 = n5041 & ~n18002 ;
  assign n18004 = ~n18000 & n18003 ;
  assign n18007 = ( n3010 & ~n13570 ) | ( n3010 & n13895 ) | ( ~n13570 & n13895 ) ;
  assign n18005 = n1474 & n3182 ;
  assign n18006 = n18005 ^ n8844 ^ n8313 ;
  assign n18008 = n18007 ^ n18006 ^ n9181 ;
  assign n18009 = n18008 ^ n17847 ^ 1'b0 ;
  assign n18010 = n3288 & n18009 ;
  assign n18011 = n10266 ^ n5031 ^ n1968 ;
  assign n18012 = ( n4162 & ~n9526 ) | ( n4162 & n12539 ) | ( ~n9526 & n12539 ) ;
  assign n18013 = n9117 ^ n6150 ^ n983 ;
  assign n18014 = ( n1203 & n6019 ) | ( n1203 & ~n18013 ) | ( n6019 & ~n18013 ) ;
  assign n18015 = n18014 ^ n7414 ^ n1065 ;
  assign n18016 = n18015 ^ n14584 ^ n7004 ;
  assign n18017 = n13275 & ~n16460 ;
  assign n18023 = n6447 ^ n4390 ^ n2438 ;
  assign n18024 = n18023 ^ n11589 ^ 1'b0 ;
  assign n18018 = ( n8411 & ~n9005 ) | ( n8411 & n12504 ) | ( ~n9005 & n12504 ) ;
  assign n18019 = n18018 ^ n15895 ^ n5170 ;
  assign n18020 = n13768 ^ n5435 ^ n2604 ;
  assign n18021 = n18020 ^ n14348 ^ 1'b0 ;
  assign n18022 = ~n18019 & n18021 ;
  assign n18025 = n18024 ^ n18022 ^ n8233 ;
  assign n18026 = n7686 ^ n4976 ^ n2685 ;
  assign n18027 = ( n5573 & n6512 ) | ( n5573 & n9091 ) | ( n6512 & n9091 ) ;
  assign n18028 = ( n4469 & n6423 ) | ( n4469 & n18027 ) | ( n6423 & n18027 ) ;
  assign n18029 = n14370 ^ n10594 ^ n1274 ;
  assign n18030 = n256 | n6040 ;
  assign n18031 = n15898 ^ n14699 ^ n5949 ;
  assign n18032 = n10877 ^ n2706 ^ x86 ;
  assign n18033 = n8188 & n13041 ;
  assign n18034 = n18032 & n18033 ;
  assign n18035 = ( n18030 & ~n18031 ) | ( n18030 & n18034 ) | ( ~n18031 & n18034 ) ;
  assign n18036 = n17982 ^ n9131 ^ n7044 ;
  assign n18037 = ~n1400 & n10029 ;
  assign n18038 = n18036 & n18037 ;
  assign n18039 = n6794 ^ n4823 ^ n4809 ;
  assign n18040 = n18039 ^ n9566 ^ n8755 ;
  assign n18041 = n16578 & ~n18040 ;
  assign n18042 = n18041 ^ n4363 ^ 1'b0 ;
  assign n18043 = n8741 ^ n8632 ^ 1'b0 ;
  assign n18044 = n4544 & ~n18043 ;
  assign n18045 = ( ~n896 & n3040 ) | ( ~n896 & n6706 ) | ( n3040 & n6706 ) ;
  assign n18046 = ( n6540 & n18044 ) | ( n6540 & ~n18045 ) | ( n18044 & ~n18045 ) ;
  assign n18047 = ( ~n14709 & n15839 ) | ( ~n14709 & n18046 ) | ( n15839 & n18046 ) ;
  assign n18048 = n9186 ^ n8056 ^ n459 ;
  assign n18049 = n589 & ~n18048 ;
  assign n18050 = ( n2743 & n3173 ) | ( n2743 & n4205 ) | ( n3173 & n4205 ) ;
  assign n18051 = ( n13796 & n16613 ) | ( n13796 & n18050 ) | ( n16613 & n18050 ) ;
  assign n18053 = n1041 & n1326 ;
  assign n18054 = n16949 | n18053 ;
  assign n18052 = n1922 & ~n4403 ;
  assign n18055 = n18054 ^ n18052 ^ 1'b0 ;
  assign n18056 = n472 ^ n466 ^ x13 ;
  assign n18057 = n9498 & ~n17898 ;
  assign n18058 = n16771 & n18057 ;
  assign n18059 = ( ~n595 & n18056 ) | ( ~n595 & n18058 ) | ( n18056 & n18058 ) ;
  assign n18060 = n16778 ^ n5034 ^ 1'b0 ;
  assign n18061 = n7991 | n10770 ;
  assign n18062 = n14740 ^ n5425 ^ n876 ;
  assign n18063 = n10294 ^ n3617 ^ 1'b0 ;
  assign n18064 = ~n11594 & n18063 ;
  assign n18065 = n1554 & n10137 ;
  assign n18066 = n14018 & n18065 ;
  assign n18067 = n1160 | n18066 ;
  assign n18068 = n17480 | n18067 ;
  assign n18069 = n1994 & ~n3836 ;
  assign n18070 = ( n5185 & ~n11686 ) | ( n5185 & n18069 ) | ( ~n11686 & n18069 ) ;
  assign n18071 = n11603 | n18070 ;
  assign n18072 = ( ~n18064 & n18068 ) | ( ~n18064 & n18071 ) | ( n18068 & n18071 ) ;
  assign n18073 = ( n6464 & n18062 ) | ( n6464 & ~n18072 ) | ( n18062 & ~n18072 ) ;
  assign n18080 = n5342 ^ n5319 ^ n3671 ;
  assign n18075 = n1753 ^ n502 ^ 1'b0 ;
  assign n18076 = ( ~n222 & n579 ) | ( ~n222 & n18075 ) | ( n579 & n18075 ) ;
  assign n18077 = n18076 ^ n7294 ^ n7113 ;
  assign n18078 = ( n1694 & n3840 ) | ( n1694 & n18077 ) | ( n3840 & n18077 ) ;
  assign n18074 = n8940 ^ n7660 ^ 1'b0 ;
  assign n18079 = n18078 ^ n18074 ^ n16018 ;
  assign n18081 = n18080 ^ n18079 ^ 1'b0 ;
  assign n18082 = n9769 ^ n4666 ^ n2755 ;
  assign n18083 = ~n711 & n8120 ;
  assign n18084 = n4257 ^ n2548 ^ n1121 ;
  assign n18085 = n249 & ~n18084 ;
  assign n18086 = n6335 & n18085 ;
  assign n18087 = ( ~n12951 & n18083 ) | ( ~n12951 & n18086 ) | ( n18083 & n18086 ) ;
  assign n18088 = ( n243 & n18082 ) | ( n243 & n18087 ) | ( n18082 & n18087 ) ;
  assign n18089 = n2405 | n11543 ;
  assign n18090 = n4034 | n6661 ;
  assign n18091 = n5020 & ~n18090 ;
  assign n18092 = ( n9767 & ~n9861 ) | ( n9767 & n11335 ) | ( ~n9861 & n11335 ) ;
  assign n18093 = n18092 ^ n4387 ^ 1'b0 ;
  assign n18094 = n304 & ~n2238 ;
  assign n18095 = ~n5958 & n18094 ;
  assign n18096 = n1209 & ~n18095 ;
  assign n18097 = n4907 & n18096 ;
  assign n18098 = n18097 ^ n4113 ^ 1'b0 ;
  assign n18099 = ~n6158 & n18098 ;
  assign n18100 = ~n11212 & n18099 ;
  assign n18101 = ( n11200 & ~n14277 ) | ( n11200 & n18100 ) | ( ~n14277 & n18100 ) ;
  assign n18102 = n195 | n1423 ;
  assign n18103 = n6021 | n18102 ;
  assign n18104 = ( ~n10315 & n17695 ) | ( ~n10315 & n18103 ) | ( n17695 & n18103 ) ;
  assign n18105 = ( n457 & ~n1113 ) | ( n457 & n4639 ) | ( ~n1113 & n4639 ) ;
  assign n18106 = n18105 ^ n2795 ^ n2015 ;
  assign n18107 = ( x113 & n2737 ) | ( x113 & ~n18106 ) | ( n2737 & ~n18106 ) ;
  assign n18108 = ( n6223 & n13809 ) | ( n6223 & n18107 ) | ( n13809 & n18107 ) ;
  assign n18109 = n18108 ^ n4496 ^ 1'b0 ;
  assign n18110 = ( n3724 & n5268 ) | ( n3724 & n18109 ) | ( n5268 & n18109 ) ;
  assign n18111 = n6722 ^ n2692 ^ n2220 ;
  assign n18112 = ( n4214 & n7113 ) | ( n4214 & ~n18111 ) | ( n7113 & ~n18111 ) ;
  assign n18113 = n11711 ^ n3584 ^ 1'b0 ;
  assign n18114 = ( n3759 & ~n6361 ) | ( n3759 & n8403 ) | ( ~n6361 & n8403 ) ;
  assign n18115 = ( n3719 & n4085 ) | ( n3719 & ~n15728 ) | ( n4085 & ~n15728 ) ;
  assign n18119 = n9745 ^ n4480 ^ 1'b0 ;
  assign n18116 = n3928 ^ n1733 ^ 1'b0 ;
  assign n18117 = n1319 | n18116 ;
  assign n18118 = n18117 ^ n13045 ^ n2468 ;
  assign n18120 = n18119 ^ n18118 ^ n2845 ;
  assign n18121 = n10483 ^ n6630 ^ 1'b0 ;
  assign n18122 = n16031 & n18121 ;
  assign n18129 = n831 | n16327 ;
  assign n18123 = ( n2230 & n4497 ) | ( n2230 & n4600 ) | ( n4497 & n4600 ) ;
  assign n18124 = ( n2167 & n4920 ) | ( n2167 & n18123 ) | ( n4920 & n18123 ) ;
  assign n18125 = n6123 ^ n3455 ^ 1'b0 ;
  assign n18126 = n389 | n18125 ;
  assign n18127 = n869 & ~n18126 ;
  assign n18128 = n18124 & n18127 ;
  assign n18130 = n18129 ^ n18128 ^ n5443 ;
  assign n18131 = n18130 ^ n13336 ^ n8242 ;
  assign n18132 = n6913 ^ n1998 ^ n1122 ;
  assign n18133 = ( n3416 & ~n3460 ) | ( n3416 & n18132 ) | ( ~n3460 & n18132 ) ;
  assign n18134 = n5345 & ~n12398 ;
  assign n18135 = n18134 ^ n15527 ^ 1'b0 ;
  assign n18136 = n1948 | n18135 ;
  assign n18137 = n18136 ^ n12599 ^ 1'b0 ;
  assign n18138 = n7039 ^ n6223 ^ n3953 ;
  assign n18139 = n14761 & ~n18138 ;
  assign n18140 = n11177 | n18139 ;
  assign n18141 = n18140 ^ n11954 ^ 1'b0 ;
  assign n18142 = n16264 ^ n5219 ^ 1'b0 ;
  assign n18143 = n12221 & ~n18142 ;
  assign n18144 = ( n1835 & n15054 ) | ( n1835 & ~n16278 ) | ( n15054 & ~n16278 ) ;
  assign n18145 = n18144 ^ n12550 ^ n10412 ;
  assign n18146 = ( ~n3278 & n11370 ) | ( ~n3278 & n12833 ) | ( n11370 & n12833 ) ;
  assign n18147 = n10594 ^ n9351 ^ n1250 ;
  assign n18148 = n18147 ^ n7274 ^ n1830 ;
  assign n18149 = n18148 ^ n8434 ^ n3605 ;
  assign n18150 = ( n2426 & n14293 ) | ( n2426 & n18149 ) | ( n14293 & n18149 ) ;
  assign n18151 = n573 & ~n8152 ;
  assign n18152 = ~n14551 & n18151 ;
  assign n18153 = ( n2470 & n8653 ) | ( n2470 & ~n8842 ) | ( n8653 & ~n8842 ) ;
  assign n18154 = n17122 ^ n3318 ^ 1'b0 ;
  assign n18155 = n18154 ^ n10102 ^ n4283 ;
  assign n18156 = ( n18152 & ~n18153 ) | ( n18152 & n18155 ) | ( ~n18153 & n18155 ) ;
  assign n18157 = n15355 ^ n5763 ^ 1'b0 ;
  assign n18158 = ~n661 & n18157 ;
  assign n18159 = n18158 ^ n13048 ^ n7578 ;
  assign n18160 = n17362 ^ n3775 ^ n1440 ;
  assign n18161 = ( n748 & ~n18159 ) | ( n748 & n18160 ) | ( ~n18159 & n18160 ) ;
  assign n18162 = n4030 ^ n1632 ^ x22 ;
  assign n18163 = ( ~n2644 & n8881 ) | ( ~n2644 & n9216 ) | ( n8881 & n9216 ) ;
  assign n18164 = n5367 ^ n3008 ^ n2977 ;
  assign n18165 = n18164 ^ x36 ^ 1'b0 ;
  assign n18166 = n17953 & ~n18165 ;
  assign n18167 = ( n6848 & n18163 ) | ( n6848 & ~n18166 ) | ( n18163 & ~n18166 ) ;
  assign n18168 = ( n3270 & n10984 ) | ( n3270 & n18167 ) | ( n10984 & n18167 ) ;
  assign n18169 = n5493 & ~n18168 ;
  assign n18170 = n18169 ^ n1583 ^ 1'b0 ;
  assign n18172 = ( ~n1137 & n4564 ) | ( ~n1137 & n6720 ) | ( n4564 & n6720 ) ;
  assign n18171 = n14535 ^ n4962 ^ n1648 ;
  assign n18173 = n18172 ^ n18171 ^ n8741 ;
  assign n18174 = ( n2853 & n10162 ) | ( n2853 & n18173 ) | ( n10162 & n18173 ) ;
  assign n18175 = ( ~n5388 & n10053 ) | ( ~n5388 & n18174 ) | ( n10053 & n18174 ) ;
  assign n18176 = n15213 ^ n6582 ^ n404 ;
  assign n18178 = n12368 ^ n11825 ^ n6240 ;
  assign n18177 = n16357 ^ n12299 ^ n3801 ;
  assign n18179 = n18178 ^ n18177 ^ n1585 ;
  assign n18180 = n18179 ^ n12599 ^ n8906 ;
  assign n18181 = n5527 | n13051 ;
  assign n18182 = n18181 ^ n9691 ^ 1'b0 ;
  assign n18183 = n4754 ^ n2492 ^ 1'b0 ;
  assign n18184 = n13365 & ~n18183 ;
  assign n18185 = ~n1536 & n3197 ;
  assign n18186 = n18184 & ~n18185 ;
  assign n18187 = n5516 & n18186 ;
  assign n18188 = ( ~n4855 & n7636 ) | ( ~n4855 & n13768 ) | ( n7636 & n13768 ) ;
  assign n18189 = ( ~n644 & n10237 ) | ( ~n644 & n16771 ) | ( n10237 & n16771 ) ;
  assign n18190 = n17740 ^ n8860 ^ 1'b0 ;
  assign n18191 = n18190 ^ n9421 ^ n8316 ;
  assign n18192 = n13781 ^ n10864 ^ n5556 ;
  assign n18193 = n18192 ^ n6872 ^ n3319 ;
  assign n18197 = n8337 ^ n4264 ^ n228 ;
  assign n18198 = n6423 | n18197 ;
  assign n18199 = ~n5109 & n10306 ;
  assign n18200 = ~n18198 & n18199 ;
  assign n18194 = n5329 ^ n5279 ^ n4122 ;
  assign n18195 = ( n2395 & n2697 ) | ( n2395 & ~n18194 ) | ( n2697 & ~n18194 ) ;
  assign n18196 = n18195 ^ n4360 ^ n3518 ;
  assign n18201 = n18200 ^ n18196 ^ n11023 ;
  assign n18202 = ( n1285 & n4860 ) | ( n1285 & ~n10868 ) | ( n4860 & ~n10868 ) ;
  assign n18203 = n8142 ^ n2897 ^ n2879 ;
  assign n18206 = n7157 ^ n2702 ^ n817 ;
  assign n18207 = n2511 & n18206 ;
  assign n18208 = ( n1171 & n8731 ) | ( n1171 & ~n18207 ) | ( n8731 & ~n18207 ) ;
  assign n18209 = ( ~n3590 & n8609 ) | ( ~n3590 & n18208 ) | ( n8609 & n18208 ) ;
  assign n18204 = ~n725 & n5735 ;
  assign n18205 = n6899 & ~n18204 ;
  assign n18210 = n18209 ^ n18205 ^ n9268 ;
  assign n18211 = ( n2168 & ~n2548 ) | ( n2168 & n12862 ) | ( ~n2548 & n12862 ) ;
  assign n18212 = ( x28 & n5055 ) | ( x28 & ~n18211 ) | ( n5055 & ~n18211 ) ;
  assign n18213 = n18212 ^ n11892 ^ n3879 ;
  assign n18214 = n18213 ^ n4601 ^ 1'b0 ;
  assign n18215 = ( n18203 & n18210 ) | ( n18203 & ~n18214 ) | ( n18210 & ~n18214 ) ;
  assign n18225 = n3444 ^ n3240 ^ n2068 ;
  assign n18220 = n9276 ^ n7654 ^ n6770 ;
  assign n18221 = n18220 ^ n4477 ^ n2558 ;
  assign n18222 = ( ~n3796 & n11965 ) | ( ~n3796 & n18221 ) | ( n11965 & n18221 ) ;
  assign n18223 = ( n2688 & ~n13865 ) | ( n2688 & n18222 ) | ( ~n13865 & n18222 ) ;
  assign n18224 = ( n6447 & ~n13652 ) | ( n6447 & n18223 ) | ( ~n13652 & n18223 ) ;
  assign n18217 = ( n8338 & n12075 ) | ( n8338 & ~n12983 ) | ( n12075 & ~n12983 ) ;
  assign n18216 = n1982 & ~n1998 ;
  assign n18218 = n18217 ^ n18216 ^ 1'b0 ;
  assign n18219 = ( n1849 & n14055 ) | ( n1849 & n18218 ) | ( n14055 & n18218 ) ;
  assign n18226 = n18225 ^ n18224 ^ n18219 ;
  assign n18227 = n11015 ^ n8192 ^ n3825 ;
  assign n18228 = ( n3498 & n4422 ) | ( n3498 & ~n13524 ) | ( n4422 & ~n13524 ) ;
  assign n18232 = n10053 ^ n5166 ^ n1447 ;
  assign n18229 = n9131 ^ n6139 ^ n258 ;
  assign n18230 = n16799 ^ n8661 ^ 1'b0 ;
  assign n18231 = ~n18229 & n18230 ;
  assign n18233 = n18232 ^ n18231 ^ n17557 ;
  assign n18234 = n1243 & ~n8469 ;
  assign n18235 = n2494 | n14958 ;
  assign n18236 = ( n3626 & n18234 ) | ( n3626 & ~n18235 ) | ( n18234 & ~n18235 ) ;
  assign n18237 = ( n242 & ~n7086 ) | ( n242 & n18236 ) | ( ~n7086 & n18236 ) ;
  assign n18238 = n14270 ^ n5551 ^ n5005 ;
  assign n18239 = n18238 ^ n5554 ^ 1'b0 ;
  assign n18240 = n18239 ^ n12661 ^ n8306 ;
  assign n18241 = n18240 ^ n6401 ^ 1'b0 ;
  assign n18242 = n11865 ^ n3508 ^ 1'b0 ;
  assign n18243 = n2353 | n11285 ;
  assign n18244 = n18243 ^ n6040 ^ 1'b0 ;
  assign n18245 = n18244 ^ n17655 ^ 1'b0 ;
  assign n18246 = ( ~n1352 & n3067 ) | ( ~n1352 & n10266 ) | ( n3067 & n10266 ) ;
  assign n18247 = ~n4121 & n11595 ;
  assign n18248 = ~n3876 & n18247 ;
  assign n18249 = n18248 ^ n9932 ^ n4091 ;
  assign n18250 = n18249 ^ n4885 ^ n345 ;
  assign n18251 = ~n14329 & n18250 ;
  assign n18254 = n13378 ^ n3617 ^ 1'b0 ;
  assign n18255 = ~n9148 & n18254 ;
  assign n18252 = n13617 ^ n7956 ^ n160 ;
  assign n18253 = ~n9710 & n18252 ;
  assign n18256 = n18255 ^ n18253 ^ 1'b0 ;
  assign n18257 = n18256 ^ n12781 ^ n9552 ;
  assign n18258 = n3637 & n10379 ;
  assign n18259 = n10073 ^ n3028 ^ n2845 ;
  assign n18260 = ( ~n15828 & n18258 ) | ( ~n15828 & n18259 ) | ( n18258 & n18259 ) ;
  assign n18261 = n18260 ^ n15469 ^ n11502 ;
  assign n18262 = x84 & n6777 ;
  assign n18263 = ~n7660 & n18262 ;
  assign n18264 = n18263 ^ n10856 ^ n10010 ;
  assign n18265 = n18264 ^ n4167 ^ n333 ;
  assign n18266 = n5338 & ~n9903 ;
  assign n18267 = n18266 ^ n11480 ^ 1'b0 ;
  assign n18268 = n18267 ^ n12152 ^ n10438 ;
  assign n18269 = ( n2909 & n17869 ) | ( n2909 & n18268 ) | ( n17869 & n18268 ) ;
  assign n18272 = n5333 | n13034 ;
  assign n18273 = n5443 & ~n18272 ;
  assign n18274 = n5562 ^ n4914 ^ n1645 ;
  assign n18275 = ( n9447 & ~n12575 ) | ( n9447 & n18274 ) | ( ~n12575 & n18274 ) ;
  assign n18276 = ( n10827 & n18273 ) | ( n10827 & n18275 ) | ( n18273 & n18275 ) ;
  assign n18270 = n8285 ^ n5648 ^ n2358 ;
  assign n18271 = n16574 & ~n18270 ;
  assign n18277 = n18276 ^ n18271 ^ 1'b0 ;
  assign n18279 = ( n1188 & n4337 ) | ( n1188 & ~n17234 ) | ( n4337 & ~n17234 ) ;
  assign n18280 = ( n11354 & n13394 ) | ( n11354 & n18279 ) | ( n13394 & n18279 ) ;
  assign n18281 = n11304 ^ n10085 ^ n3340 ;
  assign n18282 = ( ~n6241 & n15873 ) | ( ~n6241 & n18281 ) | ( n15873 & n18281 ) ;
  assign n18283 = ( n13613 & n18280 ) | ( n13613 & ~n18282 ) | ( n18280 & ~n18282 ) ;
  assign n18278 = n14721 & n15998 ;
  assign n18284 = n18283 ^ n18278 ^ 1'b0 ;
  assign n18285 = ( n1478 & ~n6535 ) | ( n1478 & n9994 ) | ( ~n6535 & n9994 ) ;
  assign n18286 = ( n1212 & ~n1604 ) | ( n1212 & n15861 ) | ( ~n1604 & n15861 ) ;
  assign n18287 = ( n4322 & ~n7264 ) | ( n4322 & n15854 ) | ( ~n7264 & n15854 ) ;
  assign n18288 = ( n4982 & ~n10849 ) | ( n4982 & n16209 ) | ( ~n10849 & n16209 ) ;
  assign n18289 = n18288 ^ n14358 ^ n2259 ;
  assign n18290 = n1803 & ~n12842 ;
  assign n18291 = n18290 ^ n13345 ^ 1'b0 ;
  assign n18292 = n13160 ^ n11699 ^ n11675 ;
  assign n18293 = n14541 ^ n3791 ^ n3142 ;
  assign n18294 = n18292 & n18293 ;
  assign n18295 = ~n603 & n12695 ;
  assign n18296 = n7029 & n18295 ;
  assign n18297 = n6950 & n7849 ;
  assign n18298 = n18297 ^ n15116 ^ 1'b0 ;
  assign n18299 = n2849 & n18298 ;
  assign n18300 = ( n4663 & ~n18296 ) | ( n4663 & n18299 ) | ( ~n18296 & n18299 ) ;
  assign n18301 = ( ~n560 & n3186 ) | ( ~n560 & n17232 ) | ( n3186 & n17232 ) ;
  assign n18302 = ( ~n7143 & n12177 ) | ( ~n7143 & n18301 ) | ( n12177 & n18301 ) ;
  assign n18303 = n16521 ^ n1010 ^ x24 ;
  assign n18304 = n18303 ^ n6738 ^ n579 ;
  assign n18305 = ( ~n2533 & n17470 ) | ( ~n2533 & n18304 ) | ( n17470 & n18304 ) ;
  assign n18306 = ( n3996 & n6793 ) | ( n3996 & ~n9657 ) | ( n6793 & ~n9657 ) ;
  assign n18307 = ( ~n6032 & n13010 ) | ( ~n6032 & n18306 ) | ( n13010 & n18306 ) ;
  assign n18308 = n1158 & n18307 ;
  assign n18309 = n18308 ^ n9967 ^ 1'b0 ;
  assign n18310 = ~n4292 & n10406 ;
  assign n18311 = n18310 ^ n3716 ^ 1'b0 ;
  assign n18312 = n18311 ^ n17594 ^ n6013 ;
  assign n18313 = n18312 ^ n9398 ^ n7124 ;
  assign n18314 = ( n2064 & n5404 ) | ( n2064 & ~n11152 ) | ( n5404 & ~n11152 ) ;
  assign n18315 = ( n11132 & ~n13117 ) | ( n11132 & n18314 ) | ( ~n13117 & n18314 ) ;
  assign n18316 = ( n2644 & n9259 ) | ( n2644 & ~n14329 ) | ( n9259 & ~n14329 ) ;
  assign n18317 = ( ~n5219 & n5818 ) | ( ~n5219 & n12059 ) | ( n5818 & n12059 ) ;
  assign n18318 = ( n3876 & n4762 ) | ( n3876 & n18317 ) | ( n4762 & n18317 ) ;
  assign n18319 = n18318 ^ n17127 ^ n7771 ;
  assign n18320 = ( n14817 & ~n18316 ) | ( n14817 & n18319 ) | ( ~n18316 & n18319 ) ;
  assign n18321 = ( n233 & n8766 ) | ( n233 & n17374 ) | ( n8766 & n17374 ) ;
  assign n18322 = n15697 ^ n12506 ^ 1'b0 ;
  assign n18323 = n16150 ^ n4428 ^ 1'b0 ;
  assign n18324 = n18323 ^ n9405 ^ 1'b0 ;
  assign n18325 = ( n1732 & ~n2508 ) | ( n1732 & n8920 ) | ( ~n2508 & n8920 ) ;
  assign n18330 = n2392 & n11537 ;
  assign n18326 = n8577 ^ n4156 ^ 1'b0 ;
  assign n18327 = n5795 & ~n18326 ;
  assign n18328 = n18327 ^ n14745 ^ n14559 ;
  assign n18329 = n18328 ^ n6059 ^ n878 ;
  assign n18331 = n18330 ^ n18329 ^ 1'b0 ;
  assign n18332 = ( n2406 & n18325 ) | ( n2406 & n18331 ) | ( n18325 & n18331 ) ;
  assign n18333 = n16390 ^ n6016 ^ n5415 ;
  assign n18335 = n2135 & ~n2433 ;
  assign n18336 = n9455 | n18335 ;
  assign n18334 = ( n2000 & ~n4079 ) | ( n2000 & n15887 ) | ( ~n4079 & n15887 ) ;
  assign n18337 = n18336 ^ n18334 ^ n6884 ;
  assign n18338 = n4017 & ~n18337 ;
  assign n18339 = ~n2070 & n18338 ;
  assign n18340 = n3451 | n18339 ;
  assign n18341 = n15276 | n18340 ;
  assign n18342 = n17809 ^ n2806 ^ 1'b0 ;
  assign n18343 = n18342 ^ n4058 ^ 1'b0 ;
  assign n18344 = ( n3748 & ~n4108 ) | ( n3748 & n5576 ) | ( ~n4108 & n5576 ) ;
  assign n18345 = ( ~n1045 & n12018 ) | ( ~n1045 & n18344 ) | ( n12018 & n18344 ) ;
  assign n18346 = ( n223 & n5662 ) | ( n223 & ~n6626 ) | ( n5662 & ~n6626 ) ;
  assign n18347 = ( n1767 & n6827 ) | ( n1767 & ~n18346 ) | ( n6827 & ~n18346 ) ;
  assign n18348 = n5970 | n9080 ;
  assign n18349 = ( ~n8883 & n9941 ) | ( ~n8883 & n18348 ) | ( n9941 & n18348 ) ;
  assign n18350 = n18349 ^ n15928 ^ n1024 ;
  assign n18351 = n1626 ^ n857 ^ 1'b0 ;
  assign n18352 = ( n567 & n14819 ) | ( n567 & n18351 ) | ( n14819 & n18351 ) ;
  assign n18353 = ( n7486 & n9222 ) | ( n7486 & ~n18352 ) | ( n9222 & ~n18352 ) ;
  assign n18354 = ( n14187 & n18350 ) | ( n14187 & ~n18353 ) | ( n18350 & ~n18353 ) ;
  assign n18355 = ( n18345 & n18347 ) | ( n18345 & n18354 ) | ( n18347 & n18354 ) ;
  assign n18356 = n18355 ^ n10091 ^ n8309 ;
  assign n18357 = n13113 ^ n3838 ^ n244 ;
  assign n18358 = n8303 ^ n5100 ^ n2634 ;
  assign n18359 = n18117 ^ n12187 ^ n12083 ;
  assign n18360 = ( n18357 & n18358 ) | ( n18357 & n18359 ) | ( n18358 & n18359 ) ;
  assign n18361 = n12650 & ~n14239 ;
  assign n18362 = n991 & n1711 ;
  assign n18363 = n18362 ^ n1538 ^ 1'b0 ;
  assign n18364 = n18363 ^ n6115 ^ 1'b0 ;
  assign n18366 = n17329 ^ n12802 ^ n10143 ;
  assign n18365 = ~n14217 & n16139 ;
  assign n18367 = n18366 ^ n18365 ^ n4557 ;
  assign n18368 = n18367 ^ n15577 ^ n9717 ;
  assign n18369 = n18368 ^ n12030 ^ n7841 ;
  assign n18375 = ( n5038 & n8399 ) | ( n5038 & n12217 ) | ( n8399 & n12217 ) ;
  assign n18376 = ~n16909 & n18375 ;
  assign n18372 = n12521 ^ n6396 ^ 1'b0 ;
  assign n18373 = n3301 & ~n18372 ;
  assign n18370 = ( n3940 & ~n8963 ) | ( n3940 & n18357 ) | ( ~n8963 & n18357 ) ;
  assign n18371 = ( n3685 & n4450 ) | ( n3685 & n18370 ) | ( n4450 & n18370 ) ;
  assign n18374 = n18373 ^ n18371 ^ n2960 ;
  assign n18377 = n18376 ^ n18374 ^ n15250 ;
  assign n18378 = ~n5444 & n18377 ;
  assign n18380 = n3434 & ~n5464 ;
  assign n18381 = n18380 ^ n15405 ^ 1'b0 ;
  assign n18379 = ( ~n4249 & n9094 ) | ( ~n4249 & n11545 ) | ( n9094 & n11545 ) ;
  assign n18382 = n18381 ^ n18379 ^ n7932 ;
  assign n18383 = n17594 ^ n3625 ^ 1'b0 ;
  assign n18384 = ~n6302 & n18383 ;
  assign n18385 = ~n2371 & n18384 ;
  assign n18388 = ( ~n2094 & n9345 ) | ( ~n2094 & n12842 ) | ( n9345 & n12842 ) ;
  assign n18386 = n14387 ^ n8455 ^ n5290 ;
  assign n18387 = n18386 ^ n1902 ^ n1499 ;
  assign n18389 = n18388 ^ n18387 ^ n12979 ;
  assign n18390 = ( n442 & ~n1084 ) | ( n442 & n8773 ) | ( ~n1084 & n8773 ) ;
  assign n18391 = n18390 ^ n14250 ^ 1'b0 ;
  assign n18392 = ~n16348 & n18391 ;
  assign n18393 = n8203 ^ n1949 ^ n1409 ;
  assign n18394 = n16527 ^ n7634 ^ 1'b0 ;
  assign n18395 = n18393 & n18394 ;
  assign n18405 = n1401 & ~n2932 ;
  assign n18406 = n11157 ^ n6641 ^ 1'b0 ;
  assign n18407 = ~n18405 & n18406 ;
  assign n18408 = n18407 ^ n4236 ^ 1'b0 ;
  assign n18403 = n7449 ^ n4502 ^ 1'b0 ;
  assign n18404 = n18403 ^ n14811 ^ 1'b0 ;
  assign n18396 = n14547 ^ n5959 ^ n2200 ;
  assign n18398 = ( x66 & n3146 ) | ( x66 & ~n15340 ) | ( n3146 & ~n15340 ) ;
  assign n18397 = n14284 ^ n4798 ^ x105 ;
  assign n18399 = n18398 ^ n18397 ^ n12469 ;
  assign n18400 = n7812 ^ n5163 ^ n1548 ;
  assign n18401 = n8620 & ~n18400 ;
  assign n18402 = ( n18396 & ~n18399 ) | ( n18396 & n18401 ) | ( ~n18399 & n18401 ) ;
  assign n18409 = n18408 ^ n18404 ^ n18402 ;
  assign n18410 = n17414 ^ n11516 ^ n9409 ;
  assign n18411 = n9665 ^ n5303 ^ n357 ;
  assign n18412 = n1550 ^ n289 ^ 1'b0 ;
  assign n18413 = n18411 & n18412 ;
  assign n18414 = n18413 ^ n15191 ^ 1'b0 ;
  assign n18415 = n18414 ^ n17530 ^ n12245 ;
  assign n18416 = n10994 ^ n3116 ^ n1263 ;
  assign n18417 = n18416 ^ n3319 ^ 1'b0 ;
  assign n18419 = ( n1883 & n9919 ) | ( n1883 & ~n13708 ) | ( n9919 & ~n13708 ) ;
  assign n18418 = n4729 ^ n2026 ^ 1'b0 ;
  assign n18420 = n18419 ^ n18418 ^ n3966 ;
  assign n18421 = ( n1338 & n1834 ) | ( n1338 & n13913 ) | ( n1834 & n13913 ) ;
  assign n18422 = n13715 ^ n6228 ^ n3103 ;
  assign n18423 = n18422 ^ n14638 ^ 1'b0 ;
  assign n18424 = ( ~n2450 & n5285 ) | ( ~n2450 & n12366 ) | ( n5285 & n12366 ) ;
  assign n18425 = n18424 ^ n15714 ^ n11674 ;
  assign n18426 = ( n716 & n12323 ) | ( n716 & n18425 ) | ( n12323 & n18425 ) ;
  assign n18427 = n16875 | n18426 ;
  assign n18428 = n18423 | n18427 ;
  assign n18429 = n10244 ^ n9761 ^ 1'b0 ;
  assign n18430 = ~n12407 & n18429 ;
  assign n18431 = ( n3429 & n11898 ) | ( n3429 & ~n15216 ) | ( n11898 & ~n15216 ) ;
  assign n18432 = n6130 ^ n3566 ^ 1'b0 ;
  assign n18433 = n17709 & ~n18432 ;
  assign n18434 = n18433 ^ n13813 ^ n4225 ;
  assign n18435 = n7333 ^ n6925 ^ n3689 ;
  assign n18436 = n4065 ^ n3631 ^ n1089 ;
  assign n18437 = ( ~n7963 & n18435 ) | ( ~n7963 & n18436 ) | ( n18435 & n18436 ) ;
  assign n18438 = ( ~n229 & n6425 ) | ( ~n229 & n18437 ) | ( n6425 & n18437 ) ;
  assign n18439 = n18438 ^ n14130 ^ n8533 ;
  assign n18440 = n6691 ^ n2813 ^ n648 ;
  assign n18441 = n18440 ^ n5351 ^ 1'b0 ;
  assign n18442 = ( n6042 & n7561 ) | ( n6042 & ~n8672 ) | ( n7561 & ~n8672 ) ;
  assign n18443 = n9407 ^ n6180 ^ n6111 ;
  assign n18444 = n18443 ^ n2150 ^ 1'b0 ;
  assign n18445 = ~n13405 & n18444 ;
  assign n18446 = ( n748 & ~n3502 ) | ( n748 & n5352 ) | ( ~n3502 & n5352 ) ;
  assign n18447 = n18446 ^ n9367 ^ n439 ;
  assign n18448 = ( ~n6712 & n9412 ) | ( ~n6712 & n18447 ) | ( n9412 & n18447 ) ;
  assign n18449 = n18448 ^ n14275 ^ n12002 ;
  assign n18450 = ( n1950 & ~n11768 ) | ( n1950 & n15013 ) | ( ~n11768 & n15013 ) ;
  assign n18451 = n18296 ^ n8160 ^ n908 ;
  assign n18452 = ( n460 & n10814 ) | ( n460 & n18451 ) | ( n10814 & n18451 ) ;
  assign n18453 = ( ~n18449 & n18450 ) | ( ~n18449 & n18452 ) | ( n18450 & n18452 ) ;
  assign n18454 = ~n3629 & n11868 ;
  assign n18455 = ~n12936 & n18454 ;
  assign n18456 = ( ~n2558 & n8463 ) | ( ~n2558 & n18455 ) | ( n8463 & n18455 ) ;
  assign n18457 = ( n15169 & n17581 ) | ( n15169 & n18456 ) | ( n17581 & n18456 ) ;
  assign n18460 = n9958 ^ n4035 ^ n3403 ;
  assign n18458 = n10065 ^ n7908 ^ n5326 ;
  assign n18459 = n18458 ^ n15519 ^ n3794 ;
  assign n18461 = n18460 ^ n18459 ^ n9564 ;
  assign n18462 = n17600 ^ n11093 ^ n394 ;
  assign n18463 = n7122 ^ n4956 ^ 1'b0 ;
  assign n18464 = n4106 & ~n18463 ;
  assign n18465 = ( n17852 & n18462 ) | ( n17852 & ~n18464 ) | ( n18462 & ~n18464 ) ;
  assign n18466 = n2825 & ~n5645 ;
  assign n18467 = n8689 & n18466 ;
  assign n18468 = n7831 ^ n1981 ^ n743 ;
  assign n18469 = n18468 ^ n10736 ^ n9898 ;
  assign n18470 = ( n3215 & ~n9436 ) | ( n3215 & n18469 ) | ( ~n9436 & n18469 ) ;
  assign n18471 = ( n2591 & n18467 ) | ( n2591 & ~n18470 ) | ( n18467 & ~n18470 ) ;
  assign n18472 = n5700 ^ n4538 ^ 1'b0 ;
  assign n18473 = n3010 & ~n18472 ;
  assign n18474 = ~n7804 & n15822 ;
  assign n18475 = ( n2477 & n13077 ) | ( n2477 & n13787 ) | ( n13077 & n13787 ) ;
  assign n18476 = n18475 ^ n17756 ^ n7771 ;
  assign n18477 = n16416 ^ n15660 ^ n11982 ;
  assign n18478 = n14021 ^ n11601 ^ n8106 ;
  assign n18479 = n7525 ^ n2190 ^ 1'b0 ;
  assign n18480 = n18479 ^ n4104 ^ 1'b0 ;
  assign n18481 = n8850 | n18480 ;
  assign n18482 = n2640 & n3429 ;
  assign n18483 = n2019 & n18482 ;
  assign n18484 = n18483 ^ n17854 ^ 1'b0 ;
  assign n18485 = n12341 & n18484 ;
  assign n18486 = n4476 & n9487 ;
  assign n18487 = ( n18403 & n18485 ) | ( n18403 & n18486 ) | ( n18485 & n18486 ) ;
  assign n18488 = ( n5344 & n15134 ) | ( n5344 & ~n18487 ) | ( n15134 & ~n18487 ) ;
  assign n18489 = n11173 ^ n10472 ^ 1'b0 ;
  assign n18490 = ~n985 & n18489 ;
  assign n18491 = n18490 ^ n10171 ^ n8924 ;
  assign n18492 = ( n379 & n5117 ) | ( n379 & ~n18491 ) | ( n5117 & ~n18491 ) ;
  assign n18493 = n18492 ^ n6130 ^ n5276 ;
  assign n18494 = n2837 ^ n1940 ^ x21 ;
  assign n18495 = ( n1019 & ~n3568 ) | ( n1019 & n18494 ) | ( ~n3568 & n18494 ) ;
  assign n18496 = ( n475 & ~n14429 ) | ( n475 & n18495 ) | ( ~n14429 & n18495 ) ;
  assign n18497 = ~n5334 & n14375 ;
  assign n18498 = n1544 & n18497 ;
  assign n18499 = ~n6521 & n10136 ;
  assign n18500 = n18499 ^ n3499 ^ 1'b0 ;
  assign n18501 = n18500 ^ n8936 ^ n1678 ;
  assign n18502 = n15739 & n18501 ;
  assign n18503 = n18502 ^ n8936 ^ 1'b0 ;
  assign n18504 = n3771 | n18503 ;
  assign n18505 = ( ~n4332 & n4482 ) | ( ~n4332 & n17027 ) | ( n4482 & n17027 ) ;
  assign n18506 = n2914 ^ n1249 ^ n334 ;
  assign n18507 = ( n12955 & n15144 ) | ( n12955 & n18506 ) | ( n15144 & n18506 ) ;
  assign n18508 = n18507 ^ n4364 ^ 1'b0 ;
  assign n18509 = ( n3959 & n5657 ) | ( n3959 & ~n7198 ) | ( n5657 & ~n7198 ) ;
  assign n18510 = n9561 | n18509 ;
  assign n18511 = ( n5702 & n7392 ) | ( n5702 & n18510 ) | ( n7392 & n18510 ) ;
  assign n18512 = n18511 ^ n4919 ^ n4918 ;
  assign n18513 = n12031 ^ n1160 ^ n179 ;
  assign n18514 = ( n6423 & n7967 ) | ( n6423 & n18513 ) | ( n7967 & n18513 ) ;
  assign n18515 = ( n3204 & n9344 ) | ( n3204 & ~n18514 ) | ( n9344 & ~n18514 ) ;
  assign n18516 = n18515 ^ n10706 ^ n743 ;
  assign n18517 = ( ~n4207 & n12217 ) | ( ~n4207 & n15531 ) | ( n12217 & n15531 ) ;
  assign n18518 = n18517 ^ n12872 ^ n5383 ;
  assign n18519 = n13596 ^ n8629 ^ n1239 ;
  assign n18520 = n9717 ^ n8004 ^ n3923 ;
  assign n18521 = n14464 ^ n2866 ^ 1'b0 ;
  assign n18522 = n9104 & ~n18521 ;
  assign n18523 = n8694 ^ n8253 ^ n2997 ;
  assign n18524 = n18523 ^ n15801 ^ n5838 ;
  assign n18525 = n3050 & ~n3478 ;
  assign n18526 = ~n2484 & n13664 ;
  assign n18527 = n18526 ^ n15150 ^ n9632 ;
  assign n18528 = n12988 ^ n8552 ^ 1'b0 ;
  assign n18529 = n4210 & n18528 ;
  assign n18530 = ~n4761 & n18529 ;
  assign n18531 = ~n6575 & n18530 ;
  assign n18532 = ( n5736 & n18527 ) | ( n5736 & ~n18531 ) | ( n18527 & ~n18531 ) ;
  assign n18533 = ( n7730 & n9965 ) | ( n7730 & n13141 ) | ( n9965 & n13141 ) ;
  assign n18534 = ~n868 & n1954 ;
  assign n18535 = ( n1897 & n7564 ) | ( n1897 & n18534 ) | ( n7564 & n18534 ) ;
  assign n18536 = n18535 ^ n7051 ^ n6889 ;
  assign n18537 = n8547 | n18536 ;
  assign n18538 = n18537 ^ n278 ^ 1'b0 ;
  assign n18541 = ( n1257 & n7254 ) | ( n1257 & n9218 ) | ( n7254 & n9218 ) ;
  assign n18539 = n11810 & n12695 ;
  assign n18540 = n18539 ^ n6778 ^ 1'b0 ;
  assign n18542 = n18541 ^ n18540 ^ 1'b0 ;
  assign n18543 = n12231 ^ n11687 ^ n7730 ;
  assign n18545 = n4463 ^ n3579 ^ 1'b0 ;
  assign n18544 = n9777 & ~n10390 ;
  assign n18546 = n18545 ^ n18544 ^ 1'b0 ;
  assign n18547 = n2196 | n3936 ;
  assign n18548 = n1939 & ~n18547 ;
  assign n18549 = n18548 ^ n5950 ^ 1'b0 ;
  assign n18550 = n18546 & n18549 ;
  assign n18551 = ( n1000 & n13962 ) | ( n1000 & ~n18550 ) | ( n13962 & ~n18550 ) ;
  assign n18552 = ( n1927 & ~n13960 ) | ( n1927 & n16827 ) | ( ~n13960 & n16827 ) ;
  assign n18558 = n2202 & ~n7763 ;
  assign n18557 = ( ~n558 & n3905 ) | ( ~n558 & n15784 ) | ( n3905 & n15784 ) ;
  assign n18559 = n18558 ^ n18557 ^ 1'b0 ;
  assign n18560 = n18559 ^ n12930 ^ n1169 ;
  assign n18561 = n18560 ^ n16332 ^ n3794 ;
  assign n18553 = n16098 ^ n10445 ^ n2455 ;
  assign n18554 = n6626 ^ n2022 ^ n179 ;
  assign n18555 = ( n3511 & n15568 ) | ( n3511 & ~n18554 ) | ( n15568 & ~n18554 ) ;
  assign n18556 = ~n18553 & n18555 ;
  assign n18562 = n18561 ^ n18556 ^ 1'b0 ;
  assign n18564 = n13870 ^ n4966 ^ n3210 ;
  assign n18563 = n17917 ^ n16889 ^ n13856 ;
  assign n18565 = n18564 ^ n18563 ^ n12897 ;
  assign n18566 = n2239 & ~n4287 ;
  assign n18567 = n18566 ^ n6268 ^ 1'b0 ;
  assign n18568 = ( n421 & n697 ) | ( n421 & ~n17026 ) | ( n697 & ~n17026 ) ;
  assign n18569 = n1322 | n18568 ;
  assign n18570 = n12005 & ~n18569 ;
  assign n18571 = n335 & ~n4013 ;
  assign n18572 = n18571 ^ n2231 ^ 1'b0 ;
  assign n18573 = ~n2484 & n18572 ;
  assign n18574 = n18573 ^ n6446 ^ n141 ;
  assign n18575 = n18574 ^ n16152 ^ x101 ;
  assign n18576 = n437 & n4191 ;
  assign n18577 = n8856 & n18576 ;
  assign n18578 = ( n2666 & n13025 ) | ( n2666 & ~n18577 ) | ( n13025 & ~n18577 ) ;
  assign n18579 = n10347 ^ n2985 ^ 1'b0 ;
  assign n18580 = ( n6050 & ~n16388 ) | ( n6050 & n18579 ) | ( ~n16388 & n18579 ) ;
  assign n18581 = n12118 ^ n1246 ^ 1'b0 ;
  assign n18582 = n18581 ^ n17037 ^ 1'b0 ;
  assign n18583 = n6579 & ~n18582 ;
  assign n18584 = ( n11871 & ~n11944 ) | ( n11871 & n14140 ) | ( ~n11944 & n14140 ) ;
  assign n18585 = ( n8148 & ~n10701 ) | ( n8148 & n18584 ) | ( ~n10701 & n18584 ) ;
  assign n18588 = n9458 ^ n6869 ^ n4055 ;
  assign n18589 = ~n1087 & n18588 ;
  assign n18586 = n2780 & ~n9376 ;
  assign n18587 = n18586 ^ n6158 ^ 1'b0 ;
  assign n18590 = n18589 ^ n18587 ^ n15523 ;
  assign n18591 = n18585 | n18590 ;
  assign n18592 = n18591 ^ n7888 ^ 1'b0 ;
  assign n18593 = n14449 ^ n3634 ^ n1351 ;
  assign n18594 = ( n4778 & n5963 ) | ( n4778 & ~n13786 ) | ( n5963 & ~n13786 ) ;
  assign n18595 = ( n4398 & ~n8524 ) | ( n4398 & n14353 ) | ( ~n8524 & n14353 ) ;
  assign n18596 = n8496 ^ n6640 ^ n4834 ;
  assign n18597 = n12050 ^ n2988 ^ n739 ;
  assign n18598 = ( n18595 & n18596 ) | ( n18595 & ~n18597 ) | ( n18596 & ~n18597 ) ;
  assign n18601 = ( n4924 & n12092 ) | ( n4924 & n17442 ) | ( n12092 & n17442 ) ;
  assign n18602 = n2895 & n18601 ;
  assign n18603 = ~n2367 & n18602 ;
  assign n18599 = ( n176 & n1453 ) | ( n176 & ~n4000 ) | ( n1453 & ~n4000 ) ;
  assign n18600 = ( n4118 & n12051 ) | ( n4118 & n18599 ) | ( n12051 & n18599 ) ;
  assign n18604 = n18603 ^ n18600 ^ n14936 ;
  assign n18605 = n4078 ^ n2418 ^ n2260 ;
  assign n18613 = n12852 ^ n1586 ^ n1340 ;
  assign n18614 = n18613 ^ n6198 ^ n1743 ;
  assign n18610 = ( n5744 & n9153 ) | ( n5744 & n14738 ) | ( n9153 & n14738 ) ;
  assign n18606 = ( n7897 & n7993 ) | ( n7897 & ~n12672 ) | ( n7993 & ~n12672 ) ;
  assign n18607 = n18606 ^ n16321 ^ 1'b0 ;
  assign n18608 = n1340 & n18607 ;
  assign n18609 = ~n14325 & n18608 ;
  assign n18611 = n18610 ^ n18609 ^ 1'b0 ;
  assign n18612 = n7736 & n18611 ;
  assign n18615 = n18614 ^ n18612 ^ 1'b0 ;
  assign n18616 = ( n195 & n1244 ) | ( n195 & n1897 ) | ( n1244 & n1897 ) ;
  assign n18617 = n18616 ^ n658 ^ 1'b0 ;
  assign n18618 = n18617 ^ n8313 ^ n2493 ;
  assign n18619 = n5349 | n10140 ;
  assign n18620 = ( n1642 & ~n18618 ) | ( n1642 & n18619 ) | ( ~n18618 & n18619 ) ;
  assign n18626 = n18213 ^ n1505 ^ n609 ;
  assign n18621 = n3363 ^ n701 ^ n285 ;
  assign n18622 = n7514 & ~n16025 ;
  assign n18623 = n18622 ^ n6992 ^ 1'b0 ;
  assign n18624 = n805 | n18623 ;
  assign n18625 = n18621 & ~n18624 ;
  assign n18627 = n18626 ^ n18625 ^ n17298 ;
  assign n18628 = n13604 ^ n5692 ^ n4079 ;
  assign n18629 = n3064 & ~n5923 ;
  assign n18630 = ( n1281 & n18628 ) | ( n1281 & ~n18629 ) | ( n18628 & ~n18629 ) ;
  assign n18631 = ( n2156 & ~n3984 ) | ( n2156 & n14489 ) | ( ~n3984 & n14489 ) ;
  assign n18632 = ( n8885 & n10834 ) | ( n8885 & ~n18631 ) | ( n10834 & ~n18631 ) ;
  assign n18633 = n10825 ^ n6481 ^ n5421 ;
  assign n18634 = ( n9459 & ~n17511 ) | ( n9459 & n18633 ) | ( ~n17511 & n18633 ) ;
  assign n18635 = ( n5481 & n10968 ) | ( n5481 & n18634 ) | ( n10968 & n18634 ) ;
  assign n18636 = ( n1842 & n4024 ) | ( n1842 & ~n7784 ) | ( n4024 & ~n7784 ) ;
  assign n18637 = n17742 ^ n16237 ^ n9752 ;
  assign n18638 = ~n18636 & n18637 ;
  assign n18639 = ~n5556 & n18638 ;
  assign n18640 = ( n3384 & n8638 ) | ( n3384 & n13945 ) | ( n8638 & n13945 ) ;
  assign n18641 = ( ~n3615 & n4661 ) | ( ~n3615 & n14455 ) | ( n4661 & n14455 ) ;
  assign n18642 = ( n3917 & ~n9656 ) | ( n3917 & n18288 ) | ( ~n9656 & n18288 ) ;
  assign n18643 = ( ~n7111 & n18641 ) | ( ~n7111 & n18642 ) | ( n18641 & n18642 ) ;
  assign n18644 = n18643 ^ n15816 ^ n6834 ;
  assign n18645 = n5554 ^ n1634 ^ n972 ;
  assign n18646 = n18645 ^ n13918 ^ 1'b0 ;
  assign n18647 = n18646 ^ n16893 ^ n10511 ;
  assign n18648 = ( n135 & n2117 ) | ( n135 & n16113 ) | ( n2117 & n16113 ) ;
  assign n18649 = n1527 | n15600 ;
  assign n18650 = n7543 | n18649 ;
  assign n18651 = n16481 ^ n14176 ^ n10747 ;
  assign n18652 = ( n4381 & ~n4410 ) | ( n4381 & n9821 ) | ( ~n4410 & n9821 ) ;
  assign n18653 = n3008 & n3346 ;
  assign n18654 = ~n18652 & n18653 ;
  assign n18655 = ( n6322 & n10126 ) | ( n6322 & ~n18654 ) | ( n10126 & ~n18654 ) ;
  assign n18656 = n12734 ^ n4210 ^ n953 ;
  assign n18657 = n14839 & ~n18656 ;
  assign n18658 = n18657 ^ n11811 ^ n8942 ;
  assign n18659 = n7264 ^ n4129 ^ n1068 ;
  assign n18660 = n5287 | n15651 ;
  assign n18661 = ( n11380 & n18659 ) | ( n11380 & ~n18660 ) | ( n18659 & ~n18660 ) ;
  assign n18662 = ( n2105 & ~n3689 ) | ( n2105 & n11185 ) | ( ~n3689 & n11185 ) ;
  assign n18663 = n526 | n2328 ;
  assign n18664 = n4060 & ~n18663 ;
  assign n18665 = n18664 ^ n15028 ^ n11633 ;
  assign n18666 = n11037 ^ n10740 ^ 1'b0 ;
  assign n18667 = n4989 & ~n18666 ;
  assign n18668 = ( ~n6476 & n18665 ) | ( ~n6476 & n18667 ) | ( n18665 & n18667 ) ;
  assign n18669 = n14039 ^ n11994 ^ n5527 ;
  assign n18675 = n5935 ^ n183 ^ 1'b0 ;
  assign n18676 = n18675 ^ n9183 ^ n1572 ;
  assign n18677 = ( ~n208 & n4309 ) | ( ~n208 & n18676 ) | ( n4309 & n18676 ) ;
  assign n18673 = n14229 ^ n2120 ^ 1'b0 ;
  assign n18671 = ( n4354 & n4964 ) | ( n4354 & n6236 ) | ( n4964 & n6236 ) ;
  assign n18672 = n18671 ^ n10562 ^ n771 ;
  assign n18670 = n6416 ^ n6034 ^ x14 ;
  assign n18674 = n18673 ^ n18672 ^ n18670 ;
  assign n18678 = n18677 ^ n18674 ^ 1'b0 ;
  assign n18679 = n18669 & ~n18678 ;
  assign n18680 = n5970 ^ n5562 ^ n363 ;
  assign n18681 = n7386 ^ n7086 ^ n3190 ;
  assign n18682 = ( n7830 & n9789 ) | ( n7830 & n18681 ) | ( n9789 & n18681 ) ;
  assign n18683 = n18682 ^ n8672 ^ 1'b0 ;
  assign n18684 = n18680 | n18683 ;
  assign n18685 = n3168 & n3311 ;
  assign n18686 = n4940 ^ n2119 ^ n727 ;
  assign n18687 = ( ~n7767 & n18685 ) | ( ~n7767 & n18686 ) | ( n18685 & n18686 ) ;
  assign n18688 = n5004 & ~n8445 ;
  assign n18689 = n18688 ^ n8125 ^ 1'b0 ;
  assign n18690 = n18689 ^ n13560 ^ 1'b0 ;
  assign n18691 = n6073 ^ n5885 ^ 1'b0 ;
  assign n18692 = n18691 ^ n16977 ^ x124 ;
  assign n18693 = n15469 & n18652 ;
  assign n18694 = ~n3262 & n18693 ;
  assign n18695 = n18083 & ~n18694 ;
  assign n18696 = n6422 & n18695 ;
  assign n18697 = n18696 ^ n10096 ^ n6479 ;
  assign n18698 = ( n2644 & n6626 ) | ( n2644 & n6676 ) | ( n6626 & n6676 ) ;
  assign n18699 = n18698 ^ n5710 ^ 1'b0 ;
  assign n18700 = n1019 | n18031 ;
  assign n18701 = n18700 ^ n623 ^ 1'b0 ;
  assign n18704 = ~n7164 & n9413 ;
  assign n18702 = n5970 & ~n11921 ;
  assign n18703 = n1198 & n18702 ;
  assign n18705 = n18704 ^ n18703 ^ 1'b0 ;
  assign n18706 = n18701 | n18705 ;
  assign n18707 = ~n2309 & n12492 ;
  assign n18708 = ~n1122 & n18707 ;
  assign n18709 = n18708 ^ n14245 ^ n3920 ;
  assign n18710 = n12781 ^ n925 ^ 1'b0 ;
  assign n18711 = n18710 ^ n13780 ^ n1765 ;
  assign n18712 = n18711 ^ n6741 ^ n6331 ;
  assign n18713 = n18712 ^ n18001 ^ n7625 ;
  assign n18714 = ~n1588 & n15780 ;
  assign n18715 = n18714 ^ n14281 ^ 1'b0 ;
  assign n18716 = n18715 ^ n12577 ^ n2819 ;
  assign n18717 = n628 | n6336 ;
  assign n18718 = x66 | n18717 ;
  assign n18719 = n18718 ^ n14112 ^ n3695 ;
  assign n18720 = n7198 ^ n5034 ^ n3832 ;
  assign n18723 = n7417 & n8793 ;
  assign n18721 = n6829 & n11010 ;
  assign n18722 = ~n3949 & n18721 ;
  assign n18724 = n18723 ^ n18722 ^ 1'b0 ;
  assign n18725 = ~n18720 & n18724 ;
  assign n18726 = x73 & ~n18599 ;
  assign n18727 = n18726 ^ n13272 ^ 1'b0 ;
  assign n18728 = n15316 ^ n5921 ^ n5642 ;
  assign n18729 = n18728 ^ n5120 ^ 1'b0 ;
  assign n18730 = n9496 | n18729 ;
  assign n18731 = n18730 ^ n11812 ^ n4453 ;
  assign n18732 = n11718 ^ x42 ^ 1'b0 ;
  assign n18733 = n2828 & ~n18732 ;
  assign n18734 = n18733 ^ n13609 ^ 1'b0 ;
  assign n18735 = n18734 ^ n10675 ^ n5328 ;
  assign n18736 = n2444 ^ n2338 ^ x127 ;
  assign n18737 = n18736 ^ n17140 ^ 1'b0 ;
  assign n18738 = ( n3441 & n4580 ) | ( n3441 & ~n18737 ) | ( n4580 & ~n18737 ) ;
  assign n18741 = ( n877 & ~n9269 ) | ( n877 & n9964 ) | ( ~n9269 & n9964 ) ;
  assign n18739 = ( n11369 & n12859 ) | ( n11369 & ~n13299 ) | ( n12859 & ~n13299 ) ;
  assign n18740 = ( n6036 & n15458 ) | ( n6036 & ~n18739 ) | ( n15458 & ~n18739 ) ;
  assign n18742 = n18741 ^ n18740 ^ n16642 ;
  assign n18743 = n3907 ^ n3196 ^ n3085 ;
  assign n18744 = ( n2242 & n3863 ) | ( n2242 & n5204 ) | ( n3863 & n5204 ) ;
  assign n18745 = n18743 & n18744 ;
  assign n18746 = ( n3319 & n12176 ) | ( n3319 & ~n13147 ) | ( n12176 & ~n13147 ) ;
  assign n18747 = ( n14552 & n16410 ) | ( n14552 & ~n18746 ) | ( n16410 & ~n18746 ) ;
  assign n18748 = n10328 ^ n2782 ^ n1944 ;
  assign n18749 = ( ~n1129 & n7861 ) | ( ~n1129 & n18748 ) | ( n7861 & n18748 ) ;
  assign n18750 = n3513 & n11417 ;
  assign n18752 = n11225 ^ n9594 ^ n5138 ;
  assign n18751 = n12240 ^ n2274 ^ n452 ;
  assign n18753 = n18752 ^ n18751 ^ n1656 ;
  assign n18754 = ( n1158 & n3423 ) | ( n1158 & n8615 ) | ( n3423 & n8615 ) ;
  assign n18755 = n18754 ^ n8670 ^ n5474 ;
  assign n18756 = n18755 ^ n15691 ^ n14612 ;
  assign n18757 = n17496 & n18756 ;
  assign n18758 = n5543 ^ n4647 ^ 1'b0 ;
  assign n18759 = n6422 | n18758 ;
  assign n18760 = n3968 | n18759 ;
  assign n18761 = n8350 & ~n18760 ;
  assign n18762 = n1181 | n1797 ;
  assign n18763 = n2740 & ~n18762 ;
  assign n18764 = n18763 ^ n13420 ^ n1788 ;
  assign n18765 = n4399 ^ n2402 ^ 1'b0 ;
  assign n18766 = n18765 ^ n16436 ^ n6980 ;
  assign n18767 = ( n10947 & n11761 ) | ( n10947 & ~n18766 ) | ( n11761 & ~n18766 ) ;
  assign n18768 = ( n2289 & ~n5471 ) | ( n2289 & n9957 ) | ( ~n5471 & n9957 ) ;
  assign n18771 = n7156 ^ n3341 ^ n2455 ;
  assign n18772 = ( n1369 & n12277 ) | ( n1369 & ~n18771 ) | ( n12277 & ~n18771 ) ;
  assign n18770 = n528 & n8320 ;
  assign n18769 = ( n275 & n1856 ) | ( n275 & n18712 ) | ( n1856 & n18712 ) ;
  assign n18773 = n18772 ^ n18770 ^ n18769 ;
  assign n18774 = n18773 ^ n3459 ^ 1'b0 ;
  assign n18775 = n17452 & ~n18774 ;
  assign n18776 = ( n357 & n1880 ) | ( n357 & n9947 ) | ( n1880 & n9947 ) ;
  assign n18777 = n9645 ^ n3656 ^ 1'b0 ;
  assign n18778 = ~n18776 & n18777 ;
  assign n18779 = n10158 ^ n7631 ^ n2011 ;
  assign n18780 = n18779 ^ n9012 ^ n8665 ;
  assign n18781 = n6417 & n16883 ;
  assign n18782 = n18781 ^ x31 ^ 1'b0 ;
  assign n18783 = n18782 ^ n17806 ^ 1'b0 ;
  assign n18784 = n18783 ^ n8692 ^ n7742 ;
  assign n18785 = n10376 ^ n4585 ^ n2461 ;
  assign n18786 = n1898 ^ n526 ^ n401 ;
  assign n18787 = n18786 ^ n6641 ^ n735 ;
  assign n18788 = ( ~n506 & n18785 ) | ( ~n506 & n18787 ) | ( n18785 & n18787 ) ;
  assign n18790 = n13152 ^ n6731 ^ n2391 ;
  assign n18789 = ( n584 & n9308 ) | ( n584 & n12504 ) | ( n9308 & n12504 ) ;
  assign n18791 = n18790 ^ n18789 ^ n11297 ;
  assign n18792 = n18656 ^ n15408 ^ n10269 ;
  assign n18793 = n18792 ^ n13833 ^ 1'b0 ;
  assign n18795 = n9501 ^ n6637 ^ n1949 ;
  assign n18794 = n15169 | n17039 ;
  assign n18796 = n18795 ^ n18794 ^ 1'b0 ;
  assign n18797 = n3162 ^ n3096 ^ n2440 ;
  assign n18798 = n18797 ^ n9964 ^ n7045 ;
  assign n18799 = ( ~n417 & n1107 ) | ( ~n417 & n18798 ) | ( n1107 & n18798 ) ;
  assign n18805 = n12790 ^ n11396 ^ n7421 ;
  assign n18800 = n2676 ^ n1803 ^ n1129 ;
  assign n18802 = ( x5 & n8870 ) | ( x5 & ~n11883 ) | ( n8870 & ~n11883 ) ;
  assign n18801 = ( n879 & n4469 ) | ( n879 & n10621 ) | ( n4469 & n10621 ) ;
  assign n18803 = n18802 ^ n18801 ^ n13034 ;
  assign n18804 = ( n6720 & n18800 ) | ( n6720 & n18803 ) | ( n18800 & n18803 ) ;
  assign n18806 = n18805 ^ n18804 ^ 1'b0 ;
  assign n18807 = n18799 & n18806 ;
  assign n18808 = n1902 | n3368 ;
  assign n18809 = n18808 ^ n2536 ^ 1'b0 ;
  assign n18810 = ( n4459 & n9656 ) | ( n4459 & n18809 ) | ( n9656 & n18809 ) ;
  assign n18811 = n17191 ^ n12117 ^ n7083 ;
  assign n18812 = ( n3267 & ~n12472 ) | ( n3267 & n18811 ) | ( ~n12472 & n18811 ) ;
  assign n18813 = n1800 & n9691 ;
  assign n18814 = n18813 ^ n15134 ^ n13136 ;
  assign n18815 = ~n1290 & n8879 ;
  assign n18816 = n18815 ^ n7266 ^ 1'b0 ;
  assign n18817 = ( n2549 & n6095 ) | ( n2549 & ~n12299 ) | ( n6095 & ~n12299 ) ;
  assign n18818 = ( n1615 & n18816 ) | ( n1615 & ~n18817 ) | ( n18816 & ~n18817 ) ;
  assign n18819 = n18818 ^ n11764 ^ n2940 ;
  assign n18820 = ( n4788 & n17594 ) | ( n4788 & n18819 ) | ( n17594 & n18819 ) ;
  assign n18821 = n3994 ^ n3010 ^ n208 ;
  assign n18822 = ( ~n662 & n1792 ) | ( ~n662 & n9797 ) | ( n1792 & n9797 ) ;
  assign n18823 = ( n5650 & n10598 ) | ( n5650 & n18822 ) | ( n10598 & n18822 ) ;
  assign n18824 = n7083 ^ n1368 ^ 1'b0 ;
  assign n18825 = ~n18823 & n18824 ;
  assign n18826 = ~n18821 & n18825 ;
  assign n18827 = n18826 ^ n17527 ^ n8524 ;
  assign n18828 = ( ~n1903 & n6983 ) | ( ~n1903 & n9964 ) | ( n6983 & n9964 ) ;
  assign n18829 = ( n8662 & ~n14963 ) | ( n8662 & n18828 ) | ( ~n14963 & n18828 ) ;
  assign n18830 = n18829 ^ n6115 ^ 1'b0 ;
  assign n18831 = n7760 & n18830 ;
  assign n18832 = n8032 ^ n2351 ^ n366 ;
  assign n18833 = ( ~n919 & n11795 ) | ( ~n919 & n18832 ) | ( n11795 & n18832 ) ;
  assign n18834 = n18833 ^ n5892 ^ n5831 ;
  assign n18835 = ( n1169 & n13681 ) | ( n1169 & ~n18834 ) | ( n13681 & ~n18834 ) ;
  assign n18837 = n13526 ^ n4861 ^ n2174 ;
  assign n18838 = n18206 & n18837 ;
  assign n18836 = n11260 | n17423 ;
  assign n18839 = n18838 ^ n18836 ^ 1'b0 ;
  assign n18840 = n8897 & n12087 ;
  assign n18841 = ( n2596 & n18839 ) | ( n2596 & n18840 ) | ( n18839 & n18840 ) ;
  assign n18842 = n6008 | n14053 ;
  assign n18843 = n9392 | n18842 ;
  assign n18844 = n4764 ^ n287 ^ x89 ;
  assign n18845 = x49 & n18844 ;
  assign n18846 = n18845 ^ n15234 ^ 1'b0 ;
  assign n18847 = n8775 | n11391 ;
  assign n18848 = n18847 ^ n13303 ^ n388 ;
  assign n18849 = ( n2944 & ~n3436 ) | ( n2944 & n14868 ) | ( ~n3436 & n14868 ) ;
  assign n18850 = n18849 ^ n17233 ^ n12623 ;
  assign n18851 = ( n18846 & ~n18848 ) | ( n18846 & n18850 ) | ( ~n18848 & n18850 ) ;
  assign n18852 = ( ~n1008 & n18843 ) | ( ~n1008 & n18851 ) | ( n18843 & n18851 ) ;
  assign n18853 = n8709 ^ n7826 ^ n1565 ;
  assign n18854 = n18853 ^ n6654 ^ n3047 ;
  assign n18855 = n13879 ^ n7781 ^ n373 ;
  assign n18856 = ( n11155 & n18854 ) | ( n11155 & n18855 ) | ( n18854 & n18855 ) ;
  assign n18857 = n2827 & n10333 ;
  assign n18858 = n18857 ^ n6636 ^ 1'b0 ;
  assign n18859 = ~n12683 & n18414 ;
  assign n18860 = ~n2069 & n18859 ;
  assign n18861 = n1476 & ~n4342 ;
  assign n18862 = n18860 & n18861 ;
  assign n18863 = n5485 & n9127 ;
  assign n18864 = n18863 ^ n4744 ^ 1'b0 ;
  assign n18865 = n18864 ^ n18776 ^ n9429 ;
  assign n18866 = n18865 ^ n14839 ^ n4069 ;
  assign n18867 = ( n4853 & ~n10887 ) | ( n4853 & n18866 ) | ( ~n10887 & n18866 ) ;
  assign n18868 = n6696 & ~n6841 ;
  assign n18869 = n18867 & n18868 ;
  assign n18870 = n14864 ^ n9491 ^ n2102 ;
  assign n18871 = ( n2196 & n11880 ) | ( n2196 & n13798 ) | ( n11880 & n13798 ) ;
  assign n18872 = n18870 | n18871 ;
  assign n18873 = n18068 ^ n14982 ^ n4624 ;
  assign n18874 = n14716 ^ n10388 ^ n7922 ;
  assign n18875 = ( n8632 & n12101 ) | ( n8632 & ~n15840 ) | ( n12101 & ~n15840 ) ;
  assign n18876 = n18875 ^ n9611 ^ 1'b0 ;
  assign n18877 = ( n2660 & ~n6197 ) | ( n2660 & n11181 ) | ( ~n6197 & n11181 ) ;
  assign n18878 = n18877 ^ n10465 ^ 1'b0 ;
  assign n18879 = ( ~n601 & n2949 ) | ( ~n601 & n18878 ) | ( n2949 & n18878 ) ;
  assign n18880 = ( ~x33 & n4329 ) | ( ~x33 & n18879 ) | ( n4329 & n18879 ) ;
  assign n18881 = ( n6926 & ~n13283 ) | ( n6926 & n14089 ) | ( ~n13283 & n14089 ) ;
  assign n18882 = n2071 ^ n1944 ^ n776 ;
  assign n18883 = n18882 ^ n10664 ^ n4308 ;
  assign n18884 = n1494 | n2306 ;
  assign n18885 = n5220 & ~n18884 ;
  assign n18886 = n18885 ^ n5346 ^ 1'b0 ;
  assign n18890 = n14742 ^ n9183 ^ n3049 ;
  assign n18887 = n4141 ^ n3272 ^ 1'b0 ;
  assign n18888 = ~n2933 & n18887 ;
  assign n18889 = n10562 & n18888 ;
  assign n18891 = n18890 ^ n18889 ^ 1'b0 ;
  assign n18892 = x66 & n6169 ;
  assign n18893 = n18892 ^ n4106 ^ n688 ;
  assign n18894 = n6360 | n13143 ;
  assign n18895 = n18893 | n18894 ;
  assign n18896 = ~n6809 & n13915 ;
  assign n18897 = n18896 ^ n479 ^ 1'b0 ;
  assign n18898 = n18897 ^ n10059 ^ 1'b0 ;
  assign n18899 = ( n3584 & ~n6173 ) | ( n3584 & n18898 ) | ( ~n6173 & n18898 ) ;
  assign n18900 = n5802 ^ n5747 ^ n3391 ;
  assign n18903 = n7460 ^ n2312 ^ 1'b0 ;
  assign n18904 = ( n6621 & ~n7602 ) | ( n6621 & n18903 ) | ( ~n7602 & n18903 ) ;
  assign n18905 = ~n8581 & n8805 ;
  assign n18906 = n18905 ^ n5011 ^ 1'b0 ;
  assign n18907 = n18904 & n18906 ;
  assign n18901 = n12950 ^ n6863 ^ 1'b0 ;
  assign n18902 = n18606 & ~n18901 ;
  assign n18908 = n18907 ^ n18902 ^ n16804 ;
  assign n18909 = n13206 ^ n6894 ^ 1'b0 ;
  assign n18910 = n3047 & ~n4734 ;
  assign n18911 = n9610 ^ n9005 ^ n8265 ;
  assign n18912 = n18911 ^ n18485 ^ n934 ;
  assign n18913 = n13810 ^ n9178 ^ n4187 ;
  assign n18914 = n1009 & n8748 ;
  assign n18915 = n18914 ^ n16283 ^ n10181 ;
  assign n18916 = n5956 | n12937 ;
  assign n18917 = n9075 & ~n18916 ;
  assign n18918 = n16608 | n18917 ;
  assign n18919 = ( ~n2342 & n3118 ) | ( ~n2342 & n4162 ) | ( n3118 & n4162 ) ;
  assign n18920 = ( ~n3112 & n11134 ) | ( ~n3112 & n18919 ) | ( n11134 & n18919 ) ;
  assign n18922 = ( n2724 & n2845 ) | ( n2724 & ~n10892 ) | ( n2845 & ~n10892 ) ;
  assign n18921 = ( n2135 & n2285 ) | ( n2135 & ~n18786 ) | ( n2285 & ~n18786 ) ;
  assign n18923 = n18922 ^ n18921 ^ n7540 ;
  assign n18924 = n18920 | n18923 ;
  assign n18925 = n6210 & n7798 ;
  assign n18926 = n15762 ^ n8087 ^ n6995 ;
  assign n18929 = ( ~n1721 & n2496 ) | ( ~n1721 & n18864 ) | ( n2496 & n18864 ) ;
  assign n18928 = ( n543 & n6801 ) | ( n543 & ~n14034 ) | ( n6801 & ~n14034 ) ;
  assign n18930 = n18929 ^ n18928 ^ n3636 ;
  assign n18927 = n11869 ^ n11624 ^ n7140 ;
  assign n18931 = n18930 ^ n18927 ^ n159 ;
  assign n18932 = n7956 | n9400 ;
  assign n18933 = n18046 ^ n15641 ^ n7737 ;
  assign n18934 = ( ~n3816 & n5744 ) | ( ~n3816 & n12162 ) | ( n5744 & n12162 ) ;
  assign n18935 = n18934 ^ n11224 ^ 1'b0 ;
  assign n18936 = n4172 & ~n18935 ;
  assign n18937 = n18936 ^ n8336 ^ n1156 ;
  assign n18938 = ( ~n1557 & n14407 ) | ( ~n1557 & n18937 ) | ( n14407 & n18937 ) ;
  assign n18939 = n18938 ^ n10170 ^ n5734 ;
  assign n18940 = n13235 ^ n11718 ^ n9932 ;
  assign n18941 = ( n2725 & n16471 ) | ( n2725 & n18940 ) | ( n16471 & n18940 ) ;
  assign n18942 = ( n6389 & ~n8176 ) | ( n6389 & n18941 ) | ( ~n8176 & n18941 ) ;
  assign n18943 = n7933 ^ n5085 ^ n611 ;
  assign n18944 = n18943 ^ n15876 ^ x94 ;
  assign n18945 = n18944 ^ n11153 ^ n728 ;
  assign n18946 = ( ~n11359 & n18197 ) | ( ~n11359 & n18945 ) | ( n18197 & n18945 ) ;
  assign n18947 = ( n287 & ~n4921 ) | ( n287 & n13061 ) | ( ~n4921 & n13061 ) ;
  assign n18948 = ( n598 & n11519 ) | ( n598 & n13722 ) | ( n11519 & n13722 ) ;
  assign n18949 = n18948 ^ n15837 ^ 1'b0 ;
  assign n18950 = n18949 ^ n9913 ^ n8525 ;
  assign n18951 = n5364 ^ n3145 ^ 1'b0 ;
  assign n18952 = ~n18177 & n18951 ;
  assign n18953 = n9814 & n13103 ;
  assign n18954 = n18953 ^ n1623 ^ 1'b0 ;
  assign n18955 = n15441 & n16823 ;
  assign n18956 = n18955 ^ n15099 ^ 1'b0 ;
  assign n18957 = ~n16570 & n18956 ;
  assign n18958 = ( n1626 & n6637 ) | ( n1626 & ~n10035 ) | ( n6637 & ~n10035 ) ;
  assign n18959 = ( n4496 & ~n5609 ) | ( n4496 & n18958 ) | ( ~n5609 & n18958 ) ;
  assign n18960 = n6442 & ~n16620 ;
  assign n18961 = n4472 & n18960 ;
  assign n18962 = n2393 & n9478 ;
  assign n18963 = n18962 ^ n17864 ^ 1'b0 ;
  assign n18964 = ( ~n2755 & n16100 ) | ( ~n2755 & n18056 ) | ( n16100 & n18056 ) ;
  assign n18965 = n17137 ^ n5424 ^ n858 ;
  assign n18966 = n13150 ^ n6096 ^ 1'b0 ;
  assign n18967 = ( n3907 & n5868 ) | ( n3907 & ~n5954 ) | ( n5868 & ~n5954 ) ;
  assign n18968 = ( n3023 & n3927 ) | ( n3023 & n18967 ) | ( n3927 & n18967 ) ;
  assign n18969 = ( n1611 & ~n8213 ) | ( n1611 & n8784 ) | ( ~n8213 & n8784 ) ;
  assign n18970 = ( n6566 & n18968 ) | ( n6566 & n18969 ) | ( n18968 & n18969 ) ;
  assign n18971 = n18970 ^ n8333 ^ n8310 ;
  assign n18972 = ~n4553 & n17355 ;
  assign n18973 = n18972 ^ n12885 ^ 1'b0 ;
  assign n18974 = ( n1517 & n18535 ) | ( n1517 & ~n18973 ) | ( n18535 & ~n18973 ) ;
  assign n18975 = ( n842 & n2082 ) | ( n842 & n11015 ) | ( n2082 & n11015 ) ;
  assign n18979 = n17646 ^ n12440 ^ n6450 ;
  assign n18976 = ( n577 & n1773 ) | ( n577 & n2859 ) | ( n1773 & n2859 ) ;
  assign n18977 = n6700 ^ n5319 ^ n2061 ;
  assign n18978 = ( n3306 & n18976 ) | ( n3306 & ~n18977 ) | ( n18976 & ~n18977 ) ;
  assign n18980 = n18979 ^ n18978 ^ n13978 ;
  assign n18981 = n9594 & ~n18032 ;
  assign n18982 = n4648 & n18981 ;
  assign n18983 = ( n16592 & ~n16855 ) | ( n16592 & n18982 ) | ( ~n16855 & n18982 ) ;
  assign n18984 = n12809 ^ n1860 ^ 1'b0 ;
  assign n18985 = n18984 ^ n4144 ^ n4018 ;
  assign n18986 = n6622 ^ n3428 ^ 1'b0 ;
  assign n18987 = n18986 ^ n6620 ^ n731 ;
  assign n18988 = n11942 & ~n16213 ;
  assign n18989 = ~n18987 & n18988 ;
  assign n18990 = n8449 ^ n549 ^ 1'b0 ;
  assign n18991 = n2386 & ~n18990 ;
  assign n18992 = n11937 ^ n2789 ^ n2656 ;
  assign n18993 = n8071 | n18992 ;
  assign n18994 = n18993 ^ n9719 ^ 1'b0 ;
  assign n18995 = n9290 ^ n7597 ^ 1'b0 ;
  assign n18996 = n9274 | n18995 ;
  assign n18998 = ( ~n745 & n1314 ) | ( ~n745 & n11566 ) | ( n1314 & n11566 ) ;
  assign n18999 = ( ~n6024 & n11883 ) | ( ~n6024 & n18998 ) | ( n11883 & n18998 ) ;
  assign n19000 = ( n10465 & ~n12760 ) | ( n10465 & n18999 ) | ( ~n12760 & n18999 ) ;
  assign n18997 = n13725 ^ n5362 ^ 1'b0 ;
  assign n19001 = n19000 ^ n18997 ^ n6845 ;
  assign n19002 = n19001 ^ n18335 ^ n245 ;
  assign n19003 = n8858 ^ n8673 ^ n4428 ;
  assign n19004 = ( ~n8537 & n13763 ) | ( ~n8537 & n19003 ) | ( n13763 & n19003 ) ;
  assign n19005 = n3464 ^ n2511 ^ 1'b0 ;
  assign n19006 = ( n10039 & n14384 ) | ( n10039 & ~n15235 ) | ( n14384 & ~n15235 ) ;
  assign n19008 = n8288 ^ n8161 ^ n4116 ;
  assign n19007 = n10049 ^ n9639 ^ 1'b0 ;
  assign n19009 = n19008 ^ n19007 ^ n3923 ;
  assign n19010 = n10952 ^ n9324 ^ n7175 ;
  assign n19011 = ( n12914 & n12976 ) | ( n12914 & n19010 ) | ( n12976 & n19010 ) ;
  assign n19012 = n12570 ^ n6654 ^ n5720 ;
  assign n19013 = ( n6392 & ~n7906 ) | ( n6392 & n9610 ) | ( ~n7906 & n9610 ) ;
  assign n19014 = n1282 & n1508 ;
  assign n19015 = n19014 ^ n1131 ^ 1'b0 ;
  assign n19016 = n11136 ^ n6116 ^ n2639 ;
  assign n19017 = n16906 ^ n10782 ^ n4011 ;
  assign n19018 = ( n6344 & ~n18423 ) | ( n6344 & n19017 ) | ( ~n18423 & n19017 ) ;
  assign n19019 = ( ~n11396 & n19016 ) | ( ~n11396 & n19018 ) | ( n19016 & n19018 ) ;
  assign n19020 = ( n7902 & n14703 ) | ( n7902 & ~n19019 ) | ( n14703 & ~n19019 ) ;
  assign n19021 = n11476 & n19020 ;
  assign n19022 = ~n19015 & n19021 ;
  assign n19023 = ( n7235 & n19013 ) | ( n7235 & ~n19022 ) | ( n19013 & ~n19022 ) ;
  assign n19024 = n17058 ^ n14680 ^ n10331 ;
  assign n19025 = n19024 ^ n6161 ^ 1'b0 ;
  assign n19026 = n6642 | n19025 ;
  assign n19027 = n19026 ^ n13404 ^ n8522 ;
  assign n19028 = n19027 ^ n13919 ^ n1656 ;
  assign n19029 = ( n9973 & n10035 ) | ( n9973 & n10253 ) | ( n10035 & n10253 ) ;
  assign n19030 = n11276 ^ n695 ^ 1'b0 ;
  assign n19031 = ~n19029 & n19030 ;
  assign n19032 = ( n8307 & n13524 ) | ( n8307 & ~n13770 ) | ( n13524 & ~n13770 ) ;
  assign n19033 = n8441 ^ n7255 ^ n3350 ;
  assign n19034 = n1710 & n10376 ;
  assign n19035 = n19034 ^ n6517 ^ n2438 ;
  assign n19036 = n5430 & n16220 ;
  assign n19037 = n19036 ^ n2900 ^ 1'b0 ;
  assign n19038 = n4203 & n12763 ;
  assign n19039 = n19038 ^ n383 ^ 1'b0 ;
  assign n19040 = ( n1833 & ~n16367 ) | ( n1833 & n16553 ) | ( ~n16367 & n16553 ) ;
  assign n19041 = ~n7536 & n19040 ;
  assign n19042 = n7171 & ~n12742 ;
  assign n19043 = n13368 ^ n3619 ^ 1'b0 ;
  assign n19044 = n6102 ^ n3328 ^ 1'b0 ;
  assign n19045 = n19044 ^ n9827 ^ n2156 ;
  assign n19046 = ( n4341 & n8350 ) | ( n4341 & n19045 ) | ( n8350 & n19045 ) ;
  assign n19047 = n1396 & n9145 ;
  assign n19048 = ~n13140 & n19047 ;
  assign n19049 = n642 & n19048 ;
  assign n19050 = ( ~n12812 & n16767 ) | ( ~n12812 & n16787 ) | ( n16767 & n16787 ) ;
  assign n19051 = ( n202 & n3353 ) | ( n202 & ~n5838 ) | ( n3353 & ~n5838 ) ;
  assign n19052 = ( n440 & n3204 ) | ( n440 & n9368 ) | ( n3204 & n9368 ) ;
  assign n19053 = ( n12452 & n19051 ) | ( n12452 & n19052 ) | ( n19051 & n19052 ) ;
  assign n19054 = ( n2842 & n10195 ) | ( n2842 & ~n16842 ) | ( n10195 & ~n16842 ) ;
  assign n19055 = n15230 ^ n14687 ^ n1958 ;
  assign n19056 = ( n11175 & n12208 ) | ( n11175 & ~n19055 ) | ( n12208 & ~n19055 ) ;
  assign n19057 = n19056 ^ n11595 ^ n1478 ;
  assign n19058 = ~n6102 & n10987 ;
  assign n19059 = n19058 ^ n12993 ^ 1'b0 ;
  assign n19067 = ( n1314 & ~n3904 ) | ( n1314 & n18159 ) | ( ~n3904 & n18159 ) ;
  assign n19060 = n15517 ^ n13192 ^ n6153 ;
  assign n19061 = ( n7284 & n10376 ) | ( n7284 & ~n12307 ) | ( n10376 & ~n12307 ) ;
  assign n19062 = ( n3551 & n5777 ) | ( n3551 & ~n19061 ) | ( n5777 & ~n19061 ) ;
  assign n19063 = n19060 & n19062 ;
  assign n19064 = ~n1148 & n19063 ;
  assign n19065 = n9690 ^ n7407 ^ 1'b0 ;
  assign n19066 = n19064 | n19065 ;
  assign n19068 = n19067 ^ n19066 ^ 1'b0 ;
  assign n19069 = n6144 | n19068 ;
  assign n19070 = ~n14946 & n19069 ;
  assign n19071 = n4726 & n19070 ;
  assign n19072 = ( ~n379 & n3546 ) | ( ~n379 & n9048 ) | ( n3546 & n9048 ) ;
  assign n19073 = ( n13682 & ~n17739 ) | ( n13682 & n18139 ) | ( ~n17739 & n18139 ) ;
  assign n19074 = n17074 ^ n16743 ^ n1335 ;
  assign n19075 = n19074 ^ n16958 ^ n4340 ;
  assign n19076 = ( ~n12598 & n19073 ) | ( ~n12598 & n19075 ) | ( n19073 & n19075 ) ;
  assign n19077 = n7657 | n11958 ;
  assign n19078 = n19077 ^ n15272 ^ 1'b0 ;
  assign n19079 = n6255 & n19078 ;
  assign n19080 = n19079 ^ n9488 ^ n6055 ;
  assign n19081 = n13636 ^ n4224 ^ 1'b0 ;
  assign n19082 = n12872 & ~n19081 ;
  assign n19084 = n7393 ^ n1393 ^ 1'b0 ;
  assign n19083 = n17318 ^ n13144 ^ n3892 ;
  assign n19085 = n19084 ^ n19083 ^ n5043 ;
  assign n19086 = ( n3815 & n7108 ) | ( n3815 & n19085 ) | ( n7108 & n19085 ) ;
  assign n19088 = ( n1711 & n6044 ) | ( n1711 & n15188 ) | ( n6044 & n15188 ) ;
  assign n19087 = n16892 ^ n16566 ^ n14478 ;
  assign n19089 = n19088 ^ n19087 ^ n3959 ;
  assign n19090 = n11662 ^ n4651 ^ n739 ;
  assign n19091 = n10736 ^ n6146 ^ n3590 ;
  assign n19092 = ( n4175 & n12033 ) | ( n4175 & ~n19091 ) | ( n12033 & ~n19091 ) ;
  assign n19093 = ( n4283 & ~n12377 ) | ( n4283 & n19092 ) | ( ~n12377 & n19092 ) ;
  assign n19094 = ( ~n19045 & n19090 ) | ( ~n19045 & n19093 ) | ( n19090 & n19093 ) ;
  assign n19095 = ( n2294 & n2408 ) | ( n2294 & n7742 ) | ( n2408 & n7742 ) ;
  assign n19096 = ( n5959 & n7290 ) | ( n5959 & n19095 ) | ( n7290 & n19095 ) ;
  assign n19097 = n8607 ^ n4832 ^ n1115 ;
  assign n19098 = n1058 & ~n19097 ;
  assign n19099 = n1027 | n19020 ;
  assign n19100 = n19099 ^ n18696 ^ n10425 ;
  assign n19101 = n19098 & n19100 ;
  assign n19102 = ( n4667 & ~n7585 ) | ( n4667 & n17681 ) | ( ~n7585 & n17681 ) ;
  assign n19103 = n5475 | n19102 ;
  assign n19104 = n9243 ^ n4803 ^ n2673 ;
  assign n19105 = n336 & ~n19104 ;
  assign n19106 = n19105 ^ n12420 ^ 1'b0 ;
  assign n19107 = n14941 & n19106 ;
  assign n19108 = ( ~n1351 & n5747 ) | ( ~n1351 & n7180 ) | ( n5747 & n7180 ) ;
  assign n19109 = n8653 & ~n10788 ;
  assign n19110 = n19108 & n19109 ;
  assign n19111 = ( ~n11107 & n11462 ) | ( ~n11107 & n17102 ) | ( n11462 & n17102 ) ;
  assign n19112 = n4991 ^ n3652 ^ n3174 ;
  assign n19113 = n19112 ^ n6736 ^ n6330 ;
  assign n19114 = ( n6029 & n9579 ) | ( n6029 & n17574 ) | ( n9579 & n17574 ) ;
  assign n19115 = ~n4083 & n4433 ;
  assign n19116 = n10534 | n12217 ;
  assign n19117 = n19116 ^ n16291 ^ 1'b0 ;
  assign n19118 = n4128 & ~n12139 ;
  assign n19119 = n19118 ^ n11013 ^ 1'b0 ;
  assign n19121 = n9739 ^ n3765 ^ 1'b0 ;
  assign n19122 = n19121 ^ n15995 ^ n14107 ;
  assign n19123 = ( n1373 & n9690 ) | ( n1373 & ~n19122 ) | ( n9690 & ~n19122 ) ;
  assign n19120 = n7140 ^ n2420 ^ n1153 ;
  assign n19124 = n19123 ^ n19120 ^ n11750 ;
  assign n19126 = ~n733 & n3119 ;
  assign n19125 = n460 & ~n2140 ;
  assign n19127 = n19126 ^ n19125 ^ n10166 ;
  assign n19128 = ( n10043 & n17236 ) | ( n10043 & ~n19127 ) | ( n17236 & ~n19127 ) ;
  assign n19129 = n19128 ^ n8317 ^ n4080 ;
  assign n19130 = n11620 ^ n3238 ^ 1'b0 ;
  assign n19131 = ( n13696 & n13991 ) | ( n13696 & n16606 ) | ( n13991 & n16606 ) ;
  assign n19132 = n17820 ^ n13519 ^ 1'b0 ;
  assign n19134 = ( n1628 & n9271 ) | ( n1628 & n11087 ) | ( n9271 & n11087 ) ;
  assign n19133 = n2926 & n7168 ;
  assign n19135 = n19134 ^ n19133 ^ n3968 ;
  assign n19136 = ( ~n758 & n14011 ) | ( ~n758 & n15651 ) | ( n14011 & n15651 ) ;
  assign n19137 = n19136 ^ n14886 ^ n6636 ;
  assign n19138 = ( ~n251 & n3899 ) | ( ~n251 & n10166 ) | ( n3899 & n10166 ) ;
  assign n19139 = n19138 ^ n15121 ^ n13997 ;
  assign n19140 = x122 & ~n7007 ;
  assign n19141 = ~n2106 & n19140 ;
  assign n19142 = ( n916 & ~n7451 ) | ( n916 & n19141 ) | ( ~n7451 & n19141 ) ;
  assign n19143 = n5636 & ~n19142 ;
  assign n19144 = n4659 & n19143 ;
  assign n19145 = ( n232 & ~n2664 ) | ( n232 & n6657 ) | ( ~n2664 & n6657 ) ;
  assign n19146 = ( n1084 & n11116 ) | ( n1084 & n19145 ) | ( n11116 & n19145 ) ;
  assign n19147 = n19146 ^ n3051 ^ 1'b0 ;
  assign n19148 = n18722 | n19147 ;
  assign n19149 = n10351 & ~n11416 ;
  assign n19150 = ~n293 & n19149 ;
  assign n19151 = ( ~n10799 & n18677 ) | ( ~n10799 & n19150 ) | ( n18677 & n19150 ) ;
  assign n19152 = n7736 ^ n4426 ^ 1'b0 ;
  assign n19153 = ( ~n2549 & n6197 ) | ( ~n2549 & n19152 ) | ( n6197 & n19152 ) ;
  assign n19154 = ( n2800 & ~n6216 ) | ( n2800 & n6239 ) | ( ~n6216 & n6239 ) ;
  assign n19155 = ( n770 & n4874 ) | ( n770 & n19154 ) | ( n4874 & n19154 ) ;
  assign n19156 = ( n8406 & n12922 ) | ( n8406 & ~n19155 ) | ( n12922 & ~n19155 ) ;
  assign n19168 = n10105 ^ n9009 ^ n233 ;
  assign n19167 = ( ~n6088 & n11087 ) | ( ~n6088 & n12966 ) | ( n11087 & n12966 ) ;
  assign n19158 = ( ~n1861 & n3552 ) | ( ~n1861 & n5241 ) | ( n3552 & n5241 ) ;
  assign n19159 = n6771 ^ n3916 ^ 1'b0 ;
  assign n19160 = n19158 & n19159 ;
  assign n19161 = ( n1694 & ~n6896 ) | ( n1694 & n19160 ) | ( ~n6896 & n19160 ) ;
  assign n19162 = ( n4121 & ~n10270 ) | ( n4121 & n19161 ) | ( ~n10270 & n19161 ) ;
  assign n19163 = n3937 | n4561 ;
  assign n19164 = n19162 | n19163 ;
  assign n19165 = n19164 ^ n6489 ^ 1'b0 ;
  assign n19157 = n17052 ^ n5257 ^ n4093 ;
  assign n19166 = n19165 ^ n19157 ^ n17031 ;
  assign n19169 = n19168 ^ n19167 ^ n19166 ;
  assign n19170 = n10483 ^ n1582 ^ 1'b0 ;
  assign n19171 = n6875 & n19170 ;
  assign n19172 = n19171 ^ n13817 ^ 1'b0 ;
  assign n19173 = n4742 & ~n19172 ;
  assign n19174 = ( n4451 & n9084 ) | ( n4451 & ~n19173 ) | ( n9084 & ~n19173 ) ;
  assign n19175 = n5055 | n12420 ;
  assign n19176 = n14145 & ~n19175 ;
  assign n19177 = n14868 ^ n4583 ^ n1484 ;
  assign n19178 = ( n430 & ~n1153 ) | ( n430 & n19177 ) | ( ~n1153 & n19177 ) ;
  assign n19179 = n19178 ^ n17505 ^ n6449 ;
  assign n19180 = n7673 ^ n3725 ^ 1'b0 ;
  assign n19181 = n9565 | n19180 ;
  assign n19182 = n1933 ^ n1277 ^ 1'b0 ;
  assign n19183 = n12218 & n19182 ;
  assign n19184 = ( ~n7383 & n10207 ) | ( ~n7383 & n19183 ) | ( n10207 & n19183 ) ;
  assign n19185 = n19181 & ~n19184 ;
  assign n19186 = ( ~n1504 & n11018 ) | ( ~n1504 & n18403 ) | ( n11018 & n18403 ) ;
  assign n19187 = n9787 ^ n4333 ^ n232 ;
  assign n19188 = ( n6409 & n19186 ) | ( n6409 & ~n19187 ) | ( n19186 & ~n19187 ) ;
  assign n19189 = ( ~n6084 & n12230 ) | ( ~n6084 & n13557 ) | ( n12230 & n13557 ) ;
  assign n19190 = n19189 ^ n13886 ^ n12786 ;
  assign n19191 = n19190 ^ n18779 ^ n9434 ;
  assign n19192 = n14711 ^ n9620 ^ 1'b0 ;
  assign n19193 = n13090 ^ n6712 ^ n6470 ;
  assign n19194 = n17781 ^ n8491 ^ 1'b0 ;
  assign n19195 = ~n13609 & n19194 ;
  assign n19196 = ( n6628 & n19193 ) | ( n6628 & ~n19195 ) | ( n19193 & ~n19195 ) ;
  assign n19197 = ( ~n6210 & n8195 ) | ( ~n6210 & n9351 ) | ( n8195 & n9351 ) ;
  assign n19201 = n4330 & ~n9660 ;
  assign n19202 = n19201 ^ n13469 ^ n4838 ;
  assign n19198 = n8721 | n9816 ;
  assign n19199 = n4291 & ~n19198 ;
  assign n19200 = ( x122 & n6698 ) | ( x122 & n19199 ) | ( n6698 & n19199 ) ;
  assign n19203 = n19202 ^ n19200 ^ n1638 ;
  assign n19204 = ( ~n1745 & n7310 ) | ( ~n1745 & n15331 ) | ( n7310 & n15331 ) ;
  assign n19205 = n3498 ^ n3230 ^ 1'b0 ;
  assign n19206 = n17262 | n19205 ;
  assign n19207 = ~n5686 & n12268 ;
  assign n19208 = n19207 ^ n18938 ^ 1'b0 ;
  assign n19209 = n19208 ^ n17812 ^ n9195 ;
  assign n19210 = ( n19204 & ~n19206 ) | ( n19204 & n19209 ) | ( ~n19206 & n19209 ) ;
  assign n19216 = ( ~n4586 & n12784 ) | ( ~n4586 & n13209 ) | ( n12784 & n13209 ) ;
  assign n19217 = n19216 ^ n7515 ^ n520 ;
  assign n19218 = n19217 ^ n7907 ^ n1609 ;
  assign n19211 = n6091 ^ n4286 ^ 1'b0 ;
  assign n19212 = n18718 ^ n266 ^ 1'b0 ;
  assign n19213 = n19211 & ~n19212 ;
  assign n19214 = n19213 ^ n1139 ^ 1'b0 ;
  assign n19215 = n15826 & n19214 ;
  assign n19219 = n19218 ^ n19215 ^ n1385 ;
  assign n19220 = n10675 & ~n14137 ;
  assign n19221 = n19220 ^ n10970 ^ 1'b0 ;
  assign n19222 = n19221 ^ n9754 ^ n1467 ;
  assign n19223 = n9682 ^ n2938 ^ 1'b0 ;
  assign n19224 = ~n17162 & n19223 ;
  assign n19225 = ( ~n1759 & n10840 ) | ( ~n1759 & n12469 ) | ( n10840 & n12469 ) ;
  assign n19226 = n9662 ^ n1172 ^ n736 ;
  assign n19227 = ~n6336 & n19226 ;
  assign n19228 = ~n15769 & n19227 ;
  assign n19229 = ( ~n9620 & n19225 ) | ( ~n9620 & n19228 ) | ( n19225 & n19228 ) ;
  assign n19230 = ( n6733 & ~n10998 ) | ( n6733 & n15638 ) | ( ~n10998 & n15638 ) ;
  assign n19231 = n3479 | n19230 ;
  assign n19232 = n19231 ^ n11545 ^ 1'b0 ;
  assign n19233 = ( n4671 & n15036 ) | ( n4671 & n19232 ) | ( n15036 & n19232 ) ;
  assign n19234 = n13448 ^ n11487 ^ n3220 ;
  assign n19235 = n19234 ^ n1146 ^ n720 ;
  assign n19236 = ( x21 & ~n5421 ) | ( x21 & n18494 ) | ( ~n5421 & n18494 ) ;
  assign n19237 = n9871 ^ n6212 ^ n559 ;
  assign n19238 = ( n6090 & ~n14987 ) | ( n6090 & n19237 ) | ( ~n14987 & n19237 ) ;
  assign n19239 = n19238 ^ n14434 ^ n10552 ;
  assign n19240 = n19236 & ~n19239 ;
  assign n19241 = n8482 & n19240 ;
  assign n19242 = ( n1987 & n4133 ) | ( n1987 & n19241 ) | ( n4133 & n19241 ) ;
  assign n19243 = n12797 ^ n6526 ^ n4560 ;
  assign n19244 = ~n12504 & n19243 ;
  assign n19245 = n19244 ^ n175 ^ 1'b0 ;
  assign n19246 = ( ~n192 & n5477 ) | ( ~n192 & n19245 ) | ( n5477 & n19245 ) ;
  assign n19247 = n13223 ^ n9581 ^ n8184 ;
  assign n19248 = n10362 | n19247 ;
  assign n19253 = ~n9336 & n11345 ;
  assign n19254 = n19253 ^ n17764 ^ n4948 ;
  assign n19249 = ( n1805 & n3042 ) | ( n1805 & ~n3899 ) | ( n3042 & ~n3899 ) ;
  assign n19250 = n19249 ^ n2661 ^ 1'b0 ;
  assign n19251 = n5546 ^ n4166 ^ 1'b0 ;
  assign n19252 = ~n19250 & n19251 ;
  assign n19255 = n19254 ^ n19252 ^ 1'b0 ;
  assign n19256 = n15000 & n19255 ;
  assign n19257 = ( n3174 & ~n19248 ) | ( n3174 & n19256 ) | ( ~n19248 & n19256 ) ;
  assign n19258 = n18397 ^ n14864 ^ n5042 ;
  assign n19259 = ( n3218 & n7503 ) | ( n3218 & ~n19258 ) | ( n7503 & ~n19258 ) ;
  assign n19260 = ( ~n6782 & n15697 ) | ( ~n6782 & n19259 ) | ( n15697 & n19259 ) ;
  assign n19261 = ( ~n3178 & n4412 ) | ( ~n3178 & n15651 ) | ( n4412 & n15651 ) ;
  assign n19262 = ( n4271 & ~n5399 ) | ( n4271 & n13836 ) | ( ~n5399 & n13836 ) ;
  assign n19265 = n7310 ^ n2515 ^ n158 ;
  assign n19263 = n3244 & n3908 ;
  assign n19264 = ( ~n2120 & n9260 ) | ( ~n2120 & n19263 ) | ( n9260 & n19263 ) ;
  assign n19266 = n19265 ^ n19264 ^ n14002 ;
  assign n19267 = ( n1034 & ~n6759 ) | ( n1034 & n19266 ) | ( ~n6759 & n19266 ) ;
  assign n19268 = ( n778 & ~n16266 ) | ( n778 & n19267 ) | ( ~n16266 & n19267 ) ;
  assign n19269 = n1830 | n4955 ;
  assign n19270 = ( n584 & n1804 ) | ( n584 & ~n11194 ) | ( n1804 & ~n11194 ) ;
  assign n19271 = n5787 | n16235 ;
  assign n19272 = n19270 | n19271 ;
  assign n19273 = n15067 ^ n9120 ^ n6870 ;
  assign n19274 = ( n3046 & n6124 ) | ( n3046 & n19273 ) | ( n6124 & n19273 ) ;
  assign n19278 = n8549 ^ n4812 ^ 1'b0 ;
  assign n19279 = n2208 | n19278 ;
  assign n19276 = ( n3403 & ~n4042 ) | ( n3403 & n7699 ) | ( ~n4042 & n7699 ) ;
  assign n19275 = n18821 ^ n14277 ^ n3669 ;
  assign n19277 = n19276 ^ n19275 ^ n16042 ;
  assign n19280 = n19279 ^ n19277 ^ n9942 ;
  assign n19284 = ( n1087 & n6930 ) | ( n1087 & ~n8292 ) | ( n6930 & ~n8292 ) ;
  assign n19285 = n5800 ^ n339 ^ 1'b0 ;
  assign n19286 = ~n19284 & n19285 ;
  assign n19287 = ( n3597 & ~n6646 ) | ( n3597 & n19286 ) | ( ~n6646 & n19286 ) ;
  assign n19282 = ( n558 & ~n4271 ) | ( n558 & n9587 ) | ( ~n4271 & n9587 ) ;
  assign n19283 = ( n2593 & n6985 ) | ( n2593 & ~n19282 ) | ( n6985 & ~n19282 ) ;
  assign n19281 = n19062 ^ n13015 ^ n11750 ;
  assign n19288 = n19287 ^ n19283 ^ n19281 ;
  assign n19290 = ( n11240 & ~n11845 ) | ( n11240 & n12000 ) | ( ~n11845 & n12000 ) ;
  assign n19289 = n6022 & n13057 ;
  assign n19291 = n19290 ^ n19289 ^ 1'b0 ;
  assign n19292 = n4111 & n14931 ;
  assign n19293 = n19292 ^ x70 ^ 1'b0 ;
  assign n19294 = ( n3984 & n7370 ) | ( n3984 & ~n19293 ) | ( n7370 & ~n19293 ) ;
  assign n19295 = ( ~n1712 & n4651 ) | ( ~n1712 & n8628 ) | ( n4651 & n8628 ) ;
  assign n19296 = n19294 & n19295 ;
  assign n19297 = ~n8087 & n19296 ;
  assign n19298 = n2973 ^ n2795 ^ n2360 ;
  assign n19299 = n19298 ^ n15922 ^ n11707 ;
  assign n19300 = n7253 ^ n3000 ^ n654 ;
  assign n19301 = ( n4662 & n7991 ) | ( n4662 & ~n19300 ) | ( n7991 & ~n19300 ) ;
  assign n19302 = n13800 ^ n10875 ^ n10687 ;
  assign n19303 = n15247 & ~n19302 ;
  assign n19304 = ~n3502 & n11737 ;
  assign n19305 = ~n4691 & n19304 ;
  assign n19306 = n12803 ^ n12018 ^ n7300 ;
  assign n19307 = ( n10008 & n13729 ) | ( n10008 & ~n15802 ) | ( n13729 & ~n15802 ) ;
  assign n19308 = n19307 ^ n12003 ^ n9948 ;
  assign n19309 = ( n345 & ~n10901 ) | ( n345 & n12874 ) | ( ~n10901 & n12874 ) ;
  assign n19310 = ( n801 & n1316 ) | ( n801 & n2492 ) | ( n1316 & n2492 ) ;
  assign n19311 = n19310 ^ n12178 ^ n7503 ;
  assign n19312 = ( ~n4765 & n12602 ) | ( ~n4765 & n18050 ) | ( n12602 & n18050 ) ;
  assign n19313 = ( ~n3316 & n19311 ) | ( ~n3316 & n19312 ) | ( n19311 & n19312 ) ;
  assign n19314 = n6511 ^ n4519 ^ 1'b0 ;
  assign n19315 = n19314 ^ n14407 ^ n6389 ;
  assign n19319 = n5763 & n8545 ;
  assign n19317 = n18490 ^ n6960 ^ n509 ;
  assign n19316 = n17209 ^ n6426 ^ n5808 ;
  assign n19318 = n19317 ^ n19316 ^ n3865 ;
  assign n19320 = n19319 ^ n19318 ^ n4798 ;
  assign n19321 = ( n375 & n7991 ) | ( n375 & n9919 ) | ( n7991 & n9919 ) ;
  assign n19322 = n15099 ^ n9285 ^ n8382 ;
  assign n19323 = n12496 ^ n5252 ^ 1'b0 ;
  assign n19324 = ( n9469 & n10308 ) | ( n9469 & n19323 ) | ( n10308 & n19323 ) ;
  assign n19325 = ( n18393 & n19322 ) | ( n18393 & n19324 ) | ( n19322 & n19324 ) ;
  assign n19326 = n19321 & ~n19325 ;
  assign n19327 = n19326 ^ n15369 ^ 1'b0 ;
  assign n19328 = ( n6729 & ~n8737 ) | ( n6729 & n18244 ) | ( ~n8737 & n18244 ) ;
  assign n19331 = n5485 ^ n3240 ^ n621 ;
  assign n19332 = n19331 ^ n18844 ^ n4857 ;
  assign n19333 = n19332 ^ n4999 ^ n2314 ;
  assign n19329 = n10321 ^ n1847 ^ 1'b0 ;
  assign n19330 = n14904 & ~n19329 ;
  assign n19334 = n19333 ^ n19330 ^ n9585 ;
  assign n19335 = n8737 ^ n7009 ^ n4283 ;
  assign n19340 = x82 & ~n7226 ;
  assign n19341 = n19340 ^ n4723 ^ 1'b0 ;
  assign n19342 = n19341 ^ n4476 ^ n969 ;
  assign n19337 = n3232 & ~n16715 ;
  assign n19338 = n19337 ^ n15029 ^ 1'b0 ;
  assign n19339 = n19338 ^ n4121 ^ n1084 ;
  assign n19336 = ( n7468 & n10771 ) | ( n7468 & ~n15974 ) | ( n10771 & ~n15974 ) ;
  assign n19343 = n19342 ^ n19339 ^ n19336 ;
  assign n19344 = n16586 ^ n16543 ^ 1'b0 ;
  assign n19345 = n8896 & n19344 ;
  assign n19346 = n616 & ~n17920 ;
  assign n19347 = n19346 ^ n6524 ^ 1'b0 ;
  assign n19348 = n278 & ~n3711 ;
  assign n19349 = ( ~n1054 & n19347 ) | ( ~n1054 & n19348 ) | ( n19347 & n19348 ) ;
  assign n19350 = n15289 ^ n9735 ^ x44 ;
  assign n19351 = ( n7469 & ~n9732 ) | ( n7469 & n18652 ) | ( ~n9732 & n18652 ) ;
  assign n19352 = n13544 ^ n9139 ^ n3964 ;
  assign n19353 = n19352 ^ n10891 ^ n6813 ;
  assign n19355 = n8002 ^ n7436 ^ n2909 ;
  assign n19354 = ~n8102 & n11276 ;
  assign n19356 = n19355 ^ n19354 ^ 1'b0 ;
  assign n19357 = n19353 | n19356 ;
  assign n19358 = n8559 & ~n19357 ;
  assign n19359 = n4688 & n11925 ;
  assign n19360 = n19359 ^ n9285 ^ n5017 ;
  assign n19361 = n10814 ^ n9023 ^ 1'b0 ;
  assign n19362 = n19361 ^ n13275 ^ n10819 ;
  assign n19365 = ~n2735 & n3818 ;
  assign n19366 = ( n834 & n7605 ) | ( n834 & n19365 ) | ( n7605 & n19365 ) ;
  assign n19367 = ( n3754 & n9191 ) | ( n3754 & n19366 ) | ( n9191 & n19366 ) ;
  assign n19363 = ( n929 & ~n1658 ) | ( n929 & n5983 ) | ( ~n1658 & n5983 ) ;
  assign n19364 = ( n2513 & n11244 ) | ( n2513 & n19363 ) | ( n11244 & n19363 ) ;
  assign n19368 = n19367 ^ n19364 ^ n5293 ;
  assign n19369 = n8182 ^ n7031 ^ n3522 ;
  assign n19370 = n9737 ^ n2847 ^ 1'b0 ;
  assign n19371 = ~n19369 & n19370 ;
  assign n19372 = ~n4439 & n19371 ;
  assign n19373 = ( n3851 & n8123 ) | ( n3851 & n8413 ) | ( n8123 & n8413 ) ;
  assign n19375 = n11538 ^ n5215 ^ n1079 ;
  assign n19376 = n19375 ^ n14665 ^ n4016 ;
  assign n19374 = ( n1612 & n4810 ) | ( n1612 & ~n18217 ) | ( n4810 & ~n18217 ) ;
  assign n19377 = n19376 ^ n19374 ^ n7036 ;
  assign n19378 = n15803 | n19377 ;
  assign n19379 = ~n2485 & n9957 ;
  assign n19380 = n19379 ^ n18370 ^ n12615 ;
  assign n19381 = n19380 ^ n10229 ^ n9304 ;
  assign n19382 = ~n499 & n4538 ;
  assign n19383 = n19382 ^ n2252 ^ 1'b0 ;
  assign n19384 = n10839 & n19383 ;
  assign n19386 = n8705 ^ n7160 ^ 1'b0 ;
  assign n19387 = n1660 | n19386 ;
  assign n19385 = n3546 & ~n6360 ;
  assign n19388 = n19387 ^ n19385 ^ n11162 ;
  assign n19389 = ~n9518 & n15174 ;
  assign n19390 = n19389 ^ n4693 ^ 1'b0 ;
  assign n19391 = n11935 ^ n2555 ^ n2257 ;
  assign n19392 = ( n742 & n2960 ) | ( n742 & ~n9581 ) | ( n2960 & ~n9581 ) ;
  assign n19393 = n19391 & n19392 ;
  assign n19394 = n19390 & n19393 ;
  assign n19395 = n19394 ^ n8321 ^ x37 ;
  assign n19396 = n17885 ^ n15891 ^ n1397 ;
  assign n19397 = ( ~n3116 & n18669 ) | ( ~n3116 & n18821 ) | ( n18669 & n18821 ) ;
  assign n19398 = ( n5520 & n12354 ) | ( n5520 & n19397 ) | ( n12354 & n19397 ) ;
  assign n19399 = n17982 ^ n3766 ^ 1'b0 ;
  assign n19403 = n14211 ^ n12751 ^ n12239 ;
  assign n19400 = n9834 | n11480 ;
  assign n19401 = n16758 | n19400 ;
  assign n19402 = n19401 ^ n8594 ^ 1'b0 ;
  assign n19404 = n19403 ^ n19402 ^ n13857 ;
  assign n19405 = n11484 ^ n5231 ^ n1717 ;
  assign n19406 = n19405 ^ n1917 ^ 1'b0 ;
  assign n19407 = n19406 ^ n7668 ^ n2623 ;
  assign n19408 = n19407 ^ n11994 ^ 1'b0 ;
  assign n19409 = n19408 ^ n13736 ^ n1574 ;
  assign n19411 = n11048 ^ n11005 ^ n1220 ;
  assign n19412 = n18198 & ~n19411 ;
  assign n19410 = n6881 ^ n3972 ^ n1402 ;
  assign n19413 = n19412 ^ n19410 ^ 1'b0 ;
  assign n19414 = ~n3719 & n19413 ;
  assign n19415 = n5244 & ~n8316 ;
  assign n19416 = n9284 | n11980 ;
  assign n19417 = n3384 | n19416 ;
  assign n19418 = n19417 ^ n10318 ^ n6874 ;
  assign n19419 = n19418 ^ n17328 ^ n10014 ;
  assign n19420 = n17427 ^ n10633 ^ n3644 ;
  assign n19421 = ~n398 & n4532 ;
  assign n19422 = n19421 ^ n17442 ^ 1'b0 ;
  assign n19423 = ~n2704 & n5042 ;
  assign n19424 = ~n3513 & n19423 ;
  assign n19425 = ( n3429 & n7821 ) | ( n3429 & n19424 ) | ( n7821 & n19424 ) ;
  assign n19426 = ( n564 & n4144 ) | ( n564 & n19425 ) | ( n4144 & n19425 ) ;
  assign n19427 = n19426 ^ n11137 ^ n7537 ;
  assign n19428 = n19427 ^ n7406 ^ 1'b0 ;
  assign n19430 = n9763 ^ n3361 ^ n2789 ;
  assign n19429 = ~n4374 & n15826 ;
  assign n19431 = n19430 ^ n19429 ^ 1'b0 ;
  assign n19434 = n4147 & ~n12138 ;
  assign n19432 = n16466 ^ n9384 ^ n2493 ;
  assign n19433 = ( ~n16340 & n16686 ) | ( ~n16340 & n19432 ) | ( n16686 & n19432 ) ;
  assign n19435 = n19434 ^ n19433 ^ 1'b0 ;
  assign n19436 = x82 & n19435 ;
  assign n19437 = n7091 ^ n6050 ^ n4069 ;
  assign n19438 = ( ~n5966 & n17652 ) | ( ~n5966 & n19437 ) | ( n17652 & n19437 ) ;
  assign n19440 = ( n1576 & n1685 ) | ( n1576 & ~n13144 ) | ( n1685 & ~n13144 ) ;
  assign n19439 = ~n9837 & n13553 ;
  assign n19441 = n19440 ^ n19439 ^ n12231 ;
  assign n19442 = n7546 | n16133 ;
  assign n19443 = n13271 ^ n6717 ^ 1'b0 ;
  assign n19444 = ( n12502 & ~n15735 ) | ( n12502 & n19443 ) | ( ~n15735 & n19443 ) ;
  assign n19445 = ( n10564 & n19442 ) | ( n10564 & n19444 ) | ( n19442 & n19444 ) ;
  assign n19446 = ( ~n6255 & n12240 ) | ( ~n6255 & n12664 ) | ( n12240 & n12664 ) ;
  assign n19447 = n13966 ^ n12296 ^ n6281 ;
  assign n19451 = n6656 | n7057 ;
  assign n19452 = n19451 ^ n1802 ^ 1'b0 ;
  assign n19448 = ( ~n1564 & n1862 ) | ( ~n1564 & n5716 ) | ( n1862 & n5716 ) ;
  assign n19449 = n19448 ^ n16644 ^ n5600 ;
  assign n19450 = ~n3246 & n19449 ;
  assign n19453 = n19452 ^ n19450 ^ 1'b0 ;
  assign n19454 = n2314 & ~n19453 ;
  assign n19460 = n644 & n11422 ;
  assign n19461 = ~n5098 & n19460 ;
  assign n19456 = n6401 ^ n2504 ^ 1'b0 ;
  assign n19457 = n19456 ^ n18732 ^ n10792 ;
  assign n19455 = n1392 ^ n186 ^ 1'b0 ;
  assign n19458 = n19457 ^ n19455 ^ n12615 ;
  assign n19459 = ( n184 & n8719 ) | ( n184 & n19458 ) | ( n8719 & n19458 ) ;
  assign n19462 = n19461 ^ n19459 ^ n10256 ;
  assign n19466 = n7479 ^ n599 ^ 1'b0 ;
  assign n19463 = n7867 ^ n3220 ^ n1441 ;
  assign n19464 = ( n10863 & n13847 ) | ( n10863 & ~n19463 ) | ( n13847 & ~n19463 ) ;
  assign n19465 = n9380 & ~n19464 ;
  assign n19467 = n19466 ^ n19465 ^ n1131 ;
  assign n19468 = n11081 ^ n6766 ^ 1'b0 ;
  assign n19469 = n19468 ^ n18353 ^ n14493 ;
  assign n19471 = n8071 ^ n5424 ^ n2069 ;
  assign n19470 = n18977 ^ n6720 ^ n5381 ;
  assign n19472 = n19471 ^ n19470 ^ n6143 ;
  assign n19473 = ( n2612 & ~n16436 ) | ( n2612 & n18708 ) | ( ~n16436 & n18708 ) ;
  assign n19474 = n6708 ^ n912 ^ 1'b0 ;
  assign n19475 = n12079 | n19474 ;
  assign n19476 = n6967 & n18190 ;
  assign n19477 = n19476 ^ n14686 ^ n9663 ;
  assign n19478 = n4748 & n19477 ;
  assign n19479 = n19478 ^ n2450 ^ 1'b0 ;
  assign n19480 = ( ~n3552 & n6345 ) | ( ~n3552 & n18771 ) | ( n6345 & n18771 ) ;
  assign n19481 = n3846 & n5033 ;
  assign n19482 = n19481 ^ n5446 ^ n4920 ;
  assign n19483 = n19482 ^ n10562 ^ n6749 ;
  assign n19487 = n9550 | n10622 ;
  assign n19484 = n2313 | n15225 ;
  assign n19485 = n19484 ^ n325 ^ 1'b0 ;
  assign n19486 = n8988 | n19485 ;
  assign n19488 = n19487 ^ n19486 ^ n15447 ;
  assign n19489 = n11646 ^ n10962 ^ n1668 ;
  assign n19490 = n14608 ^ n5735 ^ n765 ;
  assign n19491 = n15015 & n19490 ;
  assign n19492 = ~n11872 & n19491 ;
  assign n19493 = ( n2776 & ~n12205 ) | ( n2776 & n19492 ) | ( ~n12205 & n19492 ) ;
  assign n19494 = n7757 ^ n5405 ^ n1312 ;
  assign n19495 = ( n422 & n5455 ) | ( n422 & ~n15019 ) | ( n5455 & ~n15019 ) ;
  assign n19496 = n19495 ^ n1042 ^ 1'b0 ;
  assign n19497 = n19494 & ~n19496 ;
  assign n19498 = n19493 & ~n19497 ;
  assign n19499 = n11194 ^ n1453 ^ 1'b0 ;
  assign n19500 = n19499 ^ n18037 ^ 1'b0 ;
  assign n19501 = n1176 & ~n19434 ;
  assign n19502 = n19501 ^ n4122 ^ 1'b0 ;
  assign n19503 = ( ~n1918 & n5500 ) | ( ~n1918 & n18597 ) | ( n5500 & n18597 ) ;
  assign n19504 = ( n4488 & n7195 ) | ( n4488 & ~n9579 ) | ( n7195 & ~n9579 ) ;
  assign n19505 = ( ~n2254 & n13189 ) | ( ~n2254 & n19504 ) | ( n13189 & n19504 ) ;
  assign n19506 = ( ~n4506 & n19003 ) | ( ~n4506 & n19505 ) | ( n19003 & n19505 ) ;
  assign n19507 = ~n245 & n5486 ;
  assign n19508 = ~n5894 & n19507 ;
  assign n19509 = ( n5828 & ~n6162 ) | ( n5828 & n19508 ) | ( ~n6162 & n19508 ) ;
  assign n19510 = n9638 ^ n9308 ^ n3020 ;
  assign n19511 = n19510 ^ n13389 ^ n4514 ;
  assign n19512 = n15157 ^ n3541 ^ 1'b0 ;
  assign n19513 = n11810 ^ n10467 ^ 1'b0 ;
  assign n19514 = n19512 & ~n19513 ;
  assign n19515 = n10772 & ~n18376 ;
  assign n19516 = n19515 ^ n6820 ^ n4877 ;
  assign n19517 = n11342 ^ n5014 ^ n1007 ;
  assign n19518 = n5726 ^ n5381 ^ n2697 ;
  assign n19519 = n19518 ^ n9530 ^ n5574 ;
  assign n19520 = ( ~n1483 & n19517 ) | ( ~n1483 & n19519 ) | ( n19517 & n19519 ) ;
  assign n19521 = n2882 & n6671 ;
  assign n19522 = n19521 ^ n16998 ^ n5264 ;
  assign n19523 = ( n2487 & n11479 ) | ( n2487 & n19522 ) | ( n11479 & n19522 ) ;
  assign n19527 = n19145 ^ n17435 ^ n1065 ;
  assign n19524 = ~n2527 & n2903 ;
  assign n19525 = n4856 ^ n1929 ^ n252 ;
  assign n19526 = ( n15678 & ~n19524 ) | ( n15678 & n19525 ) | ( ~n19524 & n19525 ) ;
  assign n19528 = n19527 ^ n19526 ^ n3881 ;
  assign n19529 = n12666 ^ n9530 ^ n6134 ;
  assign n19532 = n16634 ^ n7417 ^ 1'b0 ;
  assign n19530 = ( n8142 & ~n10849 ) | ( n8142 & n14554 ) | ( ~n10849 & n14554 ) ;
  assign n19531 = n19530 ^ n5696 ^ 1'b0 ;
  assign n19533 = n19532 ^ n19531 ^ n13920 ;
  assign n19534 = n4985 ^ n3619 ^ n2964 ;
  assign n19535 = n469 | n18424 ;
  assign n19536 = n6749 & ~n19535 ;
  assign n19537 = n15009 ^ n14994 ^ 1'b0 ;
  assign n19538 = ~n8138 & n19537 ;
  assign n19539 = n12936 ^ n11604 ^ n4268 ;
  assign n19540 = n19539 ^ n12547 ^ n12168 ;
  assign n19541 = ( n5904 & n6618 ) | ( n5904 & n19540 ) | ( n6618 & n19540 ) ;
  assign n19542 = n11257 ^ n3054 ^ n2502 ;
  assign n19543 = n19542 ^ n18103 ^ n765 ;
  assign n19544 = n6050 ^ n5288 ^ n4662 ;
  assign n19545 = n19544 ^ n7593 ^ 1'b0 ;
  assign n19546 = n16031 ^ n1968 ^ 1'b0 ;
  assign n19547 = n6505 & n19546 ;
  assign n19548 = ( ~n19045 & n19545 ) | ( ~n19045 & n19547 ) | ( n19545 & n19547 ) ;
  assign n19549 = n9703 ^ n8329 ^ n6698 ;
  assign n19550 = ( ~n7952 & n15784 ) | ( ~n7952 & n19549 ) | ( n15784 & n19549 ) ;
  assign n19551 = n18479 ^ n16587 ^ n15272 ;
  assign n19555 = n8721 | n9815 ;
  assign n19556 = n6733 & ~n19555 ;
  assign n19557 = n19556 ^ n5389 ^ n3377 ;
  assign n19552 = n9541 ^ n6649 ^ 1'b0 ;
  assign n19553 = n5772 | n19552 ;
  assign n19554 = n19553 ^ n1627 ^ n1452 ;
  assign n19558 = n19557 ^ n19554 ^ n2656 ;
  assign n19559 = ( n4173 & n4287 ) | ( n4173 & n4530 ) | ( n4287 & n4530 ) ;
  assign n19560 = ( n8189 & n16654 ) | ( n8189 & n19559 ) | ( n16654 & n19559 ) ;
  assign n19561 = n4813 ^ n224 ^ 1'b0 ;
  assign n19562 = n717 & n19561 ;
  assign n19563 = n447 | n19562 ;
  assign n19564 = n19563 ^ n17751 ^ 1'b0 ;
  assign n19568 = n17389 | n19228 ;
  assign n19569 = n19568 ^ n17756 ^ 1'b0 ;
  assign n19566 = n4708 ^ n4326 ^ n2116 ;
  assign n19565 = n10913 ^ n6516 ^ n6441 ;
  assign n19567 = n19566 ^ n19565 ^ n10796 ;
  assign n19570 = n19569 ^ n19567 ^ n1410 ;
  assign n19571 = n11858 ^ n10664 ^ 1'b0 ;
  assign n19572 = n17814 | n19571 ;
  assign n19573 = n19570 & ~n19572 ;
  assign n19574 = ( n374 & n11161 ) | ( n374 & ~n15976 ) | ( n11161 & ~n15976 ) ;
  assign n19575 = ( n9296 & ~n11216 ) | ( n9296 & n19574 ) | ( ~n11216 & n19574 ) ;
  assign n19576 = n7134 & n18610 ;
  assign n19577 = n19576 ^ n2788 ^ 1'b0 ;
  assign n19578 = n19577 ^ n3272 ^ n470 ;
  assign n19579 = n9146 & n9639 ;
  assign n19580 = ~n173 & n6950 ;
  assign n19581 = ( x12 & n7003 ) | ( x12 & ~n19580 ) | ( n7003 & ~n19580 ) ;
  assign n19582 = n13402 ^ n5920 ^ n3174 ;
  assign n19583 = n19582 ^ n14531 ^ 1'b0 ;
  assign n19584 = n413 | n15768 ;
  assign n19585 = n19583 | n19584 ;
  assign n19586 = ~n954 & n4505 ;
  assign n19587 = n10740 & n19586 ;
  assign n19588 = n5478 & ~n19587 ;
  assign n19589 = n11553 & n13027 ;
  assign n19590 = ( n3830 & n6110 ) | ( n3830 & n16768 ) | ( n6110 & n16768 ) ;
  assign n19591 = ( n2933 & ~n3909 ) | ( n2933 & n4737 ) | ( ~n3909 & n4737 ) ;
  assign n19592 = ( ~n6520 & n19590 ) | ( ~n6520 & n19591 ) | ( n19590 & n19591 ) ;
  assign n19593 = ( n4189 & n13279 ) | ( n4189 & n17958 ) | ( n13279 & n17958 ) ;
  assign n19594 = n419 & ~n9653 ;
  assign n19597 = n2450 & n4222 ;
  assign n19598 = ~n5714 & n19597 ;
  assign n19599 = ( n2737 & ~n9511 ) | ( n2737 & n11515 ) | ( ~n9511 & n11515 ) ;
  assign n19600 = ( n15049 & n19598 ) | ( n15049 & ~n19599 ) | ( n19598 & ~n19599 ) ;
  assign n19595 = n4379 ^ n2006 ^ n1264 ;
  assign n19596 = n19595 ^ n18440 ^ n795 ;
  assign n19601 = n19600 ^ n19596 ^ n164 ;
  assign n19602 = n14768 ^ n14403 ^ 1'b0 ;
  assign n19603 = n8607 ^ n8568 ^ n1103 ;
  assign n19604 = ~n1756 & n19603 ;
  assign n19605 = n4162 & n19604 ;
  assign n19606 = n7406 | n19605 ;
  assign n19607 = n15513 ^ n10417 ^ n9729 ;
  assign n19608 = n11526 ^ n4644 ^ 1'b0 ;
  assign n19609 = n3074 | n19608 ;
  assign n19610 = n14166 ^ n3539 ^ 1'b0 ;
  assign n19611 = n6974 & ~n19610 ;
  assign n19612 = ~n2230 & n19611 ;
  assign n19613 = n19609 & n19612 ;
  assign n19614 = ( n16768 & ~n18448 ) | ( n16768 & n19613 ) | ( ~n18448 & n19613 ) ;
  assign n19615 = n19298 ^ n2709 ^ n1791 ;
  assign n19616 = n19615 ^ n8989 ^ n2628 ;
  assign n19617 = ( n12414 & n12812 ) | ( n12414 & n19616 ) | ( n12812 & n19616 ) ;
  assign n19618 = ( n6753 & n8084 ) | ( n6753 & ~n8325 ) | ( n8084 & ~n8325 ) ;
  assign n19619 = n6443 & ~n19618 ;
  assign n19620 = n15519 & n19619 ;
  assign n19621 = ( n584 & n6942 ) | ( n584 & ~n13560 ) | ( n6942 & ~n13560 ) ;
  assign n19623 = ( n1089 & n1467 ) | ( n1089 & ~n8293 ) | ( n1467 & ~n8293 ) ;
  assign n19622 = n10765 & ~n13452 ;
  assign n19624 = n19623 ^ n19622 ^ 1'b0 ;
  assign n19625 = n12688 | n19624 ;
  assign n19626 = n19621 | n19625 ;
  assign n19627 = ( n1444 & n3385 ) | ( n1444 & ~n9023 ) | ( n3385 & ~n9023 ) ;
  assign n19628 = ~n11359 & n19627 ;
  assign n19629 = n8611 ^ n6467 ^ n5412 ;
  assign n19630 = n19629 ^ n14432 ^ n3156 ;
  assign n19631 = ~n16076 & n18111 ;
  assign n19632 = ( ~n3767 & n9485 ) | ( ~n3767 & n19631 ) | ( n9485 & n19631 ) ;
  assign n19633 = n1232 & ~n14610 ;
  assign n19636 = n4923 ^ n4413 ^ n2719 ;
  assign n19634 = ~n3867 & n13247 ;
  assign n19635 = ( n735 & ~n3385 ) | ( n735 & n19634 ) | ( ~n3385 & n19634 ) ;
  assign n19637 = n19636 ^ n19635 ^ n10799 ;
  assign n19638 = ~n4633 & n16563 ;
  assign n19639 = n19638 ^ n8858 ^ 1'b0 ;
  assign n19640 = n19639 ^ n12093 ^ n8380 ;
  assign n19641 = n2036 ^ n1762 ^ n339 ;
  assign n19642 = n19457 ^ n14940 ^ n445 ;
  assign n19643 = ( ~n14477 & n19641 ) | ( ~n14477 & n19642 ) | ( n19641 & n19642 ) ;
  assign n19644 = ( n1061 & n6767 ) | ( n1061 & ~n9981 ) | ( n6767 & ~n9981 ) ;
  assign n19645 = n4321 ^ n1898 ^ 1'b0 ;
  assign n19646 = n19645 ^ n725 ^ 1'b0 ;
  assign n19647 = ~n4085 & n19646 ;
  assign n19648 = n19647 ^ n3147 ^ n2889 ;
  assign n19649 = ( n4948 & n8188 ) | ( n4948 & n19648 ) | ( n8188 & n19648 ) ;
  assign n19651 = n6013 & n15852 ;
  assign n19650 = ( n7730 & ~n11397 ) | ( n7730 & n17433 ) | ( ~n11397 & n17433 ) ;
  assign n19652 = n19651 ^ n19650 ^ n2612 ;
  assign n19653 = ( n1767 & n3172 ) | ( n1767 & ~n17354 ) | ( n3172 & ~n17354 ) ;
  assign n19662 = ( n1858 & n3984 ) | ( n1858 & ~n13084 ) | ( n3984 & ~n13084 ) ;
  assign n19657 = ( n1998 & n3153 ) | ( n1998 & ~n8349 ) | ( n3153 & ~n8349 ) ;
  assign n19658 = n6689 ^ n4486 ^ 1'b0 ;
  assign n19659 = n8801 & ~n19658 ;
  assign n19660 = ( ~n7657 & n19657 ) | ( ~n7657 & n19659 ) | ( n19657 & n19659 ) ;
  assign n19654 = ( ~n2088 & n5841 ) | ( ~n2088 & n15463 ) | ( n5841 & n15463 ) ;
  assign n19655 = n19654 ^ n10013 ^ 1'b0 ;
  assign n19656 = ( n4236 & n16019 ) | ( n4236 & n19655 ) | ( n16019 & n19655 ) ;
  assign n19661 = n19660 ^ n19656 ^ n1360 ;
  assign n19663 = n19662 ^ n19661 ^ x110 ;
  assign n19664 = n1431 | n13870 ;
  assign n19665 = n19664 ^ n6956 ^ 1'b0 ;
  assign n19666 = ( ~n3518 & n19440 ) | ( ~n3518 & n19665 ) | ( n19440 & n19665 ) ;
  assign n19667 = n19666 ^ n10376 ^ n426 ;
  assign n19668 = ( n2055 & n13274 ) | ( n2055 & n15317 ) | ( n13274 & n15317 ) ;
  assign n19669 = n3904 & ~n19668 ;
  assign n19670 = ( n3484 & ~n4143 ) | ( n3484 & n12696 ) | ( ~n4143 & n12696 ) ;
  assign n19671 = ( n6681 & n14747 ) | ( n6681 & ~n16792 ) | ( n14747 & ~n16792 ) ;
  assign n19672 = ( n1927 & n15314 ) | ( n1927 & ~n19671 ) | ( n15314 & ~n19671 ) ;
  assign n19673 = n19672 ^ n9088 ^ n275 ;
  assign n19676 = ~n6318 & n12658 ;
  assign n19677 = ~n247 & n19676 ;
  assign n19674 = n11927 ^ n3948 ^ n2653 ;
  assign n19675 = ( ~n6614 & n10343 ) | ( ~n6614 & n19674 ) | ( n10343 & n19674 ) ;
  assign n19678 = n19677 ^ n19675 ^ n3096 ;
  assign n19679 = n18671 ^ n8259 ^ 1'b0 ;
  assign n19681 = n3580 & ~n3655 ;
  assign n19680 = ~n5549 & n6042 ;
  assign n19682 = n19681 ^ n19680 ^ 1'b0 ;
  assign n19683 = n6586 ^ n3566 ^ n1104 ;
  assign n19684 = n19683 ^ n10207 ^ n6060 ;
  assign n19685 = n19684 ^ n10109 ^ 1'b0 ;
  assign n19686 = ~n15571 & n19685 ;
  assign n19687 = n19686 ^ n5653 ^ 1'b0 ;
  assign n19688 = n11795 ^ n11745 ^ n7712 ;
  assign n19689 = ~n3884 & n14608 ;
  assign n19690 = ~n16827 & n19689 ;
  assign n19691 = n17305 | n19690 ;
  assign n19692 = ( n8446 & ~n19688 ) | ( n8446 & n19691 ) | ( ~n19688 & n19691 ) ;
  assign n19693 = ~n633 & n2229 ;
  assign n19694 = n19693 ^ n13312 ^ 1'b0 ;
  assign n19695 = ( n2680 & n8611 ) | ( n2680 & ~n19694 ) | ( n8611 & ~n19694 ) ;
  assign n19696 = n19695 ^ n13410 ^ n2209 ;
  assign n19697 = ( n4771 & n13384 ) | ( n4771 & ~n14388 ) | ( n13384 & ~n14388 ) ;
  assign n19707 = ( n2388 & n2670 ) | ( n2388 & n5319 ) | ( n2670 & n5319 ) ;
  assign n19706 = n16281 ^ n5922 ^ n1466 ;
  assign n19700 = ( ~n860 & n5800 ) | ( ~n860 & n7164 ) | ( n5800 & n7164 ) ;
  assign n19701 = ( n561 & n7176 ) | ( n561 & n15908 ) | ( n7176 & n15908 ) ;
  assign n19702 = n19701 ^ n3918 ^ n2958 ;
  assign n19703 = ( n4451 & n13387 ) | ( n4451 & n19702 ) | ( n13387 & n19702 ) ;
  assign n19704 = ( n4017 & n19700 ) | ( n4017 & ~n19703 ) | ( n19700 & ~n19703 ) ;
  assign n19698 = n16745 ^ n1333 ^ 1'b0 ;
  assign n19699 = n16227 & ~n19698 ;
  assign n19705 = n19704 ^ n19699 ^ 1'b0 ;
  assign n19708 = n19707 ^ n19706 ^ n19705 ;
  assign n19709 = n6534 & n7502 ;
  assign n19710 = ~n19708 & n19709 ;
  assign n19711 = n17458 ^ n1672 ^ 1'b0 ;
  assign n19712 = n3596 | n19711 ;
  assign n19713 = ( n1290 & n7651 ) | ( n1290 & n8900 ) | ( n7651 & n8900 ) ;
  assign n19714 = n7514 | n19713 ;
  assign n19715 = ~n4406 & n7575 ;
  assign n19716 = ~n19714 & n19715 ;
  assign n19717 = n3164 ^ n1247 ^ 1'b0 ;
  assign n19718 = ~n1312 & n3692 ;
  assign n19719 = n1743 & n19718 ;
  assign n19720 = n19719 ^ n10915 ^ 1'b0 ;
  assign n19723 = n12101 ^ n6250 ^ n4303 ;
  assign n19724 = ~n11847 & n19723 ;
  assign n19721 = ( n159 & ~n3702 ) | ( n159 & n9413 ) | ( ~n3702 & n9413 ) ;
  assign n19722 = n19721 ^ n4543 ^ 1'b0 ;
  assign n19725 = n19724 ^ n19722 ^ n6006 ;
  assign n19726 = n6567 ^ n3782 ^ 1'b0 ;
  assign n19727 = n10382 & n19726 ;
  assign n19728 = n5813 ^ n2313 ^ n1820 ;
  assign n19729 = ( n2829 & ~n11647 ) | ( n2829 & n19728 ) | ( ~n11647 & n19728 ) ;
  assign n19730 = ( n7683 & n19727 ) | ( n7683 & ~n19729 ) | ( n19727 & ~n19729 ) ;
  assign n19731 = n10610 ^ n9036 ^ n4289 ;
  assign n19732 = n1354 & n10359 ;
  assign n19733 = n19731 & n19732 ;
  assign n19734 = n19733 ^ n15484 ^ n11436 ;
  assign n19735 = n4940 & ~n7852 ;
  assign n19736 = n18664 ^ n6972 ^ n2480 ;
  assign n19737 = n17991 | n19736 ;
  assign n19738 = n19735 & ~n19737 ;
  assign n19739 = n19738 ^ n14876 ^ n3246 ;
  assign n19740 = n10000 & ~n19739 ;
  assign n19741 = n19740 ^ n231 ^ 1'b0 ;
  assign n19743 = ( ~n794 & n13200 ) | ( ~n794 & n19091 ) | ( n13200 & n19091 ) ;
  assign n19744 = ( ~n8773 & n18577 ) | ( ~n8773 & n19743 ) | ( n18577 & n19743 ) ;
  assign n19742 = n875 | n12328 ;
  assign n19745 = n19744 ^ n19742 ^ 1'b0 ;
  assign n19746 = ( n968 & ~n17634 ) | ( n968 & n18961 ) | ( ~n17634 & n18961 ) ;
  assign n19749 = n11152 ^ n6214 ^ n466 ;
  assign n19747 = ~n804 & n7614 ;
  assign n19748 = n19747 ^ n3141 ^ 1'b0 ;
  assign n19750 = n19749 ^ n19748 ^ n5348 ;
  assign n19751 = n19750 ^ n6469 ^ 1'b0 ;
  assign n19752 = ( ~n12438 & n16709 ) | ( ~n12438 & n19751 ) | ( n16709 & n19751 ) ;
  assign n19753 = n17432 ^ n10528 ^ n7327 ;
  assign n19754 = n7192 & n18211 ;
  assign n19757 = ~n3569 & n6764 ;
  assign n19755 = n3307 ^ n278 ^ 1'b0 ;
  assign n19756 = ( n2046 & ~n15532 ) | ( n2046 & n19755 ) | ( ~n15532 & n19755 ) ;
  assign n19758 = n19757 ^ n19756 ^ n576 ;
  assign n19759 = n13300 ^ n12158 ^ 1'b0 ;
  assign n19760 = ~n1427 & n19759 ;
  assign n19761 = n19760 ^ n569 ^ 1'b0 ;
  assign n19762 = ( n12715 & n19758 ) | ( n12715 & n19761 ) | ( n19758 & n19761 ) ;
  assign n19763 = ( n3095 & n14877 ) | ( n3095 & n19762 ) | ( n14877 & n19762 ) ;
  assign n19764 = ( n6116 & n19754 ) | ( n6116 & ~n19763 ) | ( n19754 & ~n19763 ) ;
  assign n19765 = n11677 | n13384 ;
  assign n19766 = x119 & n8166 ;
  assign n19767 = n5772 & n19766 ;
  assign n19768 = n19767 ^ n17150 ^ n5892 ;
  assign n19769 = n19768 ^ n14592 ^ n10252 ;
  assign n19770 = n9885 ^ n5507 ^ 1'b0 ;
  assign n19771 = n8610 | n19770 ;
  assign n19772 = n19771 ^ n1745 ^ 1'b0 ;
  assign n19773 = n1844 | n2987 ;
  assign n19774 = ( n430 & ~n2741 ) | ( n430 & n19773 ) | ( ~n2741 & n19773 ) ;
  assign n19775 = ( n5697 & n10071 ) | ( n5697 & ~n19774 ) | ( n10071 & ~n19774 ) ;
  assign n19776 = ( n1466 & n3422 ) | ( n1466 & ~n3909 ) | ( n3422 & ~n3909 ) ;
  assign n19777 = n718 | n15447 ;
  assign n19778 = n19776 & ~n19777 ;
  assign n19779 = n16248 ^ n8042 ^ n7769 ;
  assign n19780 = ( n6067 & n19778 ) | ( n6067 & n19779 ) | ( n19778 & n19779 ) ;
  assign n19781 = ( ~n3112 & n4331 ) | ( ~n3112 & n19780 ) | ( n4331 & n19780 ) ;
  assign n19784 = ( ~n1189 & n4201 ) | ( ~n1189 & n12205 ) | ( n4201 & n12205 ) ;
  assign n19782 = n10504 ^ n5572 ^ n1377 ;
  assign n19783 = ( ~n2788 & n9035 ) | ( ~n2788 & n19782 ) | ( n9035 & n19782 ) ;
  assign n19785 = n19784 ^ n19783 ^ n701 ;
  assign n19786 = ( n14779 & ~n17058 ) | ( n14779 & n19785 ) | ( ~n17058 & n19785 ) ;
  assign n19787 = n4855 ^ n3392 ^ n2834 ;
  assign n19788 = n19787 ^ n6371 ^ 1'b0 ;
  assign n19789 = n233 & ~n7004 ;
  assign n19790 = n19789 ^ n3386 ^ 1'b0 ;
  assign n19791 = n19788 | n19790 ;
  assign n19792 = n6392 & ~n11247 ;
  assign n19793 = n19792 ^ n17644 ^ 1'b0 ;
  assign n19799 = n2847 & ~n3754 ;
  assign n19800 = n1115 & n19799 ;
  assign n19801 = ( ~n12036 & n15247 ) | ( ~n12036 & n19800 ) | ( n15247 & n19800 ) ;
  assign n19794 = ( n1365 & n6917 ) | ( n1365 & ~n6933 ) | ( n6917 & ~n6933 ) ;
  assign n19795 = ( ~n3119 & n3949 ) | ( ~n3119 & n19794 ) | ( n3949 & n19794 ) ;
  assign n19796 = n19795 ^ n18943 ^ n2943 ;
  assign n19797 = n17976 ^ n5123 ^ n2835 ;
  assign n19798 = n19796 & ~n19797 ;
  assign n19802 = n19801 ^ n19798 ^ 1'b0 ;
  assign n19803 = ( n7427 & n8330 ) | ( n7427 & n10046 ) | ( n8330 & n10046 ) ;
  assign n19804 = n19803 ^ n11375 ^ 1'b0 ;
  assign n19805 = ( n3664 & n5001 ) | ( n3664 & ~n6292 ) | ( n5001 & ~n6292 ) ;
  assign n19806 = n19805 ^ n10041 ^ n9458 ;
  assign n19807 = ( n6057 & n8346 ) | ( n6057 & n19806 ) | ( n8346 & n19806 ) ;
  assign n19808 = n1631 | n3110 ;
  assign n19809 = ( ~n11656 & n12112 ) | ( ~n11656 & n19808 ) | ( n12112 & n19808 ) ;
  assign n19810 = ( ~n13696 & n14780 ) | ( ~n13696 & n18657 ) | ( n14780 & n18657 ) ;
  assign n19813 = ( n669 & n1409 ) | ( n669 & n4365 ) | ( n1409 & n4365 ) ;
  assign n19812 = ( n926 & n4030 ) | ( n926 & ~n7034 ) | ( n4030 & ~n7034 ) ;
  assign n19811 = ( n9191 & n14443 ) | ( n9191 & ~n16038 ) | ( n14443 & ~n16038 ) ;
  assign n19814 = n19813 ^ n19812 ^ n19811 ;
  assign n19815 = ( ~n4410 & n9391 ) | ( ~n4410 & n14574 ) | ( n9391 & n14574 ) ;
  assign n19818 = ( n6021 & n7697 ) | ( n6021 & n11457 ) | ( n7697 & n11457 ) ;
  assign n19816 = n13607 ^ n8152 ^ n5474 ;
  assign n19817 = ( n3876 & ~n16357 ) | ( n3876 & n19816 ) | ( ~n16357 & n19816 ) ;
  assign n19819 = n19818 ^ n19817 ^ n19112 ;
  assign n19820 = n10927 ^ n4403 ^ n1910 ;
  assign n19821 = n19820 ^ n12082 ^ n2839 ;
  assign n19822 = ~n566 & n2686 ;
  assign n19823 = ( ~n5506 & n6014 ) | ( ~n5506 & n19822 ) | ( n6014 & n19822 ) ;
  assign n19824 = n19823 ^ n1896 ^ 1'b0 ;
  assign n19825 = n19824 ^ n10933 ^ n254 ;
  assign n19826 = ( n2570 & ~n2571 ) | ( n2570 & n19825 ) | ( ~n2571 & n19825 ) ;
  assign n19827 = n5164 & n10636 ;
  assign n19828 = ( n3423 & n5871 ) | ( n3423 & n12504 ) | ( n5871 & n12504 ) ;
  assign n19829 = ( n4958 & ~n7985 ) | ( n4958 & n18039 ) | ( ~n7985 & n18039 ) ;
  assign n19830 = ( n12953 & ~n19828 ) | ( n12953 & n19829 ) | ( ~n19828 & n19829 ) ;
  assign n19831 = n2610 ^ n1742 ^ n1326 ;
  assign n19832 = n15253 ^ n14122 ^ n3900 ;
  assign n19833 = ( n3856 & n19831 ) | ( n3856 & n19832 ) | ( n19831 & n19832 ) ;
  assign n19837 = n12384 ^ n9797 ^ n2831 ;
  assign n19834 = n5668 ^ n1874 ^ 1'b0 ;
  assign n19835 = n8599 & n19834 ;
  assign n19836 = n19835 ^ n8787 ^ n517 ;
  assign n19838 = n19837 ^ n19836 ^ 1'b0 ;
  assign n19839 = ( n1387 & n2947 ) | ( n1387 & ~n2977 ) | ( n2947 & ~n2977 ) ;
  assign n19840 = ( n4042 & n11504 ) | ( n4042 & n19839 ) | ( n11504 & n19839 ) ;
  assign n19841 = n18898 ^ n4604 ^ 1'b0 ;
  assign n19842 = n19841 ^ n19544 ^ n7315 ;
  assign n19843 = n19842 ^ n16685 ^ n14387 ;
  assign n19844 = ( n2156 & n3263 ) | ( n2156 & n18811 ) | ( n3263 & n18811 ) ;
  assign n19845 = n7604 ^ n5977 ^ n3485 ;
  assign n19846 = ( n6510 & n12553 ) | ( n6510 & ~n14800 ) | ( n12553 & ~n14800 ) ;
  assign n19847 = n19846 ^ n9905 ^ n381 ;
  assign n19848 = n763 & n2739 ;
  assign n19849 = n19848 ^ n564 ^ 1'b0 ;
  assign n19852 = ~n2912 & n12293 ;
  assign n19853 = ~n16993 & n19852 ;
  assign n19850 = ~n12496 & n15613 ;
  assign n19851 = n19850 ^ n8541 ^ n4926 ;
  assign n19854 = n19853 ^ n19851 ^ n11470 ;
  assign n19855 = n13511 & n19854 ;
  assign n19856 = n19855 ^ n5474 ^ 1'b0 ;
  assign n19857 = ( ~n1778 & n5809 ) | ( ~n1778 & n7148 ) | ( n5809 & n7148 ) ;
  assign n19858 = n19857 ^ n5320 ^ 1'b0 ;
  assign n19863 = ( ~n1918 & n5487 ) | ( ~n1918 & n14864 ) | ( n5487 & n14864 ) ;
  assign n19862 = n12981 ^ n9935 ^ n2875 ;
  assign n19859 = n7456 ^ n1284 ^ n1239 ;
  assign n19860 = n13017 & n19859 ;
  assign n19861 = ( n6060 & n10234 ) | ( n6060 & ~n19860 ) | ( n10234 & ~n19860 ) ;
  assign n19864 = n19863 ^ n19862 ^ n19861 ;
  assign n19867 = n2016 & n7364 ;
  assign n19865 = ~n2502 & n11380 ;
  assign n19866 = n19865 ^ n7447 ^ n2391 ;
  assign n19868 = n19867 ^ n19866 ^ n14205 ;
  assign n19870 = ( n1139 & n4728 ) | ( n1139 & n7458 ) | ( n4728 & n7458 ) ;
  assign n19869 = n18168 ^ n9942 ^ 1'b0 ;
  assign n19871 = n19870 ^ n19869 ^ 1'b0 ;
  assign n19876 = n11279 ^ n9932 ^ n1457 ;
  assign n19877 = n19876 ^ n6443 ^ n4421 ;
  assign n19878 = ~n5498 & n19877 ;
  assign n19872 = n9332 ^ n4478 ^ n2530 ;
  assign n19873 = n8604 ^ n4396 ^ n834 ;
  assign n19874 = n19872 | n19873 ;
  assign n19875 = n8885 | n19874 ;
  assign n19879 = n19878 ^ n19875 ^ n6198 ;
  assign n19880 = n11179 ^ n6292 ^ n5008 ;
  assign n19885 = ( ~x6 & n6701 ) | ( ~x6 & n11276 ) | ( n6701 & n11276 ) ;
  assign n19881 = n16521 ^ n10962 ^ n4118 ;
  assign n19882 = n19881 ^ n11415 ^ n2000 ;
  assign n19883 = n6464 ^ n930 ^ 1'b0 ;
  assign n19884 = n19882 | n19883 ;
  assign n19886 = n19885 ^ n19884 ^ 1'b0 ;
  assign n19891 = n5634 ^ n3722 ^ n499 ;
  assign n19888 = ( n1303 & ~n5410 ) | ( n1303 & n9191 ) | ( ~n5410 & n9191 ) ;
  assign n19889 = ~n4744 & n19888 ;
  assign n19887 = ( n336 & n8100 ) | ( n336 & ~n13639 ) | ( n8100 & ~n13639 ) ;
  assign n19890 = n19889 ^ n19887 ^ n6256 ;
  assign n19892 = n19891 ^ n19890 ^ n6793 ;
  assign n19893 = ( n5306 & ~n10646 ) | ( n5306 & n12773 ) | ( ~n10646 & n12773 ) ;
  assign n19898 = n3872 ^ n935 ^ 1'b0 ;
  assign n19899 = n2145 & ~n19898 ;
  assign n19900 = ( ~x83 & n4676 ) | ( ~x83 & n19899 ) | ( n4676 & n19899 ) ;
  assign n19901 = n13781 ^ n6447 ^ n6280 ;
  assign n19902 = n19901 ^ n16281 ^ n5146 ;
  assign n19903 = ( n4838 & n19900 ) | ( n4838 & n19902 ) | ( n19900 & n19902 ) ;
  assign n19895 = n5903 & n7975 ;
  assign n19896 = n19895 ^ n783 ^ 1'b0 ;
  assign n19897 = n4087 | n19896 ;
  assign n19904 = n19903 ^ n19897 ^ 1'b0 ;
  assign n19894 = n15483 ^ n7257 ^ 1'b0 ;
  assign n19905 = n19904 ^ n19894 ^ n17558 ;
  assign n19906 = ( n4156 & n8056 ) | ( n4156 & n12337 ) | ( n8056 & n12337 ) ;
  assign n19907 = n4463 & n19906 ;
  assign n19908 = n10356 & ~n18190 ;
  assign n19909 = n19908 ^ n11735 ^ 1'b0 ;
  assign n19910 = n668 & ~n6921 ;
  assign n19911 = n19910 ^ n14249 ^ n4606 ;
  assign n19912 = n16746 ^ n12594 ^ n4459 ;
  assign n19913 = n19911 & n19912 ;
  assign n19914 = n15364 & n15785 ;
  assign n19918 = n766 & ~n6026 ;
  assign n19919 = n19918 ^ n1775 ^ 1'b0 ;
  assign n19920 = ( ~n10960 & n14974 ) | ( ~n10960 & n19919 ) | ( n14974 & n19919 ) ;
  assign n19915 = n3258 & ~n8081 ;
  assign n19916 = n4061 ^ n2733 ^ n1716 ;
  assign n19917 = ( ~n8757 & n19915 ) | ( ~n8757 & n19916 ) | ( n19915 & n19916 ) ;
  assign n19921 = n19920 ^ n19917 ^ n17125 ;
  assign n19926 = n995 | n16747 ;
  assign n19922 = ~n2468 & n4622 ;
  assign n19923 = n19922 ^ n6797 ^ n6045 ;
  assign n19924 = n19923 ^ n4516 ^ 1'b0 ;
  assign n19925 = ~n13981 & n19924 ;
  assign n19927 = n19926 ^ n19925 ^ n4569 ;
  assign n19928 = n11207 ^ n3691 ^ 1'b0 ;
  assign n19929 = ~n12355 & n18388 ;
  assign n19930 = n18212 ^ n5604 ^ n2918 ;
  assign n19931 = n19930 ^ n7614 ^ n875 ;
  assign n19932 = ( n4301 & n5825 ) | ( n4301 & n19931 ) | ( n5825 & n19931 ) ;
  assign n19933 = n2893 ^ x105 ^ 1'b0 ;
  assign n19934 = n5809 & ~n19933 ;
  assign n19936 = n14177 ^ n5367 ^ n2039 ;
  assign n19935 = ( ~n3136 & n4822 ) | ( ~n3136 & n10659 ) | ( n4822 & n10659 ) ;
  assign n19937 = n19936 ^ n19935 ^ n19016 ;
  assign n19938 = ( n9153 & ~n11046 ) | ( n9153 & n19937 ) | ( ~n11046 & n19937 ) ;
  assign n19939 = n5980 ^ n4558 ^ 1'b0 ;
  assign n19940 = n18316 | n19939 ;
  assign n19941 = ( ~n3110 & n19161 ) | ( ~n3110 & n19940 ) | ( n19161 & n19940 ) ;
  assign n19942 = n19941 ^ n19109 ^ n11847 ;
  assign n19943 = n18292 ^ n6985 ^ n2036 ;
  assign n19944 = n5551 ^ n2573 ^ n2222 ;
  assign n19945 = n10115 | n13371 ;
  assign n19946 = n11093 | n19945 ;
  assign n19947 = n411 | n1784 ;
  assign n19948 = ( n9455 & ~n19946 ) | ( n9455 & n19947 ) | ( ~n19946 & n19947 ) ;
  assign n19949 = n2375 & ~n19833 ;
  assign n19950 = n19949 ^ n5173 ^ 1'b0 ;
  assign n19951 = n17244 ^ n6664 ^ 1'b0 ;
  assign n19952 = n513 & n19951 ;
  assign n19954 = ( ~n12694 & n14027 ) | ( ~n12694 & n14391 ) | ( n14027 & n14391 ) ;
  assign n19953 = ~n7385 & n11226 ;
  assign n19955 = n19954 ^ n19953 ^ 1'b0 ;
  assign n19956 = n10331 | n10866 ;
  assign n19957 = n19956 ^ n7007 ^ 1'b0 ;
  assign n19958 = n19957 ^ n18940 ^ 1'b0 ;
  assign n19959 = n13729 ^ n1000 ^ 1'b0 ;
  assign n19960 = ( ~n17260 & n19958 ) | ( ~n17260 & n19959 ) | ( n19958 & n19959 ) ;
  assign n19961 = n12112 ^ n8809 ^ n454 ;
  assign n19962 = n11528 ^ n8996 ^ n2866 ;
  assign n19963 = ( n15420 & n17515 ) | ( n15420 & ~n19962 ) | ( n17515 & ~n19962 ) ;
  assign n19964 = ( n11871 & n14703 ) | ( n11871 & ~n18884 ) | ( n14703 & ~n18884 ) ;
  assign n19965 = ( n1253 & n7924 ) | ( n1253 & n12570 ) | ( n7924 & n12570 ) ;
  assign n19966 = n19965 ^ n3532 ^ 1'b0 ;
  assign n19967 = n19964 & ~n19966 ;
  assign n19968 = n10273 ^ n7079 ^ 1'b0 ;
  assign n19969 = n8008 & ~n19968 ;
  assign n19970 = n19969 ^ n10616 ^ 1'b0 ;
  assign n19971 = ( n157 & n7111 ) | ( n157 & ~n11569 ) | ( n7111 & ~n11569 ) ;
  assign n19973 = n4175 ^ n3540 ^ n2676 ;
  assign n19974 = n4617 & ~n19973 ;
  assign n19975 = n19974 ^ n1662 ^ 1'b0 ;
  assign n19976 = ( n8599 & n14420 ) | ( n8599 & n19975 ) | ( n14420 & n19975 ) ;
  assign n19977 = ( n2623 & ~n11213 ) | ( n2623 & n19976 ) | ( ~n11213 & n19976 ) ;
  assign n19972 = n15683 ^ n13548 ^ n9197 ;
  assign n19978 = n19977 ^ n19972 ^ n12859 ;
  assign n19979 = n17674 ^ n8678 ^ n6469 ;
  assign n19980 = n8449 ^ n2879 ^ n2131 ;
  assign n19981 = n19980 ^ n13424 ^ n545 ;
  assign n19982 = n19981 ^ n18628 ^ 1'b0 ;
  assign n19983 = ~n5437 & n19982 ;
  assign n19984 = n18435 ^ n2529 ^ n2392 ;
  assign n19985 = n19984 ^ n5014 ^ n720 ;
  assign n19986 = ( n3649 & ~n8527 ) | ( n3649 & n16313 ) | ( ~n8527 & n16313 ) ;
  assign n19987 = n11358 | n19986 ;
  assign n19988 = n19985 & ~n19987 ;
  assign n19989 = ~n1852 & n3732 ;
  assign n19990 = n19989 ^ n442 ^ 1'b0 ;
  assign n19991 = x41 & n9433 ;
  assign n19992 = ~n5667 & n19991 ;
  assign n19993 = n6400 & n19992 ;
  assign n19994 = n19993 ^ n12040 ^ n1670 ;
  assign n19995 = ( n6976 & n19990 ) | ( n6976 & ~n19994 ) | ( n19990 & ~n19994 ) ;
  assign n19996 = ( n2530 & n9947 ) | ( n2530 & n19995 ) | ( n9947 & n19995 ) ;
  assign n19997 = n6301 ^ n5693 ^ n4163 ;
  assign n19998 = n9520 ^ n8595 ^ 1'b0 ;
  assign n19999 = x28 & ~n19998 ;
  assign n20000 = ( n10205 & n19997 ) | ( n10205 & ~n19999 ) | ( n19997 & ~n19999 ) ;
  assign n20001 = n4581 ^ n2878 ^ 1'b0 ;
  assign n20002 = n1908 | n20001 ;
  assign n20003 = ( n4520 & n10798 ) | ( n4520 & ~n20002 ) | ( n10798 & ~n20002 ) ;
  assign n20004 = ( n3257 & n14498 ) | ( n3257 & n18330 ) | ( n14498 & n18330 ) ;
  assign n20005 = ( n5951 & n13120 ) | ( n5951 & ~n20004 ) | ( n13120 & ~n20004 ) ;
  assign n20006 = ( n3432 & ~n14897 ) | ( n3432 & n14940 ) | ( ~n14897 & n14940 ) ;
  assign n20007 = ( n5664 & n11158 ) | ( n5664 & n20006 ) | ( n11158 & n20006 ) ;
  assign n20008 = n19009 ^ n4070 ^ 1'b0 ;
  assign n20009 = ~n4541 & n20008 ;
  assign n20010 = n11928 & n19177 ;
  assign n20011 = n20010 ^ n15133 ^ 1'b0 ;
  assign n20012 = n3805 ^ n3785 ^ n3283 ;
  assign n20013 = n4494 ^ n2274 ^ n229 ;
  assign n20014 = ( n10526 & ~n19167 ) | ( n10526 & n20013 ) | ( ~n19167 & n20013 ) ;
  assign n20015 = n20014 ^ n4366 ^ 1'b0 ;
  assign n20016 = n10348 ^ n3049 ^ n155 ;
  assign n20017 = n20016 ^ n6637 ^ 1'b0 ;
  assign n20018 = ( n10410 & n13663 ) | ( n10410 & n16427 ) | ( n13663 & n16427 ) ;
  assign n20019 = ( n12932 & ~n20017 ) | ( n12932 & n20018 ) | ( ~n20017 & n20018 ) ;
  assign n20020 = n5332 & n17937 ;
  assign n20021 = n1577 ^ x21 ^ 1'b0 ;
  assign n20022 = n17556 & n20021 ;
  assign n20023 = ~n3140 & n6150 ;
  assign n20024 = ~n4513 & n20023 ;
  assign n20025 = n8182 | n20024 ;
  assign n20026 = n17809 ^ n6038 ^ n3135 ;
  assign n20027 = n14653 ^ n8438 ^ n8129 ;
  assign n20029 = ( n4671 & n8225 ) | ( n4671 & n15429 ) | ( n8225 & n15429 ) ;
  assign n20028 = n15690 ^ n11081 ^ 1'b0 ;
  assign n20030 = n20029 ^ n20028 ^ 1'b0 ;
  assign n20031 = n4773 | n20030 ;
  assign n20032 = n20031 ^ n4697 ^ n4291 ;
  assign n20033 = n3707 | n7321 ;
  assign n20034 = n4998 | n20033 ;
  assign n20035 = n20034 ^ n13513 ^ 1'b0 ;
  assign n20036 = n10739 ^ n9134 ^ 1'b0 ;
  assign n20037 = n2742 & n20036 ;
  assign n20038 = n20037 ^ n1878 ^ 1'b0 ;
  assign n20039 = n588 & n8684 ;
  assign n20040 = n20039 ^ n9903 ^ 1'b0 ;
  assign n20041 = n20040 ^ n17209 ^ n10059 ;
  assign n20042 = n14478 ^ n11568 ^ 1'b0 ;
  assign n20043 = n20041 | n20042 ;
  assign n20044 = n9161 & n14887 ;
  assign n20045 = n20044 ^ n5884 ^ 1'b0 ;
  assign n20046 = n5977 & n8671 ;
  assign n20047 = n20045 & n20046 ;
  assign n20048 = n3691 ^ n2642 ^ n1016 ;
  assign n20049 = ( ~n2232 & n11216 ) | ( ~n2232 & n20048 ) | ( n11216 & n20048 ) ;
  assign n20050 = ( n6873 & ~n12126 ) | ( n6873 & n20049 ) | ( ~n12126 & n20049 ) ;
  assign n20051 = ( n5106 & n9829 ) | ( n5106 & n20050 ) | ( n9829 & n20050 ) ;
  assign n20052 = n1009 & n20051 ;
  assign n20058 = ( ~n370 & n5800 ) | ( ~n370 & n6087 ) | ( n5800 & n6087 ) ;
  assign n20055 = n8925 ^ n1342 ^ 1'b0 ;
  assign n20056 = n6102 | n20055 ;
  assign n20053 = ( n9083 & n11279 ) | ( n9083 & n17632 ) | ( n11279 & n17632 ) ;
  assign n20054 = n20053 ^ n7902 ^ n1445 ;
  assign n20057 = n20056 ^ n20054 ^ n11249 ;
  assign n20059 = n20058 ^ n20057 ^ n13958 ;
  assign n20061 = n10832 ^ n6184 ^ x94 ;
  assign n20060 = n18304 ^ n15301 ^ n7146 ;
  assign n20062 = n20061 ^ n20060 ^ n19968 ;
  assign n20063 = n13489 ^ n9064 ^ 1'b0 ;
  assign n20064 = ( ~n6350 & n6852 ) | ( ~n6350 & n12708 ) | ( n6852 & n12708 ) ;
  assign n20065 = ( n6202 & n7704 ) | ( n6202 & n20064 ) | ( n7704 & n20064 ) ;
  assign n20067 = ( n355 & n4331 ) | ( n355 & n6369 ) | ( n4331 & n6369 ) ;
  assign n20068 = ( ~n5787 & n5837 ) | ( ~n5787 & n20067 ) | ( n5837 & n20067 ) ;
  assign n20066 = ( n926 & ~n3977 ) | ( n926 & n11108 ) | ( ~n3977 & n11108 ) ;
  assign n20069 = n20068 ^ n20066 ^ 1'b0 ;
  assign n20070 = n18608 & ~n20069 ;
  assign n20071 = ~n15581 & n20070 ;
  assign n20072 = n997 | n14153 ;
  assign n20073 = n20072 ^ n4640 ^ 1'b0 ;
  assign n20074 = n11794 ^ n7344 ^ 1'b0 ;
  assign n20075 = n4786 | n20074 ;
  assign n20076 = n20075 ^ n11153 ^ n2392 ;
  assign n20077 = n11598 & n20076 ;
  assign n20079 = n314 & ~n5256 ;
  assign n20080 = n20079 ^ n7329 ^ 1'b0 ;
  assign n20078 = ( n4291 & ~n6065 ) | ( n4291 & n10358 ) | ( ~n6065 & n10358 ) ;
  assign n20081 = n20080 ^ n20078 ^ n15582 ;
  assign n20082 = ( ~n315 & n6628 ) | ( ~n315 & n13052 ) | ( n6628 & n13052 ) ;
  assign n20083 = ~n12745 & n20082 ;
  assign n20093 = ( n247 & n3182 ) | ( n247 & ~n7450 ) | ( n3182 & ~n7450 ) ;
  assign n20094 = ( ~n2351 & n10504 ) | ( ~n2351 & n11054 ) | ( n10504 & n11054 ) ;
  assign n20095 = n752 & n17675 ;
  assign n20096 = ( n20093 & n20094 ) | ( n20093 & n20095 ) | ( n20094 & n20095 ) ;
  assign n20090 = n6267 ^ n3299 ^ n1474 ;
  assign n20091 = ( n693 & n13428 ) | ( n693 & ~n20090 ) | ( n13428 & ~n20090 ) ;
  assign n20092 = n20091 ^ n16822 ^ 1'b0 ;
  assign n20084 = n12145 ^ n10504 ^ n2910 ;
  assign n20085 = ~n2920 & n11595 ;
  assign n20086 = n6384 & n20085 ;
  assign n20087 = n4828 & n7616 ;
  assign n20088 = n20087 ^ n15654 ^ n3171 ;
  assign n20089 = ( n20084 & n20086 ) | ( n20084 & ~n20088 ) | ( n20086 & ~n20088 ) ;
  assign n20097 = n20096 ^ n20092 ^ n20089 ;
  assign n20098 = ( n9307 & ~n13616 ) | ( n9307 & n18460 ) | ( ~n13616 & n18460 ) ;
  assign n20099 = n20098 ^ n8154 ^ n2494 ;
  assign n20100 = n20099 ^ n13621 ^ n2158 ;
  assign n20101 = ( n8543 & n11663 ) | ( n8543 & n13798 ) | ( n11663 & n13798 ) ;
  assign n20102 = ( n11557 & n15591 ) | ( n11557 & ~n20101 ) | ( n15591 & ~n20101 ) ;
  assign n20103 = n20102 ^ n14871 ^ n5757 ;
  assign n20105 = n7999 & n14806 ;
  assign n20104 = n1988 | n6211 ;
  assign n20106 = n20105 ^ n20104 ^ n12536 ;
  assign n20107 = ( n7111 & n9443 ) | ( n7111 & n11867 ) | ( n9443 & n11867 ) ;
  assign n20108 = n14568 ^ n8586 ^ 1'b0 ;
  assign n20109 = n19743 & n20108 ;
  assign n20110 = n7399 | n7861 ;
  assign n20113 = ( n6400 & ~n7268 ) | ( n6400 & n18681 ) | ( ~n7268 & n18681 ) ;
  assign n20111 = n7645 & ~n17710 ;
  assign n20112 = n5579 & n20111 ;
  assign n20114 = n20113 ^ n20112 ^ n13803 ;
  assign n20115 = n6915 | n9227 ;
  assign n20116 = ( n728 & n18015 ) | ( n728 & n20115 ) | ( n18015 & n20115 ) ;
  assign n20117 = n3774 & ~n11752 ;
  assign n20118 = n20117 ^ n16369 ^ 1'b0 ;
  assign n20119 = ( n4603 & ~n14202 ) | ( n4603 & n20118 ) | ( ~n14202 & n20118 ) ;
  assign n20120 = n496 & n2343 ;
  assign n20121 = ~n13695 & n20120 ;
  assign n20122 = ( n6338 & n16767 ) | ( n6338 & n18178 ) | ( n16767 & n18178 ) ;
  assign n20123 = ~n9722 & n16306 ;
  assign n20124 = n20122 & n20123 ;
  assign n20125 = ( n18749 & ~n20121 ) | ( n18749 & n20124 ) | ( ~n20121 & n20124 ) ;
  assign n20126 = n18381 ^ n2242 ^ n1657 ;
  assign n20127 = ( n2330 & n5905 ) | ( n2330 & n20126 ) | ( n5905 & n20126 ) ;
  assign n20128 = ~n7633 & n12872 ;
  assign n20129 = n20127 & n20128 ;
  assign n20130 = ~n830 & n7410 ;
  assign n20131 = n20130 ^ n2589 ^ 1'b0 ;
  assign n20132 = n15726 ^ n2471 ^ 1'b0 ;
  assign n20133 = n15201 | n20132 ;
  assign n20134 = n18387 ^ n15902 ^ 1'b0 ;
  assign n20135 = n10343 ^ n5871 ^ n2737 ;
  assign n20136 = ( n6691 & n8261 ) | ( n6691 & n20135 ) | ( n8261 & n20135 ) ;
  assign n20137 = ( n10106 & n19485 ) | ( n10106 & ~n20136 ) | ( n19485 & ~n20136 ) ;
  assign n20138 = n15257 ^ n6966 ^ n6724 ;
  assign n20139 = n18670 ^ n12125 ^ n7942 ;
  assign n20140 = n547 & ~n2083 ;
  assign n20141 = ( ~n5963 & n11891 ) | ( ~n5963 & n18759 ) | ( n11891 & n18759 ) ;
  assign n20142 = ( n5493 & n5749 ) | ( n5493 & n6681 ) | ( n5749 & n6681 ) ;
  assign n20143 = ( n3759 & n17141 ) | ( n3759 & n20142 ) | ( n17141 & n20142 ) ;
  assign n20144 = ( n1444 & n8398 ) | ( n1444 & n20143 ) | ( n8398 & n20143 ) ;
  assign n20145 = ( n20140 & ~n20141 ) | ( n20140 & n20144 ) | ( ~n20141 & n20144 ) ;
  assign n20146 = n15774 ^ n12858 ^ 1'b0 ;
  assign n20147 = n577 ^ n354 ^ 1'b0 ;
  assign n20148 = n1225 & ~n20147 ;
  assign n20149 = n20148 ^ n7766 ^ n3166 ;
  assign n20150 = n17574 ^ n3423 ^ 1'b0 ;
  assign n20151 = n20150 ^ n12364 ^ n2380 ;
  assign n20152 = ( n4530 & n8839 ) | ( n4530 & ~n11094 ) | ( n8839 & ~n11094 ) ;
  assign n20153 = n14839 ^ n6089 ^ n5440 ;
  assign n20154 = n14702 ^ n13678 ^ n6356 ;
  assign n20155 = n280 & ~n4292 ;
  assign n20156 = n20155 ^ n16168 ^ 1'b0 ;
  assign n20157 = n5544 ^ n263 ^ 1'b0 ;
  assign n20158 = n20157 ^ n15160 ^ n4043 ;
  assign n20160 = ( ~n1604 & n5490 ) | ( ~n1604 & n7794 ) | ( n5490 & n7794 ) ;
  assign n20159 = ( n4728 & n8569 ) | ( n4728 & n19318 ) | ( n8569 & n19318 ) ;
  assign n20161 = n20160 ^ n20159 ^ n7850 ;
  assign n20162 = ~n12442 & n18196 ;
  assign n20163 = n8127 & n20162 ;
  assign n20164 = ~n5872 & n20163 ;
  assign n20165 = n10008 ^ n9545 ^ 1'b0 ;
  assign n20166 = ~n5436 & n20165 ;
  assign n20167 = n20166 ^ n6875 ^ n1356 ;
  assign n20168 = ( n7471 & n14348 ) | ( n7471 & ~n20167 ) | ( n14348 & ~n20167 ) ;
  assign n20171 = n2458 & n3425 ;
  assign n20169 = n9181 ^ n5318 ^ n2062 ;
  assign n20170 = ( n8517 & n18024 ) | ( n8517 & n20169 ) | ( n18024 & n20169 ) ;
  assign n20172 = n20171 ^ n20170 ^ n11568 ;
  assign n20173 = n3800 ^ n3518 ^ x73 ;
  assign n20179 = n7984 ^ n5027 ^ 1'b0 ;
  assign n20174 = n3210 & n5446 ;
  assign n20175 = n4752 & ~n20174 ;
  assign n20176 = n875 & n20175 ;
  assign n20177 = n12101 | n20176 ;
  assign n20178 = n12650 & n20177 ;
  assign n20180 = n20179 ^ n20178 ^ 1'b0 ;
  assign n20181 = ( n7597 & n20173 ) | ( n7597 & n20180 ) | ( n20173 & n20180 ) ;
  assign n20182 = n9412 ^ n2905 ^ n773 ;
  assign n20183 = ( n5050 & n14088 ) | ( n5050 & n14366 ) | ( n14088 & n14366 ) ;
  assign n20184 = n17708 ^ n4032 ^ n1674 ;
  assign n20185 = n20184 ^ n19204 ^ n2982 ;
  assign n20186 = ( n5293 & ~n14992 ) | ( n5293 & n15417 ) | ( ~n14992 & n15417 ) ;
  assign n20187 = n20186 ^ n7187 ^ x97 ;
  assign n20188 = ( n7531 & n9443 ) | ( n7531 & n15078 ) | ( n9443 & n15078 ) ;
  assign n20189 = n20188 ^ n6727 ^ n4809 ;
  assign n20190 = ( ~n963 & n20187 ) | ( ~n963 & n20189 ) | ( n20187 & n20189 ) ;
  assign n20192 = ( n987 & n3067 ) | ( n987 & n11949 ) | ( n3067 & n11949 ) ;
  assign n20191 = n4473 | n18928 ;
  assign n20193 = n20192 ^ n20191 ^ 1'b0 ;
  assign n20195 = ~n413 & n1639 ;
  assign n20196 = ~n17263 & n20195 ;
  assign n20194 = ( ~n680 & n4556 ) | ( ~n680 & n5559 ) | ( n4556 & n5559 ) ;
  assign n20197 = n20196 ^ n20194 ^ n14682 ;
  assign n20198 = n8425 | n20197 ;
  assign n20199 = n15746 & ~n20198 ;
  assign n20202 = ( n1344 & n2603 ) | ( n1344 & n4059 ) | ( n2603 & n4059 ) ;
  assign n20200 = n15132 ^ n14608 ^ n584 ;
  assign n20201 = ( n3546 & n13243 ) | ( n3546 & ~n20200 ) | ( n13243 & ~n20200 ) ;
  assign n20203 = n20202 ^ n20201 ^ n8658 ;
  assign n20204 = n730 & ~n9826 ;
  assign n20205 = n20204 ^ n2985 ^ n166 ;
  assign n20206 = ( n181 & ~n9352 ) | ( n181 & n20205 ) | ( ~n9352 & n20205 ) ;
  assign n20207 = ( n2355 & n3594 ) | ( n2355 & ~n9814 ) | ( n3594 & ~n9814 ) ;
  assign n20208 = n20207 ^ n19903 ^ n10897 ;
  assign n20209 = ( n1667 & n3882 ) | ( n1667 & n11909 ) | ( n3882 & n11909 ) ;
  assign n20210 = n15739 | n20209 ;
  assign n20211 = n3136 & ~n20210 ;
  assign n20212 = n19471 ^ n953 ^ 1'b0 ;
  assign n20213 = ~n20211 & n20212 ;
  assign n20214 = n11925 ^ n10606 ^ n2272 ;
  assign n20215 = ( n935 & ~n6467 ) | ( n935 & n20214 ) | ( ~n6467 & n20214 ) ;
  assign n20216 = n20215 ^ n17245 ^ 1'b0 ;
  assign n20217 = n4286 | n20216 ;
  assign n20218 = n20217 ^ n18914 ^ n1216 ;
  assign n20220 = n1973 | n5410 ;
  assign n20219 = n20024 ^ n7103 ^ x68 ;
  assign n20221 = n20220 ^ n20219 ^ n7020 ;
  assign n20222 = ( n1470 & ~n8478 ) | ( n1470 & n20221 ) | ( ~n8478 & n20221 ) ;
  assign n20223 = ( ~n7462 & n10463 ) | ( ~n7462 & n17086 ) | ( n10463 & n17086 ) ;
  assign n20227 = ( n3741 & ~n12508 ) | ( n3741 & n14303 ) | ( ~n12508 & n14303 ) ;
  assign n20224 = ( ~n3061 & n3648 ) | ( ~n3061 & n5113 ) | ( n3648 & n5113 ) ;
  assign n20225 = n20224 ^ n9219 ^ n1448 ;
  assign n20226 = ( n6676 & n19727 ) | ( n6676 & n20225 ) | ( n19727 & n20225 ) ;
  assign n20228 = n20227 ^ n20226 ^ 1'b0 ;
  assign n20229 = ~n8958 & n20228 ;
  assign n20230 = ( ~n993 & n13657 ) | ( ~n993 & n15993 ) | ( n13657 & n15993 ) ;
  assign n20231 = n12367 ^ n3322 ^ n2201 ;
  assign n20232 = ( n7973 & ~n12337 ) | ( n7973 & n20231 ) | ( ~n12337 & n20231 ) ;
  assign n20233 = n17740 ^ n15804 ^ n5265 ;
  assign n20234 = n20233 ^ n7078 ^ n2703 ;
  assign n20235 = n20234 ^ n257 ^ 1'b0 ;
  assign n20237 = ( ~n2411 & n7003 ) | ( ~n2411 & n9667 ) | ( n7003 & n9667 ) ;
  assign n20238 = n20237 ^ n18005 ^ 1'b0 ;
  assign n20236 = n5051 & ~n10779 ;
  assign n20239 = n20238 ^ n20236 ^ 1'b0 ;
  assign n20240 = n20239 ^ n11112 ^ n4564 ;
  assign n20241 = n12968 ^ n1456 ^ 1'b0 ;
  assign n20242 = ~n15969 & n20241 ;
  assign n20243 = n5557 & n7383 ;
  assign n20244 = n6586 & n20243 ;
  assign n20245 = n1092 & n20244 ;
  assign n20246 = n1114 | n14076 ;
  assign n20247 = n20245 | n20246 ;
  assign n20248 = n16701 | n19050 ;
  assign n20249 = n4465 & ~n20248 ;
  assign n20250 = ( n514 & n1493 ) | ( n514 & ~n3276 ) | ( n1493 & ~n3276 ) ;
  assign n20251 = ( ~x108 & n3990 ) | ( ~x108 & n8639 ) | ( n3990 & n8639 ) ;
  assign n20252 = n20251 ^ n4640 ^ 1'b0 ;
  assign n20253 = n11995 & n20252 ;
  assign n20254 = ( n5271 & n20250 ) | ( n5271 & ~n20253 ) | ( n20250 & ~n20253 ) ;
  assign n20255 = n4830 ^ n2849 ^ n1725 ;
  assign n20256 = n20255 ^ n19731 ^ n17195 ;
  assign n20257 = n11904 ^ n2856 ^ n1778 ;
  assign n20258 = n20257 ^ n7075 ^ n5304 ;
  assign n20259 = n20258 ^ n2377 ^ n747 ;
  assign n20263 = n4896 ^ n4187 ^ 1'b0 ;
  assign n20264 = n14532 & n20263 ;
  assign n20265 = ( ~x127 & n10328 ) | ( ~x127 & n20264 ) | ( n10328 & n20264 ) ;
  assign n20266 = ( n9302 & ~n12407 ) | ( n9302 & n20265 ) | ( ~n12407 & n20265 ) ;
  assign n20267 = ( ~n8508 & n11771 ) | ( ~n8508 & n12997 ) | ( n11771 & n12997 ) ;
  assign n20268 = n12284 | n20267 ;
  assign n20269 = n20266 & n20268 ;
  assign n20270 = n20269 ^ n14483 ^ 1'b0 ;
  assign n20260 = n19800 ^ n17792 ^ n1077 ;
  assign n20261 = n20260 ^ n9960 ^ n5029 ;
  assign n20262 = n20261 ^ n9754 ^ n2647 ;
  assign n20271 = n20270 ^ n20262 ^ n15769 ;
  assign n20272 = n10543 ^ n9974 ^ n4157 ;
  assign n20273 = ( n4968 & n5700 ) | ( n4968 & ~n8406 ) | ( n5700 & ~n8406 ) ;
  assign n20274 = n20273 ^ n5772 ^ 1'b0 ;
  assign n20275 = n20272 & ~n20274 ;
  assign n20276 = ( ~n10082 & n12583 ) | ( ~n10082 & n20275 ) | ( n12583 & n20275 ) ;
  assign n20277 = n19018 ^ n7031 ^ n135 ;
  assign n20278 = n2900 | n6310 ;
  assign n20279 = n20278 ^ n3767 ^ 1'b0 ;
  assign n20280 = ( n218 & n6707 ) | ( n218 & ~n20279 ) | ( n6707 & ~n20279 ) ;
  assign n20281 = ( n10936 & n19099 ) | ( n10936 & n20280 ) | ( n19099 & n20280 ) ;
  assign n20282 = n3865 & n6630 ;
  assign n20283 = n20282 ^ n7077 ^ 1'b0 ;
  assign n20284 = n20283 ^ n5145 ^ n698 ;
  assign n20285 = n9989 & ~n12993 ;
  assign n20286 = n20284 & n20285 ;
  assign n20287 = ( n4796 & n15058 ) | ( n4796 & n17938 ) | ( n15058 & n17938 ) ;
  assign n20288 = n20287 ^ n13924 ^ n7817 ;
  assign n20289 = n7511 | n16035 ;
  assign n20290 = ( n4382 & ~n16058 ) | ( n4382 & n18034 ) | ( ~n16058 & n18034 ) ;
  assign n20292 = n13365 ^ n9445 ^ n2294 ;
  assign n20293 = n20292 ^ n4767 ^ 1'b0 ;
  assign n20294 = n16897 & n20293 ;
  assign n20291 = n15090 ^ n4786 ^ n4505 ;
  assign n20295 = n20294 ^ n20291 ^ n12814 ;
  assign n20296 = n20295 ^ n6209 ^ n4529 ;
  assign n20297 = ( n1077 & ~n3657 ) | ( n1077 & n4437 ) | ( ~n3657 & n4437 ) ;
  assign n20298 = ( n2712 & n8214 ) | ( n2712 & ~n20297 ) | ( n8214 & ~n20297 ) ;
  assign n20299 = x127 & n2386 ;
  assign n20300 = ~n2903 & n20299 ;
  assign n20301 = n15968 | n20300 ;
  assign n20302 = n13376 & ~n20301 ;
  assign n20303 = n20302 ^ n13521 ^ n612 ;
  assign n20304 = n15804 ^ n14363 ^ n6091 ;
  assign n20305 = ( n7282 & n10795 ) | ( n7282 & ~n20304 ) | ( n10795 & ~n20304 ) ;
  assign n20306 = ( n256 & ~n4055 ) | ( n256 & n14483 ) | ( ~n4055 & n14483 ) ;
  assign n20307 = ( n4299 & ~n18558 ) | ( n4299 & n20306 ) | ( ~n18558 & n20306 ) ;
  assign n20308 = ( ~n4174 & n16129 ) | ( ~n4174 & n20307 ) | ( n16129 & n20307 ) ;
  assign n20309 = n20308 ^ n13960 ^ 1'b0 ;
  assign n20310 = n9195 ^ n9114 ^ n7206 ;
  assign n20311 = ( n1977 & n5424 ) | ( n1977 & ~n8344 ) | ( n5424 & ~n8344 ) ;
  assign n20312 = n20311 ^ n13612 ^ n2560 ;
  assign n20313 = ( ~n1200 & n6403 ) | ( ~n1200 & n14487 ) | ( n6403 & n14487 ) ;
  assign n20314 = n16820 & ~n20313 ;
  assign n20315 = ( n5319 & ~n20312 ) | ( n5319 & n20314 ) | ( ~n20312 & n20314 ) ;
  assign n20316 = n9768 ^ n6757 ^ n2123 ;
  assign n20317 = ( n1014 & n14881 ) | ( n1014 & ~n17096 ) | ( n14881 & ~n17096 ) ;
  assign n20318 = n17285 ^ n12151 ^ n2215 ;
  assign n20319 = ~n10822 & n14528 ;
  assign n20320 = n20319 ^ n9579 ^ 1'b0 ;
  assign n20322 = n9865 ^ n2804 ^ n1567 ;
  assign n20321 = ~n16778 & n17637 ;
  assign n20323 = n20322 ^ n20321 ^ 1'b0 ;
  assign n20324 = n19524 ^ n3222 ^ 1'b0 ;
  assign n20327 = n10458 ^ n1051 ^ 1'b0 ;
  assign n20328 = n5047 & ~n20327 ;
  assign n20325 = n14453 ^ n327 ^ 1'b0 ;
  assign n20326 = ~n7173 & n20325 ;
  assign n20329 = n20328 ^ n20326 ^ n18048 ;
  assign n20330 = ( n5682 & ~n8894 ) | ( n5682 & n9061 ) | ( ~n8894 & n9061 ) ;
  assign n20331 = n13997 & ~n20330 ;
  assign n20332 = n10772 & ~n19408 ;
  assign n20333 = n1545 | n11281 ;
  assign n20334 = n20333 ^ n10392 ^ 1'b0 ;
  assign n20335 = ( n581 & ~n1942 ) | ( n581 & n3087 ) | ( ~n1942 & n3087 ) ;
  assign n20336 = n5608 | n20335 ;
  assign n20337 = ( x62 & n10155 ) | ( x62 & n20336 ) | ( n10155 & n20336 ) ;
  assign n20338 = n16434 | n18937 ;
  assign n20339 = n20338 ^ n15478 ^ n14524 ;
  assign n20340 = n4329 & ~n11905 ;
  assign n20341 = n20340 ^ n14996 ^ 1'b0 ;
  assign n20342 = n16780 | n20341 ;
  assign n20344 = n4441 & n16408 ;
  assign n20345 = n20344 ^ n10614 ^ 1'b0 ;
  assign n20343 = n863 & ~n12112 ;
  assign n20346 = n20345 ^ n20343 ^ 1'b0 ;
  assign n20347 = n20346 ^ n17869 ^ n4444 ;
  assign n20348 = ( ~n750 & n9582 ) | ( ~n750 & n12320 ) | ( n9582 & n12320 ) ;
  assign n20349 = n16094 & n20348 ;
  assign n20350 = n15797 ^ n9322 ^ 1'b0 ;
  assign n20351 = n10733 ^ n7824 ^ n2429 ;
  assign n20352 = n20351 ^ n2771 ^ x99 ;
  assign n20353 = ( ~n9254 & n20350 ) | ( ~n9254 & n20352 ) | ( n20350 & n20352 ) ;
  assign n20354 = ( n14211 & n17249 ) | ( n14211 & n20353 ) | ( n17249 & n20353 ) ;
  assign n20355 = ( ~n5880 & n8577 ) | ( ~n5880 & n8864 ) | ( n8577 & n8864 ) ;
  assign n20356 = n5286 ^ n1385 ^ n519 ;
  assign n20357 = ~n19306 & n20356 ;
  assign n20358 = n9281 ^ n7385 ^ 1'b0 ;
  assign n20359 = ( n7047 & n7102 ) | ( n7047 & n19727 ) | ( n7102 & n19727 ) ;
  assign n20360 = ( n19846 & n20358 ) | ( n19846 & ~n20359 ) | ( n20358 & ~n20359 ) ;
  assign n20361 = n11883 ^ n4066 ^ 1'b0 ;
  assign n20362 = n934 & n20361 ;
  assign n20363 = n10181 ^ n6894 ^ 1'b0 ;
  assign n20364 = ( n6514 & n10622 ) | ( n6514 & ~n20363 ) | ( n10622 & ~n20363 ) ;
  assign n20366 = ( n2615 & n6551 ) | ( n2615 & n7791 ) | ( n6551 & n7791 ) ;
  assign n20365 = ~n10234 & n15931 ;
  assign n20367 = n20366 ^ n20365 ^ 1'b0 ;
  assign n20368 = n7134 ^ n6616 ^ n875 ;
  assign n20369 = ( n6934 & n15741 ) | ( n6934 & ~n20368 ) | ( n15741 & ~n20368 ) ;
  assign n20370 = ( n434 & ~n12521 ) | ( n434 & n15065 ) | ( ~n12521 & n15065 ) ;
  assign n20373 = n13383 ^ n1958 ^ n879 ;
  assign n20371 = n13347 ^ n5774 ^ n4452 ;
  assign n20372 = ( ~n444 & n10012 ) | ( ~n444 & n20371 ) | ( n10012 & n20371 ) ;
  assign n20374 = n20373 ^ n20372 ^ 1'b0 ;
  assign n20375 = n2706 & ~n4433 ;
  assign n20376 = n20375 ^ n4224 ^ n2862 ;
  assign n20377 = n20376 ^ n14041 ^ n4069 ;
  assign n20378 = n18944 ^ n18722 ^ n3604 ;
  assign n20379 = n20016 ^ n7935 ^ n2536 ;
  assign n20380 = ( n6253 & ~n12417 ) | ( n6253 & n20379 ) | ( ~n12417 & n20379 ) ;
  assign n20381 = n20380 ^ n17467 ^ n8423 ;
  assign n20382 = n20381 ^ n18999 ^ n14625 ;
  assign n20383 = n2845 ^ n2437 ^ 1'b0 ;
  assign n20384 = n4889 | n20383 ;
  assign n20385 = n17740 ^ n3315 ^ n2501 ;
  assign n20386 = n20385 ^ n17352 ^ n1182 ;
  assign n20387 = n20386 ^ n10508 ^ 1'b0 ;
  assign n20388 = ~n20384 & n20387 ;
  assign n20389 = ( n5720 & n9271 ) | ( n5720 & n15191 ) | ( n9271 & n15191 ) ;
  assign n20390 = n20389 ^ n8785 ^ n1398 ;
  assign n20391 = n15742 ^ n13713 ^ n9179 ;
  assign n20392 = n6156 & n6708 ;
  assign n20393 = ~n13136 & n20392 ;
  assign n20394 = ( n4754 & ~n7820 ) | ( n4754 & n20393 ) | ( ~n7820 & n20393 ) ;
  assign n20395 = ( n1440 & n14750 ) | ( n1440 & ~n20394 ) | ( n14750 & ~n20394 ) ;
  assign n20396 = ( ~n7124 & n15667 ) | ( ~n7124 & n18056 ) | ( n15667 & n18056 ) ;
  assign n20397 = n20396 ^ n6512 ^ n1517 ;
  assign n20398 = ( n4549 & n16459 ) | ( n4549 & n19980 ) | ( n16459 & n19980 ) ;
  assign n20399 = n17853 ^ n12883 ^ n5506 ;
  assign n20400 = n6052 & ~n11178 ;
  assign n20401 = n20400 ^ n8709 ^ 1'b0 ;
  assign n20402 = n20401 ^ n12105 ^ n8061 ;
  assign n20403 = n20402 ^ n17574 ^ n13465 ;
  assign n20404 = ( n4124 & n8457 ) | ( n4124 & n8676 ) | ( n8457 & n8676 ) ;
  assign n20406 = ( n1120 & n1374 ) | ( n1120 & ~n6480 ) | ( n1374 & ~n6480 ) ;
  assign n20405 = n6894 & n8854 ;
  assign n20407 = n20406 ^ n20405 ^ 1'b0 ;
  assign n20408 = n3697 ^ n3140 ^ n2806 ;
  assign n20409 = ( ~n7643 & n9801 ) | ( ~n7643 & n20408 ) | ( n9801 & n20408 ) ;
  assign n20410 = ( n1026 & n11376 ) | ( n1026 & ~n20409 ) | ( n11376 & ~n20409 ) ;
  assign n20411 = n11084 ^ n10283 ^ n8406 ;
  assign n20412 = n20411 ^ n20258 ^ n7894 ;
  assign n20413 = ( n5967 & ~n16213 ) | ( n5967 & n19731 ) | ( ~n16213 & n19731 ) ;
  assign n20418 = ( n898 & n4795 ) | ( n898 & n12382 ) | ( n4795 & n12382 ) ;
  assign n20414 = n15109 ^ n7478 ^ n2687 ;
  assign n20415 = n20414 ^ n14504 ^ n5826 ;
  assign n20416 = n20415 ^ n16912 ^ n10464 ;
  assign n20417 = ~n2429 & n20416 ;
  assign n20419 = n20418 ^ n20417 ^ n5610 ;
  assign n20420 = n20419 ^ n3228 ^ 1'b0 ;
  assign n20421 = ( ~n5556 & n18269 ) | ( ~n5556 & n20420 ) | ( n18269 & n20420 ) ;
  assign n20423 = ( n2716 & n3689 ) | ( n2716 & ~n12934 ) | ( n3689 & ~n12934 ) ;
  assign n20422 = ( n1465 & ~n6459 ) | ( n1465 & n8858 ) | ( ~n6459 & n8858 ) ;
  assign n20424 = n20423 ^ n20422 ^ n15647 ;
  assign n20425 = n20424 ^ n18878 ^ n13309 ;
  assign n20426 = n20425 ^ n3967 ^ x66 ;
  assign n20427 = n15301 ^ n13253 ^ n1723 ;
  assign n20428 = n17362 ^ n6420 ^ n1684 ;
  assign n20429 = n19045 & n20428 ;
  assign n20430 = n5538 ^ n4384 ^ 1'b0 ;
  assign n20431 = n3256 & ~n20430 ;
  assign n20432 = ( ~n596 & n4941 ) | ( ~n596 & n13532 ) | ( n4941 & n13532 ) ;
  assign n20433 = n10449 & ~n11802 ;
  assign n20434 = ( n6681 & n13453 ) | ( n6681 & ~n20433 ) | ( n13453 & ~n20433 ) ;
  assign n20435 = n20432 & ~n20434 ;
  assign n20436 = n20435 ^ n12036 ^ n3514 ;
  assign n20437 = n13750 ^ n4392 ^ n1760 ;
  assign n20438 = ( n5125 & n5794 ) | ( n5125 & ~n7931 ) | ( n5794 & ~n7931 ) ;
  assign n20439 = n20437 & ~n20438 ;
  assign n20440 = ( n9669 & n12659 ) | ( n9669 & ~n17812 ) | ( n12659 & ~n17812 ) ;
  assign n20441 = ~n18368 & n20440 ;
  assign n20444 = n13946 ^ n6065 ^ 1'b0 ;
  assign n20445 = n18390 | n20444 ;
  assign n20442 = ~n2664 & n7303 ;
  assign n20443 = ( ~n4976 & n5899 ) | ( ~n4976 & n20442 ) | ( n5899 & n20442 ) ;
  assign n20446 = n20445 ^ n20443 ^ n3286 ;
  assign n20447 = n20446 ^ n1015 ^ 1'b0 ;
  assign n20448 = n17233 ^ n8641 ^ n871 ;
  assign n20449 = n11670 ^ n9462 ^ n242 ;
  assign n20450 = n20449 ^ n19545 ^ n15888 ;
  assign n20451 = ( n1561 & n4510 ) | ( n1561 & ~n11182 ) | ( n4510 & ~n11182 ) ;
  assign n20452 = n16956 ^ n5730 ^ n2836 ;
  assign n20453 = n20451 | n20452 ;
  assign n20454 = n19073 ^ n14572 ^ n1430 ;
  assign n20455 = n2476 & ~n2756 ;
  assign n20456 = n12447 & n20455 ;
  assign n20457 = n20456 ^ n9881 ^ n4184 ;
  assign n20458 = n12852 ^ n6421 ^ n3267 ;
  assign n20462 = ( ~n1174 & n8470 ) | ( ~n1174 & n11055 ) | ( n8470 & n11055 ) ;
  assign n20461 = n7113 & ~n7685 ;
  assign n20459 = ( x110 & n1180 ) | ( x110 & n14668 ) | ( n1180 & n14668 ) ;
  assign n20460 = n20459 ^ n11281 ^ n7754 ;
  assign n20463 = n20462 ^ n20461 ^ n20460 ;
  assign n20464 = x119 & ~n7973 ;
  assign n20465 = n6658 & n19947 ;
  assign n20466 = ~n2329 & n3878 ;
  assign n20467 = ( n2511 & ~n3478 ) | ( n2511 & n4487 ) | ( ~n3478 & n4487 ) ;
  assign n20468 = n5390 & ~n20467 ;
  assign n20469 = ( n7287 & n15264 ) | ( n7287 & ~n20468 ) | ( n15264 & ~n20468 ) ;
  assign n20470 = n20469 ^ n4058 ^ 1'b0 ;
  assign n20471 = n20466 & ~n20470 ;
  assign n20472 = ( n2481 & n7071 ) | ( n2481 & ~n12308 ) | ( n7071 & ~n12308 ) ;
  assign n20473 = ( n2530 & n2674 ) | ( n2530 & ~n4346 ) | ( n2674 & ~n4346 ) ;
  assign n20474 = ( n1631 & n6654 ) | ( n1631 & ~n20473 ) | ( n6654 & ~n20473 ) ;
  assign n20475 = ( ~n8149 & n17105 ) | ( ~n8149 & n17234 ) | ( n17105 & n17234 ) ;
  assign n20476 = ( ~n3605 & n10834 ) | ( ~n3605 & n20475 ) | ( n10834 & n20475 ) ;
  assign n20477 = ~n7737 & n19574 ;
  assign n20478 = n7733 | n20477 ;
  assign n20479 = n18229 & ~n20478 ;
  assign n20480 = n17257 ^ n17010 ^ n3020 ;
  assign n20481 = ( ~x39 & n4012 ) | ( ~x39 & n12722 ) | ( n4012 & n12722 ) ;
  assign n20482 = ( n5121 & ~n15683 ) | ( n5121 & n20481 ) | ( ~n15683 & n20481 ) ;
  assign n20483 = n18229 ^ n15295 ^ n13101 ;
  assign n20485 = ( n2683 & ~n5398 ) | ( n2683 & n18849 ) | ( ~n5398 & n18849 ) ;
  assign n20484 = ( ~n4124 & n6357 ) | ( ~n4124 & n14353 ) | ( n6357 & n14353 ) ;
  assign n20486 = n20485 ^ n20484 ^ n19424 ;
  assign n20487 = ( ~n8251 & n19375 ) | ( ~n8251 & n19822 ) | ( n19375 & n19822 ) ;
  assign n20488 = ~n12021 & n14840 ;
  assign n20489 = n15768 & n20488 ;
  assign n20490 = x119 & n1897 ;
  assign n20491 = ( n10225 & ~n10993 ) | ( n10225 & n20490 ) | ( ~n10993 & n20490 ) ;
  assign n20492 = n20491 ^ n2012 ^ 1'b0 ;
  assign n20493 = n16862 ^ n10736 ^ 1'b0 ;
  assign n20494 = n7113 & ~n20493 ;
  assign n20495 = n20494 ^ n3488 ^ 1'b0 ;
  assign n20496 = ( ~n2045 & n2334 ) | ( ~n2045 & n5839 ) | ( n2334 & n5839 ) ;
  assign n20497 = ( n10618 & n13706 ) | ( n10618 & ~n13809 ) | ( n13706 & ~n13809 ) ;
  assign n20498 = ( ~n2344 & n20496 ) | ( ~n2344 & n20497 ) | ( n20496 & n20497 ) ;
  assign n20499 = ~n8878 & n12872 ;
  assign n20500 = n20499 ^ n14249 ^ 1'b0 ;
  assign n20501 = ( ~n8531 & n9575 ) | ( ~n8531 & n20500 ) | ( n9575 & n20500 ) ;
  assign n20502 = n17809 ^ n11393 ^ 1'b0 ;
  assign n20503 = x16 & n20502 ;
  assign n20507 = n5186 ^ n1710 ^ 1'b0 ;
  assign n20508 = ( n5704 & n10511 ) | ( n5704 & n20507 ) | ( n10511 & n20507 ) ;
  assign n20504 = n18311 ^ n12631 ^ n12333 ;
  assign n20505 = n3150 & ~n20504 ;
  assign n20506 = n20505 ^ n16047 ^ 1'b0 ;
  assign n20509 = n20508 ^ n20506 ^ n4828 ;
  assign n20510 = n13205 ^ n6630 ^ n2950 ;
  assign n20511 = ( n8385 & ~n13484 ) | ( n8385 & n20510 ) | ( ~n13484 & n20510 ) ;
  assign n20512 = n20511 ^ n3905 ^ 1'b0 ;
  assign n20513 = ~n20509 & n20512 ;
  assign n20514 = n16787 ^ n7505 ^ 1'b0 ;
  assign n20515 = ~n17306 & n20514 ;
  assign n20516 = ~n813 & n15452 ;
  assign n20517 = n20516 ^ n2877 ^ 1'b0 ;
  assign n20518 = n18596 ^ n16144 ^ n11759 ;
  assign n20519 = ( n2422 & n20517 ) | ( n2422 & n20518 ) | ( n20517 & n20518 ) ;
  assign n20520 = ( n1876 & n4333 ) | ( n1876 & n17496 ) | ( n4333 & n17496 ) ;
  assign n20521 = ( n9311 & n20519 ) | ( n9311 & ~n20520 ) | ( n20519 & ~n20520 ) ;
  assign n20522 = ( ~n2206 & n7974 ) | ( ~n2206 & n19762 ) | ( n7974 & n19762 ) ;
  assign n20523 = ( n282 & n11138 ) | ( n282 & ~n11375 ) | ( n11138 & ~n11375 ) ;
  assign n20524 = ( n10587 & n13787 ) | ( n10587 & ~n20523 ) | ( n13787 & ~n20523 ) ;
  assign n20525 = n20524 ^ n5581 ^ 1'b0 ;
  assign n20526 = n15879 ^ n5666 ^ n5375 ;
  assign n20527 = ~n7042 & n11048 ;
  assign n20528 = n20527 ^ n12958 ^ 1'b0 ;
  assign n20530 = ( n1684 & n10601 ) | ( n1684 & n10648 ) | ( n10601 & n10648 ) ;
  assign n20529 = n809 & ~n7340 ;
  assign n20531 = n20530 ^ n20529 ^ n2857 ;
  assign n20532 = n13003 ^ n11321 ^ n547 ;
  assign n20533 = n20532 ^ n19775 ^ n15837 ;
  assign n20534 = n12366 ^ n4032 ^ 1'b0 ;
  assign n20535 = n2504 | n7633 ;
  assign n20536 = n3016 & n20535 ;
  assign n20537 = ( ~n10755 & n20534 ) | ( ~n10755 & n20536 ) | ( n20534 & n20536 ) ;
  assign n20538 = n19439 ^ n13950 ^ n11937 ;
  assign n20539 = n9649 ^ n344 ^ 1'b0 ;
  assign n20540 = ( n889 & n3671 ) | ( n889 & ~n4830 ) | ( n3671 & ~n4830 ) ;
  assign n20541 = n9502 & ~n18092 ;
  assign n20542 = n20541 ^ n11330 ^ 1'b0 ;
  assign n20543 = ( n20539 & ~n20540 ) | ( n20539 & n20542 ) | ( ~n20540 & n20542 ) ;
  assign n20544 = n12025 ^ n1304 ^ n164 ;
  assign n20545 = ~n4627 & n18679 ;
  assign n20546 = n16172 & n20545 ;
  assign n20548 = n14893 ^ n6577 ^ 1'b0 ;
  assign n20547 = ( n4698 & ~n8479 ) | ( n4698 & n9777 ) | ( ~n8479 & n9777 ) ;
  assign n20549 = n20548 ^ n20547 ^ n3542 ;
  assign n20550 = n20549 ^ n16637 ^ 1'b0 ;
  assign n20551 = n19485 | n20550 ;
  assign n20552 = ( n580 & n4714 ) | ( n580 & n20040 ) | ( n4714 & n20040 ) ;
  assign n20553 = n17158 | n19958 ;
  assign n20554 = n20553 ^ n13980 ^ 1'b0 ;
  assign n20555 = ( n13907 & ~n17316 ) | ( n13907 & n20554 ) | ( ~n17316 & n20554 ) ;
  assign n20556 = n20555 ^ n9372 ^ n4384 ;
  assign n20560 = n3066 | n6466 ;
  assign n20557 = ( ~n6722 & n13613 ) | ( ~n6722 & n19683 ) | ( n13613 & n19683 ) ;
  assign n20558 = n2336 & n9913 ;
  assign n20559 = n20557 & n20558 ;
  assign n20561 = n20560 ^ n20559 ^ n10467 ;
  assign n20562 = n16428 ^ n16074 ^ n5950 ;
  assign n20563 = n20562 ^ n5310 ^ x65 ;
  assign n20565 = n13205 ^ n3034 ^ n1581 ;
  assign n20564 = n11737 ^ n7904 ^ n7817 ;
  assign n20566 = n20565 ^ n20564 ^ n9975 ;
  assign n20567 = n5948 ^ n215 ^ 1'b0 ;
  assign n20568 = n11801 & ~n20567 ;
  assign n20569 = n20568 ^ n6460 ^ 1'b0 ;
  assign n20570 = n16553 | n20569 ;
  assign n20574 = ( n2335 & ~n2802 ) | ( n2335 & n14490 ) | ( ~n2802 & n14490 ) ;
  assign n20571 = n1641 & n9061 ;
  assign n20572 = n20571 ^ n13822 ^ 1'b0 ;
  assign n20573 = n171 & n20572 ;
  assign n20575 = n20574 ^ n20573 ^ 1'b0 ;
  assign n20576 = ( n457 & n6664 ) | ( n457 & ~n7269 ) | ( n6664 & ~n7269 ) ;
  assign n20577 = ( n268 & n3345 ) | ( n268 & ~n20576 ) | ( n3345 & ~n20576 ) ;
  assign n20578 = n3150 & n7429 ;
  assign n20579 = n5056 & n20578 ;
  assign n20580 = ( n1718 & n6415 ) | ( n1718 & n20579 ) | ( n6415 & n20579 ) ;
  assign n20581 = ( n8071 & n19108 ) | ( n8071 & ~n20580 ) | ( n19108 & ~n20580 ) ;
  assign n20582 = ( ~n1990 & n8904 ) | ( ~n1990 & n20581 ) | ( n8904 & n20581 ) ;
  assign n20583 = n1992 ^ n804 ^ 1'b0 ;
  assign n20584 = n2039 | n20583 ;
  assign n20585 = n20584 ^ n2732 ^ n2294 ;
  assign n20586 = ( n1694 & n4408 ) | ( n1694 & n20585 ) | ( n4408 & n20585 ) ;
  assign n20587 = n14143 ^ n9476 ^ n2708 ;
  assign n20588 = n3084 ^ n163 ^ 1'b0 ;
  assign n20589 = ~n209 & n20588 ;
  assign n20590 = ~n14126 & n20589 ;
  assign n20591 = n20590 ^ n13983 ^ 1'b0 ;
  assign n20592 = n9187 ^ n7582 ^ 1'b0 ;
  assign n20593 = n20591 | n20592 ;
  assign n20594 = n15234 & n17200 ;
  assign n20595 = n20593 & n20594 ;
  assign n20596 = ( n3455 & ~n20587 ) | ( n3455 & n20595 ) | ( ~n20587 & n20595 ) ;
  assign n20597 = n2898 ^ n1004 ^ 1'b0 ;
  assign n20598 = ~n11263 & n20597 ;
  assign n20599 = ~n16281 & n20598 ;
  assign n20600 = n20599 ^ n16441 ^ n6113 ;
  assign n20601 = n6818 & n9854 ;
  assign n20602 = n902 & n9994 ;
  assign n20603 = ~n980 & n20602 ;
  assign n20604 = ( n7634 & n7738 ) | ( n7634 & ~n20603 ) | ( n7738 & ~n20603 ) ;
  assign n20605 = ( n7984 & n14651 ) | ( n7984 & ~n16948 ) | ( n14651 & ~n16948 ) ;
  assign n20606 = n3566 | n15792 ;
  assign n20607 = n1806 & ~n20606 ;
  assign n20608 = ( n4783 & ~n20605 ) | ( n4783 & n20607 ) | ( ~n20605 & n20607 ) ;
  assign n20609 = n3378 ^ n2016 ^ 1'b0 ;
  assign n20610 = n20609 ^ n18179 ^ n4604 ;
  assign n20611 = n16507 ^ n13355 ^ n11785 ;
  assign n20612 = n3777 & n12936 ;
  assign n20613 = ~n12942 & n20612 ;
  assign n20614 = n7571 ^ n6956 ^ n5901 ;
  assign n20615 = n2328 | n10939 ;
  assign n20616 = ( n19064 & ~n20614 ) | ( n19064 & n20615 ) | ( ~n20614 & n20615 ) ;
  assign n20617 = n17353 ^ n10723 ^ 1'b0 ;
  assign n20618 = ~n20616 & n20617 ;
  assign n20619 = ( n11257 & n13028 ) | ( n11257 & n14464 ) | ( n13028 & n14464 ) ;
  assign n20620 = ( n2232 & n2893 ) | ( n2232 & ~n4900 ) | ( n2893 & ~n4900 ) ;
  assign n20621 = n20620 ^ n14178 ^ 1'b0 ;
  assign n20622 = n11341 & ~n20621 ;
  assign n20623 = ( n1421 & ~n20619 ) | ( n1421 & n20622 ) | ( ~n20619 & n20622 ) ;
  assign n20624 = ~n8344 & n17941 ;
  assign n20625 = ( n623 & ~n9510 ) | ( n623 & n9622 ) | ( ~n9510 & n9622 ) ;
  assign n20626 = ( n1495 & ~n13721 ) | ( n1495 & n20625 ) | ( ~n13721 & n20625 ) ;
  assign n20627 = ( n7468 & n20624 ) | ( n7468 & ~n20626 ) | ( n20624 & ~n20626 ) ;
  assign n20628 = ( n12835 & n18121 ) | ( n12835 & n20627 ) | ( n18121 & n20627 ) ;
  assign n20629 = ( ~n1629 & n7903 ) | ( ~n1629 & n15690 ) | ( n7903 & n15690 ) ;
  assign n20630 = ( ~n9614 & n12087 ) | ( ~n9614 & n13809 ) | ( n12087 & n13809 ) ;
  assign n20631 = ( ~n11807 & n12429 ) | ( ~n11807 & n20630 ) | ( n12429 & n20630 ) ;
  assign n20632 = n11087 ^ n8641 ^ n8341 ;
  assign n20633 = n20632 ^ n9367 ^ n9235 ;
  assign n20634 = n20631 & ~n20633 ;
  assign n20635 = ~n1999 & n11486 ;
  assign n20636 = n9051 & n20635 ;
  assign n20637 = n14974 & ~n20636 ;
  assign n20638 = n2696 & n20637 ;
  assign n20639 = ( n3075 & ~n4368 ) | ( n3075 & n20638 ) | ( ~n4368 & n20638 ) ;
  assign n20640 = n17326 ^ n13106 ^ n9167 ;
  assign n20641 = ( n5036 & n8407 ) | ( n5036 & ~n14307 ) | ( n8407 & ~n14307 ) ;
  assign n20642 = n20641 ^ n2045 ^ n829 ;
  assign n20643 = n2068 & n14034 ;
  assign n20644 = ( n15638 & ~n15921 ) | ( n15638 & n20643 ) | ( ~n15921 & n20643 ) ;
  assign n20645 = ( n8144 & n13854 ) | ( n8144 & ~n20644 ) | ( n13854 & ~n20644 ) ;
  assign n20646 = ( x111 & ~n2225 ) | ( x111 & n3968 ) | ( ~n2225 & n3968 ) ;
  assign n20647 = n20646 ^ n11312 ^ n5192 ;
  assign n20648 = n20647 ^ n5815 ^ n3322 ;
  assign n20649 = ( n1170 & ~n4221 ) | ( n1170 & n20648 ) | ( ~n4221 & n20648 ) ;
  assign n20650 = n16287 ^ n13307 ^ n7660 ;
  assign n20651 = n1466 | n13616 ;
  assign n20652 = x127 | n20651 ;
  assign n20653 = n20652 ^ n15225 ^ n3262 ;
  assign n20657 = n14820 ^ n2982 ^ n2107 ;
  assign n20654 = n5006 ^ n4207 ^ 1'b0 ;
  assign n20655 = n9646 & ~n20654 ;
  assign n20656 = n20655 ^ n7183 ^ 1'b0 ;
  assign n20658 = n20657 ^ n20656 ^ n5171 ;
  assign n20659 = ( n1445 & n2854 ) | ( n1445 & n9988 ) | ( n2854 & n9988 ) ;
  assign n20660 = ( n10202 & ~n14332 ) | ( n10202 & n20659 ) | ( ~n14332 & n20659 ) ;
  assign n20661 = n12324 & ~n12504 ;
  assign n20662 = n5568 ^ n3564 ^ x56 ;
  assign n20663 = ~n2049 & n20662 ;
  assign n20664 = n2402 & ~n10688 ;
  assign n20665 = n3109 ^ n395 ^ 1'b0 ;
  assign n20666 = ( n8061 & ~n15266 ) | ( n8061 & n20665 ) | ( ~n15266 & n20665 ) ;
  assign n20667 = n20666 ^ n539 ^ 1'b0 ;
  assign n20668 = n20667 ^ n7718 ^ n7549 ;
  assign n20669 = ( n5648 & n10355 ) | ( n5648 & ~n10685 ) | ( n10355 & ~n10685 ) ;
  assign n20670 = n20669 ^ n8589 ^ n2050 ;
  assign n20671 = ( n624 & n4043 ) | ( n624 & n7325 ) | ( n4043 & n7325 ) ;
  assign n20672 = n11895 ^ n10758 ^ n3977 ;
  assign n20673 = n7925 | n19947 ;
  assign n20674 = n20673 ^ n3213 ^ 1'b0 ;
  assign n20675 = ( n15832 & n20672 ) | ( n15832 & n20674 ) | ( n20672 & n20674 ) ;
  assign n20676 = ( n1352 & n4235 ) | ( n1352 & n9423 ) | ( n4235 & n9423 ) ;
  assign n20677 = n20676 ^ n14063 ^ 1'b0 ;
  assign n20678 = n20015 | n20677 ;
  assign n20679 = ( n8803 & n9094 ) | ( n8803 & ~n17854 ) | ( n9094 & ~n17854 ) ;
  assign n20680 = n5035 ^ n3331 ^ n2687 ;
  assign n20681 = n20680 ^ n4458 ^ n4034 ;
  assign n20682 = ( n1927 & n5869 ) | ( n1927 & n20681 ) | ( n5869 & n20681 ) ;
  assign n20683 = n15449 ^ n7661 ^ n3015 ;
  assign n20684 = ( ~n4401 & n20682 ) | ( ~n4401 & n20683 ) | ( n20682 & n20683 ) ;
  assign n20685 = n4559 | n16521 ;
  assign n20686 = n20685 ^ n13162 ^ n5224 ;
  assign n20690 = ( n215 & ~n2230 ) | ( n215 & n3716 ) | ( ~n2230 & n3716 ) ;
  assign n20687 = n2984 ^ n521 ^ 1'b0 ;
  assign n20688 = n4519 & n20687 ;
  assign n20689 = ( n1970 & ~n10876 ) | ( n1970 & n20688 ) | ( ~n10876 & n20688 ) ;
  assign n20691 = n20690 ^ n20689 ^ n8743 ;
  assign n20692 = ( n4418 & n10645 ) | ( n4418 & ~n10827 ) | ( n10645 & ~n10827 ) ;
  assign n20693 = n20692 ^ n18634 ^ 1'b0 ;
  assign n20694 = n19997 & n20693 ;
  assign n20695 = n4939 & n10332 ;
  assign n20696 = ~n2450 & n20695 ;
  assign n20697 = ( n457 & n2429 ) | ( n457 & ~n20696 ) | ( n2429 & ~n20696 ) ;
  assign n20698 = ( n5484 & ~n10142 ) | ( n5484 & n20697 ) | ( ~n10142 & n20697 ) ;
  assign n20699 = n2893 | n20698 ;
  assign n20700 = n20699 ^ n20624 ^ 1'b0 ;
  assign n20701 = ( n1503 & n15954 ) | ( n1503 & ~n19109 ) | ( n15954 & ~n19109 ) ;
  assign n20702 = n19300 ^ n10075 ^ n6255 ;
  assign n20703 = n19812 ^ n8039 ^ n1724 ;
  assign n20704 = n20703 ^ n16022 ^ n2108 ;
  assign n20705 = ( n9391 & ~n9423 ) | ( n9391 & n15739 ) | ( ~n9423 & n15739 ) ;
  assign n20706 = n10170 & ~n20705 ;
  assign n20707 = n20706 ^ n1805 ^ 1'b0 ;
  assign n20708 = n20707 ^ n17513 ^ n13273 ;
  assign n20709 = ( n7453 & n11613 ) | ( n7453 & ~n20708 ) | ( n11613 & ~n20708 ) ;
  assign n20710 = n8414 ^ n3650 ^ n2704 ;
  assign n20711 = ( n7926 & ~n15930 ) | ( n7926 & n20710 ) | ( ~n15930 & n20710 ) ;
  assign n20712 = ( n11921 & n18936 ) | ( n11921 & n20711 ) | ( n18936 & n20711 ) ;
  assign n20713 = ( ~n8010 & n12460 ) | ( ~n8010 & n20712 ) | ( n12460 & n20712 ) ;
  assign n20714 = n360 | n20713 ;
  assign n20715 = n6019 ^ n2083 ^ n507 ;
  assign n20716 = n16046 ^ n9663 ^ 1'b0 ;
  assign n20717 = n20715 & n20716 ;
  assign n20718 = n1481 ^ n1361 ^ 1'b0 ;
  assign n20719 = ~n2198 & n19924 ;
  assign n20720 = ~n20718 & n20719 ;
  assign n20721 = ( n1607 & ~n11605 ) | ( n1607 & n20720 ) | ( ~n11605 & n20720 ) ;
  assign n20722 = n20717 & ~n20721 ;
  assign n20723 = n20722 ^ n13918 ^ 1'b0 ;
  assign n20724 = n13416 ^ n9212 ^ 1'b0 ;
  assign n20725 = n2662 | n20724 ;
  assign n20726 = n15741 ^ n1617 ^ 1'b0 ;
  assign n20727 = n2383 & ~n20726 ;
  assign n20728 = ~n8468 & n9117 ;
  assign n20729 = n20728 ^ n10511 ^ 1'b0 ;
  assign n20730 = n20729 ^ n9611 ^ n6236 ;
  assign n20731 = ( n5892 & ~n6480 ) | ( n5892 & n7830 ) | ( ~n6480 & n7830 ) ;
  assign n20732 = n2643 & n4848 ;
  assign n20733 = ~n20731 & n20732 ;
  assign n20734 = ~n5167 & n20733 ;
  assign n20735 = ( n10046 & n11128 ) | ( n10046 & n12967 ) | ( n11128 & n12967 ) ;
  assign n20736 = n9594 ^ n4243 ^ n1515 ;
  assign n20737 = n20736 ^ x92 ^ 1'b0 ;
  assign n20739 = n1455 & n13316 ;
  assign n20740 = n20739 ^ n3485 ^ 1'b0 ;
  assign n20738 = n12885 ^ n5667 ^ n4598 ;
  assign n20741 = n20740 ^ n20738 ^ n5476 ;
  assign n20743 = ( n4240 & ~n4861 ) | ( n4240 & n12060 ) | ( ~n4861 & n12060 ) ;
  assign n20744 = n6731 ^ n2902 ^ 1'b0 ;
  assign n20745 = ( n14774 & n20743 ) | ( n14774 & ~n20744 ) | ( n20743 & ~n20744 ) ;
  assign n20746 = ~n10480 & n20745 ;
  assign n20747 = n13341 & n20746 ;
  assign n20742 = n1042 & n13857 ;
  assign n20748 = n20747 ^ n20742 ^ 1'b0 ;
  assign n20749 = n17470 ^ n14833 ^ n9186 ;
  assign n20750 = ( n10587 & n15603 ) | ( n10587 & ~n20749 ) | ( n15603 & ~n20749 ) ;
  assign n20751 = n6562 ^ n3424 ^ n382 ;
  assign n20752 = n20751 ^ n11845 ^ n2495 ;
  assign n20753 = ( n4830 & n10022 ) | ( n4830 & n10519 ) | ( n10022 & n10519 ) ;
  assign n20754 = ( n1411 & ~n2664 ) | ( n1411 & n11812 ) | ( ~n2664 & n11812 ) ;
  assign n20755 = ( n6698 & n20753 ) | ( n6698 & ~n20754 ) | ( n20753 & ~n20754 ) ;
  assign n20756 = ( ~n6301 & n7721 ) | ( ~n6301 & n18771 ) | ( n7721 & n18771 ) ;
  assign n20757 = n20756 ^ n1526 ^ 1'b0 ;
  assign n20758 = ~n483 & n4577 ;
  assign n20760 = n8467 ^ n1731 ^ 1'b0 ;
  assign n20759 = ~n4259 & n16058 ;
  assign n20761 = n20760 ^ n20759 ^ 1'b0 ;
  assign n20762 = n13102 ^ n3487 ^ n3432 ;
  assign n20763 = ( ~n163 & n827 ) | ( ~n163 & n20762 ) | ( n827 & n20762 ) ;
  assign n20764 = n8165 ^ n5446 ^ 1'b0 ;
  assign n20765 = n20764 ^ n12824 ^ n5864 ;
  assign n20766 = ( ~n4760 & n13334 ) | ( ~n4760 & n19040 ) | ( n13334 & n19040 ) ;
  assign n20767 = n11959 ^ n10982 ^ n1398 ;
  assign n20768 = n2767 & ~n3987 ;
  assign n20769 = n7080 & n20768 ;
  assign n20770 = n20769 ^ n3773 ^ 1'b0 ;
  assign n20771 = n20767 | n20770 ;
  assign n20772 = n13378 ^ n11304 ^ 1'b0 ;
  assign n20773 = ~n5533 & n20772 ;
  assign n20774 = ( ~n1889 & n4668 ) | ( ~n1889 & n7344 ) | ( n4668 & n7344 ) ;
  assign n20775 = n5446 & n18821 ;
  assign n20776 = n20775 ^ n8212 ^ n5588 ;
  assign n20777 = ( n1170 & n13604 ) | ( n1170 & ~n20776 ) | ( n13604 & ~n20776 ) ;
  assign n20778 = ( n1007 & n20774 ) | ( n1007 & ~n20777 ) | ( n20774 & ~n20777 ) ;
  assign n20779 = ~n737 & n8554 ;
  assign n20780 = n20779 ^ n1690 ^ 1'b0 ;
  assign n20781 = ( n5544 & n6478 ) | ( n5544 & ~n7321 ) | ( n6478 & ~n7321 ) ;
  assign n20782 = ( ~n1051 & n20780 ) | ( ~n1051 & n20781 ) | ( n20780 & n20781 ) ;
  assign n20788 = n8698 ^ n1501 ^ n1131 ;
  assign n20789 = n20788 ^ n6621 ^ n2127 ;
  assign n20786 = ( n159 & n6418 ) | ( n159 & n6983 ) | ( n6418 & n6983 ) ;
  assign n20787 = n20786 ^ n150 ^ 1'b0 ;
  assign n20783 = ( n1278 & ~n11909 ) | ( n1278 & n17668 ) | ( ~n11909 & n17668 ) ;
  assign n20784 = ( ~n3115 & n6383 ) | ( ~n3115 & n6413 ) | ( n6383 & n6413 ) ;
  assign n20785 = ( n10651 & n20783 ) | ( n10651 & n20784 ) | ( n20783 & n20784 ) ;
  assign n20790 = n20789 ^ n20787 ^ n20785 ;
  assign n20791 = n12491 & ~n20790 ;
  assign n20792 = ( n1892 & ~n8547 ) | ( n1892 & n9885 ) | ( ~n8547 & n9885 ) ;
  assign n20793 = n4039 & n20792 ;
  assign n20794 = n3056 & n12435 ;
  assign n20795 = ~n13271 & n20794 ;
  assign n20796 = n8647 ^ n5489 ^ n1715 ;
  assign n20797 = n18443 ^ n15869 ^ n4257 ;
  assign n20798 = n20796 & ~n20797 ;
  assign n20799 = n20795 & n20798 ;
  assign n20800 = ( ~n9279 & n12963 ) | ( ~n9279 & n18802 ) | ( n12963 & n18802 ) ;
  assign n20801 = ( n2719 & n12710 ) | ( n2719 & ~n19167 ) | ( n12710 & ~n19167 ) ;
  assign n20802 = ( n2093 & n3876 ) | ( n2093 & n19580 ) | ( n3876 & n19580 ) ;
  assign n20803 = n20802 ^ n8461 ^ n6169 ;
  assign n20804 = n5645 | n15175 ;
  assign n20805 = n20804 ^ n9927 ^ 1'b0 ;
  assign n20806 = n20805 ^ n13722 ^ n745 ;
  assign n20807 = n2528 ^ n235 ^ 1'b0 ;
  assign n20808 = ( n6119 & n18851 ) | ( n6119 & ~n20807 ) | ( n18851 & ~n20807 ) ;
  assign n20809 = ( n1218 & n1432 ) | ( n1218 & ~n16647 ) | ( n1432 & ~n16647 ) ;
  assign n20810 = n20809 ^ n20184 ^ n2819 ;
  assign n20811 = n20810 ^ n11766 ^ n5351 ;
  assign n20812 = n16030 ^ n964 ^ 1'b0 ;
  assign n20813 = n3056 | n8414 ;
  assign n20814 = n20813 ^ n13615 ^ n12321 ;
  assign n20815 = ( ~n6801 & n10925 ) | ( ~n6801 & n20814 ) | ( n10925 & n20814 ) ;
  assign n20816 = ( n12053 & n20812 ) | ( n12053 & ~n20815 ) | ( n20812 & ~n20815 ) ;
  assign n20817 = n6231 ^ n4016 ^ 1'b0 ;
  assign n20818 = n20817 ^ n2144 ^ n247 ;
  assign n20819 = ( ~n10314 & n20131 ) | ( ~n10314 & n20818 ) | ( n20131 & n20818 ) ;
  assign n20820 = n15242 ^ n8109 ^ n7128 ;
  assign n20821 = n20820 ^ n19181 ^ n9291 ;
  assign n20822 = n8983 ^ n5273 ^ n2411 ;
  assign n20823 = ( n1449 & ~n16668 ) | ( n1449 & n17031 ) | ( ~n16668 & n17031 ) ;
  assign n20824 = ( n10171 & ~n20822 ) | ( n10171 & n20823 ) | ( ~n20822 & n20823 ) ;
  assign n20825 = n20401 ^ n18613 ^ n2210 ;
  assign n20829 = n7881 & ~n10040 ;
  assign n20826 = n15266 ^ n9754 ^ 1'b0 ;
  assign n20827 = n5816 | n20826 ;
  assign n20828 = n20827 ^ n17519 ^ n7198 ;
  assign n20830 = n20829 ^ n20828 ^ 1'b0 ;
  assign n20831 = n10170 & ~n14641 ;
  assign n20832 = n745 & ~n10706 ;
  assign n20833 = ~n14538 & n17417 ;
  assign n20834 = n20833 ^ n14187 ^ n991 ;
  assign n20835 = n20834 ^ n709 ^ 1'b0 ;
  assign n20836 = n4532 & n20835 ;
  assign n20837 = n15838 ^ n6852 ^ n1920 ;
  assign n20838 = ( n6530 & n6880 ) | ( n6530 & ~n14197 ) | ( n6880 & ~n14197 ) ;
  assign n20839 = n20820 ^ n20143 ^ n4899 ;
  assign n20840 = ( n1899 & ~n2944 ) | ( n1899 & n9276 ) | ( ~n2944 & n9276 ) ;
  assign n20841 = ( n20838 & n20839 ) | ( n20838 & ~n20840 ) | ( n20839 & ~n20840 ) ;
  assign n20842 = n6094 ^ n5346 ^ n4989 ;
  assign n20843 = n5597 & ~n14920 ;
  assign n20844 = n20843 ^ n4232 ^ 1'b0 ;
  assign n20845 = n4909 | n20844 ;
  assign n20846 = n5078 & ~n10866 ;
  assign n20847 = n20846 ^ n567 ^ 1'b0 ;
  assign n20848 = n17430 ^ n17085 ^ n6087 ;
  assign n20849 = n16617 ^ n854 ^ 1'b0 ;
  assign n20850 = n4584 & n20849 ;
  assign n20851 = ( n939 & ~n9335 ) | ( n939 & n20850 ) | ( ~n9335 & n20850 ) ;
  assign n20852 = ( n5399 & n5406 ) | ( n5399 & n18363 ) | ( n5406 & n18363 ) ;
  assign n20853 = ~n7164 & n13917 ;
  assign n20854 = n20853 ^ n2868 ^ 1'b0 ;
  assign n20855 = n20764 ^ n3518 ^ n826 ;
  assign n20856 = ( n6966 & n15769 ) | ( n6966 & n20855 ) | ( n15769 & n20855 ) ;
  assign n20857 = n5587 ^ n1797 ^ n1268 ;
  assign n20858 = n20467 ^ n10722 ^ n1901 ;
  assign n20859 = ( n962 & ~n5843 ) | ( n962 & n20858 ) | ( ~n5843 & n20858 ) ;
  assign n20860 = ( ~n20469 & n20825 ) | ( ~n20469 & n20859 ) | ( n20825 & n20859 ) ;
  assign n20861 = n13887 ^ n2640 ^ 1'b0 ;
  assign n20862 = n816 & ~n20861 ;
  assign n20863 = n7450 ^ n6048 ^ n1513 ;
  assign n20864 = n18795 ^ n10912 ^ n1866 ;
  assign n20865 = n20864 ^ n12362 ^ n4439 ;
  assign n20866 = ( n8577 & n20863 ) | ( n8577 & ~n20865 ) | ( n20863 & ~n20865 ) ;
  assign n20867 = ( n7345 & n20862 ) | ( n7345 & ~n20866 ) | ( n20862 & ~n20866 ) ;
  assign n20868 = ~n786 & n10638 ;
  assign n20869 = ( n1940 & ~n19674 ) | ( n1940 & n20868 ) | ( ~n19674 & n20868 ) ;
  assign n20870 = n19920 ^ n14202 ^ 1'b0 ;
  assign n20871 = n20869 & n20870 ;
  assign n20872 = n20871 ^ n15459 ^ n10247 ;
  assign n20875 = n16038 ^ n5981 ^ n1776 ;
  assign n20874 = n14053 ^ n11896 ^ n3746 ;
  assign n20876 = n20875 ^ n20874 ^ n1137 ;
  assign n20873 = ( x26 & n2147 ) | ( x26 & n5248 ) | ( n2147 & n5248 ) ;
  assign n20877 = n20876 ^ n20873 ^ n13424 ;
  assign n20878 = n685 | n10244 ;
  assign n20879 = n9383 & ~n20878 ;
  assign n20880 = n15026 ^ n2735 ^ n1249 ;
  assign n20881 = ~n18795 & n20880 ;
  assign n20882 = ( n4208 & n11048 ) | ( n4208 & n19706 ) | ( n11048 & n19706 ) ;
  assign n20883 = ( n10744 & ~n11076 ) | ( n10744 & n20265 ) | ( ~n11076 & n20265 ) ;
  assign n20884 = ( n15019 & ~n20882 ) | ( n15019 & n20883 ) | ( ~n20882 & n20883 ) ;
  assign n20885 = ( ~n4834 & n5229 ) | ( ~n4834 & n8785 ) | ( n5229 & n8785 ) ;
  assign n20886 = n20885 ^ n5547 ^ n3773 ;
  assign n20887 = n3268 ^ n318 ^ n145 ;
  assign n20888 = n20887 ^ n19915 ^ n14875 ;
  assign n20889 = ( n5943 & ~n12075 ) | ( n5943 & n20888 ) | ( ~n12075 & n20888 ) ;
  assign n20890 = ( n3147 & n3469 ) | ( n3147 & n8460 ) | ( n3469 & n8460 ) ;
  assign n20891 = n20890 ^ n10610 ^ n8731 ;
  assign n20892 = ( n17016 & n18045 ) | ( n17016 & ~n18218 ) | ( n18045 & ~n18218 ) ;
  assign n20893 = n7775 | n10192 ;
  assign n20894 = n20893 ^ n10344 ^ 1'b0 ;
  assign n20895 = n1046 | n20894 ;
  assign n20896 = ( n4459 & n10678 ) | ( n4459 & n13396 ) | ( n10678 & n13396 ) ;
  assign n20897 = n2305 & n20896 ;
  assign n20898 = n20897 ^ n14646 ^ 1'b0 ;
  assign n20899 = n14592 & ~n20898 ;
  assign n20900 = n8058 ^ n6219 ^ n3262 ;
  assign n20901 = n20900 ^ n5332 ^ n4788 ;
  assign n20903 = ( n3447 & n13716 ) | ( n3447 & n18561 ) | ( n13716 & n18561 ) ;
  assign n20902 = n17609 ^ n16818 ^ n7378 ;
  assign n20904 = n20903 ^ n20902 ^ n10869 ;
  assign n20905 = ( ~n237 & n2260 ) | ( ~n237 & n20904 ) | ( n2260 & n20904 ) ;
  assign n20906 = ( n4127 & n5243 ) | ( n4127 & n7177 ) | ( n5243 & n7177 ) ;
  assign n20907 = ( ~n7933 & n10631 ) | ( ~n7933 & n20906 ) | ( n10631 & n20906 ) ;
  assign n20908 = ( n4963 & n14875 ) | ( n4963 & n20907 ) | ( n14875 & n20907 ) ;
  assign n20909 = ( n849 & n7917 ) | ( n849 & ~n12999 ) | ( n7917 & ~n12999 ) ;
  assign n20910 = ( ~n3257 & n4528 ) | ( ~n3257 & n14649 ) | ( n4528 & n14649 ) ;
  assign n20911 = n19812 & n20910 ;
  assign n20912 = n20911 ^ n16171 ^ 1'b0 ;
  assign n20913 = n20912 ^ n9439 ^ n8211 ;
  assign n20914 = n20913 ^ n11189 ^ n398 ;
  assign n20915 = n1902 | n9265 ;
  assign n20916 = n20915 ^ n6495 ^ 1'b0 ;
  assign n20917 = n10235 ^ n3324 ^ 1'b0 ;
  assign n20918 = ( n7644 & n9210 ) | ( n7644 & ~n19000 ) | ( n9210 & ~n19000 ) ;
  assign n20919 = ( ~n20916 & n20917 ) | ( ~n20916 & n20918 ) | ( n20917 & n20918 ) ;
  assign n20920 = ( n2458 & n7260 ) | ( n2458 & n19093 ) | ( n7260 & n19093 ) ;
  assign n20921 = n6130 & n8883 ;
  assign n20923 = ( n1875 & n6671 ) | ( n1875 & ~n10786 ) | ( n6671 & ~n10786 ) ;
  assign n20922 = ( n5138 & n5721 ) | ( n5138 & ~n14055 ) | ( n5721 & ~n14055 ) ;
  assign n20924 = n20923 ^ n20922 ^ n2025 ;
  assign n20925 = n12755 & ~n20924 ;
  assign n20926 = n20921 & n20925 ;
  assign n20927 = n6242 | n9476 ;
  assign n20928 = n20927 ^ n8762 ^ 1'b0 ;
  assign n20931 = n17234 ^ n6335 ^ n2594 ;
  assign n20929 = n7031 ^ n4092 ^ 1'b0 ;
  assign n20930 = n12229 & ~n20929 ;
  assign n20932 = n20931 ^ n20930 ^ n1865 ;
  assign n20933 = n14911 ^ n3031 ^ n900 ;
  assign n20937 = ( ~n1604 & n1740 ) | ( ~n1604 & n2081 ) | ( n1740 & n2081 ) ;
  assign n20934 = n15739 ^ n15592 ^ n6610 ;
  assign n20935 = n10292 & n20934 ;
  assign n20936 = n2599 & n20935 ;
  assign n20938 = n20937 ^ n20936 ^ n17713 ;
  assign n20939 = ( ~n6277 & n20933 ) | ( ~n6277 & n20938 ) | ( n20933 & n20938 ) ;
  assign n20940 = n2950 | n19226 ;
  assign n20941 = n20940 ^ n18099 ^ n4363 ;
  assign n20942 = ( n8809 & n17729 ) | ( n8809 & ~n18550 ) | ( n17729 & ~n18550 ) ;
  assign n20943 = n12297 ^ n7154 ^ n258 ;
  assign n20948 = n4541 ^ n681 ^ 1'b0 ;
  assign n20949 = n18743 & n20948 ;
  assign n20950 = n20949 ^ n1395 ^ n1084 ;
  assign n20947 = n14644 ^ n6857 ^ n6581 ;
  assign n20951 = n20950 ^ n20947 ^ 1'b0 ;
  assign n20952 = ~n6801 & n20951 ;
  assign n20944 = n1165 & ~n1813 ;
  assign n20945 = n4954 & n20944 ;
  assign n20946 = n20945 ^ n3618 ^ n2047 ;
  assign n20953 = n20952 ^ n20946 ^ n17857 ;
  assign n20954 = n8164 ^ n4421 ^ n1081 ;
  assign n20955 = n20954 ^ n11755 ^ n11250 ;
  assign n20956 = n16346 ^ n5495 ^ n3977 ;
  assign n20957 = n14680 ^ n5543 ^ n696 ;
  assign n20958 = ( n6024 & n13995 ) | ( n6024 & n20957 ) | ( n13995 & n20957 ) ;
  assign n20959 = ( ~n9084 & n20956 ) | ( ~n9084 & n20958 ) | ( n20956 & n20958 ) ;
  assign n20960 = n20959 ^ n12749 ^ n5526 ;
  assign n20961 = n6729 ^ n1231 ^ x58 ;
  assign n20962 = n3624 ^ n3213 ^ 1'b0 ;
  assign n20963 = n5394 | n20962 ;
  assign n20964 = n20963 ^ n6676 ^ n6186 ;
  assign n20965 = n12537 ^ n4336 ^ n3539 ;
  assign n20966 = ( ~n8958 & n20964 ) | ( ~n8958 & n20965 ) | ( n20964 & n20965 ) ;
  assign n20967 = ~n379 & n3564 ;
  assign n20968 = n20967 ^ n11492 ^ 1'b0 ;
  assign n20969 = n16575 & n16820 ;
  assign n20970 = ~n7028 & n20969 ;
  assign n20971 = n6407 ^ n4583 ^ n890 ;
  assign n20972 = n1812 & ~n20971 ;
  assign n20973 = ( n5672 & n8592 ) | ( n5672 & n20972 ) | ( n8592 & n20972 ) ;
  assign n20974 = n20973 ^ n18468 ^ n16648 ;
  assign n20975 = ( n6503 & n9863 ) | ( n6503 & n11832 ) | ( n9863 & n11832 ) ;
  assign n20976 = n13448 ^ n4760 ^ n3161 ;
  assign n20977 = n10681 | n19228 ;
  assign n20978 = n20977 ^ n7792 ^ n2393 ;
  assign n20979 = ( n5998 & n7831 ) | ( n5998 & ~n15084 ) | ( n7831 & ~n15084 ) ;
  assign n20980 = n20979 ^ n18626 ^ n14595 ;
  assign n20981 = n20980 ^ n11766 ^ 1'b0 ;
  assign n20982 = n8036 | n20981 ;
  assign n20983 = ( n2907 & n5474 ) | ( n2907 & ~n13663 ) | ( n5474 & ~n13663 ) ;
  assign n20984 = n20983 ^ n1263 ^ 1'b0 ;
  assign n20985 = n7979 ^ n7303 ^ n6598 ;
  assign n20986 = ( n514 & ~n2688 ) | ( n514 & n4167 ) | ( ~n2688 & n4167 ) ;
  assign n20987 = ( n5731 & n8793 ) | ( n5731 & ~n20986 ) | ( n8793 & ~n20986 ) ;
  assign n20988 = n1893 & n20987 ;
  assign n20989 = n20988 ^ n2427 ^ 1'b0 ;
  assign n20990 = n20989 ^ n6411 ^ n5227 ;
  assign n20991 = ( n1662 & n20985 ) | ( n1662 & n20990 ) | ( n20985 & n20990 ) ;
  assign n20992 = n20984 | n20991 ;
  assign n20993 = ( ~n773 & n2029 ) | ( ~n773 & n2092 ) | ( n2029 & n2092 ) ;
  assign n20994 = n20993 ^ n3000 ^ n2084 ;
  assign n20995 = ~n5564 & n19723 ;
  assign n20996 = ~n2004 & n20995 ;
  assign n20997 = n17973 ^ n16479 ^ n8178 ;
  assign n20998 = ( ~n9662 & n20996 ) | ( ~n9662 & n20997 ) | ( n20996 & n20997 ) ;
  assign n20999 = ( n4633 & n20994 ) | ( n4633 & n20998 ) | ( n20994 & n20998 ) ;
  assign n21005 = n17006 ^ n7039 ^ n2531 ;
  assign n21003 = n9083 ^ n6987 ^ n450 ;
  assign n21004 = n21003 ^ n12040 ^ n3667 ;
  assign n21000 = n6513 ^ n6000 ^ 1'b0 ;
  assign n21001 = n21000 ^ n1456 ^ n688 ;
  assign n21002 = n21001 ^ n13763 ^ n2441 ;
  assign n21006 = n21005 ^ n21004 ^ n21002 ;
  assign n21007 = n6818 ^ n3135 ^ n523 ;
  assign n21008 = n8193 ^ n3030 ^ 1'b0 ;
  assign n21009 = n4934 | n7633 ;
  assign n21010 = n21008 & ~n21009 ;
  assign n21011 = n14524 ^ n4434 ^ n1244 ;
  assign n21012 = n9977 ^ n9738 ^ n4213 ;
  assign n21013 = ( n8711 & ~n9125 ) | ( n8711 & n21012 ) | ( ~n9125 & n21012 ) ;
  assign n21014 = ( n10693 & ~n15429 ) | ( n10693 & n20469 ) | ( ~n15429 & n20469 ) ;
  assign n21015 = n20245 ^ n18789 ^ n5436 ;
  assign n21016 = n20769 ^ n3893 ^ n2554 ;
  assign n21017 = ( ~n13828 & n19872 ) | ( ~n13828 & n21016 ) | ( n19872 & n21016 ) ;
  assign n21018 = ( ~x42 & n2983 ) | ( ~x42 & n15340 ) | ( n2983 & n15340 ) ;
  assign n21019 = ~n12493 & n13920 ;
  assign n21020 = n21019 ^ n8112 ^ 1'b0 ;
  assign n21021 = n21018 | n21020 ;
  assign n21022 = n15759 ^ n11304 ^ n1244 ;
  assign n21023 = n21022 ^ n4676 ^ 1'b0 ;
  assign n21024 = n14063 & ~n16127 ;
  assign n21025 = n21023 & n21024 ;
  assign n21026 = n21021 | n21025 ;
  assign n21027 = n21026 ^ n4485 ^ 1'b0 ;
  assign n21028 = ( n1883 & ~n2081 ) | ( n1883 & n4400 ) | ( ~n2081 & n4400 ) ;
  assign n21029 = ( ~n1728 & n19236 ) | ( ~n1728 & n21028 ) | ( n19236 & n21028 ) ;
  assign n21030 = n21029 ^ n8111 ^ 1'b0 ;
  assign n21031 = n15817 ^ n7342 ^ n7070 ;
  assign n21032 = n21031 ^ n17891 ^ n6588 ;
  assign n21033 = n4419 ^ n2976 ^ n1797 ;
  assign n21034 = n21033 ^ n17443 ^ n6608 ;
  assign n21035 = ( x38 & ~n10181 ) | ( x38 & n15775 ) | ( ~n10181 & n15775 ) ;
  assign n21036 = n6637 ^ n1990 ^ 1'b0 ;
  assign n21037 = n21036 ^ n20500 ^ n194 ;
  assign n21038 = ( n19405 & n21035 ) | ( n19405 & n21037 ) | ( n21035 & n21037 ) ;
  assign n21039 = n10821 ^ n513 ^ n248 ;
  assign n21040 = ~n5671 & n21039 ;
  assign n21041 = n5074 ^ n4680 ^ 1'b0 ;
  assign n21042 = n4102 & n21041 ;
  assign n21043 = ( n1304 & ~n1956 ) | ( n1304 & n6466 ) | ( ~n1956 & n6466 ) ;
  assign n21044 = ( n9116 & ~n17775 ) | ( n9116 & n21043 ) | ( ~n17775 & n21043 ) ;
  assign n21045 = n16180 ^ n14492 ^ n6997 ;
  assign n21046 = ( n9121 & n13187 ) | ( n9121 & ~n17825 ) | ( n13187 & ~n17825 ) ;
  assign n21047 = n13571 ^ n13465 ^ n10133 ;
  assign n21048 = ( ~n1773 & n7241 ) | ( ~n1773 & n12871 ) | ( n7241 & n12871 ) ;
  assign n21049 = ( ~n11755 & n17077 ) | ( ~n11755 & n21048 ) | ( n17077 & n21048 ) ;
  assign n21050 = n3757 & n14545 ;
  assign n21051 = ~n21049 & n21050 ;
  assign n21052 = ( n6340 & ~n6426 ) | ( n6340 & n7824 ) | ( ~n6426 & n7824 ) ;
  assign n21054 = n19375 ^ n13402 ^ n11021 ;
  assign n21053 = n4465 | n14017 ;
  assign n21055 = n21054 ^ n21053 ^ 1'b0 ;
  assign n21056 = ( n1091 & ~n1292 ) | ( n1091 & n1969 ) | ( ~n1292 & n1969 ) ;
  assign n21057 = n1842 ^ n944 ^ 1'b0 ;
  assign n21058 = n21056 & ~n21057 ;
  assign n21059 = n9444 ^ n164 ^ 1'b0 ;
  assign n21060 = ( ~n1880 & n21058 ) | ( ~n1880 & n21059 ) | ( n21058 & n21059 ) ;
  assign n21061 = ( ~n21052 & n21055 ) | ( ~n21052 & n21060 ) | ( n21055 & n21060 ) ;
  assign n21062 = n6556 ^ n6391 ^ n3899 ;
  assign n21063 = n18800 ^ n7366 ^ 1'b0 ;
  assign n21064 = ( n2959 & ~n9652 ) | ( n2959 & n21063 ) | ( ~n9652 & n21063 ) ;
  assign n21065 = n21064 ^ n19485 ^ n17631 ;
  assign n21066 = n21065 ^ n5219 ^ n3703 ;
  assign n21067 = n7251 ^ n4477 ^ n2790 ;
  assign n21068 = ( n8685 & n19736 ) | ( n8685 & ~n21067 ) | ( n19736 & ~n21067 ) ;
  assign n21069 = ( n152 & n5217 ) | ( n152 & n15476 ) | ( n5217 & n15476 ) ;
  assign n21070 = n3885 | n7329 ;
  assign n21071 = n21069 & ~n21070 ;
  assign n21072 = n15821 ^ n1578 ^ 1'b0 ;
  assign n21073 = n21072 ^ n19865 ^ 1'b0 ;
  assign n21074 = n13511 ^ n1420 ^ 1'b0 ;
  assign n21075 = n12113 ^ n10090 ^ n2677 ;
  assign n21076 = n14193 ^ n14024 ^ n9674 ;
  assign n21077 = n3590 ^ n3042 ^ 1'b0 ;
  assign n21078 = n21077 ^ n11018 ^ n6076 ;
  assign n21079 = ( n212 & n7428 ) | ( n212 & ~n21078 ) | ( n7428 & ~n21078 ) ;
  assign n21080 = n21076 & n21079 ;
  assign n21081 = n17405 & n21080 ;
  assign n21083 = n14550 ^ n6187 ^ 1'b0 ;
  assign n21084 = n21083 ^ n4971 ^ n2228 ;
  assign n21082 = n3400 | n10408 ;
  assign n21085 = n21084 ^ n21082 ^ n13175 ;
  assign n21086 = n20780 ^ n1690 ^ 1'b0 ;
  assign n21087 = n7053 | n21086 ;
  assign n21088 = ~n17180 & n21087 ;
  assign n21089 = ( ~n1369 & n7650 ) | ( ~n1369 & n12223 ) | ( n7650 & n12223 ) ;
  assign n21090 = n21089 ^ n7516 ^ n4122 ;
  assign n21092 = n8323 ^ n5088 ^ n3042 ;
  assign n21091 = n14768 ^ n1544 ^ n1225 ;
  assign n21093 = n21092 ^ n21091 ^ x70 ;
  assign n21094 = ( n5622 & n9036 ) | ( n5622 & n21093 ) | ( n9036 & n21093 ) ;
  assign n21095 = ~n3531 & n3892 ;
  assign n21096 = ( n5494 & ~n10024 ) | ( n5494 & n21095 ) | ( ~n10024 & n21095 ) ;
  assign n21097 = ( ~n3063 & n11754 ) | ( ~n3063 & n21096 ) | ( n11754 & n21096 ) ;
  assign n21098 = ( n1027 & ~n1100 ) | ( n1027 & n21097 ) | ( ~n1100 & n21097 ) ;
  assign n21099 = n5650 & ~n8837 ;
  assign n21100 = n2220 & n21099 ;
  assign n21101 = n21100 ^ n9737 ^ 1'b0 ;
  assign n21102 = n18921 | n20997 ;
  assign n21103 = n16558 ^ n12489 ^ n5902 ;
  assign n21104 = n15268 ^ n7519 ^ 1'b0 ;
  assign n21105 = n3355 & ~n21104 ;
  assign n21106 = n8010 & ~n14001 ;
  assign n21107 = ( n855 & n7883 ) | ( n855 & ~n9335 ) | ( n7883 & ~n9335 ) ;
  assign n21118 = ( n400 & ~n3541 ) | ( n400 & n3705 ) | ( ~n3541 & n3705 ) ;
  assign n21108 = n9121 ^ n5051 ^ n1657 ;
  assign n21109 = n21108 ^ n6884 ^ n5454 ;
  assign n21110 = n2004 & ~n7678 ;
  assign n21111 = ~n21109 & n21110 ;
  assign n21112 = n12395 ^ n11635 ^ n11075 ;
  assign n21113 = ( n7772 & ~n21111 ) | ( n7772 & n21112 ) | ( ~n21111 & n21112 ) ;
  assign n21114 = ( n6130 & n6163 ) | ( n6130 & n16708 ) | ( n6163 & n16708 ) ;
  assign n21115 = ( n1231 & n5148 ) | ( n1231 & ~n7942 ) | ( n5148 & ~n7942 ) ;
  assign n21116 = ( n11366 & ~n21114 ) | ( n11366 & n21115 ) | ( ~n21114 & n21115 ) ;
  assign n21117 = ( n6835 & n21113 ) | ( n6835 & ~n21116 ) | ( n21113 & ~n21116 ) ;
  assign n21119 = n21118 ^ n21117 ^ n1356 ;
  assign n21122 = ~n5644 & n15620 ;
  assign n21120 = n8725 | n16065 ;
  assign n21121 = n19582 | n21120 ;
  assign n21123 = n21122 ^ n21121 ^ n13921 ;
  assign n21124 = n10291 ^ n7732 ^ n3832 ;
  assign n21125 = ( n3727 & n5081 ) | ( n3727 & ~n5354 ) | ( n5081 & ~n5354 ) ;
  assign n21126 = n21125 ^ n19267 ^ 1'b0 ;
  assign n21127 = ( ~n15217 & n21124 ) | ( ~n15217 & n21126 ) | ( n21124 & n21126 ) ;
  assign n21128 = n10083 ^ n4958 ^ n1677 ;
  assign n21129 = ( n8467 & ~n11433 ) | ( n8467 & n21128 ) | ( ~n11433 & n21128 ) ;
  assign n21130 = ( n8291 & ~n12156 ) | ( n8291 & n21129 ) | ( ~n12156 & n21129 ) ;
  assign n21131 = ( n3091 & ~n11258 ) | ( n3091 & n18350 ) | ( ~n11258 & n18350 ) ;
  assign n21132 = ( ~n5264 & n6459 ) | ( ~n5264 & n21131 ) | ( n6459 & n21131 ) ;
  assign n21134 = ( n5726 & n7162 ) | ( n5726 & ~n12626 ) | ( n7162 & ~n12626 ) ;
  assign n21135 = ~n12322 & n21134 ;
  assign n21136 = ~n14370 & n21135 ;
  assign n21133 = n9528 & n12289 ;
  assign n21137 = n21136 ^ n21133 ^ 1'b0 ;
  assign n21138 = n4223 ^ n3541 ^ 1'b0 ;
  assign n21144 = n10457 ^ n10385 ^ n235 ;
  assign n21141 = ~n2928 & n11829 ;
  assign n21142 = ~n10843 & n21141 ;
  assign n21139 = n13428 & ~n14458 ;
  assign n21140 = n21139 ^ n14623 ^ 1'b0 ;
  assign n21143 = n21142 ^ n21140 ^ n15206 ;
  assign n21145 = n21144 ^ n21143 ^ n8972 ;
  assign n21146 = ( x64 & n8051 ) | ( x64 & ~n17163 ) | ( n8051 & ~n17163 ) ;
  assign n21147 = ( n6962 & n9128 ) | ( n6962 & n13645 ) | ( n9128 & n13645 ) ;
  assign n21148 = n11227 ^ n4728 ^ n4166 ;
  assign n21152 = n18811 ^ n12441 ^ n8540 ;
  assign n21149 = n14768 ^ n9034 ^ 1'b0 ;
  assign n21150 = ~n5641 & n21149 ;
  assign n21151 = n8704 & n21150 ;
  assign n21153 = n21152 ^ n21151 ^ n10239 ;
  assign n21154 = n9056 ^ n337 ^ 1'b0 ;
  assign n21155 = n19391 ^ n15835 ^ 1'b0 ;
  assign n21156 = n11868 & ~n21155 ;
  assign n21158 = n5949 ^ n4105 ^ 1'b0 ;
  assign n21159 = n21158 ^ n4233 ^ n4102 ;
  assign n21157 = ( n941 & n5932 ) | ( n941 & ~n17114 ) | ( n5932 & ~n17114 ) ;
  assign n21160 = n21159 ^ n21157 ^ n16573 ;
  assign n21161 = ( ~n3272 & n4504 ) | ( ~n3272 & n12742 ) | ( n4504 & n12742 ) ;
  assign n21162 = n21161 ^ n18917 ^ n5548 ;
  assign n21163 = ( n5608 & n18426 ) | ( n5608 & ~n18703 ) | ( n18426 & ~n18703 ) ;
  assign n21164 = n3706 & ~n4270 ;
  assign n21165 = n21164 ^ n8932 ^ n8749 ;
  assign n21166 = ( n4861 & ~n7715 ) | ( n4861 & n11771 ) | ( ~n7715 & n11771 ) ;
  assign n21167 = n15535 & n21166 ;
  assign n21168 = n21167 ^ n20194 ^ 1'b0 ;
  assign n21169 = ( n3742 & n4940 ) | ( n3742 & n17496 ) | ( n4940 & n17496 ) ;
  assign n21170 = ( n4837 & n5955 ) | ( n4837 & n6107 ) | ( n5955 & n6107 ) ;
  assign n21171 = ( n3660 & ~n8218 ) | ( n3660 & n21170 ) | ( ~n8218 & n21170 ) ;
  assign n21172 = n17041 ^ n12717 ^ n11168 ;
  assign n21173 = n13383 ^ n7042 ^ n2108 ;
  assign n21181 = n2999 ^ n1302 ^ n1104 ;
  assign n21182 = n21181 ^ n8674 ^ n1625 ;
  assign n21179 = n15735 ^ n4803 ^ 1'b0 ;
  assign n21180 = n21179 ^ n19788 ^ n9244 ;
  assign n21177 = n10337 ^ n4373 ^ n1710 ;
  assign n21178 = ( n7440 & n19052 ) | ( n7440 & n21177 ) | ( n19052 & n21177 ) ;
  assign n21183 = n21182 ^ n21180 ^ n21178 ;
  assign n21174 = ( n8608 & ~n12611 ) | ( n8608 & n18798 ) | ( ~n12611 & n18798 ) ;
  assign n21175 = n21174 ^ n18039 ^ n14417 ;
  assign n21176 = n21175 ^ n11762 ^ n3572 ;
  assign n21184 = n21183 ^ n21176 ^ n15265 ;
  assign n21185 = ( n10706 & ~n18319 ) | ( n10706 & n19795 ) | ( ~n18319 & n19795 ) ;
  assign n21186 = n7593 & ~n15742 ;
  assign n21187 = n21185 & n21186 ;
  assign n21188 = n3823 & ~n8303 ;
  assign n21189 = n14264 & n21188 ;
  assign n21190 = n17507 ^ n708 ^ 1'b0 ;
  assign n21191 = n8261 & ~n21190 ;
  assign n21192 = ( ~n1998 & n10093 ) | ( ~n1998 & n15901 ) | ( n10093 & n15901 ) ;
  assign n21193 = ( ~n6641 & n13318 ) | ( ~n6641 & n21192 ) | ( n13318 & n21192 ) ;
  assign n21194 = ( n3141 & ~n4289 ) | ( n3141 & n5574 ) | ( ~n4289 & n5574 ) ;
  assign n21195 = ( n7350 & n8241 ) | ( n7350 & ~n14676 ) | ( n8241 & ~n14676 ) ;
  assign n21197 = ( n9587 & n11441 ) | ( n9587 & n14120 ) | ( n11441 & n14120 ) ;
  assign n21196 = ~n2376 & n7387 ;
  assign n21198 = n21197 ^ n21196 ^ 1'b0 ;
  assign n21199 = n19701 ^ n8709 ^ n6904 ;
  assign n21200 = n10158 | n21199 ;
  assign n21201 = ~n868 & n21200 ;
  assign n21202 = n2723 & n21201 ;
  assign n21203 = n7549 ^ n534 ^ n207 ;
  assign n21204 = n21203 ^ n3722 ^ n2244 ;
  assign n21205 = ~n1456 & n4766 ;
  assign n21206 = ~n19651 & n21205 ;
  assign n21207 = ( n3428 & n11399 ) | ( n3428 & ~n21206 ) | ( n11399 & ~n21206 ) ;
  assign n21208 = ( n574 & n2360 ) | ( n574 & n8184 ) | ( n2360 & n8184 ) ;
  assign n21209 = n21208 ^ n1022 ^ 1'b0 ;
  assign n21210 = n21209 ^ n14915 ^ n7445 ;
  assign n21211 = n18526 ^ n13847 ^ n10467 ;
  assign n21212 = n21211 ^ n19981 ^ n2084 ;
  assign n21213 = n3863 & n5328 ;
  assign n21214 = n12976 ^ n4421 ^ n2208 ;
  assign n21215 = ( n516 & ~n7381 ) | ( n516 & n7441 ) | ( ~n7381 & n7441 ) ;
  assign n21216 = n10030 ^ n710 ^ 1'b0 ;
  assign n21217 = n3126 | n21216 ;
  assign n21218 = n19827 ^ n16407 ^ 1'b0 ;
  assign n21219 = n3339 | n21218 ;
  assign n21220 = n1922 & n18526 ;
  assign n21221 = n17966 & n21220 ;
  assign n21222 = n15879 ^ n8022 ^ n3917 ;
  assign n21223 = ( ~n5142 & n5313 ) | ( ~n5142 & n21222 ) | ( n5313 & n21222 ) ;
  assign n21224 = n6572 ^ n5137 ^ n889 ;
  assign n21225 = n394 & ~n11736 ;
  assign n21226 = ( n588 & n16035 ) | ( n588 & ~n16316 ) | ( n16035 & ~n16316 ) ;
  assign n21227 = ( n7312 & n15090 ) | ( n7312 & n21226 ) | ( n15090 & n21226 ) ;
  assign n21228 = n21227 ^ n11759 ^ n1392 ;
  assign n21229 = ( n21224 & n21225 ) | ( n21224 & n21228 ) | ( n21225 & n21228 ) ;
  assign n21230 = ( n7706 & n12859 ) | ( n7706 & n15416 ) | ( n12859 & n15416 ) ;
  assign n21231 = n3188 | n11113 ;
  assign n21232 = n17668 | n21231 ;
  assign n21233 = n21232 ^ n20632 ^ n20266 ;
  assign n21234 = ( n4340 & n4433 ) | ( n4340 & n11415 ) | ( n4433 & n11415 ) ;
  assign n21235 = n21234 ^ n7453 ^ n4653 ;
  assign n21236 = n3221 ^ n784 ^ n150 ;
  assign n21237 = n7091 & n21236 ;
  assign n21238 = n4204 & n21237 ;
  assign n21239 = n21235 & n21238 ;
  assign n21240 = n9871 ^ n1412 ^ x106 ;
  assign n21241 = ( n3157 & n5274 ) | ( n3157 & ~n5630 ) | ( n5274 & ~n5630 ) ;
  assign n21242 = ( ~n15612 & n17297 ) | ( ~n15612 & n21241 ) | ( n17297 & n21241 ) ;
  assign n21243 = n14786 ^ n489 ^ 1'b0 ;
  assign n21244 = n21243 ^ n4666 ^ 1'b0 ;
  assign n21245 = n13931 ^ n10597 ^ n5691 ;
  assign n21246 = n21245 ^ n1104 ^ 1'b0 ;
  assign n21247 = n4733 | n21246 ;
  assign n21248 = n11768 & ~n21247 ;
  assign n21249 = ( n1867 & ~n12711 ) | ( n1867 & n17390 ) | ( ~n12711 & n17390 ) ;
  assign n21250 = n13053 ^ n8875 ^ n3096 ;
  assign n21251 = n21250 ^ n16820 ^ n1657 ;
  assign n21252 = ~n4726 & n11479 ;
  assign n21253 = ~n16476 & n21252 ;
  assign n21254 = n14634 ^ n12387 ^ n3380 ;
  assign n21255 = n14325 ^ n5537 ^ n2422 ;
  assign n21256 = n21255 ^ n3780 ^ n1840 ;
  assign n21257 = ( n6352 & n15242 ) | ( n6352 & n20609 ) | ( n15242 & n20609 ) ;
  assign n21258 = ( n1896 & ~n4384 ) | ( n1896 & n5413 ) | ( ~n4384 & n5413 ) ;
  assign n21259 = n14284 & n21258 ;
  assign n21260 = n4949 & n21259 ;
  assign n21261 = n4508 & n21260 ;
  assign n21262 = n1835 | n17216 ;
  assign n21263 = n7581 ^ n2430 ^ n1748 ;
  assign n21264 = ( n4165 & n15242 ) | ( n4165 & ~n21263 ) | ( n15242 & ~n21263 ) ;
  assign n21265 = ~n1604 & n21264 ;
  assign n21266 = n5479 & n21265 ;
  assign n21267 = n13491 ^ n1217 ^ 1'b0 ;
  assign n21268 = ( ~n657 & n5978 ) | ( ~n657 & n8100 ) | ( n5978 & n8100 ) ;
  assign n21269 = n15892 ^ n8482 ^ 1'b0 ;
  assign n21270 = ~n21268 & n21269 ;
  assign n21271 = n5727 & ~n21270 ;
  assign n21272 = n10953 ^ n6231 ^ n1264 ;
  assign n21273 = ( n4037 & ~n8607 ) | ( n4037 & n21272 ) | ( ~n8607 & n21272 ) ;
  assign n21274 = n14661 ^ n3581 ^ n1878 ;
  assign n21275 = n15973 ^ n15157 ^ 1'b0 ;
  assign n21276 = n13915 & ~n21275 ;
  assign n21277 = ( n5665 & n10479 ) | ( n5665 & ~n12277 ) | ( n10479 & ~n12277 ) ;
  assign n21278 = n8920 ^ n3971 ^ 1'b0 ;
  assign n21279 = ( n4344 & n5629 ) | ( n4344 & ~n21278 ) | ( n5629 & ~n21278 ) ;
  assign n21281 = n13517 ^ n9113 ^ n1324 ;
  assign n21280 = n10109 ^ n2429 ^ n1233 ;
  assign n21282 = n21281 ^ n21280 ^ n4966 ;
  assign n21283 = ~n7943 & n21282 ;
  assign n21284 = ~n8267 & n21283 ;
  assign n21285 = n9449 ^ n1573 ^ 1'b0 ;
  assign n21286 = ~n11812 & n21285 ;
  assign n21287 = ( n12833 & n18370 ) | ( n12833 & ~n21286 ) | ( n18370 & ~n21286 ) ;
  assign n21288 = n13654 ^ n8846 ^ n2114 ;
  assign n21289 = n21288 ^ n12818 ^ n1025 ;
  assign n21290 = n21289 ^ n13980 ^ 1'b0 ;
  assign n21291 = n7130 ^ n5262 ^ n2762 ;
  assign n21292 = n21291 ^ n15412 ^ n3489 ;
  assign n21293 = n21292 ^ n20993 ^ n13468 ;
  assign n21294 = ( n4568 & n6268 ) | ( n4568 & ~n11884 ) | ( n6268 & ~n11884 ) ;
  assign n21295 = n8891 ^ n3901 ^ 1'b0 ;
  assign n21296 = n3773 & ~n21295 ;
  assign n21297 = ~n5951 & n10125 ;
  assign n21298 = ~n502 & n21297 ;
  assign n21299 = n13997 ^ n12947 ^ n2457 ;
  assign n21300 = n4177 ^ n2562 ^ n2506 ;
  assign n21301 = n724 & ~n20292 ;
  assign n21302 = n21301 ^ n19656 ^ n9774 ;
  assign n21303 = n5219 | n5585 ;
  assign n21304 = n4310 & ~n21303 ;
  assign n21305 = n21304 ^ n4158 ^ 1'b0 ;
  assign n21306 = n5146 | n21305 ;
  assign n21307 = n21306 ^ n9156 ^ n6455 ;
  assign n21308 = ( x87 & n5274 ) | ( x87 & ~n21307 ) | ( n5274 & ~n21307 ) ;
  assign n21309 = ~n2635 & n4569 ;
  assign n21310 = n21309 ^ n2439 ^ 1'b0 ;
  assign n21311 = n21310 ^ n7504 ^ 1'b0 ;
  assign n21312 = ~n7865 & n21311 ;
  assign n21313 = ( n1129 & n14661 ) | ( n1129 & n21312 ) | ( n14661 & n21312 ) ;
  assign n21314 = n261 & n1422 ;
  assign n21315 = n21314 ^ n9241 ^ 1'b0 ;
  assign n21316 = ( ~n7795 & n8634 ) | ( ~n7795 & n9347 ) | ( n8634 & n9347 ) ;
  assign n21317 = ( n3150 & n15635 ) | ( n3150 & n18676 ) | ( n15635 & n18676 ) ;
  assign n21321 = ~n7910 & n10864 ;
  assign n21322 = n21321 ^ n2726 ^ 1'b0 ;
  assign n21318 = n14675 ^ n7980 ^ n4940 ;
  assign n21319 = n1680 | n20176 ;
  assign n21320 = n21318 | n21319 ;
  assign n21323 = n21322 ^ n21320 ^ n15703 ;
  assign n21324 = n11488 ^ n4168 ^ 1'b0 ;
  assign n21325 = n2933 & ~n4627 ;
  assign n21326 = n17199 ^ n8531 ^ 1'b0 ;
  assign n21327 = ~n334 & n21326 ;
  assign n21328 = n15996 ^ n10010 ^ n3226 ;
  assign n21329 = ( ~n8716 & n21327 ) | ( ~n8716 & n21328 ) | ( n21327 & n21328 ) ;
  assign n21331 = ( n612 & n3812 ) | ( n612 & ~n6391 ) | ( n3812 & ~n6391 ) ;
  assign n21330 = ( n196 & n7369 ) | ( n196 & n20991 ) | ( n7369 & n20991 ) ;
  assign n21332 = n21331 ^ n21330 ^ n20707 ;
  assign n21333 = ( n3741 & n15766 ) | ( n3741 & n16656 ) | ( n15766 & n16656 ) ;
  assign n21334 = n13645 ^ n7714 ^ n946 ;
  assign n21335 = n21334 ^ n9298 ^ n291 ;
  assign n21336 = n18307 ^ n12985 ^ n1158 ;
  assign n21337 = n21336 ^ n15476 ^ 1'b0 ;
  assign n21338 = n14347 ^ n9331 ^ n5185 ;
  assign n21339 = n21338 ^ n9995 ^ 1'b0 ;
  assign n21340 = ( n204 & n11850 ) | ( n204 & n21339 ) | ( n11850 & n21339 ) ;
  assign n21341 = n873 | n21340 ;
  assign n21342 = n8182 ^ n5306 ^ n4821 ;
  assign n21343 = n21342 ^ n16087 ^ 1'b0 ;
  assign n21344 = ~n4406 & n21343 ;
  assign n21345 = ( ~n11201 & n13387 ) | ( ~n11201 & n21344 ) | ( n13387 & n21344 ) ;
  assign n21346 = n2190 & n5351 ;
  assign n21347 = ( ~n1844 & n2405 ) | ( ~n1844 & n21346 ) | ( n2405 & n21346 ) ;
  assign n21348 = ( n576 & n1143 ) | ( n576 & n21347 ) | ( n1143 & n21347 ) ;
  assign n21349 = n21348 ^ n18244 ^ 1'b0 ;
  assign n21350 = ~n18675 & n21349 ;
  assign n21351 = ( x51 & n2077 ) | ( x51 & n21350 ) | ( n2077 & n21350 ) ;
  assign n21354 = n7351 & ~n19341 ;
  assign n21355 = n3542 & n21354 ;
  assign n21356 = n21355 ^ n19300 ^ n12689 ;
  assign n21352 = n17265 ^ n2007 ^ 1'b0 ;
  assign n21353 = n3407 & n21352 ;
  assign n21357 = n21356 ^ n21353 ^ n20820 ;
  assign n21358 = ( n7042 & n7402 ) | ( n7042 & ~n11219 ) | ( n7402 & ~n11219 ) ;
  assign n21359 = n11571 ^ n862 ^ 1'b0 ;
  assign n21360 = n479 & n21013 ;
  assign n21361 = n9721 & n21360 ;
  assign n21362 = n21361 ^ n6687 ^ 1'b0 ;
  assign n21363 = n16872 | n21362 ;
  assign n21364 = ( n8429 & n10804 ) | ( n8429 & ~n16776 ) | ( n10804 & ~n16776 ) ;
  assign n21365 = n2659 & ~n21364 ;
  assign n21366 = n21365 ^ n8713 ^ 1'b0 ;
  assign n21367 = ( n1695 & n12750 ) | ( n1695 & ~n13313 ) | ( n12750 & ~n13313 ) ;
  assign n21368 = n6209 ^ n2827 ^ n1401 ;
  assign n21369 = ( n1897 & n3477 ) | ( n1897 & n21368 ) | ( n3477 & n21368 ) ;
  assign n21370 = n10456 ^ n6971 ^ n197 ;
  assign n21371 = n13205 | n21370 ;
  assign n21372 = ( n2926 & n4123 ) | ( n2926 & n5088 ) | ( n4123 & n5088 ) ;
  assign n21373 = n21372 ^ n20440 ^ n14611 ;
  assign n21374 = ( n3559 & ~n21371 ) | ( n3559 & n21373 ) | ( ~n21371 & n21373 ) ;
  assign n21375 = n2959 | n13436 ;
  assign n21376 = n11511 ^ n242 ^ 1'b0 ;
  assign n21377 = ~n21375 & n21376 ;
  assign n21378 = n20890 ^ n16254 ^ n1263 ;
  assign n21379 = ( n1399 & n5730 ) | ( n1399 & n8155 ) | ( n5730 & n8155 ) ;
  assign n21380 = ( ~n464 & n3469 ) | ( ~n464 & n11832 ) | ( n3469 & n11832 ) ;
  assign n21381 = ( n18948 & n21379 ) | ( n18948 & ~n21380 ) | ( n21379 & ~n21380 ) ;
  assign n21382 = ( n5447 & ~n6569 ) | ( n5447 & n15467 ) | ( ~n6569 & n15467 ) ;
  assign n21383 = n5830 ^ n5000 ^ n2982 ;
  assign n21384 = n21383 ^ n14864 ^ 1'b0 ;
  assign n21385 = n12515 ^ n7139 ^ n3554 ;
  assign n21386 = n17724 ^ n10772 ^ n6617 ;
  assign n21387 = n17034 ^ n12531 ^ n5529 ;
  assign n21388 = n6787 | n21387 ;
  assign n21389 = n16012 | n21388 ;
  assign n21390 = n11764 & ~n21389 ;
  assign n21391 = n19068 ^ n9296 ^ n7727 ;
  assign n21392 = ( n18147 & n18629 ) | ( n18147 & ~n18802 ) | ( n18629 & ~n18802 ) ;
  assign n21393 = ( n588 & ~n3728 ) | ( n588 & n6027 ) | ( ~n3728 & n6027 ) ;
  assign n21394 = n21393 ^ n5786 ^ n3276 ;
  assign n21396 = n16213 ^ n5365 ^ n4802 ;
  assign n21395 = ( n2411 & n6144 ) | ( n2411 & ~n17539 ) | ( n6144 & ~n17539 ) ;
  assign n21397 = n21396 ^ n21395 ^ n13317 ;
  assign n21398 = ( n11459 & n17793 ) | ( n11459 & ~n21397 ) | ( n17793 & ~n21397 ) ;
  assign n21399 = ( ~n6071 & n13175 ) | ( ~n6071 & n18209 ) | ( n13175 & n18209 ) ;
  assign n21400 = n7168 & n20561 ;
  assign n21401 = ~n6251 & n21400 ;
  assign n21402 = n3996 | n15269 ;
  assign n21403 = n21402 ^ n11796 ^ n4552 ;
  assign n21404 = n21403 ^ n2906 ^ 1'b0 ;
  assign n21405 = n9597 ^ n3272 ^ n2660 ;
  assign n21406 = n21405 ^ n13379 ^ n11194 ;
  assign n21407 = n16407 | n16441 ;
  assign n21408 = n21407 ^ n2011 ^ 1'b0 ;
  assign n21409 = ( x72 & ~n19656 ) | ( x72 & n21408 ) | ( ~n19656 & n21408 ) ;
  assign n21410 = n6172 ^ n4445 ^ n2436 ;
  assign n21411 = x115 & ~n21410 ;
  assign n21412 = n21411 ^ n14716 ^ 1'b0 ;
  assign n21413 = n21412 ^ n1003 ^ 1'b0 ;
  assign n21414 = ~n947 & n21413 ;
  assign n21415 = n21414 ^ n6588 ^ n4585 ;
  assign n21417 = n5715 ^ n5475 ^ n2142 ;
  assign n21416 = ( ~n4804 & n5844 ) | ( ~n4804 & n17687 ) | ( n5844 & n17687 ) ;
  assign n21418 = n21417 ^ n21416 ^ 1'b0 ;
  assign n21419 = n19735 ^ n9845 ^ n7931 ;
  assign n21420 = n3462 ^ n2809 ^ n2131 ;
  assign n21421 = n16470 | n21420 ;
  assign n21422 = ( n2932 & n19900 ) | ( n2932 & n21421 ) | ( n19900 & n21421 ) ;
  assign n21423 = n21422 ^ n16879 ^ n8199 ;
  assign n21424 = n5364 ^ n2579 ^ n1243 ;
  assign n21426 = ( n3814 & n6430 ) | ( n3814 & ~n19171 ) | ( n6430 & ~n19171 ) ;
  assign n21425 = n1381 | n15123 ;
  assign n21427 = n21426 ^ n21425 ^ 1'b0 ;
  assign n21428 = ( ~n14822 & n21424 ) | ( ~n14822 & n21427 ) | ( n21424 & n21427 ) ;
  assign n21429 = n7083 & n8291 ;
  assign n21430 = n21429 ^ n11699 ^ 1'b0 ;
  assign n21431 = n18588 ^ n6272 ^ 1'b0 ;
  assign n21432 = n12763 & n21431 ;
  assign n21433 = ( n5006 & n18675 ) | ( n5006 & n20209 ) | ( n18675 & n20209 ) ;
  assign n21434 = n21433 ^ n20365 ^ n20170 ;
  assign n21435 = n14384 ^ n14242 ^ n7855 ;
  assign n21436 = n21435 ^ n13958 ^ 1'b0 ;
  assign n21437 = n6739 | n21436 ;
  assign n21438 = n21437 ^ n2140 ^ 1'b0 ;
  assign n21439 = ( x117 & n7001 ) | ( x117 & ~n10802 ) | ( n7001 & ~n10802 ) ;
  assign n21440 = n12892 ^ n10536 ^ 1'b0 ;
  assign n21441 = n10315 | n18942 ;
  assign n21442 = n21441 ^ n16642 ^ 1'b0 ;
  assign n21443 = ( n5062 & n9397 ) | ( n5062 & ~n14078 ) | ( n9397 & ~n14078 ) ;
  assign n21444 = n12597 ^ n10818 ^ n670 ;
  assign n21445 = ( n4075 & n12364 ) | ( n4075 & ~n17080 ) | ( n12364 & ~n17080 ) ;
  assign n21446 = n4764 | n21445 ;
  assign n21447 = n9563 ^ n8701 ^ n4031 ;
  assign n21448 = n3713 | n14364 ;
  assign n21449 = n21448 ^ x94 ^ 1'b0 ;
  assign n21450 = ( n9137 & n21447 ) | ( n9137 & n21449 ) | ( n21447 & n21449 ) ;
  assign n21451 = ( n633 & ~n6412 ) | ( n633 & n21450 ) | ( ~n6412 & n21450 ) ;
  assign n21452 = n15614 | n17012 ;
  assign n21453 = ( n1284 & n4838 ) | ( n1284 & ~n5948 ) | ( n4838 & ~n5948 ) ;
  assign n21454 = n21453 ^ n13548 ^ n5987 ;
  assign n21455 = n5104 ^ n1166 ^ 1'b0 ;
  assign n21456 = n21455 ^ n14296 ^ n5031 ;
  assign n21457 = n21456 ^ n10454 ^ n730 ;
  assign n21458 = ( ~n13763 & n17640 ) | ( ~n13763 & n17742 ) | ( n17640 & n17742 ) ;
  assign n21459 = ( ~n8935 & n9167 ) | ( ~n8935 & n21458 ) | ( n9167 & n21458 ) ;
  assign n21460 = n6757 | n21459 ;
  assign n21461 = n21457 & ~n21460 ;
  assign n21462 = n1388 ^ n894 ^ 1'b0 ;
  assign n21463 = n8774 ^ n2327 ^ 1'b0 ;
  assign n21464 = x26 & n21463 ;
  assign n21465 = n21464 ^ n14454 ^ 1'b0 ;
  assign n21466 = n8713 | n21465 ;
  assign n21467 = n6096 & n21466 ;
  assign n21468 = n21462 & ~n21467 ;
  assign n21469 = ~n10127 & n21468 ;
  assign n21471 = ( n2390 & n7604 ) | ( n2390 & n11840 ) | ( n7604 & n11840 ) ;
  assign n21470 = n10983 ^ n10262 ^ x86 ;
  assign n21472 = n21471 ^ n21470 ^ 1'b0 ;
  assign n21473 = ~n21469 & n21472 ;
  assign n21474 = n13113 ^ n9564 ^ n9092 ;
  assign n21475 = n11885 ^ n1440 ^ n702 ;
  assign n21476 = ( n16762 & ~n19600 ) | ( n16762 & n21475 ) | ( ~n19600 & n21475 ) ;
  assign n21477 = n8199 ^ n1710 ^ n878 ;
  assign n21478 = ( ~n390 & n8878 ) | ( ~n390 & n10650 ) | ( n8878 & n10650 ) ;
  assign n21479 = ( n4021 & ~n7641 ) | ( n4021 & n8035 ) | ( ~n7641 & n8035 ) ;
  assign n21480 = n18899 ^ n3668 ^ 1'b0 ;
  assign n21481 = ~n7687 & n21480 ;
  assign n21484 = n10054 ^ n6097 ^ n934 ;
  assign n21482 = ( ~n4323 & n5922 ) | ( ~n4323 & n18045 ) | ( n5922 & n18045 ) ;
  assign n21483 = n7999 | n21482 ;
  assign n21485 = n21484 ^ n21483 ^ 1'b0 ;
  assign n21488 = n7021 ^ n1659 ^ n1215 ;
  assign n21489 = n4668 ^ n1294 ^ 1'b0 ;
  assign n21490 = n11084 ^ n9025 ^ n1984 ;
  assign n21491 = ( n14901 & n21489 ) | ( n14901 & ~n21490 ) | ( n21489 & ~n21490 ) ;
  assign n21492 = n21488 & n21491 ;
  assign n21493 = n21492 ^ n8856 ^ 1'b0 ;
  assign n21486 = n12368 ^ n1765 ^ 1'b0 ;
  assign n21487 = n21486 ^ n10749 ^ n2570 ;
  assign n21494 = n21493 ^ n21487 ^ n1744 ;
  assign n21495 = n14382 ^ n13058 ^ n11333 ;
  assign n21496 = ( n2189 & n5668 ) | ( n2189 & n21495 ) | ( n5668 & n21495 ) ;
  assign n21497 = n17764 ^ n11604 ^ n6378 ;
  assign n21498 = n21497 ^ n4425 ^ n1944 ;
  assign n21499 = n5262 & ~n15340 ;
  assign n21500 = n3622 & n21499 ;
  assign n21501 = n15898 ^ n15033 ^ n276 ;
  assign n21502 = n17576 ^ n16185 ^ n14244 ;
  assign n21503 = n5465 ^ n1367 ^ n314 ;
  assign n21504 = ( n9378 & n21502 ) | ( n9378 & ~n21503 ) | ( n21502 & ~n21503 ) ;
  assign n21505 = ( ~n2438 & n8986 ) | ( ~n2438 & n16105 ) | ( n8986 & n16105 ) ;
  assign n21506 = n19093 ^ n15121 ^ n9810 ;
  assign n21507 = n21506 ^ n16874 ^ 1'b0 ;
  assign n21508 = n18273 ^ n10158 ^ n9023 ;
  assign n21509 = ( n1252 & n7914 ) | ( n1252 & n21508 ) | ( n7914 & n21508 ) ;
  assign n21510 = n21509 ^ n1678 ^ 1'b0 ;
  assign n21511 = n5068 & ~n21510 ;
  assign n21512 = n21511 ^ n10881 ^ 1'b0 ;
  assign n21513 = n1701 & ~n9757 ;
  assign n21514 = n17257 & ~n21513 ;
  assign n21515 = n20964 & n21514 ;
  assign n21516 = n6073 ^ n5748 ^ 1'b0 ;
  assign n21517 = n18460 ^ n5730 ^ n5063 ;
  assign n21518 = ( n13156 & n21516 ) | ( n13156 & ~n21517 ) | ( n21516 & ~n21517 ) ;
  assign n21519 = n6285 | n10467 ;
  assign n21524 = n10693 ^ n4816 ^ n793 ;
  assign n21520 = n2110 | n13463 ;
  assign n21521 = n9477 & ~n21520 ;
  assign n21522 = x113 & ~n21521 ;
  assign n21523 = n21522 ^ n1588 ^ 1'b0 ;
  assign n21525 = n21524 ^ n21523 ^ n12075 ;
  assign n21526 = ( n469 & n21519 ) | ( n469 & ~n21525 ) | ( n21519 & ~n21525 ) ;
  assign n21527 = ( x50 & n4277 ) | ( x50 & ~n7842 ) | ( n4277 & ~n7842 ) ;
  assign n21528 = ( ~n2792 & n3798 ) | ( ~n2792 & n6766 ) | ( n3798 & n6766 ) ;
  assign n21529 = n21528 ^ n7730 ^ n6956 ;
  assign n21530 = n18943 ^ n10606 ^ n3968 ;
  assign n21531 = n13827 ^ n7873 ^ n4948 ;
  assign n21532 = ( ~n5498 & n11894 ) | ( ~n5498 & n21531 ) | ( n11894 & n21531 ) ;
  assign n21533 = n21532 ^ n17074 ^ n3191 ;
  assign n21534 = ( n13935 & n17725 ) | ( n13935 & n19624 ) | ( n17725 & n19624 ) ;
  assign n21535 = n16505 ^ n7266 ^ n5713 ;
  assign n21536 = n21535 ^ n4378 ^ n4275 ;
  assign n21537 = ( ~n16680 & n18130 ) | ( ~n16680 & n21536 ) | ( n18130 & n21536 ) ;
  assign n21538 = n16541 ^ n8122 ^ n7249 ;
  assign n21539 = ( ~n3117 & n6963 ) | ( ~n3117 & n21538 ) | ( n6963 & n21538 ) ;
  assign n21540 = n7300 | n21539 ;
  assign n21541 = n5601 | n21540 ;
  assign n21542 = n2405 & ~n2726 ;
  assign n21543 = n18957 | n21542 ;
  assign n21544 = n21543 ^ n13610 ^ 1'b0 ;
  assign n21545 = n21199 ^ n9221 ^ 1'b0 ;
  assign n21546 = n17930 ^ n8300 ^ n3461 ;
  assign n21547 = ( n10581 & n16316 ) | ( n10581 & ~n21495 ) | ( n16316 & ~n21495 ) ;
  assign n21548 = ( ~n1317 & n15326 ) | ( ~n1317 & n18545 ) | ( n15326 & n18545 ) ;
  assign n21549 = ( n2041 & n21528 ) | ( n2041 & n21548 ) | ( n21528 & n21548 ) ;
  assign n21550 = n8743 ^ n4494 ^ 1'b0 ;
  assign n21551 = n21550 ^ n20813 ^ n10013 ;
  assign n21552 = n13184 ^ n2983 ^ n2009 ;
  assign n21553 = ( n4553 & n7098 ) | ( n4553 & ~n21552 ) | ( n7098 & ~n21552 ) ;
  assign n21554 = ( n6809 & n13620 ) | ( n6809 & ~n21553 ) | ( n13620 & ~n21553 ) ;
  assign n21555 = n14444 ^ n10181 ^ n8403 ;
  assign n21556 = n7397 ^ n1745 ^ 1'b0 ;
  assign n21557 = n21555 & n21556 ;
  assign n21558 = ( n6325 & n8308 ) | ( n6325 & n21557 ) | ( n8308 & n21557 ) ;
  assign n21559 = n4025 ^ n3870 ^ n3422 ;
  assign n21560 = n21559 ^ n8199 ^ n3588 ;
  assign n21561 = ( n10424 & n16071 ) | ( n10424 & ~n21560 ) | ( n16071 & ~n21560 ) ;
  assign n21562 = n21561 ^ n18884 ^ n15012 ;
  assign n21563 = ~n7022 & n15689 ;
  assign n21564 = n4876 & n10575 ;
  assign n21565 = ( n7581 & n21563 ) | ( n7581 & ~n21564 ) | ( n21563 & ~n21564 ) ;
  assign n21566 = n10238 ^ n7323 ^ n506 ;
  assign n21567 = n5493 ^ n263 ^ 1'b0 ;
  assign n21568 = n21567 ^ n6098 ^ n4911 ;
  assign n21569 = n21568 ^ n20871 ^ n11394 ;
  assign n21570 = n4723 & n14302 ;
  assign n21571 = ~n2528 & n21570 ;
  assign n21573 = n5934 | n10760 ;
  assign n21574 = n6021 | n21573 ;
  assign n21572 = ( ~n252 & n9548 ) | ( ~n252 & n9670 ) | ( n9548 & n9670 ) ;
  assign n21575 = n21574 ^ n21572 ^ n12357 ;
  assign n21576 = n10143 ^ n8355 ^ n543 ;
  assign n21577 = n14045 ^ n753 ^ n212 ;
  assign n21578 = n9272 ^ n8156 ^ 1'b0 ;
  assign n21579 = n12939 ^ n9760 ^ n6411 ;
  assign n21580 = n21579 ^ n7560 ^ n6218 ;
  assign n21581 = n12026 ^ n7618 ^ n683 ;
  assign n21582 = ( n4294 & ~n21122 ) | ( n4294 & n21581 ) | ( ~n21122 & n21581 ) ;
  assign n21583 = n12167 ^ n12098 ^ x64 ;
  assign n21584 = ( ~n5477 & n8863 ) | ( ~n5477 & n21583 ) | ( n8863 & n21583 ) ;
  assign n21585 = ( ~n16283 & n21582 ) | ( ~n16283 & n21584 ) | ( n21582 & n21584 ) ;
  assign n21586 = n21585 ^ n11258 ^ 1'b0 ;
  assign n21587 = n5049 & ~n16746 ;
  assign n21588 = n21587 ^ n3651 ^ 1'b0 ;
  assign n21601 = ( n1898 & n2038 ) | ( n1898 & ~n3115 ) | ( n2038 & ~n3115 ) ;
  assign n21589 = n21453 ^ n13731 ^ n10572 ;
  assign n21595 = n5273 & ~n7319 ;
  assign n21596 = n21595 ^ n20196 ^ n15780 ;
  assign n21597 = n21596 ^ n9254 ^ 1'b0 ;
  assign n21598 = n21597 ^ n10526 ^ n4410 ;
  assign n21590 = ~n4463 & n11648 ;
  assign n21591 = n21590 ^ n2299 ^ 1'b0 ;
  assign n21592 = ( n7119 & n9189 ) | ( n7119 & n21591 ) | ( n9189 & n21591 ) ;
  assign n21593 = n17911 ^ n15409 ^ 1'b0 ;
  assign n21594 = n21592 & n21593 ;
  assign n21599 = n21598 ^ n21594 ^ 1'b0 ;
  assign n21600 = n21589 & n21599 ;
  assign n21602 = n21601 ^ n21600 ^ n6456 ;
  assign n21606 = ( n1766 & ~n4691 ) | ( n1766 & n6808 ) | ( ~n4691 & n6808 ) ;
  assign n21603 = n12342 ^ n5174 ^ n4041 ;
  assign n21604 = ~n17742 & n21603 ;
  assign n21605 = ~n4419 & n21604 ;
  assign n21607 = n21606 ^ n21605 ^ n19796 ;
  assign n21608 = ~n8588 & n19490 ;
  assign n21609 = n19228 ^ n8737 ^ n1588 ;
  assign n21610 = ( n2976 & n8898 ) | ( n2976 & n21609 ) | ( n8898 & n21609 ) ;
  assign n21611 = n21610 ^ n13833 ^ n417 ;
  assign n21612 = ( n17740 & n20424 ) | ( n17740 & ~n21611 ) | ( n20424 & ~n21611 ) ;
  assign n21613 = ( n11356 & n16241 ) | ( n11356 & n18867 ) | ( n16241 & n18867 ) ;
  assign n21614 = n13385 & ~n17755 ;
  assign n21615 = n7441 ^ n3268 ^ 1'b0 ;
  assign n21616 = ~n19225 & n21615 ;
  assign n21617 = n4730 ^ n2943 ^ n1078 ;
  assign n21618 = ~n11271 & n21617 ;
  assign n21619 = n12293 ^ n3093 ^ n1872 ;
  assign n21620 = ( n2165 & n10231 ) | ( n2165 & n21619 ) | ( n10231 & n21619 ) ;
  assign n21624 = n4320 ^ n4107 ^ 1'b0 ;
  assign n21625 = n12336 & n21624 ;
  assign n21626 = ( n7678 & n15486 ) | ( n7678 & n21625 ) | ( n15486 & n21625 ) ;
  assign n21621 = n12742 | n16782 ;
  assign n21622 = n21621 ^ n3177 ^ 1'b0 ;
  assign n21623 = n15458 & ~n21622 ;
  assign n21627 = n21626 ^ n21623 ^ 1'b0 ;
  assign n21628 = n21627 ^ n20280 ^ 1'b0 ;
  assign n21629 = n9474 ^ n9064 ^ n9035 ;
  assign n21630 = n648 & n21629 ;
  assign n21631 = n10303 ^ n1639 ^ 1'b0 ;
  assign n21632 = n8413 & n21631 ;
  assign n21633 = n4223 & ~n21632 ;
  assign n21634 = n21633 ^ n18838 ^ 1'b0 ;
  assign n21635 = n3316 | n16776 ;
  assign n21636 = n14213 | n21635 ;
  assign n21637 = ~n20580 & n21636 ;
  assign n21638 = n21637 ^ n19582 ^ 1'b0 ;
  assign n21641 = n7582 ^ n1136 ^ x105 ;
  assign n21642 = n21641 ^ n13334 ^ n830 ;
  assign n21639 = n9544 ^ n5860 ^ 1'b0 ;
  assign n21640 = ~n15010 & n21639 ;
  assign n21643 = n21642 ^ n21640 ^ n19250 ;
  assign n21644 = n17715 ^ n4175 ^ n4092 ;
  assign n21646 = x89 & ~n9022 ;
  assign n21647 = n21646 ^ n8484 ^ 1'b0 ;
  assign n21648 = n21647 ^ n8831 ^ n2676 ;
  assign n21645 = ( n263 & n399 ) | ( n263 & n16634 ) | ( n399 & n16634 ) ;
  assign n21649 = n21648 ^ n21645 ^ n15704 ;
  assign n21650 = ~n21644 & n21649 ;
  assign n21651 = ~n1612 & n21467 ;
  assign n21652 = ( ~n8895 & n9198 ) | ( ~n8895 & n15759 ) | ( n9198 & n15759 ) ;
  assign n21653 = n11827 ^ n5447 ^ 1'b0 ;
  assign n21654 = n21653 ^ n876 ^ 1'b0 ;
  assign n21655 = ~n254 & n21654 ;
  assign n21656 = n8810 ^ n4651 ^ 1'b0 ;
  assign n21657 = ( n5268 & n6291 ) | ( n5268 & n21656 ) | ( n6291 & n21656 ) ;
  assign n21658 = n21657 ^ n16127 ^ 1'b0 ;
  assign n21659 = n5160 & ~n21658 ;
  assign n21660 = n19623 ^ n18297 ^ n12854 ;
  assign n21661 = n14459 | n21660 ;
  assign n21662 = n21659 | n21661 ;
  assign n21667 = n4841 ^ n1417 ^ n834 ;
  assign n21668 = n14308 ^ n7348 ^ 1'b0 ;
  assign n21669 = n21667 & n21668 ;
  assign n21664 = ( n1949 & ~n4071 ) | ( n1949 & n20936 ) | ( ~n4071 & n20936 ) ;
  assign n21663 = ( n7453 & ~n8154 ) | ( n7453 & n19051 ) | ( ~n8154 & n19051 ) ;
  assign n21665 = n21664 ^ n21663 ^ n10772 ;
  assign n21666 = n6731 & ~n21665 ;
  assign n21670 = n21669 ^ n21666 ^ 1'b0 ;
  assign n21671 = n4168 ^ n3655 ^ n2861 ;
  assign n21672 = ( n2147 & n17500 ) | ( n2147 & ~n21671 ) | ( n17500 & ~n21671 ) ;
  assign n21673 = n12438 ^ n5761 ^ n4560 ;
  assign n21674 = ~n2850 & n19392 ;
  assign n21675 = n9920 & n21674 ;
  assign n21676 = n15446 ^ n15148 ^ 1'b0 ;
  assign n21677 = ~n9839 & n21676 ;
  assign n21678 = ( n5652 & ~n21675 ) | ( n5652 & n21677 ) | ( ~n21675 & n21677 ) ;
  assign n21679 = n375 & n16427 ;
  assign n21680 = n9816 | n13072 ;
  assign n21681 = n21680 ^ n1967 ^ 1'b0 ;
  assign n21682 = n10802 ^ n5365 ^ n2910 ;
  assign n21683 = ( n8875 & ~n9492 ) | ( n8875 & n21682 ) | ( ~n9492 & n21682 ) ;
  assign n21684 = n1550 & ~n18654 ;
  assign n21685 = ~n21683 & n21684 ;
  assign n21686 = n4139 & ~n21685 ;
  assign n21687 = ( n19394 & n21681 ) | ( n19394 & n21686 ) | ( n21681 & n21686 ) ;
  assign n21688 = ( n844 & ~n5101 ) | ( n844 & n10765 ) | ( ~n5101 & n10765 ) ;
  assign n21689 = ( n8146 & n8731 ) | ( n8146 & ~n11979 ) | ( n8731 & ~n11979 ) ;
  assign n21690 = ( n12051 & n21688 ) | ( n12051 & n21689 ) | ( n21688 & n21689 ) ;
  assign n21691 = n21690 ^ n11280 ^ n10562 ;
  assign n21695 = ( ~n3137 & n10632 ) | ( ~n3137 & n11677 ) | ( n10632 & n11677 ) ;
  assign n21692 = n3441 ^ n743 ^ n471 ;
  assign n21693 = ( ~n1794 & n11778 ) | ( ~n1794 & n21692 ) | ( n11778 & n21692 ) ;
  assign n21694 = ~n16041 & n21693 ;
  assign n21696 = n21695 ^ n21694 ^ 1'b0 ;
  assign n21697 = ~n8651 & n13050 ;
  assign n21698 = n21697 ^ n1166 ^ 1'b0 ;
  assign n21699 = n21698 ^ n7245 ^ 1'b0 ;
  assign n21700 = n7392 | n21699 ;
  assign n21701 = ~n20442 & n21700 ;
  assign n21702 = n9327 & ~n11825 ;
  assign n21703 = n21702 ^ n5266 ^ 1'b0 ;
  assign n21704 = ~n5873 & n14869 ;
  assign n21706 = n11415 ^ n6337 ^ n1539 ;
  assign n21705 = n5909 ^ n2287 ^ n940 ;
  assign n21707 = n21706 ^ n21705 ^ n689 ;
  assign n21708 = ( n8670 & ~n15349 ) | ( n8670 & n16745 ) | ( ~n15349 & n16745 ) ;
  assign n21709 = n21708 ^ n14751 ^ n12968 ;
  assign n21710 = n12366 ^ n9288 ^ n7660 ;
  assign n21712 = n16391 ^ n13018 ^ n1103 ;
  assign n21711 = n17240 ^ n12125 ^ n4788 ;
  assign n21713 = n21712 ^ n21711 ^ n2971 ;
  assign n21714 = n13603 ^ n10195 ^ 1'b0 ;
  assign n21715 = n20202 ^ n18956 ^ n14143 ;
  assign n21716 = n8613 ^ n8211 ^ n4303 ;
  assign n21717 = ( n2055 & n20863 ) | ( n2055 & ~n21716 ) | ( n20863 & ~n21716 ) ;
  assign n21718 = n4296 & ~n17594 ;
  assign n21719 = n21718 ^ n16341 ^ 1'b0 ;
  assign n21720 = n21719 ^ n11770 ^ n605 ;
  assign n21721 = n14829 ^ n8755 ^ n8710 ;
  assign n21722 = ( ~x104 & n10036 ) | ( ~x104 & n21721 ) | ( n10036 & n21721 ) ;
  assign n21723 = n3005 & ~n21722 ;
  assign n21724 = ~n10339 & n21723 ;
  assign n21726 = ( n6928 & n7620 ) | ( n6928 & ~n12367 ) | ( n7620 & ~n12367 ) ;
  assign n21727 = n21726 ^ n12947 ^ n1649 ;
  assign n21725 = n1572 & n9566 ;
  assign n21728 = n21727 ^ n21725 ^ 1'b0 ;
  assign n21729 = ( n896 & n5202 ) | ( n896 & n6550 ) | ( n5202 & n6550 ) ;
  assign n21730 = n3253 ^ n1966 ^ 1'b0 ;
  assign n21731 = ( n4723 & n7810 ) | ( n4723 & ~n20756 ) | ( n7810 & ~n20756 ) ;
  assign n21732 = n21731 ^ n1644 ^ 1'b0 ;
  assign n21733 = n21730 & ~n21732 ;
  assign n21734 = n21733 ^ n10097 ^ 1'b0 ;
  assign n21735 = ( n6762 & n18437 ) | ( n6762 & ~n21734 ) | ( n18437 & ~n21734 ) ;
  assign n21736 = ( ~n8212 & n10885 ) | ( ~n8212 & n14856 ) | ( n10885 & n14856 ) ;
  assign n21737 = ( ~n7769 & n8593 ) | ( ~n7769 & n12364 ) | ( n8593 & n12364 ) ;
  assign n21738 = n21737 ^ n18595 ^ 1'b0 ;
  assign n21739 = ( n4544 & ~n17504 ) | ( n4544 & n21738 ) | ( ~n17504 & n21738 ) ;
  assign n21740 = n2625 & n21739 ;
  assign n21741 = n21736 & n21740 ;
  assign n21742 = n21741 ^ n4577 ^ 1'b0 ;
  assign n21743 = ( ~n1549 & n8242 ) | ( ~n1549 & n12313 ) | ( n8242 & n12313 ) ;
  assign n21744 = n21743 ^ n12126 ^ 1'b0 ;
  assign n21745 = n14686 ^ n4171 ^ n4150 ;
  assign n21746 = n21745 ^ n13213 ^ 1'b0 ;
  assign n21747 = ( ~n5491 & n21610 ) | ( ~n5491 & n21746 ) | ( n21610 & n21746 ) ;
  assign n21748 = n21747 ^ n1871 ^ n1648 ;
  assign n21749 = n21748 ^ n13636 ^ n4109 ;
  assign n21750 = ( n459 & ~n5657 ) | ( n459 & n7345 ) | ( ~n5657 & n7345 ) ;
  assign n21751 = n21750 ^ n11011 ^ 1'b0 ;
  assign n21752 = ~n19629 & n21751 ;
  assign n21753 = n21752 ^ n8658 ^ 1'b0 ;
  assign n21754 = n14122 ^ n13437 ^ n1007 ;
  assign n21755 = n21754 ^ n14591 ^ n636 ;
  assign n21756 = n14687 ^ n1852 ^ 1'b0 ;
  assign n21757 = n21756 ^ n7872 ^ 1'b0 ;
  assign n21758 = ( n5610 & n20865 ) | ( n5610 & n21757 ) | ( n20865 & n21757 ) ;
  assign n21759 = ~n4160 & n7096 ;
  assign n21760 = n21759 ^ n4423 ^ 1'b0 ;
  assign n21761 = n21760 ^ n14032 ^ x20 ;
  assign n21762 = ( n5280 & n11980 ) | ( n5280 & n21761 ) | ( n11980 & n21761 ) ;
  assign n21763 = n21762 ^ n17828 ^ n586 ;
  assign n21764 = ( ~n218 & n2428 ) | ( ~n218 & n2879 ) | ( n2428 & n2879 ) ;
  assign n21765 = ( ~n10244 & n11162 ) | ( ~n10244 & n19426 ) | ( n11162 & n19426 ) ;
  assign n21766 = n21764 | n21765 ;
  assign n21767 = ( n4351 & n9810 ) | ( n4351 & ~n21375 ) | ( n9810 & ~n21375 ) ;
  assign n21768 = n21767 ^ n8985 ^ n1498 ;
  assign n21769 = n14310 | n21768 ;
  assign n21770 = n21766 | n21769 ;
  assign n21771 = n21770 ^ n19549 ^ n2891 ;
  assign n21772 = n10030 | n17943 ;
  assign n21773 = n7077 ^ n7059 ^ 1'b0 ;
  assign n21774 = n21773 ^ n11916 ^ n3115 ;
  assign n21775 = n15146 ^ n8963 ^ n4979 ;
  assign n21776 = ~n7419 & n21775 ;
  assign n21777 = n5849 | n21776 ;
  assign n21778 = n18234 ^ n12125 ^ 1'b0 ;
  assign n21779 = n21778 ^ n14989 ^ n6409 ;
  assign n21780 = n13191 ^ n7139 ^ 1'b0 ;
  assign n21781 = ( n2804 & n5484 ) | ( n2804 & n6228 ) | ( n5484 & n6228 ) ;
  assign n21782 = n21781 ^ n2947 ^ n619 ;
  assign n21783 = ( ~n9757 & n11338 ) | ( ~n9757 & n21782 ) | ( n11338 & n21782 ) ;
  assign n21784 = n19392 ^ n5432 ^ 1'b0 ;
  assign n21785 = n21784 ^ n7613 ^ n4487 ;
  assign n21786 = ( n4439 & n10296 ) | ( n4439 & n21785 ) | ( n10296 & n21785 ) ;
  assign n21787 = n5260 ^ n3302 ^ 1'b0 ;
  assign n21788 = ( n3356 & n4975 ) | ( n3356 & n21787 ) | ( n4975 & n21787 ) ;
  assign n21789 = n9622 ^ n4153 ^ n3024 ;
  assign n21790 = ( n8033 & n21788 ) | ( n8033 & n21789 ) | ( n21788 & n21789 ) ;
  assign n21791 = n20769 ^ n20304 ^ 1'b0 ;
  assign n21792 = ~n21790 & n21791 ;
  assign n21793 = ( n8512 & n8679 ) | ( n8512 & n21631 ) | ( n8679 & n21631 ) ;
  assign n21794 = n5154 ^ n2230 ^ 1'b0 ;
  assign n21795 = n12312 & ~n21794 ;
  assign n21796 = n21795 ^ n16651 ^ n7905 ;
  assign n21797 = n21796 ^ n3615 ^ 1'b0 ;
  assign n21798 = n21793 & n21797 ;
  assign n21799 = n11359 ^ n5659 ^ n354 ;
  assign n21800 = ( n5513 & n18675 ) | ( n5513 & n21799 ) | ( n18675 & n21799 ) ;
  assign n21801 = n6319 & n21800 ;
  assign n21802 = n21801 ^ n18066 ^ n13143 ;
  assign n21803 = n1922 & n2163 ;
  assign n21804 = n21803 ^ n12775 ^ 1'b0 ;
  assign n21805 = n7848 | n21804 ;
  assign n21806 = n21805 ^ n21180 ^ n15924 ;
  assign n21807 = ( n160 & ~n5230 ) | ( n160 & n8428 ) | ( ~n5230 & n8428 ) ;
  assign n21808 = ( ~n4803 & n10790 ) | ( ~n4803 & n21807 ) | ( n10790 & n21807 ) ;
  assign n21809 = ( n1134 & ~n7133 ) | ( n1134 & n19684 ) | ( ~n7133 & n19684 ) ;
  assign n21810 = ( ~n7856 & n11503 ) | ( ~n7856 & n21809 ) | ( n11503 & n21809 ) ;
  assign n21811 = n11545 ^ n5929 ^ 1'b0 ;
  assign n21812 = n21811 ^ n10223 ^ n4352 ;
  assign n21813 = n15878 ^ n12809 ^ n1207 ;
  assign n21814 = n21813 ^ n15734 ^ 1'b0 ;
  assign n21815 = ~n11435 & n21814 ;
  assign n21816 = n3766 & ~n4828 ;
  assign n21817 = n9927 & n21816 ;
  assign n21818 = n7658 ^ n4070 ^ 1'b0 ;
  assign n21819 = n2749 & n21818 ;
  assign n21820 = n21819 ^ n4336 ^ n1141 ;
  assign n21826 = n13018 ^ n11415 ^ n2146 ;
  assign n21822 = ( n3644 & n3899 ) | ( n3644 & ~n6897 ) | ( n3899 & ~n6897 ) ;
  assign n21823 = ( n674 & ~n8003 ) | ( n674 & n21822 ) | ( ~n8003 & n21822 ) ;
  assign n21824 = n9850 ^ n8300 ^ n7493 ;
  assign n21825 = n21823 | n21824 ;
  assign n21821 = ( n944 & n2874 ) | ( n944 & ~n18097 ) | ( n2874 & ~n18097 ) ;
  assign n21827 = n21826 ^ n21825 ^ n21821 ;
  assign n21828 = n13517 ^ n8803 ^ n3267 ;
  assign n21829 = n21828 ^ n10722 ^ 1'b0 ;
  assign n21830 = ( ~n7486 & n11407 ) | ( ~n7486 & n21829 ) | ( n11407 & n21829 ) ;
  assign n21832 = n21641 ^ n15516 ^ n13661 ;
  assign n21831 = n14070 ^ n959 ^ n855 ;
  assign n21833 = n21832 ^ n21831 ^ n14653 ;
  assign n21835 = n3909 | n4479 ;
  assign n21836 = n2145 | n21835 ;
  assign n21837 = n21836 ^ n4216 ^ 1'b0 ;
  assign n21834 = n508 | n9506 ;
  assign n21838 = n21837 ^ n21834 ^ 1'b0 ;
  assign n21839 = ~n4008 & n10353 ;
  assign n21840 = n21839 ^ n3331 ^ 1'b0 ;
  assign n21841 = n19366 ^ n15922 ^ n15214 ;
  assign n21842 = n11655 ^ n9819 ^ n7840 ;
  assign n21845 = n496 & ~n1004 ;
  assign n21846 = ~n588 & n21845 ;
  assign n21843 = ( n19761 & n20365 ) | ( n19761 & ~n21553 ) | ( n20365 & ~n21553 ) ;
  assign n21844 = ( n237 & n10059 ) | ( n237 & n21843 ) | ( n10059 & n21843 ) ;
  assign n21847 = n21846 ^ n21844 ^ n5984 ;
  assign n21849 = ( x105 & n261 ) | ( x105 & ~n1801 ) | ( n261 & ~n1801 ) ;
  assign n21848 = ( n7726 & ~n11071 ) | ( n7726 & n17003 ) | ( ~n11071 & n17003 ) ;
  assign n21850 = n21849 ^ n21848 ^ 1'b0 ;
  assign n21851 = ( n206 & n4941 ) | ( n206 & n17050 ) | ( n4941 & n17050 ) ;
  assign n21852 = n18527 ^ n5344 ^ 1'b0 ;
  assign n21853 = ( n13003 & n19900 ) | ( n13003 & n21852 ) | ( n19900 & n21852 ) ;
  assign n21854 = n21851 & ~n21853 ;
  assign n21855 = ( n2757 & n7260 ) | ( n2757 & ~n21854 ) | ( n7260 & ~n21854 ) ;
  assign n21856 = n8319 ^ x119 ^ 1'b0 ;
  assign n21857 = n11182 & n14545 ;
  assign n21858 = ~n20792 & n21857 ;
  assign n21859 = ~n10729 & n21858 ;
  assign n21860 = ( n1032 & n21856 ) | ( n1032 & n21859 ) | ( n21856 & n21859 ) ;
  assign n21861 = n18039 ^ n15813 ^ n7703 ;
  assign n21862 = ( n11612 & n14391 ) | ( n11612 & n21861 ) | ( n14391 & n21861 ) ;
  assign n21863 = n19752 & n20167 ;
  assign n21864 = n21863 ^ n1557 ^ 1'b0 ;
  assign n21865 = ( ~n8963 & n14428 ) | ( ~n8963 & n19154 ) | ( n14428 & n19154 ) ;
  assign n21866 = n19311 ^ n17764 ^ n8989 ;
  assign n21867 = ( n18001 & n21865 ) | ( n18001 & n21866 ) | ( n21865 & n21866 ) ;
  assign n21868 = n21867 ^ n15860 ^ n10843 ;
  assign n21869 = ~n12361 & n21868 ;
  assign n21870 = n1805 & n21869 ;
  assign n21871 = n1887 ^ n1245 ^ n1134 ;
  assign n21872 = ( n10241 & n15452 ) | ( n10241 & n21871 ) | ( n15452 & n21871 ) ;
  assign n21873 = n155 & ~n15335 ;
  assign n21874 = n21873 ^ n7513 ^ 1'b0 ;
  assign n21875 = ( ~n6386 & n21872 ) | ( ~n6386 & n21874 ) | ( n21872 & n21874 ) ;
  assign n21876 = ( n5967 & n13710 ) | ( n5967 & n16471 ) | ( n13710 & n16471 ) ;
  assign n21877 = n11011 ^ n5886 ^ 1'b0 ;
  assign n21878 = ( ~n3272 & n6793 ) | ( ~n3272 & n21877 ) | ( n6793 & n21877 ) ;
  assign n21879 = n11845 ^ n7928 ^ n6688 ;
  assign n21880 = n21879 ^ n18208 ^ n2267 ;
  assign n21881 = ( n5077 & n19284 ) | ( n5077 & n21880 ) | ( n19284 & n21880 ) ;
  assign n21882 = n8849 ^ n2405 ^ n1654 ;
  assign n21883 = ( n15059 & n15292 ) | ( n15059 & n21882 ) | ( n15292 & n21882 ) ;
  assign n21884 = n13588 ^ n13515 ^ n2973 ;
  assign n21885 = ( n2886 & n6785 ) | ( n2886 & ~n15467 ) | ( n6785 & ~n15467 ) ;
  assign n21886 = n2978 & n9354 ;
  assign n21887 = ~n13666 & n21886 ;
  assign n21888 = n10884 | n19591 ;
  assign n21889 = n7008 | n21888 ;
  assign n21890 = ( ~n8582 & n21887 ) | ( ~n8582 & n21889 ) | ( n21887 & n21889 ) ;
  assign n21891 = n9439 ^ n9354 ^ n1400 ;
  assign n21892 = ( n2330 & n7354 ) | ( n2330 & ~n16367 ) | ( n7354 & ~n16367 ) ;
  assign n21893 = n21892 ^ n19832 ^ 1'b0 ;
  assign n21894 = ( n816 & n1602 ) | ( n816 & n16993 ) | ( n1602 & n16993 ) ;
  assign n21895 = n1883 | n21894 ;
  assign n21896 = ( n17207 & ~n19857 ) | ( n17207 & n21895 ) | ( ~n19857 & n21895 ) ;
  assign n21897 = n2598 | n10925 ;
  assign n21898 = n21897 ^ n19437 ^ 1'b0 ;
  assign n21899 = n2037 ^ n1550 ^ 1'b0 ;
  assign n21900 = n12852 & n21899 ;
  assign n21901 = n18665 ^ n14432 ^ n14403 ;
  assign n21902 = n21900 & n21901 ;
  assign n21903 = ~n5005 & n21902 ;
  assign n21904 = n1152 & n3186 ;
  assign n21905 = n21904 ^ n7478 ^ 1'b0 ;
  assign n21906 = ~n2905 & n5183 ;
  assign n21907 = n21906 ^ n10922 ^ n1491 ;
  assign n21908 = n15233 ^ n10449 ^ n2309 ;
  assign n21909 = ( ~n2507 & n5183 ) | ( ~n2507 & n21908 ) | ( n5183 & n21908 ) ;
  assign n21910 = n2555 & n18357 ;
  assign n21911 = n21910 ^ n19727 ^ n15638 ;
  assign n21912 = n11733 ^ n4111 ^ 1'b0 ;
  assign n21913 = n19412 & ~n21912 ;
  assign n21914 = n15759 ^ n4998 ^ 1'b0 ;
  assign n21915 = n10875 & n21914 ;
  assign n21916 = n14876 ^ n6889 ^ n4115 ;
  assign n21917 = ( n13062 & ~n15151 ) | ( n13062 & n17473 ) | ( ~n15151 & n17473 ) ;
  assign n21918 = n21917 ^ n12893 ^ n12277 ;
  assign n21919 = ( n1065 & n3484 ) | ( n1065 & n21918 ) | ( n3484 & n21918 ) ;
  assign n21920 = n4565 ^ n428 ^ 1'b0 ;
  assign n21921 = n5824 & n21920 ;
  assign n21922 = n21921 ^ n19264 ^ n9705 ;
  assign n21923 = n4595 & ~n15989 ;
  assign n21924 = ( n4511 & n5444 ) | ( n4511 & ~n21923 ) | ( n5444 & ~n21923 ) ;
  assign n21929 = ( ~n3186 & n11077 ) | ( ~n3186 & n14051 ) | ( n11077 & n14051 ) ;
  assign n21930 = n21929 ^ n17473 ^ n8909 ;
  assign n21931 = n21930 ^ n11486 ^ n1383 ;
  assign n21928 = ( n4540 & n9695 ) | ( n4540 & n17118 ) | ( n9695 & n17118 ) ;
  assign n21925 = n18184 ^ n13649 ^ n1095 ;
  assign n21926 = ~n10598 & n21925 ;
  assign n21927 = ~n10322 & n21926 ;
  assign n21932 = n21931 ^ n21928 ^ n21927 ;
  assign n21933 = ( n12139 & n21924 ) | ( n12139 & ~n21932 ) | ( n21924 & ~n21932 ) ;
  assign n21934 = n21854 ^ n13012 ^ n6228 ;
  assign n21937 = n13610 ^ n12797 ^ n10372 ;
  assign n21935 = ( n5624 & n8724 ) | ( n5624 & ~n16485 ) | ( n8724 & ~n16485 ) ;
  assign n21936 = n21935 ^ n9668 ^ n6052 ;
  assign n21938 = n21937 ^ n21936 ^ n8109 ;
  assign n21939 = n10579 ^ n5400 ^ n5043 ;
  assign n21940 = ( n1398 & n3931 ) | ( n1398 & n21939 ) | ( n3931 & n21939 ) ;
  assign n21941 = ( n718 & ~n17715 ) | ( n718 & n21940 ) | ( ~n17715 & n21940 ) ;
  assign n21942 = n4662 ^ n4290 ^ n3026 ;
  assign n21943 = n7323 & n19157 ;
  assign n21944 = ~n21942 & n21943 ;
  assign n21945 = n4017 & n7452 ;
  assign n21946 = n21945 ^ n11865 ^ 1'b0 ;
  assign n21947 = n11285 ^ n6918 ^ n3237 ;
  assign n21949 = n19889 ^ n7890 ^ n2732 ;
  assign n21948 = n263 & ~n15576 ;
  assign n21950 = n21949 ^ n21948 ^ n1356 ;
  assign n21951 = ( n5881 & n21947 ) | ( n5881 & ~n21950 ) | ( n21947 & ~n21950 ) ;
  assign n21952 = ( n1367 & n11035 ) | ( n1367 & n13416 ) | ( n11035 & n13416 ) ;
  assign n21953 = n21952 ^ n9957 ^ 1'b0 ;
  assign n21954 = n3378 & n13692 ;
  assign n21955 = n11814 & n21954 ;
  assign n21957 = ( n4179 & n5301 ) | ( n4179 & ~n12553 ) | ( n5301 & ~n12553 ) ;
  assign n21956 = n2043 & n13915 ;
  assign n21958 = n21957 ^ n21956 ^ n4642 ;
  assign n21959 = ~n16435 & n21958 ;
  assign n21960 = n10695 ^ n6302 ^ 1'b0 ;
  assign n21962 = n5263 ^ n1549 ^ n974 ;
  assign n21961 = n11759 ^ n5301 ^ 1'b0 ;
  assign n21963 = n21962 ^ n21961 ^ n6272 ;
  assign n21964 = n2771 | n14338 ;
  assign n21965 = n10073 | n21964 ;
  assign n21966 = n21965 ^ n6917 ^ n4463 ;
  assign n21967 = n21966 ^ n5556 ^ 1'b0 ;
  assign n21968 = ~n2727 & n21967 ;
  assign n21969 = n4155 & ~n19034 ;
  assign n21970 = ~n21968 & n21969 ;
  assign n21971 = ( n21960 & ~n21963 ) | ( n21960 & n21970 ) | ( ~n21963 & n21970 ) ;
  assign n21972 = n21959 & ~n21971 ;
  assign n21973 = ~n764 & n21972 ;
  assign n21974 = ~n2132 & n7954 ;
  assign n21975 = n4179 & n21974 ;
  assign n21976 = n11571 ^ n4532 ^ n4027 ;
  assign n21977 = ( n3713 & n12260 ) | ( n3713 & ~n21976 ) | ( n12260 & ~n21976 ) ;
  assign n21979 = n4160 ^ n2862 ^ n2813 ;
  assign n21978 = n7034 ^ n6519 ^ n6104 ;
  assign n21980 = n21979 ^ n21978 ^ n4986 ;
  assign n21981 = ( ~n6312 & n13168 ) | ( ~n6312 & n21980 ) | ( n13168 & n21980 ) ;
  assign n21982 = n18728 ^ n3190 ^ 1'b0 ;
  assign n21983 = n8868 & ~n21982 ;
  assign n21984 = n20571 ^ n20565 ^ 1'b0 ;
  assign n21985 = ( n8281 & n21983 ) | ( n8281 & ~n21984 ) | ( n21983 & ~n21984 ) ;
  assign n21986 = ( n1234 & n5677 ) | ( n1234 & ~n10597 ) | ( n5677 & ~n10597 ) ;
  assign n21987 = n5488 & n20188 ;
  assign n21988 = ( n6963 & n17411 ) | ( n6963 & ~n21516 ) | ( n17411 & ~n21516 ) ;
  assign n21989 = n21988 ^ n17220 ^ n14671 ;
  assign n21990 = n21989 ^ n6018 ^ n4622 ;
  assign n21991 = n10648 | n14570 ;
  assign n21992 = n21990 | n21991 ;
  assign n21993 = n16040 ^ n5429 ^ 1'b0 ;
  assign n21994 = ( ~n9620 & n11850 ) | ( ~n9620 & n21993 ) | ( n11850 & n21993 ) ;
  assign n21995 = n15240 ^ n3762 ^ n1918 ;
  assign n21996 = n19286 ^ n17256 ^ n4712 ;
  assign n21997 = ( n1563 & n20897 ) | ( n1563 & ~n21996 ) | ( n20897 & ~n21996 ) ;
  assign n21998 = ( n2327 & n2855 ) | ( n2327 & n8930 ) | ( n2855 & n8930 ) ;
  assign n21999 = ( n15175 & ~n17410 ) | ( n15175 & n21998 ) | ( ~n17410 & n21998 ) ;
  assign n22000 = n2876 ^ n2440 ^ 1'b0 ;
  assign n22001 = ~n3115 & n22000 ;
  assign n22002 = n22001 ^ n3233 ^ n2884 ;
  assign n22003 = n2153 | n22002 ;
  assign n22004 = n13473 ^ n7117 ^ 1'b0 ;
  assign n22005 = n8013 & n22004 ;
  assign n22006 = n22005 ^ n17034 ^ n4830 ;
  assign n22007 = ( n5382 & ~n7646 ) | ( n5382 & n10173 ) | ( ~n7646 & n10173 ) ;
  assign n22008 = ( ~n1741 & n12049 ) | ( ~n1741 & n22007 ) | ( n12049 & n22007 ) ;
  assign n22009 = n22008 ^ n13165 ^ n7168 ;
  assign n22010 = n9701 & ~n14652 ;
  assign n22011 = n22010 ^ n3495 ^ 1'b0 ;
  assign n22012 = n20459 ^ n15924 ^ n4087 ;
  assign n22013 = n12894 & n22012 ;
  assign n22014 = n18867 & n22013 ;
  assign n22015 = n22014 ^ n21663 ^ n12616 ;
  assign n22016 = ( n4218 & n5629 ) | ( n4218 & ~n7130 ) | ( n5629 & ~n7130 ) ;
  assign n22017 = ( n16473 & ~n18398 ) | ( n16473 & n22016 ) | ( ~n18398 & n22016 ) ;
  assign n22019 = n10649 ^ n6280 ^ n4714 ;
  assign n22020 = ( n3880 & n5692 ) | ( n3880 & ~n22019 ) | ( n5692 & ~n22019 ) ;
  assign n22018 = n14133 ^ n2973 ^ n1800 ;
  assign n22021 = n22020 ^ n22018 ^ n5096 ;
  assign n22022 = n22021 ^ n13620 ^ n6626 ;
  assign n22023 = ( ~n18631 & n22017 ) | ( ~n18631 & n22022 ) | ( n22017 & n22022 ) ;
  assign n22024 = n18119 ^ n15199 ^ n4377 ;
  assign n22025 = n22024 ^ n6433 ^ 1'b0 ;
  assign n22026 = ( n7816 & ~n20221 ) | ( n7816 & n22025 ) | ( ~n20221 & n22025 ) ;
  assign n22027 = n19299 ^ n6548 ^ n4863 ;
  assign n22028 = ( n1131 & ~n13509 ) | ( n1131 & n19104 ) | ( ~n13509 & n19104 ) ;
  assign n22029 = ( n5027 & ~n9069 ) | ( n5027 & n22028 ) | ( ~n9069 & n22028 ) ;
  assign n22030 = n22029 ^ n12091 ^ 1'b0 ;
  assign n22031 = n20428 ^ n9100 ^ n7644 ;
  assign n22032 = n16468 ^ n2006 ^ 1'b0 ;
  assign n22033 = n1368 & n22032 ;
  assign n22036 = n8107 ^ n7344 ^ n1469 ;
  assign n22034 = ( ~n1784 & n4059 ) | ( ~n1784 & n10640 ) | ( n4059 & n10640 ) ;
  assign n22035 = n22034 ^ n20244 ^ n15408 ;
  assign n22037 = n22036 ^ n22035 ^ n15455 ;
  assign n22038 = n9527 ^ n6872 ^ n3082 ;
  assign n22039 = ~n2602 & n13596 ;
  assign n22040 = ( n3373 & n13855 ) | ( n3373 & n22039 ) | ( n13855 & n22039 ) ;
  assign n22041 = ( n2631 & n3982 ) | ( n2631 & n4677 ) | ( n3982 & n4677 ) ;
  assign n22042 = n377 & ~n8256 ;
  assign n22043 = ~n15331 & n22042 ;
  assign n22044 = n22043 ^ n4587 ^ 1'b0 ;
  assign n22045 = n11451 & n22044 ;
  assign n22046 = n11330 ^ n7805 ^ n6114 ;
  assign n22047 = ( n4178 & n12437 ) | ( n4178 & n22046 ) | ( n12437 & n22046 ) ;
  assign n22048 = n955 & n1580 ;
  assign n22049 = ~n1820 & n22048 ;
  assign n22050 = n1325 | n7848 ;
  assign n22051 = n13814 | n22050 ;
  assign n22052 = ( ~n13636 & n22049 ) | ( ~n13636 & n22051 ) | ( n22049 & n22051 ) ;
  assign n22054 = ( n507 & ~n1009 ) | ( n507 & n5325 ) | ( ~n1009 & n5325 ) ;
  assign n22053 = n20949 ^ n7856 ^ 1'b0 ;
  assign n22055 = n22054 ^ n22053 ^ n6432 ;
  assign n22056 = ( ~n4032 & n5462 ) | ( ~n4032 & n8268 ) | ( n5462 & n8268 ) ;
  assign n22057 = n10349 & ~n22056 ;
  assign n22058 = ( n3668 & n22055 ) | ( n3668 & n22057 ) | ( n22055 & n22057 ) ;
  assign n22059 = n6370 ^ n5237 ^ 1'b0 ;
  assign n22060 = n22059 ^ n20984 ^ n11883 ;
  assign n22061 = n17592 ^ n9010 ^ 1'b0 ;
  assign n22062 = n6729 & n22061 ;
  assign n22063 = ( ~n10307 & n20467 ) | ( ~n10307 & n22062 ) | ( n20467 & n22062 ) ;
  assign n22064 = n13259 ^ n13226 ^ 1'b0 ;
  assign n22065 = n22063 | n22064 ;
  assign n22066 = n16367 ^ n10329 ^ 1'b0 ;
  assign n22067 = n1768 & n22066 ;
  assign n22068 = n18612 ^ n5088 ^ n4802 ;
  assign n22069 = ~n14105 & n18525 ;
  assign n22073 = n1749 & n14552 ;
  assign n22070 = ( n6107 & n7861 ) | ( n6107 & n16295 ) | ( n7861 & n16295 ) ;
  assign n22071 = n22070 ^ n15753 ^ n8552 ;
  assign n22072 = n22071 ^ n20916 ^ n19010 ;
  assign n22074 = n22073 ^ n22072 ^ n13778 ;
  assign n22075 = ( n10130 & ~n16911 ) | ( n10130 & n19084 ) | ( ~n16911 & n19084 ) ;
  assign n22076 = n22075 ^ n9354 ^ n7469 ;
  assign n22078 = ( n6824 & n16771 ) | ( n6824 & n21685 ) | ( n16771 & n21685 ) ;
  assign n22077 = n11618 | n12101 ;
  assign n22079 = n22078 ^ n22077 ^ n6233 ;
  assign n22081 = ( n3996 & ~n7605 ) | ( n3996 & n11021 ) | ( ~n7605 & n11021 ) ;
  assign n22080 = n10404 & n16310 ;
  assign n22082 = n22081 ^ n22080 ^ n2723 ;
  assign n22083 = ( n582 & n11394 ) | ( n582 & ~n22082 ) | ( n11394 & ~n22082 ) ;
  assign n22084 = ( n276 & n8868 ) | ( n276 & n12171 ) | ( n8868 & n12171 ) ;
  assign n22085 = n22084 ^ n4836 ^ n1591 ;
  assign n22086 = ( ~n5836 & n13948 ) | ( ~n5836 & n22085 ) | ( n13948 & n22085 ) ;
  assign n22087 = ( n3660 & ~n4439 ) | ( n3660 & n6072 ) | ( ~n4439 & n6072 ) ;
  assign n22088 = n20676 ^ n7645 ^ n4036 ;
  assign n22089 = n22088 ^ n1742 ^ 1'b0 ;
  assign n22090 = ~n22087 & n22089 ;
  assign n22091 = ( n3865 & n9887 ) | ( n3865 & ~n22090 ) | ( n9887 & ~n22090 ) ;
  assign n22092 = n20790 ^ n3750 ^ 1'b0 ;
  assign n22093 = ~n19521 & n22092 ;
  assign n22094 = n21450 ^ n13706 ^ 1'b0 ;
  assign n22096 = n16513 ^ n5038 ^ n2931 ;
  assign n22097 = n22096 ^ n9272 ^ 1'b0 ;
  assign n22095 = n7092 & ~n12563 ;
  assign n22098 = n22097 ^ n22095 ^ 1'b0 ;
  assign n22100 = n20227 ^ n6156 ^ n2446 ;
  assign n22101 = n14191 & ~n19481 ;
  assign n22102 = n22101 ^ n921 ^ 1'b0 ;
  assign n22103 = ( n9829 & ~n22100 ) | ( n9829 & n22102 ) | ( ~n22100 & n22102 ) ;
  assign n22099 = n18219 ^ n12592 ^ n4840 ;
  assign n22104 = n22103 ^ n22099 ^ n21936 ;
  assign n22105 = n17821 ^ n10751 ^ 1'b0 ;
  assign n22106 = ( ~n2728 & n6582 ) | ( ~n2728 & n12635 ) | ( n6582 & n12635 ) ;
  assign n22107 = n13196 | n19869 ;
  assign n22108 = n7605 & ~n22107 ;
  assign n22109 = n16754 ^ n8777 ^ n8750 ;
  assign n22111 = n8062 ^ n6188 ^ n1278 ;
  assign n22110 = ( ~n5118 & n7929 ) | ( ~n5118 & n11758 ) | ( n7929 & n11758 ) ;
  assign n22112 = n22111 ^ n22110 ^ 1'b0 ;
  assign n22113 = n22109 | n22112 ;
  assign n22114 = n18597 ^ n1278 ^ 1'b0 ;
  assign n22115 = ( n5571 & ~n5676 ) | ( n5571 & n18083 ) | ( ~n5676 & n18083 ) ;
  assign n22116 = n7620 ^ n5524 ^ n3228 ;
  assign n22119 = n16786 ^ n9851 ^ n1064 ;
  assign n22118 = n11867 ^ n6020 ^ x119 ;
  assign n22117 = n21828 ^ n12748 ^ n8207 ;
  assign n22120 = n22119 ^ n22118 ^ n22117 ;
  assign n22121 = n8127 ^ n2978 ^ n1328 ;
  assign n22122 = ( ~n366 & n8773 ) | ( ~n366 & n22121 ) | ( n8773 & n22121 ) ;
  assign n22123 = n7400 | n22122 ;
  assign n22124 = n16164 ^ n13748 ^ n2623 ;
  assign n22125 = n4387 | n22124 ;
  assign n22126 = n14160 | n22001 ;
  assign n22127 = ( n9893 & ~n22125 ) | ( n9893 & n22126 ) | ( ~n22125 & n22126 ) ;
  assign n22128 = ~n14379 & n22127 ;
  assign n22129 = ~n1381 & n16067 ;
  assign n22130 = ~n20902 & n22129 ;
  assign n22131 = ( n12101 & n18773 ) | ( n12101 & ~n22130 ) | ( n18773 & ~n22130 ) ;
  assign n22132 = n989 | n10781 ;
  assign n22133 = n22132 ^ n15097 ^ n12910 ;
  assign n22134 = ( n5552 & ~n17498 ) | ( n5552 & n21535 ) | ( ~n17498 & n21535 ) ;
  assign n22135 = n22134 ^ n15592 ^ n5982 ;
  assign n22136 = n939 ^ n828 ^ 1'b0 ;
  assign n22137 = n946 & n22136 ;
  assign n22138 = n22137 ^ n8203 ^ n5101 ;
  assign n22143 = ( n10106 & ~n13160 ) | ( n10106 & n20105 ) | ( ~n13160 & n20105 ) ;
  assign n22144 = n22143 ^ n9396 ^ 1'b0 ;
  assign n22139 = n21781 ^ n4478 ^ 1'b0 ;
  assign n22140 = n1201 | n22139 ;
  assign n22141 = ( n887 & n946 ) | ( n887 & n13756 ) | ( n946 & n13756 ) ;
  assign n22142 = ~n22140 & n22141 ;
  assign n22145 = n22144 ^ n22142 ^ 1'b0 ;
  assign n22146 = n22138 & n22145 ;
  assign n22147 = n9216 & n22146 ;
  assign n22148 = n21745 ^ n573 ^ 1'b0 ;
  assign n22149 = n19234 ^ n14349 ^ n6149 ;
  assign n22150 = ( n9836 & ~n12429 ) | ( n9836 & n22149 ) | ( ~n12429 & n22149 ) ;
  assign n22151 = n16592 ^ n15803 ^ n6513 ;
  assign n22152 = ( n2487 & n3424 ) | ( n2487 & n4693 ) | ( n3424 & n4693 ) ;
  assign n22153 = ( ~n8368 & n22151 ) | ( ~n8368 & n22152 ) | ( n22151 & n22152 ) ;
  assign n22154 = n5447 ^ n2699 ^ 1'b0 ;
  assign n22155 = ( n1684 & n4253 ) | ( n1684 & ~n11584 ) | ( n4253 & ~n11584 ) ;
  assign n22156 = n15612 ^ n12555 ^ n656 ;
  assign n22157 = n22156 ^ n17993 ^ n6085 ;
  assign n22158 = ( n10162 & ~n22155 ) | ( n10162 & n22157 ) | ( ~n22155 & n22157 ) ;
  assign n22159 = ( n2519 & ~n15107 ) | ( n2519 & n22158 ) | ( ~n15107 & n22158 ) ;
  assign n22160 = n22159 ^ n6027 ^ n4664 ;
  assign n22161 = ( n5178 & n5208 ) | ( n5178 & n14996 ) | ( n5208 & n14996 ) ;
  assign n22162 = ( n560 & n5678 ) | ( n560 & n22161 ) | ( n5678 & n22161 ) ;
  assign n22163 = n22162 ^ n12776 ^ n8849 ;
  assign n22167 = ~n1688 & n9811 ;
  assign n22168 = n22167 ^ n1453 ^ 1'b0 ;
  assign n22169 = ( ~n762 & n4600 ) | ( ~n762 & n22168 ) | ( n4600 & n22168 ) ;
  assign n22164 = x87 & n3044 ;
  assign n22165 = n22164 ^ n3935 ^ 1'b0 ;
  assign n22166 = n22165 ^ n16152 ^ 1'b0 ;
  assign n22170 = n22169 ^ n22166 ^ n12980 ;
  assign n22171 = ( n11416 & n14439 ) | ( n11416 & ~n18108 ) | ( n14439 & ~n18108 ) ;
  assign n22172 = n17446 ^ n10445 ^ 1'b0 ;
  assign n22173 = ~n22171 & n22172 ;
  assign n22174 = n22173 ^ n21054 ^ n18405 ;
  assign n22175 = n14477 ^ n8524 ^ n3549 ;
  assign n22176 = n19091 ^ n18888 ^ n10850 ;
  assign n22177 = ( n2414 & n8503 ) | ( n2414 & ~n18633 ) | ( n8503 & ~n18633 ) ;
  assign n22178 = n10850 ^ n10456 ^ n413 ;
  assign n22179 = n5377 | n22178 ;
  assign n22180 = n22179 ^ n13952 ^ 1'b0 ;
  assign n22181 = ~n11280 & n22180 ;
  assign n22182 = n8890 ^ n8105 ^ n7071 ;
  assign n22183 = n5131 & ~n22182 ;
  assign n22184 = ~n5453 & n22183 ;
  assign n22185 = ( n4298 & n8482 ) | ( n4298 & n18168 ) | ( n8482 & n18168 ) ;
  assign n22186 = ( n12402 & n22184 ) | ( n12402 & ~n22185 ) | ( n22184 & ~n22185 ) ;
  assign n22187 = ( n3037 & n6493 ) | ( n3037 & ~n22186 ) | ( n6493 & ~n22186 ) ;
  assign n22189 = ( x60 & ~n201 ) | ( x60 & n7704 ) | ( ~n201 & n7704 ) ;
  assign n22190 = n22189 ^ n10082 ^ n8367 ;
  assign n22188 = n6226 & ~n7235 ;
  assign n22191 = n22190 ^ n22188 ^ 1'b0 ;
  assign n22192 = n5811 ^ x97 ^ 1'b0 ;
  assign n22193 = n8966 & ~n22192 ;
  assign n22194 = ( n7897 & n8345 ) | ( n7897 & ~n11722 ) | ( n8345 & ~n11722 ) ;
  assign n22195 = n6794 ^ n6703 ^ n3480 ;
  assign n22196 = n22195 ^ n5550 ^ n3979 ;
  assign n22197 = ( ~n11836 & n14169 ) | ( ~n11836 & n22196 ) | ( n14169 & n22196 ) ;
  assign n22198 = n3497 & n13945 ;
  assign n22199 = n258 & n22198 ;
  assign n22200 = n21331 ^ n12520 ^ n4355 ;
  assign n22201 = ( ~n19553 & n22199 ) | ( ~n19553 & n22200 ) | ( n22199 & n22200 ) ;
  assign n22202 = ( n11699 & ~n13491 ) | ( n11699 & n22201 ) | ( ~n13491 & n22201 ) ;
  assign n22203 = n20934 ^ n10748 ^ n6169 ;
  assign n22204 = n6210 ^ n2055 ^ 1'b0 ;
  assign n22205 = ( n21008 & n22203 ) | ( n21008 & n22204 ) | ( n22203 & n22204 ) ;
  assign n22209 = n8263 & n20571 ;
  assign n22210 = n22209 ^ n4173 ^ 1'b0 ;
  assign n22206 = n5731 ^ n4315 ^ 1'b0 ;
  assign n22207 = n1973 | n22206 ;
  assign n22208 = n22207 ^ n21653 ^ n16642 ;
  assign n22211 = n22210 ^ n22208 ^ n5121 ;
  assign n22212 = n12278 ^ n11609 ^ n3475 ;
  assign n22218 = ( n3907 & n12113 ) | ( n3907 & n12481 ) | ( n12113 & n12481 ) ;
  assign n22219 = n22218 ^ n15159 ^ 1'b0 ;
  assign n22220 = n22219 ^ n8113 ^ n6723 ;
  assign n22221 = n9743 ^ n9079 ^ n1731 ;
  assign n22222 = ( ~n8455 & n21306 ) | ( ~n8455 & n22221 ) | ( n21306 & n22221 ) ;
  assign n22223 = n22222 ^ n6370 ^ n5671 ;
  assign n22224 = ( n7405 & n22220 ) | ( n7405 & ~n22223 ) | ( n22220 & ~n22223 ) ;
  assign n22213 = n18197 ^ n16287 ^ n14011 ;
  assign n22214 = n22213 ^ n18138 ^ n16218 ;
  assign n22215 = ( ~n11855 & n16443 ) | ( ~n11855 & n16737 ) | ( n16443 & n16737 ) ;
  assign n22216 = n22215 ^ n13276 ^ n4435 ;
  assign n22217 = ( n22155 & n22214 ) | ( n22155 & n22216 ) | ( n22214 & n22216 ) ;
  assign n22225 = n22224 ^ n22217 ^ n528 ;
  assign n22231 = ~n2783 & n12191 ;
  assign n22232 = n22231 ^ n9638 ^ 1'b0 ;
  assign n22229 = ( n1398 & n5429 ) | ( n1398 & n6018 ) | ( n5429 & n6018 ) ;
  assign n22226 = ( ~n787 & n5465 ) | ( ~n787 & n8351 ) | ( n5465 & n8351 ) ;
  assign n22227 = n22226 ^ n13460 ^ n8300 ;
  assign n22228 = ( ~n5256 & n10901 ) | ( ~n5256 & n22227 ) | ( n10901 & n22227 ) ;
  assign n22230 = n22229 ^ n22228 ^ n2555 ;
  assign n22233 = n22232 ^ n22230 ^ n18734 ;
  assign n22234 = n500 | n1076 ;
  assign n22235 = n5337 & ~n22234 ;
  assign n22236 = n9134 ^ n5624 ^ 1'b0 ;
  assign n22237 = n1937 | n3519 ;
  assign n22238 = n11596 ^ n5058 ^ n1057 ;
  assign n22239 = ( n7331 & ~n21581 ) | ( n7331 & n22238 ) | ( ~n21581 & n22238 ) ;
  assign n22240 = n6886 | n22239 ;
  assign n22241 = n9498 & ~n10730 ;
  assign n22242 = n22241 ^ n1841 ^ 1'b0 ;
  assign n22243 = n13117 & ~n22242 ;
  assign n22244 = ( ~n1899 & n3820 ) | ( ~n1899 & n22243 ) | ( n3820 & n22243 ) ;
  assign n22245 = n4691 | n5878 ;
  assign n22246 = ( n13808 & ~n21789 ) | ( n13808 & n22245 ) | ( ~n21789 & n22245 ) ;
  assign n22247 = ( n20459 & n22244 ) | ( n20459 & ~n22246 ) | ( n22244 & ~n22246 ) ;
  assign n22248 = n5531 ^ n1340 ^ 1'b0 ;
  assign n22249 = ( n3591 & n10504 ) | ( n3591 & ~n22248 ) | ( n10504 & ~n22248 ) ;
  assign n22250 = ( n2696 & ~n7832 ) | ( n2696 & n8489 ) | ( ~n7832 & n8489 ) ;
  assign n22251 = n22250 ^ n14302 ^ n5015 ;
  assign n22252 = ( n4868 & n11654 ) | ( n4868 & ~n22251 ) | ( n11654 & ~n22251 ) ;
  assign n22253 = n7830 ^ n1726 ^ 1'b0 ;
  assign n22254 = ( n9358 & n20823 ) | ( n9358 & n22072 ) | ( n20823 & n22072 ) ;
  assign n22257 = n12255 ^ n3492 ^ n1275 ;
  assign n22255 = ( n856 & n2335 ) | ( n856 & ~n4009 ) | ( n2335 & ~n4009 ) ;
  assign n22256 = n22255 ^ n725 ^ 1'b0 ;
  assign n22258 = n22257 ^ n22256 ^ n18290 ;
  assign n22259 = n6364 & ~n15953 ;
  assign n22260 = n22259 ^ n20014 ^ 1'b0 ;
  assign n22261 = ( ~n4196 & n12539 ) | ( ~n4196 & n22260 ) | ( n12539 & n22260 ) ;
  assign n22263 = n7227 ^ n3697 ^ 1'b0 ;
  assign n22264 = n9514 | n22263 ;
  assign n22262 = ( n3978 & n11331 ) | ( n3978 & ~n12780 ) | ( n11331 & ~n12780 ) ;
  assign n22265 = n22264 ^ n22262 ^ n4068 ;
  assign n22266 = ( n7916 & n8903 ) | ( n7916 & ~n13537 ) | ( n8903 & ~n13537 ) ;
  assign n22267 = n21795 ^ n10136 ^ n5805 ;
  assign n22268 = n14211 ^ n466 ^ 1'b0 ;
  assign n22269 = n22267 & n22268 ;
  assign n22270 = n19250 ^ n17041 ^ 1'b0 ;
  assign n22271 = n5912 ^ n2412 ^ 1'b0 ;
  assign n22272 = n14592 & ~n22271 ;
  assign n22273 = ( n3640 & n11304 ) | ( n3640 & n22272 ) | ( n11304 & n22272 ) ;
  assign n22274 = n10371 ^ n1179 ^ n133 ;
  assign n22275 = n7458 | n22012 ;
  assign n22276 = n22275 ^ n1463 ^ 1'b0 ;
  assign n22277 = n22274 & n22276 ;
  assign n22278 = n2654 & ~n22277 ;
  assign n22279 = n22278 ^ n12354 ^ n3375 ;
  assign n22280 = ( n2342 & n8798 ) | ( n2342 & ~n22279 ) | ( n8798 & ~n22279 ) ;
  assign n22281 = n21422 ^ n11737 ^ n9402 ;
  assign n22285 = n1579 & ~n8893 ;
  assign n22286 = n13758 & n22285 ;
  assign n22283 = n1453 | n3986 ;
  assign n22282 = n12482 | n18095 ;
  assign n22284 = n22283 ^ n22282 ^ 1'b0 ;
  assign n22287 = n22286 ^ n22284 ^ n6350 ;
  assign n22288 = ( n18706 & ~n22281 ) | ( n18706 & n22287 ) | ( ~n22281 & n22287 ) ;
  assign n22290 = n14996 ^ n8755 ^ 1'b0 ;
  assign n22289 = n11430 ^ n9388 ^ n1889 ;
  assign n22291 = n22290 ^ n22289 ^ n8618 ;
  assign n22292 = n16226 ^ n8104 ^ n5454 ;
  assign n22296 = n8562 ^ n7407 ^ n6150 ;
  assign n22293 = n6252 ^ n1968 ^ n620 ;
  assign n22294 = ( n564 & n13168 ) | ( n564 & n22293 ) | ( n13168 & n22293 ) ;
  assign n22295 = n22294 ^ n19877 ^ n1251 ;
  assign n22297 = n22296 ^ n22295 ^ n5578 ;
  assign n22298 = ( n5683 & n8247 ) | ( n5683 & ~n15295 ) | ( n8247 & ~n15295 ) ;
  assign n22299 = n1374 | n7339 ;
  assign n22300 = n22298 | n22299 ;
  assign n22301 = n10136 ^ n8406 ^ n1940 ;
  assign n22302 = n22301 ^ n17300 ^ x104 ;
  assign n22303 = n22302 ^ n15613 ^ n4497 ;
  assign n22304 = n19463 ^ n12060 ^ n9741 ;
  assign n22305 = n22304 ^ n527 ^ 1'b0 ;
  assign n22306 = n22305 ^ n13915 ^ n6693 ;
  assign n22307 = ( n1174 & ~n10081 ) | ( n1174 & n21950 ) | ( ~n10081 & n21950 ) ;
  assign n22308 = ( x119 & ~n4395 ) | ( x119 & n22307 ) | ( ~n4395 & n22307 ) ;
  assign n22309 = n17034 ^ n12597 ^ n4247 ;
  assign n22310 = ( ~n2988 & n3209 ) | ( ~n2988 & n8368 ) | ( n3209 & n8368 ) ;
  assign n22311 = ( n5446 & ~n18754 ) | ( n5446 & n22310 ) | ( ~n18754 & n22310 ) ;
  assign n22312 = ( ~n13047 & n18579 ) | ( ~n13047 & n20547 ) | ( n18579 & n20547 ) ;
  assign n22313 = n22312 ^ n9484 ^ n3505 ;
  assign n22314 = ( n4295 & n13556 ) | ( n4295 & n20648 ) | ( n13556 & n20648 ) ;
  assign n22315 = ( n1004 & n1393 ) | ( n1004 & n12496 ) | ( n1393 & n12496 ) ;
  assign n22316 = ( n1116 & ~n6251 ) | ( n1116 & n14630 ) | ( ~n6251 & n14630 ) ;
  assign n22317 = ~n1068 & n10359 ;
  assign n22318 = n6761 & n22317 ;
  assign n22319 = n17336 ^ n4783 ^ n1174 ;
  assign n22320 = n22319 ^ n19810 ^ 1'b0 ;
  assign n22321 = n12893 & ~n22320 ;
  assign n22323 = n18211 ^ n3935 ^ n2603 ;
  assign n22322 = ~n16614 & n18509 ;
  assign n22324 = n22323 ^ n22322 ^ 1'b0 ;
  assign n22325 = ( n6340 & n11609 ) | ( n6340 & n15073 ) | ( n11609 & n15073 ) ;
  assign n22326 = n16094 ^ n13778 ^ x66 ;
  assign n22327 = n22326 ^ n19087 ^ n6782 ;
  assign n22332 = ( n1391 & ~n3468 ) | ( n1391 & n6409 ) | ( ~n3468 & n6409 ) ;
  assign n22328 = n13813 ^ n10844 ^ n3508 ;
  assign n22329 = ( n1451 & n3777 ) | ( n1451 & n22328 ) | ( n3777 & n22328 ) ;
  assign n22330 = n22329 ^ n6994 ^ 1'b0 ;
  assign n22331 = n4077 & n22330 ;
  assign n22333 = n22332 ^ n22331 ^ n16150 ;
  assign n22334 = n7029 ^ n3972 ^ n3938 ;
  assign n22335 = n22334 ^ n12728 ^ n8142 ;
  assign n22336 = n10990 ^ n3518 ^ n745 ;
  assign n22337 = ( n13379 & n15226 ) | ( n13379 & n22336 ) | ( n15226 & n22336 ) ;
  assign n22338 = ( ~n21682 & n22335 ) | ( ~n21682 & n22337 ) | ( n22335 & n22337 ) ;
  assign n22339 = ( n16047 & n19093 ) | ( n16047 & ~n22338 ) | ( n19093 & ~n22338 ) ;
  assign n22340 = n6205 & n13050 ;
  assign n22341 = n22340 ^ n3204 ^ 1'b0 ;
  assign n22342 = ( n5448 & n9136 ) | ( n5448 & n22341 ) | ( n9136 & n22341 ) ;
  assign n22343 = ( ~n698 & n2531 ) | ( ~n698 & n2928 ) | ( n2531 & n2928 ) ;
  assign n22344 = ( n240 & ~n7757 ) | ( n240 & n22343 ) | ( ~n7757 & n22343 ) ;
  assign n22345 = ( n8637 & n12187 ) | ( n8637 & n22344 ) | ( n12187 & n22344 ) ;
  assign n22346 = ( n686 & n1794 ) | ( n686 & n10442 ) | ( n1794 & n10442 ) ;
  assign n22347 = n20690 ^ n8753 ^ 1'b0 ;
  assign n22348 = ( ~n10371 & n22346 ) | ( ~n10371 & n22347 ) | ( n22346 & n22347 ) ;
  assign n22349 = n13128 & ~n22348 ;
  assign n22350 = n22349 ^ n19755 ^ n13559 ;
  assign n22351 = ( n1285 & n6219 ) | ( n1285 & ~n15709 ) | ( n6219 & ~n15709 ) ;
  assign n22352 = n18149 & ~n22351 ;
  assign n22353 = n22350 & n22352 ;
  assign n22354 = n4917 | n19476 ;
  assign n22355 = n1026 | n22354 ;
  assign n22356 = n16732 ^ n6071 ^ n441 ;
  assign n22357 = n15960 | n22356 ;
  assign n22358 = n22357 ^ n19493 ^ n4616 ;
  assign n22359 = n5815 | n7986 ;
  assign n22360 = n1919 & ~n22359 ;
  assign n22361 = n22360 ^ n12743 ^ 1'b0 ;
  assign n22362 = n22358 & n22361 ;
  assign n22363 = ( ~n9364 & n9413 ) | ( ~n9364 & n11071 ) | ( n9413 & n11071 ) ;
  assign n22364 = n22363 ^ n18772 ^ n4767 ;
  assign n22365 = ( ~n651 & n6469 ) | ( ~n651 & n22364 ) | ( n6469 & n22364 ) ;
  assign n22366 = n22365 ^ n19657 ^ 1'b0 ;
  assign n22367 = n16285 ^ n1464 ^ 1'b0 ;
  assign n22368 = ( ~x117 & n14015 ) | ( ~x117 & n17953 ) | ( n14015 & n17953 ) ;
  assign n22369 = n22368 ^ n9948 ^ n3107 ;
  assign n22370 = n17325 ^ n4915 ^ 1'b0 ;
  assign n22371 = n22370 ^ n11873 ^ n1857 ;
  assign n22372 = ~n3074 & n22371 ;
  assign n22373 = n22372 ^ n11447 ^ 1'b0 ;
  assign n22374 = ( n11628 & ~n12895 ) | ( n11628 & n22373 ) | ( ~n12895 & n22373 ) ;
  assign n22375 = ( ~n6290 & n16745 ) | ( ~n6290 & n21097 ) | ( n16745 & n21097 ) ;
  assign n22376 = n218 | n1822 ;
  assign n22377 = n3179 | n22376 ;
  assign n22378 = n9778 ^ n7731 ^ n643 ;
  assign n22379 = n22377 & n22378 ;
  assign n22380 = n22161 & n22379 ;
  assign n22381 = ~n333 & n987 ;
  assign n22382 = n22381 ^ n19985 ^ 1'b0 ;
  assign n22383 = ( n1050 & ~n7072 ) | ( n1050 & n10888 ) | ( ~n7072 & n10888 ) ;
  assign n22384 = n21200 ^ n12093 ^ n1361 ;
  assign n22385 = ( n846 & ~n12315 ) | ( n846 & n22384 ) | ( ~n12315 & n22384 ) ;
  assign n22386 = n22385 ^ n9754 ^ n7643 ;
  assign n22387 = ~n16023 & n22210 ;
  assign n22388 = n22387 ^ n19641 ^ 1'b0 ;
  assign n22389 = ~n1930 & n17246 ;
  assign n22390 = ( n19562 & ~n22388 ) | ( n19562 & n22389 ) | ( ~n22388 & n22389 ) ;
  assign n22391 = ( ~n5268 & n10644 ) | ( ~n5268 & n10837 ) | ( n10644 & n10837 ) ;
  assign n22392 = ( n3011 & ~n7726 ) | ( n3011 & n10089 ) | ( ~n7726 & n10089 ) ;
  assign n22393 = ( n11732 & n16983 ) | ( n11732 & ~n22392 ) | ( n16983 & ~n22392 ) ;
  assign n22394 = n16765 ^ n13382 ^ n1440 ;
  assign n22395 = n21018 ^ n4771 ^ 1'b0 ;
  assign n22396 = n22394 | n22395 ;
  assign n22397 = ( n5785 & n13316 ) | ( n5785 & ~n22347 ) | ( n13316 & ~n22347 ) ;
  assign n22400 = n7232 & ~n9581 ;
  assign n22398 = n12121 ^ n2047 ^ n943 ;
  assign n22399 = ( ~x78 & n6660 ) | ( ~x78 & n22398 ) | ( n6660 & n22398 ) ;
  assign n22401 = n22400 ^ n22399 ^ n15000 ;
  assign n22402 = n7167 & ~n15295 ;
  assign n22403 = ~n6131 & n22402 ;
  assign n22405 = n15638 ^ n12146 ^ x43 ;
  assign n22406 = n22405 ^ n16455 ^ n8647 ;
  assign n22404 = n4698 & n18083 ;
  assign n22407 = n22406 ^ n22404 ^ 1'b0 ;
  assign n22408 = ( n573 & n9399 ) | ( n573 & n22407 ) | ( n9399 & n22407 ) ;
  assign n22409 = n22408 ^ n21424 ^ n17722 ;
  assign n22410 = n7908 ^ n1833 ^ n1648 ;
  assign n22411 = ( n1766 & n5252 ) | ( n1766 & n22410 ) | ( n5252 & n22410 ) ;
  assign n22412 = n12642 ^ n6586 ^ 1'b0 ;
  assign n22413 = ~n4376 & n22412 ;
  assign n22414 = ( n17716 & ~n22411 ) | ( n17716 & n22413 ) | ( ~n22411 & n22413 ) ;
  assign n22415 = ( n22403 & n22409 ) | ( n22403 & n22414 ) | ( n22409 & n22414 ) ;
  assign n22416 = n14683 ^ n5035 ^ 1'b0 ;
  assign n22417 = n13844 | n22416 ;
  assign n22418 = n13255 ^ n1901 ^ 1'b0 ;
  assign n22421 = ( n422 & n1281 ) | ( n422 & ~n12831 ) | ( n1281 & ~n12831 ) ;
  assign n22419 = ( ~n4326 & n7071 ) | ( ~n4326 & n16847 ) | ( n7071 & n16847 ) ;
  assign n22420 = n22419 ^ n16803 ^ n6989 ;
  assign n22422 = n22421 ^ n22420 ^ n6226 ;
  assign n22423 = n7936 ^ n5744 ^ n1883 ;
  assign n22424 = n8605 ^ n4992 ^ n252 ;
  assign n22425 = ( ~n8850 & n15790 ) | ( ~n8850 & n22424 ) | ( n15790 & n22424 ) ;
  assign n22426 = ( n2461 & n3204 ) | ( n2461 & ~n8816 ) | ( n3204 & ~n8816 ) ;
  assign n22427 = ( ~n9366 & n15728 ) | ( ~n9366 & n22426 ) | ( n15728 & n22426 ) ;
  assign n22428 = n6295 | n15660 ;
  assign n22429 = n8875 | n22428 ;
  assign n22430 = n9804 & ~n22429 ;
  assign n22431 = ( n1109 & ~n5954 ) | ( n1109 & n9561 ) | ( ~n5954 & n9561 ) ;
  assign n22432 = n1143 | n3213 ;
  assign n22433 = n22432 ^ n13666 ^ 1'b0 ;
  assign n22434 = n22433 ^ n15206 ^ n10075 ;
  assign n22435 = n8989 ^ n509 ^ 1'b0 ;
  assign n22437 = ( n1688 & ~n1702 ) | ( n1688 & n8113 ) | ( ~n1702 & n8113 ) ;
  assign n22436 = ~n8018 & n9871 ;
  assign n22438 = n22437 ^ n22436 ^ n13981 ;
  assign n22439 = ( n797 & ~n3818 ) | ( n797 & n11997 ) | ( ~n3818 & n11997 ) ;
  assign n22440 = x54 & n22439 ;
  assign n22441 = n22440 ^ n2831 ^ 1'b0 ;
  assign n22442 = n22441 ^ n11377 ^ n9549 ;
  assign n22443 = n9250 ^ n4855 ^ 1'b0 ;
  assign n22444 = n22442 & ~n22443 ;
  assign n22445 = n12071 ^ n3470 ^ 1'b0 ;
  assign n22446 = ( n4020 & n19840 ) | ( n4020 & ~n22445 ) | ( n19840 & ~n22445 ) ;
  assign n22447 = n8087 ^ n7564 ^ n6524 ;
  assign n22448 = n22447 ^ n6569 ^ n4196 ;
  assign n22449 = ( n5614 & ~n18585 ) | ( n5614 & n22448 ) | ( ~n18585 & n22448 ) ;
  assign n22450 = ( n5560 & n8475 ) | ( n5560 & ~n10394 ) | ( n8475 & ~n10394 ) ;
  assign n22451 = ( n2457 & n6219 ) | ( n2457 & n22450 ) | ( n6219 & n22450 ) ;
  assign n22452 = n1682 & n9638 ;
  assign n22453 = ( ~n1390 & n22220 ) | ( ~n1390 & n22452 ) | ( n22220 & n22452 ) ;
  assign n22454 = n22453 ^ n4603 ^ n3973 ;
  assign n22456 = n9383 ^ n2918 ^ 1'b0 ;
  assign n22455 = n13027 ^ n8303 ^ 1'b0 ;
  assign n22457 = n22456 ^ n22455 ^ n16694 ;
  assign n22458 = n4443 & ~n18998 ;
  assign n22459 = n22458 ^ n6829 ^ 1'b0 ;
  assign n22460 = ( n2381 & ~n7780 ) | ( n2381 & n22459 ) | ( ~n7780 & n22459 ) ;
  assign n22461 = n10783 ^ n4213 ^ n2286 ;
  assign n22462 = ( n14664 & ~n22460 ) | ( n14664 & n22461 ) | ( ~n22460 & n22461 ) ;
  assign n22463 = n17511 ^ n12812 ^ n6582 ;
  assign n22464 = ( n20580 & n20717 ) | ( n20580 & ~n22463 ) | ( n20717 & ~n22463 ) ;
  assign n22465 = ( n3733 & ~n3995 ) | ( n3733 & n19973 ) | ( ~n3995 & n19973 ) ;
  assign n22466 = n22465 ^ n5723 ^ 1'b0 ;
  assign n22467 = ( n416 & ~n3357 ) | ( n416 & n11864 ) | ( ~n3357 & n11864 ) ;
  assign n22468 = ( n17728 & ~n17899 ) | ( n17728 & n22467 ) | ( ~n17899 & n22467 ) ;
  assign n22469 = n5431 ^ n4838 ^ 1'b0 ;
  assign n22470 = ~n22468 & n22469 ;
  assign n22471 = n22470 ^ n16640 ^ 1'b0 ;
  assign n22473 = ( ~n411 & n6636 ) | ( ~n411 & n6753 ) | ( n6636 & n6753 ) ;
  assign n22472 = n10273 ^ n9579 ^ n4414 ;
  assign n22474 = n22473 ^ n22472 ^ n12159 ;
  assign n22475 = ( n11553 & n13669 ) | ( n11553 & ~n14228 ) | ( n13669 & ~n14228 ) ;
  assign n22476 = n22475 ^ n18082 ^ n1296 ;
  assign n22477 = ( n3355 & n18749 ) | ( n3355 & ~n22476 ) | ( n18749 & ~n22476 ) ;
  assign n22478 = n4628 & n15828 ;
  assign n22480 = n5905 ^ n2023 ^ 1'b0 ;
  assign n22481 = n1219 & ~n22480 ;
  assign n22479 = n22196 ^ n8345 ^ n3919 ;
  assign n22482 = n22481 ^ n22479 ^ n12369 ;
  assign n22483 = ( ~n8127 & n17825 ) | ( ~n8127 & n21782 ) | ( n17825 & n21782 ) ;
  assign n22484 = n15641 ^ n11864 ^ 1'b0 ;
  assign n22485 = n15599 & ~n22484 ;
  assign n22486 = n22485 ^ n15210 ^ 1'b0 ;
  assign n22487 = n22483 & ~n22486 ;
  assign n22488 = n20297 ^ n10080 ^ n2651 ;
  assign n22489 = n12934 ^ n10512 ^ n6891 ;
  assign n22490 = n22489 ^ n15459 ^ n4982 ;
  assign n22491 = n22490 ^ n12800 ^ n3657 ;
  assign n22492 = ( n7625 & n10365 ) | ( n7625 & n18922 ) | ( n10365 & n18922 ) ;
  assign n22493 = n916 & ~n22492 ;
  assign n22494 = n18631 ^ n11799 ^ n10491 ;
  assign n22495 = n22494 ^ n2875 ^ n1805 ;
  assign n22496 = n10158 ^ n1259 ^ 1'b0 ;
  assign n22497 = ( n5366 & ~n18654 ) | ( n5366 & n22496 ) | ( ~n18654 & n22496 ) ;
  assign n22498 = ( n4218 & n5988 ) | ( n4218 & ~n6964 ) | ( n5988 & ~n6964 ) ;
  assign n22499 = n6990 & n7538 ;
  assign n22500 = n22498 & n22499 ;
  assign n22501 = n19523 & ~n22500 ;
  assign n22502 = n12821 & n22501 ;
  assign n22503 = n1485 & n8423 ;
  assign n22504 = n5752 | n20963 ;
  assign n22505 = ( ~n5478 & n18211 ) | ( ~n5478 & n22504 ) | ( n18211 & n22504 ) ;
  assign n22506 = n17992 ^ n14167 ^ n4173 ;
  assign n22507 = ( n344 & n1521 ) | ( n344 & n13416 ) | ( n1521 & n13416 ) ;
  assign n22508 = n17227 ^ n14533 ^ n139 ;
  assign n22509 = n3909 | n9477 ;
  assign n22510 = n22508 & ~n22509 ;
  assign n22511 = ( ~n13898 & n22507 ) | ( ~n13898 & n22510 ) | ( n22507 & n22510 ) ;
  assign n22512 = n10594 ^ n3790 ^ n1987 ;
  assign n22513 = n22512 ^ n5261 ^ n1923 ;
  assign n22514 = ( n19461 & n21770 ) | ( n19461 & n22513 ) | ( n21770 & n22513 ) ;
  assign n22515 = n7978 ^ x26 ^ 1'b0 ;
  assign n22516 = n17480 & ~n22515 ;
  assign n22517 = ( n2029 & n3316 ) | ( n2029 & ~n7957 ) | ( n3316 & ~n7957 ) ;
  assign n22518 = n10765 ^ n6150 ^ n3240 ;
  assign n22519 = ( n4885 & n5543 ) | ( n4885 & ~n22518 ) | ( n5543 & ~n22518 ) ;
  assign n22520 = n22519 ^ n14414 ^ n2387 ;
  assign n22522 = n2981 | n8241 ;
  assign n22521 = n17275 ^ n15100 ^ n13341 ;
  assign n22523 = n22522 ^ n22521 ^ n5080 ;
  assign n22524 = n7841 | n21142 ;
  assign n22525 = n22524 ^ n765 ^ 1'b0 ;
  assign n22526 = ( ~n7445 & n11505 ) | ( ~n7445 & n22525 ) | ( n11505 & n22525 ) ;
  assign n22527 = n13652 ^ n10269 ^ n4966 ;
  assign n22528 = n22527 ^ n11454 ^ n586 ;
  assign n22529 = n11403 | n13734 ;
  assign n22530 = n22528 & ~n22529 ;
  assign n22531 = ( n4286 & n4488 ) | ( n4286 & ~n4692 ) | ( n4488 & ~n4692 ) ;
  assign n22532 = ( n10385 & ~n11597 ) | ( n10385 & n22531 ) | ( ~n11597 & n22531 ) ;
  assign n22533 = n22532 ^ n15293 ^ n7737 ;
  assign n22534 = n13900 ^ n3197 ^ 1'b0 ;
  assign n22535 = ( ~n7133 & n8885 ) | ( ~n7133 & n18739 ) | ( n8885 & n18739 ) ;
  assign n22536 = n22535 ^ n1950 ^ 1'b0 ;
  assign n22537 = n6170 ^ n3972 ^ n1303 ;
  assign n22538 = n11037 ^ n10935 ^ 1'b0 ;
  assign n22539 = n22538 ^ n15199 ^ n2874 ;
  assign n22540 = n15956 ^ n13066 ^ 1'b0 ;
  assign n22541 = n17851 ^ n10359 ^ 1'b0 ;
  assign n22542 = ~n3646 & n8989 ;
  assign n22543 = n22541 & n22542 ;
  assign n22544 = n1576 & ~n14089 ;
  assign n22545 = n22544 ^ n18506 ^ 1'b0 ;
  assign n22546 = n19813 ^ n18832 ^ 1'b0 ;
  assign n22547 = ~n5946 & n10525 ;
  assign n22548 = ~n22546 & n22547 ;
  assign n22549 = n12238 ^ n11338 ^ n7485 ;
  assign n22550 = n11615 ^ n9224 ^ n8120 ;
  assign n22551 = n22550 ^ n21738 ^ n10030 ;
  assign n22553 = n2716 | n6057 ;
  assign n22554 = n290 & ~n22553 ;
  assign n22552 = n15503 ^ n8630 ^ n3771 ;
  assign n22555 = n22554 ^ n22552 ^ n17729 ;
  assign n22556 = n1919 | n2030 ;
  assign n22557 = n8684 | n22556 ;
  assign n22558 = ( ~n3721 & n9985 ) | ( ~n3721 & n22557 ) | ( n9985 & n22557 ) ;
  assign n22559 = n22558 ^ n7842 ^ n1569 ;
  assign n22560 = n22232 ^ n16915 ^ n15979 ;
  assign n22561 = ( n1970 & n3569 ) | ( n1970 & n20090 ) | ( n3569 & n20090 ) ;
  assign n22562 = n12824 & n22561 ;
  assign n22563 = n22562 ^ n15165 ^ 1'b0 ;
  assign n22564 = ( n20703 & ~n21823 ) | ( n20703 & n22563 ) | ( ~n21823 & n22563 ) ;
  assign n22565 = ( n1025 & n12508 ) | ( n1025 & n17297 ) | ( n12508 & n17297 ) ;
  assign n22566 = ~n22564 & n22565 ;
  assign n22571 = n17500 ^ n3880 ^ n2512 ;
  assign n22567 = ( n1790 & n2889 ) | ( n1790 & n5452 ) | ( n2889 & n5452 ) ;
  assign n22568 = n22567 ^ n17403 ^ n13261 ;
  assign n22569 = ~n8161 & n20161 ;
  assign n22570 = n22568 & n22569 ;
  assign n22572 = n22571 ^ n22570 ^ n12605 ;
  assign n22573 = ( ~n7603 & n11758 ) | ( ~n7603 & n21619 ) | ( n11758 & n21619 ) ;
  assign n22574 = ( n3915 & n6535 ) | ( n3915 & n15722 ) | ( n6535 & n15722 ) ;
  assign n22575 = ( n5659 & ~n13097 ) | ( n5659 & n20491 ) | ( ~n13097 & n20491 ) ;
  assign n22576 = n22508 ^ n2390 ^ 1'b0 ;
  assign n22577 = n5712 & ~n22576 ;
  assign n22578 = n7600 ^ n6095 ^ 1'b0 ;
  assign n22579 = n1574 | n22578 ;
  assign n22580 = ( n2400 & ~n21263 ) | ( n2400 & n22579 ) | ( ~n21263 & n22579 ) ;
  assign n22581 = n19691 ^ n3004 ^ n1005 ;
  assign n22585 = ( x75 & n5852 ) | ( x75 & ~n11092 ) | ( n5852 & ~n11092 ) ;
  assign n22582 = ( n4205 & ~n6689 ) | ( n4205 & n17744 ) | ( ~n6689 & n17744 ) ;
  assign n22583 = n13704 & n22582 ;
  assign n22584 = ( ~n6475 & n22077 ) | ( ~n6475 & n22583 ) | ( n22077 & n22583 ) ;
  assign n22586 = n22585 ^ n22584 ^ n16018 ;
  assign n22587 = ( n3209 & n5058 ) | ( n3209 & ~n9749 ) | ( n5058 & ~n9749 ) ;
  assign n22588 = n3939 ^ n1988 ^ n1679 ;
  assign n22589 = n8679 ^ n7746 ^ n4514 ;
  assign n22590 = n22588 & n22589 ;
  assign n22591 = n22590 ^ n14869 ^ 1'b0 ;
  assign n22592 = n7894 ^ n3531 ^ 1'b0 ;
  assign n22593 = ( n287 & n520 ) | ( n287 & ~n13537 ) | ( n520 & ~n13537 ) ;
  assign n22594 = ( ~n2725 & n3652 ) | ( ~n2725 & n22593 ) | ( n3652 & n22593 ) ;
  assign n22595 = ( n10402 & ~n18541 ) | ( n10402 & n22594 ) | ( ~n18541 & n22594 ) ;
  assign n22596 = n16051 ^ n797 ^ 1'b0 ;
  assign n22597 = ~n4521 & n22596 ;
  assign n22598 = n2043 & n7254 ;
  assign n22599 = n22598 ^ n1638 ^ 1'b0 ;
  assign n22600 = ~n327 & n22599 ;
  assign n22601 = n22600 ^ n22020 ^ n6507 ;
  assign n22602 = n22601 ^ n1949 ^ 1'b0 ;
  assign n22603 = ( x87 & n8676 ) | ( x87 & n22602 ) | ( n8676 & n22602 ) ;
  assign n22604 = n22603 ^ n14269 ^ 1'b0 ;
  assign n22605 = n22597 | n22604 ;
  assign n22606 = ( n8544 & n12105 ) | ( n8544 & n13074 ) | ( n12105 & n13074 ) ;
  assign n22607 = ( ~n3836 & n7799 ) | ( ~n3836 & n10536 ) | ( n7799 & n10536 ) ;
  assign n22608 = n20933 ^ n13141 ^ 1'b0 ;
  assign n22609 = ~n2054 & n22608 ;
  assign n22610 = ( n18139 & ~n22607 ) | ( n18139 & n22609 ) | ( ~n22607 & n22609 ) ;
  assign n22611 = n14244 | n22610 ;
  assign n22612 = ( n15115 & ~n22606 ) | ( n15115 & n22611 ) | ( ~n22606 & n22611 ) ;
  assign n22613 = n11485 | n12889 ;
  assign n22614 = n19019 ^ n1481 ^ 1'b0 ;
  assign n22615 = n22613 | n22614 ;
  assign n22616 = n643 & n1401 ;
  assign n22617 = ~n18225 & n22616 ;
  assign n22618 = n22617 ^ n14368 ^ n13405 ;
  assign n22619 = n20740 ^ n16575 ^ n7067 ;
  assign n22620 = n6363 ^ n5757 ^ n2802 ;
  assign n22621 = n22620 ^ n10099 ^ n3996 ;
  assign n22622 = n22621 ^ n10171 ^ n4289 ;
  assign n22623 = ( ~n6727 & n11511 ) | ( ~n6727 & n15441 ) | ( n11511 & n15441 ) ;
  assign n22624 = ( n879 & n4388 ) | ( n879 & ~n9787 ) | ( n4388 & ~n9787 ) ;
  assign n22625 = n11678 ^ n11152 ^ n6884 ;
  assign n22626 = n12340 ^ n6498 ^ 1'b0 ;
  assign n22627 = ~n2331 & n22626 ;
  assign n22628 = n10861 ^ n10761 ^ n9423 ;
  assign n22629 = n1065 | n2740 ;
  assign n22630 = n22628 & ~n22629 ;
  assign n22631 = n13397 ^ n11402 ^ n7855 ;
  assign n22632 = n18811 ^ n4547 ^ n3621 ;
  assign n22633 = n21128 ^ n18435 ^ 1'b0 ;
  assign n22634 = n8832 ^ n8419 ^ n1464 ;
  assign n22635 = n22634 ^ n20207 ^ n19238 ;
  assign n22636 = ( n4865 & n11234 ) | ( n4865 & ~n21908 ) | ( n11234 & ~n21908 ) ;
  assign n22638 = n6370 & n10479 ;
  assign n22639 = n22638 ^ n10818 ^ n8769 ;
  assign n22637 = n11510 ^ n10545 ^ 1'b0 ;
  assign n22640 = n22639 ^ n22637 ^ n6502 ;
  assign n22641 = n13355 ^ n8627 ^ 1'b0 ;
  assign n22642 = n21179 ^ n9391 ^ 1'b0 ;
  assign n22643 = n1129 | n22642 ;
  assign n22644 = n19018 ^ n9158 ^ n5360 ;
  assign n22645 = n14406 ^ n1860 ^ 1'b0 ;
  assign n22646 = n4678 & n22645 ;
  assign n22647 = n22646 ^ n22207 ^ n6734 ;
  assign n22648 = ( n5763 & ~n11155 ) | ( n5763 & n22647 ) | ( ~n11155 & n22647 ) ;
  assign n22649 = ( n390 & n18388 ) | ( n390 & ~n22648 ) | ( n18388 & ~n22648 ) ;
  assign n22650 = ( n2356 & n10145 ) | ( n2356 & n16171 ) | ( n10145 & n16171 ) ;
  assign n22651 = ( n2041 & ~n6867 ) | ( n2041 & n7873 ) | ( ~n6867 & n7873 ) ;
  assign n22652 = n13187 ^ n4139 ^ n3650 ;
  assign n22653 = n22652 ^ n11402 ^ n3696 ;
  assign n22654 = n19323 ^ n5820 ^ 1'b0 ;
  assign n22655 = n247 & ~n22654 ;
  assign n22656 = n13705 ^ n10587 ^ n213 ;
  assign n22657 = n22656 ^ n10253 ^ n6048 ;
  assign n22658 = n716 & n14044 ;
  assign n22659 = n22658 ^ n16792 ^ 1'b0 ;
  assign n22660 = n22659 ^ n10940 ^ n7449 ;
  assign n22664 = ( n3214 & ~n5109 ) | ( n3214 & n10889 ) | ( ~n5109 & n10889 ) ;
  assign n22662 = n14922 ^ n11704 ^ n4667 ;
  assign n22661 = n4579 & ~n13931 ;
  assign n22663 = n22662 ^ n22661 ^ 1'b0 ;
  assign n22665 = n22664 ^ n22663 ^ n10399 ;
  assign n22666 = n10322 ^ n4612 ^ 1'b0 ;
  assign n22667 = n5542 ^ n2609 ^ 1'b0 ;
  assign n22668 = n9412 ^ n9176 ^ n7166 ;
  assign n22669 = ( ~n19062 & n22667 ) | ( ~n19062 & n22668 ) | ( n22667 & n22668 ) ;
  assign n22670 = ( ~n10950 & n15099 ) | ( ~n10950 & n22669 ) | ( n15099 & n22669 ) ;
  assign n22671 = ( ~n14595 & n17376 ) | ( ~n14595 & n22670 ) | ( n17376 & n22670 ) ;
  assign n22672 = n12791 | n15897 ;
  assign n22678 = n527 & ~n15341 ;
  assign n22679 = ~n15924 & n22678 ;
  assign n22676 = ( ~n9407 & n10479 ) | ( ~n9407 & n18509 ) | ( n10479 & n18509 ) ;
  assign n22673 = n11711 ^ n6393 ^ n197 ;
  assign n22674 = n22673 ^ n10942 ^ n9312 ;
  assign n22675 = n6412 | n22674 ;
  assign n22677 = n22676 ^ n22675 ^ 1'b0 ;
  assign n22680 = n22679 ^ n22677 ^ n18641 ;
  assign n22681 = ( n1578 & n5973 ) | ( n1578 & n8503 ) | ( n5973 & n8503 ) ;
  assign n22682 = ( n6158 & n9727 ) | ( n6158 & ~n18124 ) | ( n9727 & ~n18124 ) ;
  assign n22683 = n20536 ^ n11717 ^ 1'b0 ;
  assign n22684 = n17984 ^ n15263 ^ n9506 ;
  assign n22685 = n8367 | n21721 ;
  assign n22686 = n22685 ^ n20304 ^ n9495 ;
  assign n22687 = n22686 ^ n9205 ^ 1'b0 ;
  assign n22688 = n22348 ^ n20095 ^ n18710 ;
  assign n22689 = n14798 & n16495 ;
  assign n22690 = n22689 ^ n19738 ^ 1'b0 ;
  assign n22691 = n12838 & n22690 ;
  assign n22692 = ( n4637 & ~n9024 ) | ( n4637 & n17744 ) | ( ~n9024 & n17744 ) ;
  assign n22697 = n13278 ^ n8759 ^ n7655 ;
  assign n22694 = n17396 ^ n14456 ^ n7617 ;
  assign n22693 = n19587 ^ n10142 ^ 1'b0 ;
  assign n22695 = n22694 ^ n22693 ^ n10120 ;
  assign n22696 = n2502 | n22695 ;
  assign n22698 = n22697 ^ n22696 ^ 1'b0 ;
  assign n22699 = ( n4730 & n10529 ) | ( n4730 & n22698 ) | ( n10529 & n22698 ) ;
  assign n22700 = n17581 ^ n15577 ^ 1'b0 ;
  assign n22701 = n13044 | n21642 ;
  assign n22702 = n22701 ^ n13972 ^ n6281 ;
  assign n22703 = n22199 ^ n17847 ^ n16192 ;
  assign n22704 = n4929 ^ n4697 ^ n3900 ;
  assign n22705 = n22704 ^ n5429 ^ n954 ;
  assign n22706 = n22274 ^ n9903 ^ 1'b0 ;
  assign n22707 = n864 & ~n7424 ;
  assign n22708 = ( n7565 & ~n22706 ) | ( n7565 & n22707 ) | ( ~n22706 & n22707 ) ;
  assign n22709 = n7350 & ~n8614 ;
  assign n22710 = n20780 | n22709 ;
  assign n22711 = n2181 | n22710 ;
  assign n22712 = ( ~n18783 & n22708 ) | ( ~n18783 & n22711 ) | ( n22708 & n22711 ) ;
  assign n22713 = ( n1194 & n22705 ) | ( n1194 & n22712 ) | ( n22705 & n22712 ) ;
  assign n22715 = n4076 ^ n1214 ^ 1'b0 ;
  assign n22714 = n10289 ^ n8927 ^ n2348 ;
  assign n22716 = n22715 ^ n22714 ^ n3789 ;
  assign n22717 = n22716 ^ n13017 ^ n6406 ;
  assign n22718 = n10394 & ~n15041 ;
  assign n22719 = ~n10327 & n14971 ;
  assign n22720 = n22718 & n22719 ;
  assign n22721 = n21461 ^ n8816 ^ 1'b0 ;
  assign n22722 = ~n22720 & n22721 ;
  assign n22723 = n14115 ^ n5259 ^ 1'b0 ;
  assign n22724 = ( n2070 & n3531 ) | ( n2070 & ~n18574 ) | ( n3531 & ~n18574 ) ;
  assign n22725 = n22723 & ~n22724 ;
  assign n22726 = ~n19781 & n22725 ;
  assign n22727 = ( ~x49 & n18437 ) | ( ~x49 & n21281 ) | ( n18437 & n21281 ) ;
  assign n22728 = ( n5100 & ~n12751 ) | ( n5100 & n22456 ) | ( ~n12751 & n22456 ) ;
  assign n22729 = n22727 & n22728 ;
  assign n22730 = ( n11376 & n16139 ) | ( n11376 & ~n16521 ) | ( n16139 & ~n16521 ) ;
  assign n22731 = ( n2508 & n15850 ) | ( n2508 & n22730 ) | ( n15850 & n22730 ) ;
  assign n22732 = n22731 ^ n20194 ^ n17581 ;
  assign n22733 = n18319 ^ n2588 ^ 1'b0 ;
  assign n22734 = n18799 & n22733 ;
  assign n22735 = n22734 ^ n5655 ^ n2810 ;
  assign n22736 = ( ~n2881 & n6060 ) | ( ~n2881 & n10511 ) | ( n6060 & n10511 ) ;
  assign n22737 = n9475 | n22736 ;
  assign n22738 = n22737 ^ n16516 ^ 1'b0 ;
  assign n22739 = n22738 ^ n8425 ^ 1'b0 ;
  assign n22740 = n11726 & ~n22739 ;
  assign n22741 = n7532 ^ n3081 ^ n2131 ;
  assign n22742 = ( ~n7021 & n7157 ) | ( ~n7021 & n22741 ) | ( n7157 & n22741 ) ;
  assign n22743 = n22742 ^ n7969 ^ 1'b0 ;
  assign n22744 = n8538 | n22743 ;
  assign n22745 = n9296 ^ n3954 ^ n1030 ;
  assign n22746 = ( n17819 & n20808 ) | ( n17819 & ~n22745 ) | ( n20808 & ~n22745 ) ;
  assign n22747 = ( n4204 & n11754 ) | ( n4204 & n16667 ) | ( n11754 & n16667 ) ;
  assign n22748 = ( ~n2871 & n5998 ) | ( ~n2871 & n9014 ) | ( n5998 & n9014 ) ;
  assign n22749 = n10998 ^ n216 ^ 1'b0 ;
  assign n22750 = ( ~n16026 & n22508 ) | ( ~n16026 & n22749 ) | ( n22508 & n22749 ) ;
  assign n22751 = n22750 ^ n21743 ^ n2078 ;
  assign n22752 = n5889 | n17544 ;
  assign n22753 = n22752 ^ n16047 ^ 1'b0 ;
  assign n22754 = n17851 ^ n11778 ^ n6230 ;
  assign n22755 = ~n1267 & n17884 ;
  assign n22756 = n22755 ^ n17352 ^ n4326 ;
  assign n22757 = n7726 ^ n5527 ^ 1'b0 ;
  assign n22758 = n10783 | n22757 ;
  assign n22759 = ( ~n6439 & n7433 ) | ( ~n6439 & n22758 ) | ( n7433 & n22758 ) ;
  assign n22760 = n2701 | n10373 ;
  assign n22761 = n21959 | n22760 ;
  assign n22762 = n16721 ^ n13052 ^ n6188 ;
  assign n22763 = ( n11773 & n13774 ) | ( n11773 & ~n17024 ) | ( n13774 & ~n17024 ) ;
  assign n22764 = n8539 ^ n3491 ^ n2752 ;
  assign n22765 = n18234 ^ n16688 ^ n5871 ;
  assign n22766 = ( n5504 & n16416 ) | ( n5504 & n22765 ) | ( n16416 & n22765 ) ;
  assign n22767 = ( n823 & n3882 ) | ( n823 & ~n4339 ) | ( n3882 & ~n4339 ) ;
  assign n22768 = ( n12656 & ~n13108 ) | ( n12656 & n22767 ) | ( ~n13108 & n22767 ) ;
  assign n22769 = n10179 & n22768 ;
  assign n22770 = n12848 ^ n9418 ^ n2447 ;
  assign n22771 = ~n16751 & n22770 ;
  assign n22774 = n8085 & ~n18030 ;
  assign n22775 = n22774 ^ n18097 ^ 1'b0 ;
  assign n22772 = n11505 & n21998 ;
  assign n22773 = n3262 & n22772 ;
  assign n22776 = n22775 ^ n22773 ^ n20262 ;
  assign n22777 = ~n10768 & n13424 ;
  assign n22778 = ~n3901 & n22777 ;
  assign n22779 = n4881 | n10266 ;
  assign n22780 = n8171 & n22779 ;
  assign n22781 = n22780 ^ n5118 ^ 1'b0 ;
  assign n22782 = ( n3315 & n5713 ) | ( n3315 & n22706 ) | ( n5713 & n22706 ) ;
  assign n22783 = n12462 ^ n9662 ^ n760 ;
  assign n22784 = ( ~n3702 & n22782 ) | ( ~n3702 & n22783 ) | ( n22782 & n22783 ) ;
  assign n22785 = ( n4646 & ~n20689 ) | ( n4646 & n22784 ) | ( ~n20689 & n22784 ) ;
  assign n22786 = ( n2793 & n6464 ) | ( n2793 & ~n7190 ) | ( n6464 & ~n7190 ) ;
  assign n22787 = ( n1044 & n9760 ) | ( n1044 & ~n22786 ) | ( n9760 & ~n22786 ) ;
  assign n22788 = ( ~n6875 & n7616 ) | ( ~n6875 & n14906 ) | ( n7616 & n14906 ) ;
  assign n22795 = ( n3327 & n13690 ) | ( n3327 & ~n18509 ) | ( n13690 & ~n18509 ) ;
  assign n22794 = n10657 ^ n10445 ^ 1'b0 ;
  assign n22796 = n22795 ^ n22794 ^ n7086 ;
  assign n22791 = ( ~n272 & n7590 ) | ( ~n272 & n7622 ) | ( n7590 & n7622 ) ;
  assign n22789 = n14890 ^ n3586 ^ n1100 ;
  assign n22790 = n11174 | n22789 ;
  assign n22792 = n22791 ^ n22790 ^ n959 ;
  assign n22793 = n7485 | n22792 ;
  assign n22797 = n22796 ^ n22793 ^ n12595 ;
  assign n22798 = n12444 ^ n7593 ^ n1788 ;
  assign n22799 = n801 & ~n15036 ;
  assign n22800 = n22799 ^ n16093 ^ n1259 ;
  assign n22801 = n18212 ^ n7593 ^ 1'b0 ;
  assign n22802 = n7013 & ~n22801 ;
  assign n22803 = ( ~n13801 & n16991 ) | ( ~n13801 & n22638 ) | ( n16991 & n22638 ) ;
  assign n22804 = n22803 ^ n5989 ^ n159 ;
  assign n22805 = n12750 ^ n11005 ^ n9037 ;
  assign n22806 = x87 & ~n5473 ;
  assign n22807 = n5943 & n22806 ;
  assign n22808 = n18365 & ~n22436 ;
  assign n22809 = n22807 & n22808 ;
  assign n22810 = ( n1214 & n9164 ) | ( n1214 & ~n22711 ) | ( n9164 & ~n22711 ) ;
  assign n22811 = ( n21572 & n22809 ) | ( n21572 & n22810 ) | ( n22809 & n22810 ) ;
  assign n22812 = ( ~n11796 & n22805 ) | ( ~n11796 & n22811 ) | ( n22805 & n22811 ) ;
  assign n22813 = n8152 ^ n6277 ^ n3082 ;
  assign n22814 = n9594 & n20089 ;
  assign n22815 = ( n1488 & ~n2034 ) | ( n1488 & n17050 ) | ( ~n2034 & n17050 ) ;
  assign n22816 = n17677 ^ n15683 ^ n13619 ;
  assign n22817 = n6283 | n22816 ;
  assign n22818 = ( n18514 & ~n21023 ) | ( n18514 & n22817 ) | ( ~n21023 & n22817 ) ;
  assign n22819 = ( n4479 & n8716 ) | ( n4479 & ~n19805 ) | ( n8716 & ~n19805 ) ;
  assign n22820 = ( ~n5026 & n20122 ) | ( ~n5026 & n22667 ) | ( n20122 & n22667 ) ;
  assign n22821 = n22820 ^ n17909 ^ n4760 ;
  assign n22822 = ~n2799 & n4643 ;
  assign n22823 = ~n22821 & n22822 ;
  assign n22824 = n9705 | n13123 ;
  assign n22825 = x112 | n22824 ;
  assign n22826 = ( n5703 & ~n7093 ) | ( n5703 & n7470 ) | ( ~n7093 & n7470 ) ;
  assign n22827 = n9885 & n22826 ;
  assign n22828 = n22827 ^ n226 ^ 1'b0 ;
  assign n22829 = n22593 ^ n16064 ^ n12543 ;
  assign n22831 = x115 & ~n3761 ;
  assign n22832 = n22831 ^ n14176 ^ 1'b0 ;
  assign n22833 = n21681 & n22832 ;
  assign n22834 = n22833 ^ n22084 ^ 1'b0 ;
  assign n22830 = n20868 ^ n13300 ^ n12983 ;
  assign n22835 = n22834 ^ n22830 ^ n11728 ;
  assign n22836 = ( n7041 & n7641 ) | ( n7041 & ~n7917 ) | ( n7641 & ~n7917 ) ;
  assign n22837 = n5340 ^ n671 ^ n384 ;
  assign n22838 = n11196 & ~n22837 ;
  assign n22839 = ( ~n459 & n1842 ) | ( ~n459 & n4806 ) | ( n1842 & n4806 ) ;
  assign n22840 = n18327 ^ n9023 ^ 1'b0 ;
  assign n22841 = ~n22839 & n22840 ;
  assign n22842 = n21415 & n22841 ;
  assign n22843 = n234 & n22842 ;
  assign n22844 = n254 & n15575 ;
  assign n22845 = n22844 ^ n16067 ^ n6047 ;
  assign n22846 = n6687 & ~n10184 ;
  assign n22847 = ~n22845 & n22846 ;
  assign n22852 = n1342 & ~n10187 ;
  assign n22853 = n22852 ^ n9599 ^ 1'b0 ;
  assign n22850 = ( n11099 & n14153 ) | ( n11099 & n18673 ) | ( n14153 & n18673 ) ;
  assign n22849 = n21686 ^ n8729 ^ 1'b0 ;
  assign n22848 = ( ~n15243 & n15706 ) | ( ~n15243 & n17478 ) | ( n15706 & n17478 ) ;
  assign n22851 = n22850 ^ n22849 ^ n22848 ;
  assign n22854 = n22853 ^ n22851 ^ 1'b0 ;
  assign n22855 = n3255 ^ n2265 ^ n1686 ;
  assign n22856 = ( n13975 & n14308 ) | ( n13975 & ~n22855 ) | ( n14308 & ~n22855 ) ;
  assign n22857 = n22856 ^ n1911 ^ 1'b0 ;
  assign n22858 = n6356 ^ n5866 ^ n2461 ;
  assign n22859 = ( ~n1791 & n2381 ) | ( ~n1791 & n2800 ) | ( n2381 & n2800 ) ;
  assign n22860 = n22859 ^ n11674 ^ n2758 ;
  assign n22861 = n14329 ^ n8881 ^ n7974 ;
  assign n22862 = n2709 & n9300 ;
  assign n22863 = n22862 ^ n18050 ^ 1'b0 ;
  assign n22864 = ( n22860 & n22861 ) | ( n22860 & ~n22863 ) | ( n22861 & ~n22863 ) ;
  assign n22865 = ( n4852 & ~n5241 ) | ( n4852 & n22864 ) | ( ~n5241 & n22864 ) ;
  assign n22866 = n15090 ^ n10294 ^ 1'b0 ;
  assign n22867 = ( n3009 & n10242 ) | ( n3009 & ~n12814 ) | ( n10242 & ~n12814 ) ;
  assign n22868 = n22867 ^ n19380 ^ n15837 ;
  assign n22869 = n5079 ^ n840 ^ n761 ;
  assign n22870 = n22869 ^ n16434 ^ n9836 ;
  assign n22871 = ( n3669 & n8436 ) | ( n3669 & ~n14729 ) | ( n8436 & ~n14729 ) ;
  assign n22872 = ( n1447 & n5563 ) | ( n1447 & n22871 ) | ( n5563 & n22871 ) ;
  assign n22875 = ( n7297 & ~n7431 ) | ( n7297 & n8137 ) | ( ~n7431 & n8137 ) ;
  assign n22876 = ( ~n1350 & n6383 ) | ( ~n1350 & n12054 ) | ( n6383 & n12054 ) ;
  assign n22877 = ( n3166 & ~n9209 ) | ( n3166 & n22876 ) | ( ~n9209 & n22876 ) ;
  assign n22878 = n1088 & n22877 ;
  assign n22879 = ~n22875 & n22878 ;
  assign n22873 = n1182 & n4399 ;
  assign n22874 = n22873 ^ n15609 ^ 1'b0 ;
  assign n22880 = n22879 ^ n22874 ^ n14133 ;
  assign n22881 = ~n3257 & n11997 ;
  assign n22882 = n17899 ^ n13654 ^ 1'b0 ;
  assign n22883 = ~n3891 & n12150 ;
  assign n22884 = n22883 ^ n2808 ^ 1'b0 ;
  assign n22888 = n8925 | n12549 ;
  assign n22889 = n22888 ^ n1697 ^ 1'b0 ;
  assign n22890 = n22889 ^ n16540 ^ n14291 ;
  assign n22885 = n16540 ^ n7268 ^ n3432 ;
  assign n22886 = ( n5295 & ~n18560 ) | ( n5295 & n22885 ) | ( ~n18560 & n22885 ) ;
  assign n22887 = n6822 & n22886 ;
  assign n22891 = n22890 ^ n22887 ^ 1'b0 ;
  assign n22892 = n19919 ^ n19808 ^ n17806 ;
  assign n22895 = n15890 ^ n11515 ^ 1'b0 ;
  assign n22893 = ( n2060 & n6073 ) | ( n2060 & ~n7531 ) | ( n6073 & ~n7531 ) ;
  assign n22894 = ( ~n14567 & n20260 ) | ( ~n14567 & n22893 ) | ( n20260 & n22893 ) ;
  assign n22896 = n22895 ^ n22894 ^ n13909 ;
  assign n22897 = ( n3731 & n22892 ) | ( n3731 & n22896 ) | ( n22892 & n22896 ) ;
  assign n22898 = ( n5384 & n12898 ) | ( n5384 & n16213 ) | ( n12898 & n16213 ) ;
  assign n22899 = n22898 ^ n9405 ^ 1'b0 ;
  assign n22902 = n8556 ^ n4096 ^ 1'b0 ;
  assign n22903 = ~n17143 & n22902 ;
  assign n22904 = n22903 ^ n10299 ^ n2688 ;
  assign n22900 = ( ~n295 & n4557 ) | ( ~n295 & n14496 ) | ( n4557 & n14496 ) ;
  assign n22901 = ( n7006 & n7402 ) | ( n7006 & ~n22900 ) | ( n7402 & ~n22900 ) ;
  assign n22905 = n22904 ^ n22901 ^ n13795 ;
  assign n22906 = n22905 ^ n16215 ^ n2214 ;
  assign n22907 = n3774 & ~n8615 ;
  assign n22908 = n9075 & n22907 ;
  assign n22909 = n2360 & ~n4459 ;
  assign n22910 = n3106 | n22909 ;
  assign n22911 = n22910 ^ n5301 ^ 1'b0 ;
  assign n22912 = n21829 ^ n7129 ^ n6643 ;
  assign n22913 = n16405 ^ n14453 ^ n13854 ;
  assign n22914 = n22912 | n22913 ;
  assign n22915 = n22914 ^ n7160 ^ 1'b0 ;
  assign n22916 = ~n22911 & n22915 ;
  assign n22917 = ( n12730 & n22908 ) | ( n12730 & n22916 ) | ( n22908 & n22916 ) ;
  assign n22918 = n20610 ^ n17158 ^ n12031 ;
  assign n22919 = n6323 & ~n17589 ;
  assign n22921 = ( ~n2061 & n2714 ) | ( ~n2061 & n21036 ) | ( n2714 & n21036 ) ;
  assign n22920 = ( n3610 & n9347 ) | ( n3610 & ~n16072 ) | ( n9347 & ~n16072 ) ;
  assign n22922 = n22921 ^ n22920 ^ n8220 ;
  assign n22923 = n3653 & n6425 ;
  assign n22924 = ( ~n5320 & n22679 ) | ( ~n5320 & n22923 ) | ( n22679 & n22923 ) ;
  assign n22925 = n5224 | n10362 ;
  assign n22926 = n13761 ^ n1078 ^ 1'b0 ;
  assign n22927 = ~n10252 & n12233 ;
  assign n22928 = n22927 ^ n5885 ^ 1'b0 ;
  assign n22929 = n9458 ^ n3115 ^ 1'b0 ;
  assign n22930 = ~n22928 & n22929 ;
  assign n22931 = ( n10041 & n10861 ) | ( n10041 & n18822 ) | ( n10861 & n18822 ) ;
  assign n22932 = n22931 ^ n21191 ^ 1'b0 ;
  assign n22933 = n22930 & ~n22932 ;
  assign n22934 = n2651 & n8344 ;
  assign n22935 = n22934 ^ n21939 ^ 1'b0 ;
  assign n22936 = n1519 & n4407 ;
  assign n22937 = ( n4469 & n5495 ) | ( n4469 & ~n22936 ) | ( n5495 & ~n22936 ) ;
  assign n22938 = ( n3934 & n13394 ) | ( n3934 & n22937 ) | ( n13394 & n22937 ) ;
  assign n22939 = n22938 ^ n20875 ^ n17581 ;
  assign n22940 = ( ~n4620 & n5151 ) | ( ~n4620 & n6582 ) | ( n5151 & n6582 ) ;
  assign n22941 = n22081 ^ n3510 ^ 1'b0 ;
  assign n22942 = n21523 & ~n22941 ;
  assign n22943 = ( ~n573 & n22940 ) | ( ~n573 & n22942 ) | ( n22940 & n22942 ) ;
  assign n22944 = n16206 ^ n6446 ^ n4478 ;
  assign n22945 = ( n10103 & ~n22274 ) | ( n10103 & n22944 ) | ( ~n22274 & n22944 ) ;
  assign n22946 = n7094 ^ n4848 ^ n2444 ;
  assign n22947 = ( n5148 & n10770 ) | ( n5148 & ~n22555 ) | ( n10770 & ~n22555 ) ;
  assign n22948 = n5954 | n12153 ;
  assign n22949 = ~n4691 & n13139 ;
  assign n22950 = ~n22948 & n22949 ;
  assign n22951 = n8873 ^ n3661 ^ n623 ;
  assign n22952 = n1191 & n22951 ;
  assign n22953 = n22952 ^ n9668 ^ 1'b0 ;
  assign n22954 = n21560 ^ n7427 ^ 1'b0 ;
  assign n22955 = ( n2173 & n8403 ) | ( n2173 & n15583 ) | ( n8403 & n15583 ) ;
  assign n22956 = ( ~n4029 & n22954 ) | ( ~n4029 & n22955 ) | ( n22954 & n22955 ) ;
  assign n22957 = ( n10678 & n22953 ) | ( n10678 & ~n22956 ) | ( n22953 & ~n22956 ) ;
  assign n22958 = n10763 & n21356 ;
  assign n22959 = n22958 ^ n10150 ^ n2105 ;
  assign n22960 = n657 | n21958 ;
  assign n22961 = n12368 ^ n2875 ^ 1'b0 ;
  assign n22962 = n16327 & n18290 ;
  assign n22963 = n22962 ^ n8718 ^ 1'b0 ;
  assign n22964 = ~n15123 & n22963 ;
  assign n22965 = n22964 ^ n13343 ^ 1'b0 ;
  assign n22966 = ~n21456 & n22965 ;
  assign n22967 = ( n15165 & ~n19090 ) | ( n15165 & n21395 ) | ( ~n19090 & n21395 ) ;
  assign n22968 = n10875 & n22967 ;
  assign n22969 = n22968 ^ n8034 ^ 1'b0 ;
  assign n22970 = ~n9985 & n10860 ;
  assign n22971 = n22970 ^ n12866 ^ 1'b0 ;
  assign n22972 = n22971 ^ n7417 ^ 1'b0 ;
  assign n22978 = ( n3130 & n13299 ) | ( n3130 & ~n16398 ) | ( n13299 & ~n16398 ) ;
  assign n22973 = n5953 ^ n3460 ^ 1'b0 ;
  assign n22974 = n129 & ~n22973 ;
  assign n22975 = n22974 ^ n2775 ^ n519 ;
  assign n22976 = n22975 ^ n13796 ^ 1'b0 ;
  assign n22977 = n22976 ^ n20805 ^ n6117 ;
  assign n22979 = n22978 ^ n22977 ^ n18407 ;
  assign n22980 = n9288 ^ n6689 ^ n724 ;
  assign n22981 = n3777 & n22980 ;
  assign n22982 = n2277 & n22981 ;
  assign n22983 = ( n9520 & n14378 ) | ( n9520 & n22982 ) | ( n14378 & n22982 ) ;
  assign n22984 = n11279 ^ n7613 ^ n4111 ;
  assign n22985 = n22984 ^ n19312 ^ n2526 ;
  assign n22986 = n16229 ^ n13647 ^ n11752 ;
  assign n22987 = ( n2256 & n5566 ) | ( n2256 & n22986 ) | ( n5566 & n22986 ) ;
  assign n22988 = n18337 ^ n3946 ^ n1836 ;
  assign n22989 = ( n4247 & ~n19532 ) | ( n4247 & n22988 ) | ( ~n19532 & n22988 ) ;
  assign n22990 = ( n4740 & ~n17162 ) | ( n4740 & n20211 ) | ( ~n17162 & n20211 ) ;
  assign n22991 = n22990 ^ n22789 ^ 1'b0 ;
  assign n22992 = n22989 & ~n22991 ;
  assign n22993 = n14788 ^ n10210 ^ 1'b0 ;
  assign n22994 = n22993 ^ n11633 ^ n9306 ;
  assign n22995 = n4396 ^ x127 ^ x94 ;
  assign n22996 = ( n951 & n16164 ) | ( n951 & n22995 ) | ( n16164 & n22995 ) ;
  assign n22997 = ( n1261 & n1726 ) | ( n1261 & ~n8239 ) | ( n1726 & ~n8239 ) ;
  assign n22998 = ( n11808 & ~n13140 ) | ( n11808 & n22997 ) | ( ~n13140 & n22997 ) ;
  assign n22999 = n18928 ^ n17046 ^ n4452 ;
  assign n23000 = n7956 & ~n18984 ;
  assign n23001 = ( n9980 & n14250 ) | ( n9980 & ~n19369 ) | ( n14250 & ~n19369 ) ;
  assign n23002 = n903 & ~n15954 ;
  assign n23003 = n23001 & n23002 ;
  assign n23004 = ( n3959 & n10301 ) | ( n3959 & n23003 ) | ( n10301 & n23003 ) ;
  assign n23007 = n6128 ^ n4327 ^ n3573 ;
  assign n23008 = n23007 ^ n17259 ^ n4665 ;
  assign n23009 = ( ~n3697 & n5664 ) | ( ~n3697 & n23008 ) | ( n5664 & n23008 ) ;
  assign n23005 = n10657 ^ n7203 ^ n2056 ;
  assign n23006 = ( n142 & n2756 ) | ( n142 & n23005 ) | ( n2756 & n23005 ) ;
  assign n23010 = n23009 ^ n23006 ^ n5398 ;
  assign n23011 = n23010 ^ n18752 ^ n7541 ;
  assign n23012 = ~n2850 & n3990 ;
  assign n23013 = ~n17259 & n23012 ;
  assign n23014 = n23013 ^ n21340 ^ n2795 ;
  assign n23023 = ~n4121 & n7582 ;
  assign n23015 = n2872 ^ n1527 ^ 1'b0 ;
  assign n23016 = n12498 | n23015 ;
  assign n23017 = ( n1073 & n14561 ) | ( n1073 & ~n23016 ) | ( n14561 & ~n23016 ) ;
  assign n23018 = n13950 & n23017 ;
  assign n23019 = n23018 ^ n20415 ^ 1'b0 ;
  assign n23020 = ( n9421 & n13839 ) | ( n9421 & ~n23019 ) | ( n13839 & ~n23019 ) ;
  assign n23021 = ( n852 & n8412 ) | ( n852 & ~n23020 ) | ( n8412 & ~n23020 ) ;
  assign n23022 = n21756 | n23021 ;
  assign n23024 = n23023 ^ n23022 ^ n11986 ;
  assign n23025 = n11986 ^ x66 ^ 1'b0 ;
  assign n23026 = ~n16803 & n23025 ;
  assign n23027 = n8837 ^ n1425 ^ 1'b0 ;
  assign n23028 = ( ~n1679 & n9802 ) | ( ~n1679 & n23027 ) | ( n9802 & n23027 ) ;
  assign n23029 = n11856 | n23028 ;
  assign n23030 = n10472 | n13264 ;
  assign n23031 = n23030 ^ n11751 ^ 1'b0 ;
  assign n23032 = n23031 ^ n14122 ^ n9949 ;
  assign n23033 = ( x79 & n7692 ) | ( x79 & ~n23032 ) | ( n7692 & ~n23032 ) ;
  assign n23034 = n22049 ^ n12637 ^ n399 ;
  assign n23035 = ( ~n8016 & n19281 ) | ( ~n8016 & n23034 ) | ( n19281 & n23034 ) ;
  assign n23036 = n11199 ^ n4122 ^ n652 ;
  assign n23037 = ( n8646 & n20014 ) | ( n8646 & ~n21859 ) | ( n20014 & ~n21859 ) ;
  assign n23038 = n23036 & n23037 ;
  assign n23039 = n20705 ^ n15587 ^ n1368 ;
  assign n23040 = n17753 ^ n13138 ^ n11355 ;
  assign n23041 = n23040 ^ n17739 ^ n1837 ;
  assign n23042 = ( ~n7390 & n18293 ) | ( ~n7390 & n23041 ) | ( n18293 & n23041 ) ;
  assign n23043 = n16691 ^ n12827 ^ n11118 ;
  assign n23044 = n8644 ^ n5056 ^ 1'b0 ;
  assign n23047 = n3226 ^ n3131 ^ n488 ;
  assign n23048 = ~n16216 & n23047 ;
  assign n23045 = ( n9566 & n18860 ) | ( n9566 & ~n22016 ) | ( n18860 & ~n22016 ) ;
  assign n23046 = ( n14134 & ~n19359 ) | ( n14134 & n23045 ) | ( ~n19359 & n23045 ) ;
  assign n23049 = n23048 ^ n23046 ^ n12092 ;
  assign n23050 = n1039 & n17447 ;
  assign n23051 = n23050 ^ n10934 ^ n10667 ;
  assign n23052 = n12331 & n16157 ;
  assign n23053 = ( n17762 & n23051 ) | ( n17762 & n23052 ) | ( n23051 & n23052 ) ;
  assign n23054 = n19824 ^ n5586 ^ n5166 ;
  assign n23055 = n12889 | n23054 ;
  assign n23056 = n23055 ^ n5974 ^ 1'b0 ;
  assign n23057 = n6148 ^ n5142 ^ n1922 ;
  assign n23058 = n1562 & n23057 ;
  assign n23059 = n23058 ^ n15736 ^ n3729 ;
  assign n23060 = ( n8611 & n21157 ) | ( n8611 & ~n23059 ) | ( n21157 & ~n23059 ) ;
  assign n23061 = n16548 | n23060 ;
  assign n23062 = n17927 & ~n23061 ;
  assign n23063 = n159 | n8182 ;
  assign n23064 = ( n8873 & n9068 ) | ( n8873 & n13439 ) | ( n9068 & n13439 ) ;
  assign n23065 = ( n547 & ~n1258 ) | ( n547 & n15768 ) | ( ~n1258 & n15768 ) ;
  assign n23066 = n23065 ^ n22749 ^ n7473 ;
  assign n23067 = n23066 ^ n20520 ^ n17122 ;
  assign n23068 = n12996 ^ n8039 ^ n7618 ;
  assign n23069 = n21243 ^ n12159 ^ n3746 ;
  assign n23070 = n22698 | n23069 ;
  assign n23071 = n11756 ^ n2492 ^ n1950 ;
  assign n23072 = ( n2837 & n13192 ) | ( n2837 & ~n23071 ) | ( n13192 & ~n23071 ) ;
  assign n23073 = n20094 ^ n14850 ^ n6667 ;
  assign n23074 = ( n5442 & n9660 ) | ( n5442 & ~n11738 ) | ( n9660 & ~n11738 ) ;
  assign n23075 = ( n3617 & ~n6227 ) | ( n3617 & n6742 ) | ( ~n6227 & n6742 ) ;
  assign n23076 = n23075 ^ n692 ^ 1'b0 ;
  assign n23077 = ~n15326 & n23076 ;
  assign n23078 = ~n20696 & n23077 ;
  assign n23079 = n23078 ^ n3193 ^ 1'b0 ;
  assign n23080 = ( n8793 & ~n19390 ) | ( n8793 & n20676 ) | ( ~n19390 & n20676 ) ;
  assign n23081 = ( n3896 & n19062 ) | ( n3896 & n23080 ) | ( n19062 & n23080 ) ;
  assign n23082 = ( n10083 & ~n11011 ) | ( n10083 & n12519 ) | ( ~n11011 & n12519 ) ;
  assign n23083 = ( ~n8786 & n17115 ) | ( ~n8786 & n23082 ) | ( n17115 & n23082 ) ;
  assign n23085 = ( n3845 & n7860 ) | ( n3845 & n9705 ) | ( n7860 & n9705 ) ;
  assign n23086 = n23085 ^ n22018 ^ n129 ;
  assign n23084 = ( ~n5012 & n11018 ) | ( ~n5012 & n21113 ) | ( n11018 & n21113 ) ;
  assign n23087 = n23086 ^ n23084 ^ n12362 ;
  assign n23088 = n9106 ^ n3513 ^ n1742 ;
  assign n23089 = n7602 | n22617 ;
  assign n23090 = n3492 & ~n23089 ;
  assign n23091 = n23088 & ~n23090 ;
  assign n23092 = n8766 & n10878 ;
  assign n23093 = ~x25 & n23092 ;
  assign n23094 = n23093 ^ n5436 ^ n5103 ;
  assign n23095 = n23094 ^ n20598 ^ n16182 ;
  assign n23096 = n7564 ^ n4322 ^ 1'b0 ;
  assign n23097 = n4425 & n23096 ;
  assign n23098 = n11118 & n23097 ;
  assign n23099 = n15449 & n23098 ;
  assign n23100 = ( n3222 & n7039 ) | ( n3222 & n15897 ) | ( n7039 & n15897 ) ;
  assign n23101 = n605 | n23100 ;
  assign n23102 = n23041 & ~n23101 ;
  assign n23103 = ( n2988 & ~n3025 ) | ( n2988 & n9328 ) | ( ~n3025 & n9328 ) ;
  assign n23104 = n23103 ^ n3713 ^ 1'b0 ;
  assign n23105 = n23104 ^ n19015 ^ n1685 ;
  assign n23106 = n23105 ^ n15161 ^ 1'b0 ;
  assign n23110 = n2960 & n5035 ;
  assign n23111 = n7617 & n23110 ;
  assign n23107 = n13337 ^ n6608 ^ 1'b0 ;
  assign n23108 = n16011 & ~n23107 ;
  assign n23109 = n23108 ^ n20998 ^ n9026 ;
  assign n23112 = n23111 ^ n23109 ^ n22742 ;
  assign n23113 = n9320 ^ n4238 ^ 1'b0 ;
  assign n23114 = n2088 & ~n23113 ;
  assign n23115 = ( n5230 & ~n5943 ) | ( n5230 & n23114 ) | ( ~n5943 & n23114 ) ;
  assign n23116 = ~n179 & n23115 ;
  assign n23117 = n2644 & n23116 ;
  assign n23118 = n7353 & n7670 ;
  assign n23119 = n23118 ^ n8024 ^ 1'b0 ;
  assign n23120 = ( n964 & n8121 ) | ( n964 & n23119 ) | ( n8121 & n23119 ) ;
  assign n23121 = ( n10687 & ~n13271 ) | ( n10687 & n15629 ) | ( ~n13271 & n15629 ) ;
  assign n23122 = ( n4574 & n12347 ) | ( n4574 & n17361 ) | ( n12347 & n17361 ) ;
  assign n23123 = n14444 ^ n10938 ^ n543 ;
  assign n23124 = ( n3473 & ~n7756 ) | ( n3473 & n15444 ) | ( ~n7756 & n15444 ) ;
  assign n23125 = n23124 ^ n21504 ^ n15604 ;
  assign n23127 = n4577 & ~n18922 ;
  assign n23128 = ( ~n6884 & n17107 ) | ( ~n6884 & n23127 ) | ( n17107 & n23127 ) ;
  assign n23126 = n6765 | n12838 ;
  assign n23129 = n23128 ^ n23126 ^ 1'b0 ;
  assign n23130 = n13117 & ~n20095 ;
  assign n23131 = n23130 ^ n11404 ^ 1'b0 ;
  assign n23132 = n18921 ^ n18609 ^ n814 ;
  assign n23133 = n2947 & n15516 ;
  assign n23134 = n5668 ^ n317 ^ 1'b0 ;
  assign n23135 = n23134 ^ n4796 ^ n1279 ;
  assign n23138 = ( n2587 & n6715 ) | ( n2587 & ~n11929 ) | ( n6715 & ~n11929 ) ;
  assign n23136 = n11052 & n17717 ;
  assign n23137 = n9079 & n23136 ;
  assign n23139 = n23138 ^ n23137 ^ n22312 ;
  assign n23140 = ( ~n10651 & n17273 ) | ( ~n10651 & n17872 ) | ( n17273 & n17872 ) ;
  assign n23141 = n23140 ^ n11749 ^ 1'b0 ;
  assign n23142 = n6560 | n23141 ;
  assign n23143 = n23142 ^ n22668 ^ n8884 ;
  assign n23144 = n8691 & n13984 ;
  assign n23145 = n23144 ^ n6702 ^ 1'b0 ;
  assign n23146 = n6277 ^ n3642 ^ n153 ;
  assign n23147 = n5804 ^ n3104 ^ n1332 ;
  assign n23148 = ( n2858 & n3052 ) | ( n2858 & n23147 ) | ( n3052 & n23147 ) ;
  assign n23149 = n9503 | n23148 ;
  assign n23150 = ( n9236 & n23146 ) | ( n9236 & ~n23149 ) | ( n23146 & ~n23149 ) ;
  assign n23151 = n23150 ^ n22467 ^ n7456 ;
  assign n23152 = n13245 ^ n5569 ^ x7 ;
  assign n23153 = n23152 ^ n7881 ^ n4829 ;
  assign n23156 = n13066 ^ n8120 ^ n7119 ;
  assign n23157 = n23156 ^ n18220 ^ n9104 ;
  assign n23154 = ( ~n2614 & n4532 ) | ( ~n2614 & n13369 ) | ( n4532 & n13369 ) ;
  assign n23155 = ~n319 & n23154 ;
  assign n23158 = n23157 ^ n23155 ^ 1'b0 ;
  assign n23159 = ~n5576 & n12464 ;
  assign n23160 = ( n23153 & n23158 ) | ( n23153 & ~n23159 ) | ( n23158 & ~n23159 ) ;
  assign n23161 = n10013 ^ n8333 ^ 1'b0 ;
  assign n23162 = n9134 ^ n4829 ^ n4299 ;
  assign n23163 = ( n3543 & n19407 ) | ( n3543 & n23162 ) | ( n19407 & n23162 ) ;
  assign n23164 = ( n10274 & n14271 ) | ( n10274 & ~n15024 ) | ( n14271 & ~n15024 ) ;
  assign n23165 = ~n425 & n21497 ;
  assign n23166 = n23165 ^ n2091 ^ 1'b0 ;
  assign n23167 = ( ~n10008 & n11973 ) | ( ~n10008 & n17496 ) | ( n11973 & n17496 ) ;
  assign n23168 = n23167 ^ n1494 ^ 1'b0 ;
  assign n23169 = n22210 & n23168 ;
  assign n23170 = ( ~n6297 & n7034 ) | ( ~n6297 & n7516 ) | ( n7034 & n7516 ) ;
  assign n23171 = ( n6386 & n10493 ) | ( n6386 & ~n23170 ) | ( n10493 & ~n23170 ) ;
  assign n23172 = ( ~n4424 & n14654 ) | ( ~n4424 & n16358 ) | ( n14654 & n16358 ) ;
  assign n23173 = n23172 ^ n4976 ^ 1'b0 ;
  assign n23174 = n13160 ^ n1657 ^ 1'b0 ;
  assign n23175 = ( n287 & n798 ) | ( n287 & ~n23174 ) | ( n798 & ~n23174 ) ;
  assign n23176 = n19073 ^ n3316 ^ n2083 ;
  assign n23177 = n23176 ^ n9260 ^ n8944 ;
  assign n23178 = ( n7139 & n15813 ) | ( n7139 & ~n20376 ) | ( n15813 & ~n20376 ) ;
  assign n23179 = n8300 & n15721 ;
  assign n23180 = ~n23178 & n23179 ;
  assign n23181 = n23180 ^ n21475 ^ n11826 ;
  assign n23182 = n23181 ^ n14138 ^ 1'b0 ;
  assign n23183 = n2965 & ~n21782 ;
  assign n23184 = n12981 ^ n905 ^ 1'b0 ;
  assign n23185 = n21281 & n23184 ;
  assign n23186 = n4606 & n23185 ;
  assign n23187 = n17057 & n23186 ;
  assign n23188 = n23187 ^ n3226 ^ n3108 ;
  assign n23189 = ~n8207 & n22988 ;
  assign n23190 = n18652 ^ n15234 ^ n6642 ;
  assign n23191 = n23190 ^ n19545 ^ 1'b0 ;
  assign n23192 = n17412 ^ n16270 ^ n8060 ;
  assign n23193 = n9338 ^ n7173 ^ 1'b0 ;
  assign n23194 = n23193 ^ n18435 ^ n14533 ;
  assign n23195 = n23194 ^ n16831 ^ n15564 ;
  assign n23196 = n23195 ^ n8463 ^ n3722 ;
  assign n23197 = n21339 ^ n14996 ^ n8519 ;
  assign n23198 = n2983 & n4540 ;
  assign n23199 = n7165 | n23198 ;
  assign n23200 = n23197 & ~n23199 ;
  assign n23202 = n20822 ^ n2027 ^ 1'b0 ;
  assign n23201 = ~n17582 & n19685 ;
  assign n23203 = n23202 ^ n23201 ^ 1'b0 ;
  assign n23205 = ( n1762 & n11379 ) | ( n1762 & n14905 ) | ( n11379 & n14905 ) ;
  assign n23204 = n16708 ^ n8766 ^ n1481 ;
  assign n23206 = n23205 ^ n23204 ^ n1752 ;
  assign n23207 = n18686 ^ n11767 ^ n1880 ;
  assign n23208 = ~n1457 & n23207 ;
  assign n23209 = n16182 & n23208 ;
  assign n23210 = n21131 | n23209 ;
  assign n23211 = n13981 ^ n10899 ^ n6009 ;
  assign n23212 = ( ~n20341 & n20876 ) | ( ~n20341 & n23211 ) | ( n20876 & n23211 ) ;
  assign n23213 = ( n9176 & ~n9671 ) | ( n9176 & n13170 ) | ( ~n9671 & n13170 ) ;
  assign n23214 = n12172 ^ n4494 ^ n401 ;
  assign n23215 = n11417 ^ n1814 ^ 1'b0 ;
  assign n23216 = n23215 ^ n20420 ^ n14830 ;
  assign n23219 = n5017 ^ n4745 ^ n133 ;
  assign n23217 = n5645 | n5889 ;
  assign n23218 = n2447 | n23217 ;
  assign n23220 = n23219 ^ n23218 ^ n13594 ;
  assign n23221 = ( n9862 & n14318 ) | ( n9862 & n19688 ) | ( n14318 & n19688 ) ;
  assign n23222 = n23221 ^ n18553 ^ 1'b0 ;
  assign n23223 = n19265 ^ n17914 ^ n5809 ;
  assign n23224 = n14795 | n23223 ;
  assign n23225 = n12299 ^ n3655 ^ 1'b0 ;
  assign n23229 = ~n162 & n2442 ;
  assign n23226 = n22137 ^ n9152 ^ n8706 ;
  assign n23227 = n23226 ^ n1883 ^ 1'b0 ;
  assign n23228 = n23227 ^ n22830 ^ n2158 ;
  assign n23230 = n23229 ^ n23228 ^ 1'b0 ;
  assign n23231 = n5791 ^ n2551 ^ n298 ;
  assign n23232 = n6622 & n7440 ;
  assign n23233 = ~n15524 & n23232 ;
  assign n23235 = ( n2024 & n2747 ) | ( n2024 & n16241 ) | ( n2747 & n16241 ) ;
  assign n23234 = n6360 | n21240 ;
  assign n23236 = n23235 ^ n23234 ^ 1'b0 ;
  assign n23237 = ( ~n335 & n9146 ) | ( ~n335 & n11275 ) | ( n9146 & n11275 ) ;
  assign n23238 = n13168 ^ n8294 ^ 1'b0 ;
  assign n23239 = n23238 ^ n8308 ^ n3087 ;
  assign n23240 = n12609 ^ n8620 ^ 1'b0 ;
  assign n23241 = n2426 & ~n14752 ;
  assign n23242 = ~n16501 & n23241 ;
  assign n23243 = n23242 ^ n16485 ^ n9946 ;
  assign n23244 = n7207 ^ n5217 ^ n1421 ;
  assign n23245 = ~n12026 & n23244 ;
  assign n23246 = ( n858 & n11694 ) | ( n858 & ~n15853 ) | ( n11694 & ~n15853 ) ;
  assign n23247 = n23246 ^ n12645 ^ n2952 ;
  assign n23248 = n8481 | n22468 ;
  assign n23249 = n23193 & ~n23248 ;
  assign n23250 = ( n11774 & n17483 ) | ( n11774 & ~n20056 ) | ( n17483 & ~n20056 ) ;
  assign n23251 = n23250 ^ n20918 ^ n8777 ;
  assign n23252 = ( n2455 & n15337 ) | ( n2455 & ~n17648 ) | ( n15337 & ~n17648 ) ;
  assign n23253 = ~n3060 & n6593 ;
  assign n23254 = n17844 & n23253 ;
  assign n23255 = ( n9011 & n18755 ) | ( n9011 & n23254 ) | ( n18755 & n23254 ) ;
  assign n23256 = ~n7215 & n12505 ;
  assign n23257 = ~n13326 & n23256 ;
  assign n23258 = ( ~n6610 & n15813 ) | ( ~n6610 & n20132 ) | ( n15813 & n20132 ) ;
  assign n23259 = ( ~n22995 & n23257 ) | ( ~n22995 & n23258 ) | ( n23257 & n23258 ) ;
  assign n23260 = n23259 ^ n15728 ^ n9351 ;
  assign n23261 = ( n1354 & ~n3166 ) | ( n1354 & n10243 ) | ( ~n3166 & n10243 ) ;
  assign n23262 = n21424 ^ n4702 ^ 1'b0 ;
  assign n23263 = ( n5562 & n13854 ) | ( n5562 & n23262 ) | ( n13854 & n23262 ) ;
  assign n23264 = ( n1395 & n15128 ) | ( n1395 & ~n23263 ) | ( n15128 & ~n23263 ) ;
  assign n23265 = ( n3766 & ~n4429 ) | ( n3766 & n21595 ) | ( ~n4429 & n21595 ) ;
  assign n23266 = ~n2644 & n23265 ;
  assign n23267 = n23266 ^ n19347 ^ 1'b0 ;
  assign n23268 = n3053 ^ n1259 ^ 1'b0 ;
  assign n23269 = ~n1638 & n23268 ;
  assign n23271 = n12389 ^ n4672 ^ n2458 ;
  assign n23272 = n23271 ^ n6482 ^ n2248 ;
  assign n23273 = n8628 ^ n5164 ^ n1810 ;
  assign n23274 = n22518 | n23273 ;
  assign n23275 = n10292 ^ n2479 ^ n1372 ;
  assign n23276 = ( n23272 & ~n23274 ) | ( n23272 & n23275 ) | ( ~n23274 & n23275 ) ;
  assign n23270 = n19298 ^ n15846 ^ n5754 ;
  assign n23277 = n23276 ^ n23270 ^ 1'b0 ;
  assign n23278 = ( n1520 & ~n7036 ) | ( n1520 & n13002 ) | ( ~n7036 & n13002 ) ;
  assign n23279 = ( n4368 & ~n9741 ) | ( n4368 & n11234 ) | ( ~n9741 & n11234 ) ;
  assign n23280 = n13688 | n23279 ;
  assign n23281 = ( n1504 & ~n6633 ) | ( n1504 & n11189 ) | ( ~n6633 & n11189 ) ;
  assign n23282 = ( ~n12171 & n20823 ) | ( ~n12171 & n23281 ) | ( n20823 & n23281 ) ;
  assign n23283 = n7067 ^ n1028 ^ n451 ;
  assign n23284 = n4550 & ~n17492 ;
  assign n23285 = n4734 & n23284 ;
  assign n23286 = ( n3976 & ~n23283 ) | ( n3976 & n23285 ) | ( ~n23283 & n23285 ) ;
  assign n23288 = n9300 ^ n4508 ^ n1144 ;
  assign n23287 = ( n7713 & n10907 ) | ( n7713 & n19275 ) | ( n10907 & n19275 ) ;
  assign n23289 = n23288 ^ n23287 ^ n19146 ;
  assign n23291 = ( n6996 & ~n8009 ) | ( n6996 & n11487 ) | ( ~n8009 & n11487 ) ;
  assign n23290 = n8639 & n14702 ;
  assign n23292 = n23291 ^ n23290 ^ 1'b0 ;
  assign n23293 = n8234 & ~n23292 ;
  assign n23294 = n6979 & n23293 ;
  assign n23295 = n23294 ^ n18641 ^ n12277 ;
  assign n23296 = ( x119 & ~n21427 ) | ( x119 & n23295 ) | ( ~n21427 & n23295 ) ;
  assign n23297 = n9478 & n20070 ;
  assign n23298 = ~n4283 & n14848 ;
  assign n23299 = ~n149 & n23298 ;
  assign n23300 = n440 & n6931 ;
  assign n23301 = n838 & n23300 ;
  assign n23302 = ( ~n211 & n2276 ) | ( ~n211 & n23301 ) | ( n2276 & n23301 ) ;
  assign n23303 = n23302 ^ n9708 ^ 1'b0 ;
  assign n23304 = n7651 ^ n6402 ^ n3769 ;
  assign n23305 = n23303 & n23304 ;
  assign n23306 = ~n11099 & n23305 ;
  assign n23307 = ( x62 & ~n4134 ) | ( x62 & n16213 ) | ( ~n4134 & n16213 ) ;
  assign n23308 = ( ~n7513 & n9575 ) | ( ~n7513 & n23307 ) | ( n9575 & n23307 ) ;
  assign n23309 = n23308 ^ n14515 ^ n1705 ;
  assign n23310 = ( ~n5011 & n7698 ) | ( ~n5011 & n7859 ) | ( n7698 & n7859 ) ;
  assign n23311 = ( ~n12063 & n14834 ) | ( ~n12063 & n23310 ) | ( n14834 & n23310 ) ;
  assign n23312 = ( n17046 & n19850 ) | ( n17046 & n23311 ) | ( n19850 & n23311 ) ;
  assign n23313 = n17195 ^ n17070 ^ 1'b0 ;
  assign n23314 = n3589 & n23313 ;
  assign n23315 = ~n6959 & n23314 ;
  assign n23316 = ( x95 & ~n2267 ) | ( x95 & n4405 ) | ( ~n2267 & n4405 ) ;
  assign n23317 = ( n1231 & ~n2982 ) | ( n1231 & n9157 ) | ( ~n2982 & n9157 ) ;
  assign n23318 = ( n3711 & n23316 ) | ( n3711 & n23317 ) | ( n23316 & n23317 ) ;
  assign n23319 = ( n10373 & n23315 ) | ( n10373 & n23318 ) | ( n23315 & n23318 ) ;
  assign n23321 = n2879 ^ n784 ^ 1'b0 ;
  assign n23322 = ( n469 & n12228 ) | ( n469 & n23321 ) | ( n12228 & n23321 ) ;
  assign n23320 = n14957 ^ n13704 ^ n6071 ;
  assign n23323 = n23322 ^ n23320 ^ n19750 ;
  assign n23324 = ( n11514 & ~n11627 ) | ( n11514 & n12653 ) | ( ~n11627 & n12653 ) ;
  assign n23325 = n5362 ^ n2570 ^ 1'b0 ;
  assign n23326 = n23324 | n23325 ;
  assign n23327 = n12268 & ~n23326 ;
  assign n23328 = n23327 ^ n10344 ^ 1'b0 ;
  assign n23329 = ( n6660 & n7930 ) | ( n6660 & n23328 ) | ( n7930 & n23328 ) ;
  assign n23330 = ( n5316 & n10670 ) | ( n5316 & ~n21005 ) | ( n10670 & ~n21005 ) ;
  assign n23331 = n16789 ^ n8497 ^ 1'b0 ;
  assign n23332 = n23330 & ~n23331 ;
  assign n23333 = n16229 ^ n14568 ^ 1'b0 ;
  assign n23334 = n22347 & n23333 ;
  assign n23335 = ( ~n8537 & n22073 ) | ( ~n8537 & n22184 ) | ( n22073 & n22184 ) ;
  assign n23336 = n23335 ^ n900 ^ 1'b0 ;
  assign n23337 = ( n3835 & n18371 ) | ( n3835 & n23336 ) | ( n18371 & n23336 ) ;
  assign n23338 = n8801 & n15818 ;
  assign n23339 = n23338 ^ n18349 ^ n17789 ;
  assign n23342 = n8143 ^ n1853 ^ x20 ;
  assign n23340 = n7905 | n20188 ;
  assign n23341 = n7704 | n23340 ;
  assign n23343 = n23342 ^ n23341 ^ n19421 ;
  assign n23344 = n6043 ^ n2754 ^ n2355 ;
  assign n23345 = n17757 ^ n13919 ^ n7196 ;
  assign n23346 = n16593 ^ n15049 ^ n2391 ;
  assign n23347 = ( n16573 & n23345 ) | ( n16573 & ~n23346 ) | ( n23345 & ~n23346 ) ;
  assign n23348 = n15759 & ~n18517 ;
  assign n23349 = n23348 ^ n6720 ^ n1852 ;
  assign n23350 = n1494 | n7940 ;
  assign n23351 = n23350 ^ n11359 ^ 1'b0 ;
  assign n23352 = n6530 & n19607 ;
  assign n23353 = n11666 ^ n6713 ^ n3220 ;
  assign n23354 = ( n11052 & n18452 ) | ( n11052 & n23353 ) | ( n18452 & n23353 ) ;
  assign n23359 = n12380 ^ n6265 ^ 1'b0 ;
  assign n23356 = n5549 ^ n719 ^ 1'b0 ;
  assign n23357 = n13780 | n23356 ;
  assign n23355 = n5732 ^ n2398 ^ n1402 ;
  assign n23358 = n23357 ^ n23355 ^ n20363 ;
  assign n23360 = n23359 ^ n23358 ^ n5573 ;
  assign n23364 = n13768 ^ n7348 ^ n305 ;
  assign n23361 = ( n8074 & n8154 ) | ( n8074 & ~n11500 ) | ( n8154 & ~n11500 ) ;
  assign n23362 = ( ~n1093 & n3256 ) | ( ~n1093 & n9777 ) | ( n3256 & n9777 ) ;
  assign n23363 = ( ~n1305 & n23361 ) | ( ~n1305 & n23362 ) | ( n23361 & n23362 ) ;
  assign n23365 = n23364 ^ n23363 ^ n14509 ;
  assign n23366 = n4080 & n4147 ;
  assign n23367 = ~n2722 & n23366 ;
  assign n23368 = n23367 ^ n21805 ^ n20473 ;
  assign n23370 = ( ~n1103 & n3739 ) | ( ~n1103 & n13495 ) | ( n3739 & n13495 ) ;
  assign n23369 = n21572 ^ n2055 ^ 1'b0 ;
  assign n23371 = n23370 ^ n23369 ^ n10390 ;
  assign n23372 = ( n11432 & n22110 ) | ( n11432 & n23371 ) | ( n22110 & n23371 ) ;
  assign n23373 = n13480 | n19171 ;
  assign n23374 = n22282 ^ n20292 ^ 1'b0 ;
  assign n23375 = n23374 ^ n22805 ^ n1709 ;
  assign n23376 = n23375 ^ n7153 ^ 1'b0 ;
  assign n23377 = n1852 | n23376 ;
  assign n23378 = ( n13384 & n14158 ) | ( n13384 & n15905 ) | ( n14158 & n15905 ) ;
  assign n23379 = n18194 ^ n13143 ^ 1'b0 ;
  assign n23380 = ( n3810 & ~n14702 ) | ( n3810 & n23379 ) | ( ~n14702 & n23379 ) ;
  assign n23383 = ( ~n2792 & n5437 ) | ( ~n2792 & n9117 ) | ( n5437 & n9117 ) ;
  assign n23384 = ( ~n9701 & n14212 ) | ( ~n9701 & n23383 ) | ( n14212 & n23383 ) ;
  assign n23381 = ( n5296 & n17354 ) | ( n5296 & ~n19636 ) | ( n17354 & ~n19636 ) ;
  assign n23382 = ( ~n3464 & n7483 ) | ( ~n3464 & n23381 ) | ( n7483 & n23381 ) ;
  assign n23385 = n23384 ^ n23382 ^ n2970 ;
  assign n23386 = n12001 & n21871 ;
  assign n23387 = n14526 ^ n3973 ^ 1'b0 ;
  assign n23388 = ( n1299 & ~n6218 ) | ( n1299 & n23387 ) | ( ~n6218 & n23387 ) ;
  assign n23389 = n1145 ^ x89 ^ 1'b0 ;
  assign n23390 = n10280 | n23389 ;
  assign n23391 = ( ~n2655 & n9982 ) | ( ~n2655 & n23390 ) | ( n9982 & n23390 ) ;
  assign n23392 = n5458 & ~n23391 ;
  assign n23393 = n23392 ^ n2860 ^ 1'b0 ;
  assign n23394 = n9186 & ~n19710 ;
  assign n23395 = ( n6929 & n8858 ) | ( n6929 & ~n12648 ) | ( n8858 & ~n12648 ) ;
  assign n23396 = ~n19443 & n23395 ;
  assign n23397 = n23019 ^ n18854 ^ n11558 ;
  assign n23398 = ( ~n5998 & n8355 ) | ( ~n5998 & n12159 ) | ( n8355 & n12159 ) ;
  assign n23399 = n23398 ^ n11116 ^ 1'b0 ;
  assign n23400 = n14923 ^ n11986 ^ n1914 ;
  assign n23401 = ~n9735 & n10562 ;
  assign n23402 = n23401 ^ n12785 ^ n3010 ;
  assign n23406 = ~n4059 & n15635 ;
  assign n23407 = ~n1338 & n23406 ;
  assign n23403 = n18221 ^ n9947 ^ n5791 ;
  assign n23404 = ( n2214 & ~n11566 ) | ( n2214 & n23403 ) | ( ~n11566 & n23403 ) ;
  assign n23405 = n8122 & ~n23404 ;
  assign n23408 = n23407 ^ n23405 ^ 1'b0 ;
  assign n23409 = ( n2853 & n20956 ) | ( n2853 & ~n23408 ) | ( n20956 & ~n23408 ) ;
  assign n23410 = n2348 ^ n2276 ^ 1'b0 ;
  assign n23411 = ( n5072 & n5909 ) | ( n5072 & n23410 ) | ( n5909 & n23410 ) ;
  assign n23412 = ( ~n186 & n10630 ) | ( ~n186 & n11470 ) | ( n10630 & n11470 ) ;
  assign n23413 = n23412 ^ n23189 ^ n2875 ;
  assign n23414 = ( n1662 & n5488 ) | ( n1662 & ~n9929 ) | ( n5488 & ~n9929 ) ;
  assign n23415 = n23414 ^ n17313 ^ n3368 ;
  assign n23416 = n14431 ^ n7916 ^ n4918 ;
  assign n23417 = n618 & ~n23416 ;
  assign n23418 = n23417 ^ n6783 ^ n6649 ;
  assign n23419 = n18460 ^ n1254 ^ 1'b0 ;
  assign n23420 = ~n7222 & n23419 ;
  assign n23421 = n6384 ^ n1230 ^ 1'b0 ;
  assign n23422 = n23420 & n23421 ;
  assign n23423 = n19615 ^ n10197 ^ n7101 ;
  assign n23424 = n8148 ^ n5141 ^ n553 ;
  assign n23425 = n9155 & n23424 ;
  assign n23426 = n1999 | n2363 ;
  assign n23427 = n23426 ^ n13062 ^ 1'b0 ;
  assign n23428 = n4885 ^ n3757 ^ n3175 ;
  assign n23429 = ( n1387 & n10852 ) | ( n1387 & n12780 ) | ( n10852 & n12780 ) ;
  assign n23430 = ( n255 & n23428 ) | ( n255 & n23429 ) | ( n23428 & n23429 ) ;
  assign n23431 = n23430 ^ n6073 ^ 1'b0 ;
  assign n23432 = n23427 & ~n23431 ;
  assign n23433 = ( n8706 & n10036 ) | ( n8706 & n23432 ) | ( n10036 & n23432 ) ;
  assign n23434 = n16445 ^ n9673 ^ 1'b0 ;
  assign n23435 = ( ~n14103 & n16956 ) | ( ~n14103 & n23434 ) | ( n16956 & n23434 ) ;
  assign n23439 = ( ~x100 & n13168 ) | ( ~x100 & n14271 ) | ( n13168 & n14271 ) ;
  assign n23440 = n23439 ^ n7429 ^ n1183 ;
  assign n23436 = ( n5598 & n6059 ) | ( n5598 & n9324 ) | ( n6059 & n9324 ) ;
  assign n23437 = n447 | n23436 ;
  assign n23438 = n9134 | n23437 ;
  assign n23441 = n23440 ^ n23438 ^ 1'b0 ;
  assign n23442 = n16840 ^ n13396 ^ n11771 ;
  assign n23443 = x0 & n3766 ;
  assign n23444 = ~n4723 & n23443 ;
  assign n23445 = n23444 ^ n11792 ^ n1928 ;
  assign n23446 = n7235 & n23445 ;
  assign n23447 = ( n2112 & n5313 ) | ( n2112 & n12410 ) | ( n5313 & n12410 ) ;
  assign n23448 = n23447 ^ n12799 ^ n4278 ;
  assign n23449 = n4979 | n23448 ;
  assign n23450 = n11834 ^ n5410 ^ n5296 ;
  assign n23451 = n23450 ^ n17505 ^ n3937 ;
  assign n23452 = n23451 ^ n6493 ^ 1'b0 ;
  assign n23453 = n15058 | n20211 ;
  assign n23454 = n23453 ^ n14169 ^ 1'b0 ;
  assign n23455 = n23454 ^ n6080 ^ n4482 ;
  assign n23456 = n23455 ^ n11563 ^ n7225 ;
  assign n23457 = ( n4951 & ~n5622 ) | ( n4951 & n23456 ) | ( ~n5622 & n23456 ) ;
  assign n23458 = ( n6535 & ~n9408 ) | ( n6535 & n11525 ) | ( ~n9408 & n11525 ) ;
  assign n23459 = n23458 ^ n16038 ^ n14222 ;
  assign n23461 = ( n380 & n1959 ) | ( n380 & n3608 ) | ( n1959 & n3608 ) ;
  assign n23462 = n20672 ^ n4609 ^ n3066 ;
  assign n23463 = n23461 & ~n23462 ;
  assign n23460 = n6792 | n13313 ;
  assign n23464 = n23463 ^ n23460 ^ 1'b0 ;
  assign n23465 = ~n2147 & n23464 ;
  assign n23466 = ~n15634 & n19653 ;
  assign n23467 = n23466 ^ n20510 ^ 1'b0 ;
  assign n23468 = n5068 ^ n3165 ^ n1159 ;
  assign n23469 = ( n5392 & n6159 ) | ( n5392 & n8328 ) | ( n6159 & n8328 ) ;
  assign n23470 = n23469 ^ n5287 ^ n3444 ;
  assign n23471 = n5665 ^ n3996 ^ n2483 ;
  assign n23472 = ( n8380 & ~n23470 ) | ( n8380 & n23471 ) | ( ~n23470 & n23471 ) ;
  assign n23473 = n19074 ^ n16833 ^ 1'b0 ;
  assign n23474 = n23473 ^ n9331 ^ n7308 ;
  assign n23475 = ( n4375 & n7232 ) | ( n4375 & n21925 ) | ( n7232 & n21925 ) ;
  assign n23476 = n661 | n12660 ;
  assign n23478 = n11832 ^ n2759 ^ 1'b0 ;
  assign n23479 = n23478 ^ n14896 ^ 1'b0 ;
  assign n23477 = n8966 & ~n10738 ;
  assign n23480 = n23479 ^ n23477 ^ 1'b0 ;
  assign n23482 = n23301 ^ n3507 ^ n1751 ;
  assign n23481 = n9032 & ~n9441 ;
  assign n23483 = n23482 ^ n23481 ^ 1'b0 ;
  assign n23484 = n23483 ^ n21748 ^ 1'b0 ;
  assign n23485 = n15476 | n23484 ;
  assign n23486 = n23485 ^ n22995 ^ n11779 ;
  assign n23487 = n23486 ^ n16357 ^ n2642 ;
  assign n23489 = n22784 ^ n17771 ^ n5241 ;
  assign n23488 = n9597 ^ n9125 ^ 1'b0 ;
  assign n23490 = n23489 ^ n23488 ^ n16216 ;
  assign n23491 = n8721 ^ n3507 ^ n937 ;
  assign n23492 = ( n7092 & n15024 ) | ( n7092 & n23491 ) | ( n15024 & n23491 ) ;
  assign n23493 = ( n6082 & n17613 ) | ( n6082 & ~n23492 ) | ( n17613 & ~n23492 ) ;
  assign n23494 = ~n12362 & n15988 ;
  assign n23495 = ~n894 & n23494 ;
  assign n23496 = n13011 ^ n9897 ^ 1'b0 ;
  assign n23497 = n23495 | n23496 ;
  assign n23498 = n23493 & ~n23497 ;
  assign n23499 = n23498 ^ n22500 ^ n13950 ;
  assign n23500 = n6435 ^ n6180 ^ 1'b0 ;
  assign n23501 = ~n14915 & n23500 ;
  assign n23502 = n19563 ^ n14646 ^ n5935 ;
  assign n23503 = n19743 ^ n17072 ^ n3855 ;
  assign n23504 = n23503 ^ n15537 ^ n5870 ;
  assign n23505 = n11781 | n20850 ;
  assign n23506 = ( ~n4731 & n17733 ) | ( ~n4731 & n18424 ) | ( n17733 & n18424 ) ;
  assign n23507 = ( n3302 & n19672 ) | ( n3302 & n23506 ) | ( n19672 & n23506 ) ;
  assign n23508 = ( ~n8599 & n14524 ) | ( ~n8599 & n20972 ) | ( n14524 & n20972 ) ;
  assign n23509 = ~n15099 & n23508 ;
  assign n23520 = n10631 | n18840 ;
  assign n23521 = n23520 ^ n2369 ^ 1'b0 ;
  assign n23515 = n9084 ^ n4961 ^ n3296 ;
  assign n23516 = n23515 ^ n9185 ^ n8549 ;
  assign n23517 = ( n209 & ~n12071 ) | ( n209 & n23516 ) | ( ~n12071 & n23516 ) ;
  assign n23511 = n19837 ^ n16559 ^ n13872 ;
  assign n23510 = n3102 & n5036 ;
  assign n23512 = n23511 ^ n23510 ^ 1'b0 ;
  assign n23513 = n7907 & ~n23512 ;
  assign n23514 = ~n4669 & n23513 ;
  assign n23518 = n23517 ^ n23514 ^ n7452 ;
  assign n23519 = ( n5888 & n12095 ) | ( n5888 & ~n23518 ) | ( n12095 & ~n23518 ) ;
  assign n23522 = n23521 ^ n23519 ^ n20416 ;
  assign n23523 = n15427 ^ n6405 ^ n5448 ;
  assign n23524 = n8238 & n23523 ;
  assign n23525 = ( n8282 & ~n19783 ) | ( n8282 & n23524 ) | ( ~n19783 & n23524 ) ;
  assign n23526 = n23525 ^ n1562 ^ 1'b0 ;
  assign n23527 = n5664 & n9202 ;
  assign n23528 = n22638 & n23527 ;
  assign n23530 = n2888 & n3273 ;
  assign n23529 = n13646 ^ n9943 ^ n4222 ;
  assign n23531 = n23530 ^ n23529 ^ 1'b0 ;
  assign n23533 = n18194 ^ n12811 ^ n10333 ;
  assign n23532 = n16459 ^ n13528 ^ n5248 ;
  assign n23534 = n23533 ^ n23532 ^ n23148 ;
  assign n23535 = n7278 ^ n5248 ^ n1340 ;
  assign n23536 = ( n16814 & n19860 ) | ( n16814 & ~n23535 ) | ( n19860 & ~n23535 ) ;
  assign n23537 = ( n18673 & ~n22450 ) | ( n18673 & n23536 ) | ( ~n22450 & n23536 ) ;
  assign n23538 = ( n5506 & n13375 ) | ( n5506 & ~n20866 ) | ( n13375 & ~n20866 ) ;
  assign n23539 = n3568 & n4225 ;
  assign n23540 = ( ~n638 & n2831 ) | ( ~n638 & n14742 ) | ( n2831 & n14742 ) ;
  assign n23541 = ( n4728 & ~n23539 ) | ( n4728 & n23540 ) | ( ~n23539 & n23540 ) ;
  assign n23542 = ( n9391 & n16818 ) | ( n9391 & n23541 ) | ( n16818 & n23541 ) ;
  assign n23543 = ( n596 & ~n18036 ) | ( n596 & n23542 ) | ( ~n18036 & n23542 ) ;
  assign n23544 = ~n16019 & n16359 ;
  assign n23545 = ( n6067 & n8089 ) | ( n6067 & ~n23544 ) | ( n8089 & ~n23544 ) ;
  assign n23546 = n4455 ^ n3466 ^ n2577 ;
  assign n23547 = n18580 ^ n17655 ^ 1'b0 ;
  assign n23548 = ~n5283 & n23547 ;
  assign n23549 = n21002 ^ n8873 ^ 1'b0 ;
  assign n23550 = n7597 & n23549 ;
  assign n23551 = n21356 ^ n5725 ^ 1'b0 ;
  assign n23552 = ( n18930 & n19790 ) | ( n18930 & n23551 ) | ( n19790 & n23551 ) ;
  assign n23553 = n23552 ^ n9224 ^ n5574 ;
  assign n23554 = n10569 ^ n6182 ^ n4069 ;
  assign n23555 = n20261 ^ n14201 ^ n12760 ;
  assign n23556 = ( ~n23021 & n23554 ) | ( ~n23021 & n23555 ) | ( n23554 & n23555 ) ;
  assign n23557 = n6932 & n9778 ;
  assign n23558 = n23557 ^ n6565 ^ 1'b0 ;
  assign n23559 = n23558 ^ n12385 ^ n1632 ;
  assign n23560 = ( n11764 & ~n17039 ) | ( n11764 & n23559 ) | ( ~n17039 & n23559 ) ;
  assign n23561 = n1753 & ~n11307 ;
  assign n23562 = n16767 & n23561 ;
  assign n23563 = n23562 ^ n4046 ^ n1194 ;
  assign n23564 = n23202 ^ n13135 ^ 1'b0 ;
  assign n23565 = ~n23563 & n23564 ;
  assign n23566 = ( n17469 & ~n22709 ) | ( n17469 & n23565 ) | ( ~n22709 & n23565 ) ;
  assign n23567 = n17471 ^ n13226 ^ n8998 ;
  assign n23568 = n15391 ^ n6989 ^ n5308 ;
  assign n23569 = n8626 & n8685 ;
  assign n23570 = n23569 ^ n8406 ^ n7988 ;
  assign n23571 = n1471 & ~n23570 ;
  assign n23572 = n3545 & n23571 ;
  assign n23573 = n2083 | n14807 ;
  assign n23574 = n23573 ^ n15489 ^ 1'b0 ;
  assign n23575 = ( ~n3119 & n3158 ) | ( ~n3119 & n8646 ) | ( n3158 & n8646 ) ;
  assign n23576 = n3508 & n23575 ;
  assign n23577 = n14076 & n23576 ;
  assign n23578 = ( ~n2182 & n8254 ) | ( ~n2182 & n22936 ) | ( n8254 & n22936 ) ;
  assign n23579 = ( n359 & n12498 ) | ( n359 & n23578 ) | ( n12498 & n23578 ) ;
  assign n23580 = ( n14063 & n14160 ) | ( n14063 & ~n19648 ) | ( n14160 & ~n19648 ) ;
  assign n23581 = n23580 ^ n18207 ^ n3897 ;
  assign n23582 = ( ~n6252 & n14188 ) | ( ~n6252 & n14976 ) | ( n14188 & n14976 ) ;
  assign n23583 = n17263 ^ n15988 ^ n7668 ;
  assign n23584 = ( n8144 & n20902 ) | ( n8144 & n23583 ) | ( n20902 & n23583 ) ;
  assign n23585 = ( n1368 & ~n4070 ) | ( n1368 & n14318 ) | ( ~n4070 & n14318 ) ;
  assign n23586 = n23585 ^ n22755 ^ n8601 ;
  assign n23587 = n23586 ^ n8111 ^ 1'b0 ;
  assign n23588 = n13697 & n23587 ;
  assign n23590 = ( n5067 & n7855 ) | ( n5067 & ~n7889 ) | ( n7855 & ~n7889 ) ;
  assign n23591 = ( n3072 & ~n18867 ) | ( n3072 & n23590 ) | ( ~n18867 & n23590 ) ;
  assign n23589 = n1077 & n15119 ;
  assign n23592 = n23591 ^ n23589 ^ 1'b0 ;
  assign n23593 = ( n7327 & n21517 ) | ( n7327 & ~n23592 ) | ( n21517 & ~n23592 ) ;
  assign n23594 = ( n7835 & n16367 ) | ( n7835 & ~n18177 ) | ( n16367 & ~n18177 ) ;
  assign n23595 = ( n3576 & ~n3888 ) | ( n3576 & n20993 ) | ( ~n3888 & n20993 ) ;
  assign n23596 = ( n3852 & n3853 ) | ( n3852 & ~n5935 ) | ( n3853 & ~n5935 ) ;
  assign n23597 = n23596 ^ n19016 ^ n6117 ;
  assign n23598 = ( ~n8701 & n23595 ) | ( ~n8701 & n23597 ) | ( n23595 & n23597 ) ;
  assign n23599 = n7887 ^ n2412 ^ 1'b0 ;
  assign n23600 = n23599 ^ n17419 ^ 1'b0 ;
  assign n23601 = ( n826 & n7798 ) | ( n826 & ~n23600 ) | ( n7798 & ~n23600 ) ;
  assign n23602 = n23601 ^ n3820 ^ n428 ;
  assign n23603 = ( n13002 & n13727 ) | ( n13002 & n17074 ) | ( n13727 & n17074 ) ;
  assign n23604 = ( n4725 & n20482 ) | ( n4725 & ~n23603 ) | ( n20482 & ~n23603 ) ;
  assign n23610 = n18621 ^ n10788 ^ n6255 ;
  assign n23605 = ( n4451 & n7582 ) | ( n4451 & ~n21291 ) | ( n7582 & ~n21291 ) ;
  assign n23606 = n23605 ^ n14884 ^ n10148 ;
  assign n23607 = ( n905 & ~n3189 ) | ( n905 & n5394 ) | ( ~n3189 & n5394 ) ;
  assign n23608 = n15287 & n23607 ;
  assign n23609 = n23606 & n23608 ;
  assign n23611 = n23610 ^ n23609 ^ 1'b0 ;
  assign n23612 = ( n5583 & n9544 ) | ( n5583 & n10722 ) | ( n9544 & n10722 ) ;
  assign n23613 = ~n14460 & n16424 ;
  assign n23614 = n13067 & n23613 ;
  assign n23615 = n14637 | n23614 ;
  assign n23618 = ( n5800 & n16872 ) | ( n5800 & ~n19310 ) | ( n16872 & ~n19310 ) ;
  assign n23616 = n7639 ^ n6130 ^ 1'b0 ;
  assign n23617 = n23616 ^ n10990 ^ n2379 ;
  assign n23619 = n23618 ^ n23617 ^ n11648 ;
  assign n23620 = n6873 ^ n4115 ^ n3480 ;
  assign n23621 = n23620 ^ n21396 ^ n18085 ;
  assign n23622 = n6244 | n6659 ;
  assign n23623 = n5442 & ~n5951 ;
  assign n23624 = n244 & n23623 ;
  assign n23625 = n7604 & ~n8549 ;
  assign n23626 = n23625 ^ n12595 ^ 1'b0 ;
  assign n23627 = ( n421 & ~n4511 ) | ( n421 & n13103 ) | ( ~n4511 & n13103 ) ;
  assign n23628 = ( n5500 & ~n11617 ) | ( n5500 & n20445 ) | ( ~n11617 & n20445 ) ;
  assign n23629 = ( n8920 & ~n23627 ) | ( n8920 & n23628 ) | ( ~n23627 & n23628 ) ;
  assign n23630 = n23629 ^ n12632 ^ n1372 ;
  assign n23631 = ( ~n5816 & n19910 ) | ( ~n5816 & n23630 ) | ( n19910 & n23630 ) ;
  assign n23632 = ( n429 & n10872 ) | ( n429 & n15065 ) | ( n10872 & n15065 ) ;
  assign n23633 = n2249 ^ n1009 ^ 1'b0 ;
  assign n23634 = ( n23209 & n23632 ) | ( n23209 & ~n23633 ) | ( n23632 & ~n23633 ) ;
  assign n23635 = n7541 ^ n7112 ^ 1'b0 ;
  assign n23636 = n2526 & n23635 ;
  assign n23637 = ~n4264 & n23636 ;
  assign n23638 = n23637 ^ n16047 ^ 1'b0 ;
  assign n23639 = n23638 ^ n18818 ^ n5365 ;
  assign n23640 = n7119 ^ n1398 ^ 1'b0 ;
  assign n23641 = n5600 ^ n2832 ^ 1'b0 ;
  assign n23642 = ~n5038 & n23641 ;
  assign n23643 = n23642 ^ n18712 ^ n772 ;
  assign n23644 = n4534 & n18366 ;
  assign n23645 = n23644 ^ n2980 ^ 1'b0 ;
  assign n23646 = n8285 ^ n5648 ^ n5306 ;
  assign n23647 = n23646 ^ n8623 ^ n430 ;
  assign n23648 = n12146 ^ n3965 ^ n2969 ;
  assign n23649 = n23648 ^ n8057 ^ n5961 ;
  assign n23658 = ( ~n9001 & n17162 ) | ( ~n9001 & n17526 ) | ( n17162 & n17526 ) ;
  assign n23655 = n9258 ^ n6724 ^ n6138 ;
  assign n23656 = n344 & ~n23655 ;
  assign n23657 = n23656 ^ n1234 ^ 1'b0 ;
  assign n23650 = n9253 ^ n5658 ^ 1'b0 ;
  assign n23651 = n5234 & n23650 ;
  assign n23652 = n23651 ^ n10827 ^ n430 ;
  assign n23653 = n7002 ^ n3965 ^ 1'b0 ;
  assign n23654 = n23652 | n23653 ;
  assign n23659 = n23658 ^ n23657 ^ n23654 ;
  assign n23665 = n17668 ^ n5808 ^ n2599 ;
  assign n23666 = ( ~n635 & n19065 ) | ( ~n635 & n23665 ) | ( n19065 & n23665 ) ;
  assign n23660 = n18078 ^ n10610 ^ n7950 ;
  assign n23661 = n915 & ~n14686 ;
  assign n23662 = n13504 ^ n6260 ^ n5849 ;
  assign n23663 = ( n8613 & n23661 ) | ( n8613 & ~n23662 ) | ( n23661 & ~n23662 ) ;
  assign n23664 = ( n7829 & n23660 ) | ( n7829 & n23663 ) | ( n23660 & n23663 ) ;
  assign n23667 = n23666 ^ n23664 ^ n21657 ;
  assign n23670 = n5574 & n10514 ;
  assign n23671 = ( n7703 & n11038 ) | ( n7703 & ~n23670 ) | ( n11038 & ~n23670 ) ;
  assign n23668 = n1333 & n23226 ;
  assign n23669 = n14117 & n23668 ;
  assign n23672 = n23671 ^ n23669 ^ 1'b0 ;
  assign n23673 = ~n2715 & n23672 ;
  assign n23674 = ( n12470 & n19190 ) | ( n12470 & ~n23673 ) | ( n19190 & ~n23673 ) ;
  assign n23675 = n1383 & n6140 ;
  assign n23676 = ( n2494 & n5513 ) | ( n2494 & n23675 ) | ( n5513 & n23675 ) ;
  assign n23677 = ~n2512 & n5239 ;
  assign n23678 = n23677 ^ n6015 ^ 1'b0 ;
  assign n23679 = ( n4356 & ~n9264 ) | ( n4356 & n12070 ) | ( ~n9264 & n12070 ) ;
  assign n23680 = n23127 ^ n10124 ^ n7157 ;
  assign n23681 = n20294 & n21692 ;
  assign n23682 = ( ~n13844 & n21545 ) | ( ~n13844 & n23681 ) | ( n21545 & n23681 ) ;
  assign n23683 = ( n2739 & ~n11306 ) | ( n2739 & n12751 ) | ( ~n11306 & n12751 ) ;
  assign n23686 = ( n844 & n948 ) | ( n844 & n3289 ) | ( n948 & n3289 ) ;
  assign n23687 = ( n8784 & n13239 ) | ( n8784 & n23686 ) | ( n13239 & n23686 ) ;
  assign n23684 = n12084 ^ n7016 ^ n3752 ;
  assign n23685 = n23684 ^ n23311 ^ n10551 ;
  assign n23688 = n23687 ^ n23685 ^ n8386 ;
  assign n23689 = n497 & n667 ;
  assign n23690 = ~n453 & n23689 ;
  assign n23691 = n10736 & ~n23690 ;
  assign n23692 = n8692 ^ n5955 ^ n4645 ;
  assign n23693 = n23692 ^ n14209 ^ n3400 ;
  assign n23694 = n23693 ^ n18613 ^ 1'b0 ;
  assign n23695 = n5207 & ~n9482 ;
  assign n23696 = n8217 & n23695 ;
  assign n23697 = ~n1990 & n23696 ;
  assign n23698 = n13963 ^ n7578 ^ n2390 ;
  assign n23699 = n13885 ^ n7773 ^ n1535 ;
  assign n23700 = n23699 ^ n17187 ^ n9719 ;
  assign n23701 = n9292 | n15162 ;
  assign n23702 = ( n10867 & n11858 ) | ( n10867 & ~n15568 ) | ( n11858 & ~n15568 ) ;
  assign n23703 = ( n9263 & n13345 ) | ( n9263 & ~n23702 ) | ( n13345 & ~n23702 ) ;
  assign n23704 = n2486 | n6519 ;
  assign n23705 = n23704 ^ n7881 ^ 1'b0 ;
  assign n23706 = n13963 & ~n23705 ;
  assign n23707 = n7226 & n23706 ;
  assign n23708 = n17999 | n18346 ;
  assign n23709 = n11481 | n12450 ;
  assign n23710 = n23708 | n23709 ;
  assign n23711 = ( n4086 & n16967 ) | ( n4086 & ~n21718 ) | ( n16967 & ~n21718 ) ;
  assign n23712 = n23711 ^ n22579 ^ n16320 ;
  assign n23713 = n21823 ^ n13695 ^ n4899 ;
  assign n23714 = n22195 ^ n19353 ^ n5005 ;
  assign n23715 = n20605 ^ n6548 ^ x91 ;
  assign n23716 = n10062 ^ n9717 ^ n978 ;
  assign n23717 = ( n7572 & n19311 ) | ( n7572 & ~n23716 ) | ( n19311 & ~n23716 ) ;
  assign n23718 = ( n4341 & n22714 ) | ( n4341 & n23717 ) | ( n22714 & n23717 ) ;
  assign n23719 = n5375 & n23718 ;
  assign n23720 = n23719 ^ n6469 ^ n5425 ;
  assign n23721 = ( ~n2688 & n3089 ) | ( ~n2688 & n10121 ) | ( n3089 & n10121 ) ;
  assign n23722 = n12583 ^ n10406 ^ n4983 ;
  assign n23723 = n23722 ^ n15780 ^ n6442 ;
  assign n23724 = ( n798 & ~n23721 ) | ( n798 & n23723 ) | ( ~n23721 & n23723 ) ;
  assign n23725 = ( ~n6551 & n17263 ) | ( ~n6551 & n23724 ) | ( n17263 & n23724 ) ;
  assign n23726 = n23310 ^ n17115 ^ 1'b0 ;
  assign n23727 = n23725 | n23726 ;
  assign n23728 = n9185 ^ n6739 ^ n1424 ;
  assign n23729 = n12942 ^ n10764 ^ 1'b0 ;
  assign n23730 = n23729 ^ n13940 ^ 1'b0 ;
  assign n23731 = n15028 & ~n23730 ;
  assign n23732 = n6361 | n23731 ;
  assign n23733 = n23732 ^ n21104 ^ n2737 ;
  assign n23734 = ( ~n6121 & n6354 ) | ( ~n6121 & n22492 ) | ( n6354 & n22492 ) ;
  assign n23735 = ( n12881 & n18190 ) | ( n12881 & n18811 ) | ( n18190 & n18811 ) ;
  assign n23736 = ~n1705 & n21412 ;
  assign n23737 = n23735 & n23736 ;
  assign n23738 = ( ~n12032 & n23734 ) | ( ~n12032 & n23737 ) | ( n23734 & n23737 ) ;
  assign n23740 = n22975 ^ n4477 ^ 1'b0 ;
  assign n23739 = n4071 & ~n7339 ;
  assign n23741 = n23740 ^ n23739 ^ 1'b0 ;
  assign n23742 = n8081 ^ n412 ^ n202 ;
  assign n23743 = n23742 ^ n11758 ^ n517 ;
  assign n23744 = n23743 ^ n12962 ^ 1'b0 ;
  assign n23745 = n15090 ^ n11424 ^ n9928 ;
  assign n23746 = n5042 ^ n507 ^ 1'b0 ;
  assign n23747 = n23745 & ~n23746 ;
  assign n23748 = n16167 ^ n12745 ^ n6329 ;
  assign n23749 = n23748 ^ n23292 ^ n16404 ;
  assign n23750 = n23749 ^ n22686 ^ n9441 ;
  assign n23751 = ( n3866 & ~n6007 ) | ( n3866 & n9181 ) | ( ~n6007 & n9181 ) ;
  assign n23752 = n23751 ^ n4515 ^ n4244 ;
  assign n23753 = n14890 ^ n9995 ^ n9567 ;
  assign n23755 = ( n491 & ~n3450 ) | ( n491 & n9001 ) | ( ~n3450 & n9001 ) ;
  assign n23756 = n23755 ^ n2444 ^ 1'b0 ;
  assign n23754 = n451 | n2285 ;
  assign n23757 = n23756 ^ n23754 ^ 1'b0 ;
  assign n23758 = ( n1818 & n23753 ) | ( n1818 & n23757 ) | ( n23753 & n23757 ) ;
  assign n23759 = n8751 ^ n8651 ^ n2902 ;
  assign n23760 = n23759 ^ n19018 ^ 1'b0 ;
  assign n23761 = n17845 ^ n16552 ^ n14516 ;
  assign n23762 = ( n4461 & n23760 ) | ( n4461 & ~n23761 ) | ( n23760 & ~n23761 ) ;
  assign n23763 = n10358 ^ n944 ^ n598 ;
  assign n23764 = n14584 ^ n8307 ^ n5667 ;
  assign n23765 = n8383 ^ n2163 ^ 1'b0 ;
  assign n23766 = n23764 & n23765 ;
  assign n23767 = ~n23515 & n23766 ;
  assign n23768 = n23767 ^ n3912 ^ 1'b0 ;
  assign n23769 = ( n15901 & ~n23763 ) | ( n15901 & n23768 ) | ( ~n23763 & n23768 ) ;
  assign n23770 = n5763 & ~n5939 ;
  assign n23777 = ( n5885 & n15803 ) | ( n5885 & ~n20385 ) | ( n15803 & ~n20385 ) ;
  assign n23771 = n22807 ^ n11450 ^ n5598 ;
  assign n23772 = n12447 ^ n3268 ^ n3220 ;
  assign n23773 = n17492 ^ n17144 ^ n15526 ;
  assign n23774 = n9696 & ~n23773 ;
  assign n23775 = n23774 ^ n7654 ^ 1'b0 ;
  assign n23776 = ( n23771 & n23772 ) | ( n23771 & ~n23775 ) | ( n23772 & ~n23775 ) ;
  assign n23778 = n23777 ^ n23776 ^ n3237 ;
  assign n23779 = ~n23770 & n23778 ;
  assign n23780 = ( n4445 & n5450 ) | ( n4445 & ~n23779 ) | ( n5450 & ~n23779 ) ;
  assign n23781 = ~n11911 & n14342 ;
  assign n23782 = n2091 & ~n14431 ;
  assign n23783 = n23782 ^ n1039 ^ 1'b0 ;
  assign n23784 = n23781 & ~n23783 ;
  assign n23786 = n1789 & n2170 ;
  assign n23785 = n7681 | n17100 ;
  assign n23787 = n23786 ^ n23785 ^ 1'b0 ;
  assign n23788 = n11106 ^ n350 ^ 1'b0 ;
  assign n23789 = n829 & n23788 ;
  assign n23790 = ( ~n4519 & n22124 ) | ( ~n4519 & n23789 ) | ( n22124 & n23789 ) ;
  assign n23791 = ~n9416 & n12519 ;
  assign n23792 = n10845 | n23791 ;
  assign n23793 = ( n2230 & n3156 ) | ( n2230 & ~n12657 ) | ( n3156 & ~n12657 ) ;
  assign n23794 = n15902 ^ n3589 ^ 1'b0 ;
  assign n23795 = n18584 ^ n11576 ^ 1'b0 ;
  assign n23796 = n13930 ^ n3081 ^ 1'b0 ;
  assign n23797 = ( ~n3466 & n8696 ) | ( ~n3466 & n23796 ) | ( n8696 & n23796 ) ;
  assign n23798 = ( ~n15139 & n23795 ) | ( ~n15139 & n23797 ) | ( n23795 & n23797 ) ;
  assign n23804 = n14914 ^ n8416 ^ n4732 ;
  assign n23803 = ( ~n7693 & n16627 ) | ( ~n7693 & n19495 ) | ( n16627 & n19495 ) ;
  assign n23805 = n23804 ^ n23803 ^ n12099 ;
  assign n23800 = n6899 ^ n2330 ^ 1'b0 ;
  assign n23801 = ~n14738 & n23800 ;
  assign n23799 = n840 & n11368 ;
  assign n23802 = n23801 ^ n23799 ^ 1'b0 ;
  assign n23806 = n23805 ^ n23802 ^ n12943 ;
  assign n23807 = n10646 ^ n10636 ^ n2799 ;
  assign n23808 = n17631 ^ n16481 ^ n1154 ;
  assign n23809 = ( n9773 & n22281 ) | ( n9773 & ~n23808 ) | ( n22281 & ~n23808 ) ;
  assign n23810 = n21095 ^ n17470 ^ n12385 ;
  assign n23811 = ( n8931 & n12730 ) | ( n8931 & n23810 ) | ( n12730 & n23810 ) ;
  assign n23812 = n17065 ^ n12784 ^ n12328 ;
  assign n23813 = ~n12653 & n23812 ;
  assign n23814 = n14711 ^ n14574 ^ 1'b0 ;
  assign n23815 = ~n21052 & n23814 ;
  assign n23816 = n2050 & n6510 ;
  assign n23817 = n7895 & n23816 ;
  assign n23818 = n23817 ^ n7746 ^ 1'b0 ;
  assign n23822 = n6366 & n14515 ;
  assign n23823 = ~n7564 & n23822 ;
  assign n23820 = n6870 ^ n4672 ^ 1'b0 ;
  assign n23821 = ~n7153 & n23820 ;
  assign n23824 = n23823 ^ n23821 ^ n17923 ;
  assign n23819 = ~n4203 & n18132 ;
  assign n23825 = n23824 ^ n23819 ^ 1'b0 ;
  assign n23826 = n23818 & n23825 ;
  assign n23827 = ~n18668 & n23826 ;
  assign n23828 = n23827 ^ n23805 ^ 1'b0 ;
  assign n23829 = n13892 | n14970 ;
  assign n23830 = n5407 & ~n23829 ;
  assign n23837 = n22207 ^ n13264 ^ 1'b0 ;
  assign n23838 = n5550 & n23837 ;
  assign n23835 = ( n1526 & n6424 ) | ( n1526 & ~n8810 ) | ( n6424 & ~n8810 ) ;
  assign n23836 = n6292 & ~n23835 ;
  assign n23833 = ( n1800 & n3236 ) | ( n1800 & ~n15403 ) | ( n3236 & ~n15403 ) ;
  assign n23831 = ~n1744 & n8451 ;
  assign n23832 = n23831 ^ n11750 ^ n3046 ;
  assign n23834 = n23833 ^ n23832 ^ n13932 ;
  assign n23839 = n23838 ^ n23836 ^ n23834 ;
  assign n23840 = n14449 ^ n5664 ^ n4405 ;
  assign n23841 = n23840 ^ n8056 ^ n1825 ;
  assign n23842 = n23841 ^ n17904 ^ n15314 ;
  assign n23843 = ( x63 & n3283 ) | ( x63 & n10383 ) | ( n3283 & n10383 ) ;
  assign n23844 = ~n9093 & n23843 ;
  assign n23845 = ( n13491 & n19571 ) | ( n13491 & n23532 ) | ( n19571 & n23532 ) ;
  assign n23846 = n14393 ^ n12277 ^ 1'b0 ;
  assign n23847 = n23846 ^ n20813 ^ n8687 ;
  assign n23848 = ( ~n11159 & n22758 ) | ( ~n11159 & n23847 ) | ( n22758 & n23847 ) ;
  assign n23849 = ~n11727 & n14881 ;
  assign n23850 = n723 & n23849 ;
  assign n23851 = n8699 & n19442 ;
  assign n23852 = ( ~n1319 & n11459 ) | ( ~n1319 & n12924 ) | ( n11459 & n12924 ) ;
  assign n23853 = n23852 ^ n3081 ^ n3054 ;
  assign n23854 = ( n14037 & ~n23851 ) | ( n14037 & n23853 ) | ( ~n23851 & n23853 ) ;
  assign n23855 = n10330 ^ n4763 ^ n4329 ;
  assign n23856 = ( n10831 & n20517 ) | ( n10831 & n23855 ) | ( n20517 & n23855 ) ;
  assign n23857 = n23856 ^ n1304 ^ 1'b0 ;
  assign n23861 = ( n1631 & ~n1709 ) | ( n1631 & n2764 ) | ( ~n1709 & n2764 ) ;
  assign n23862 = n12799 & ~n23861 ;
  assign n23858 = n2134 & n9104 ;
  assign n23859 = n23858 ^ n2274 ^ 1'b0 ;
  assign n23860 = ~n3697 & n23859 ;
  assign n23863 = n23862 ^ n23860 ^ n23304 ;
  assign n23864 = ( ~n1554 & n7665 ) | ( ~n1554 & n12951 ) | ( n7665 & n12951 ) ;
  assign n23865 = n23864 ^ n13814 ^ n10392 ;
  assign n23866 = ( ~n16466 & n21062 ) | ( ~n16466 & n23865 ) | ( n21062 & n23865 ) ;
  assign n23867 = ( n3695 & ~n17444 ) | ( n3695 & n21115 ) | ( ~n17444 & n21115 ) ;
  assign n23868 = n21092 ^ n14535 ^ n8719 ;
  assign n23869 = ( ~n11490 & n14359 ) | ( ~n11490 & n17883 ) | ( n14359 & n17883 ) ;
  assign n23870 = n23869 ^ n4927 ^ 1'b0 ;
  assign n23871 = n1368 & ~n14725 ;
  assign n23872 = ~n23870 & n23871 ;
  assign n23873 = n21405 ^ n11402 ^ 1'b0 ;
  assign n23874 = n11810 ^ n7156 ^ n2808 ;
  assign n23875 = n16079 ^ n11661 ^ n7998 ;
  assign n23876 = n21747 ^ n8731 ^ n6260 ;
  assign n23877 = ( n10875 & ~n21690 ) | ( n10875 & n23876 ) | ( ~n21690 & n23876 ) ;
  assign n23878 = n11741 ^ n7827 ^ n6645 ;
  assign n23879 = ( n804 & n3689 ) | ( n804 & n4218 ) | ( n3689 & n4218 ) ;
  assign n23880 = n23879 ^ n12914 ^ n3997 ;
  assign n23881 = n507 & n23880 ;
  assign n23882 = n23881 ^ n1823 ^ 1'b0 ;
  assign n23883 = n17481 ^ n9382 ^ n8854 ;
  assign n23884 = ( n12313 & n20906 ) | ( n12313 & n23766 ) | ( n20906 & n23766 ) ;
  assign n23885 = ( ~n4710 & n6368 ) | ( ~n4710 & n11331 ) | ( n6368 & n11331 ) ;
  assign n23886 = ( n5315 & n13526 ) | ( n5315 & n23885 ) | ( n13526 & n23885 ) ;
  assign n23887 = n14232 ^ n11015 ^ 1'b0 ;
  assign n23888 = n14228 & ~n23887 ;
  assign n23889 = n18126 ^ n16119 ^ 1'b0 ;
  assign n23890 = ( n18534 & ~n23888 ) | ( n18534 & n23889 ) | ( ~n23888 & n23889 ) ;
  assign n23891 = ( n2444 & n4017 ) | ( n2444 & n12881 ) | ( n4017 & n12881 ) ;
  assign n23892 = ( ~n4118 & n8403 ) | ( ~n4118 & n18152 ) | ( n8403 & n18152 ) ;
  assign n23893 = n10049 & n23892 ;
  assign n23894 = ~n10264 & n23893 ;
  assign n23895 = n6426 ^ n6253 ^ 1'b0 ;
  assign n23896 = n14631 | n23895 ;
  assign n23897 = n23896 ^ n4561 ^ 1'b0 ;
  assign n23898 = ~n20202 & n23897 ;
  assign n23899 = ( n23891 & n23894 ) | ( n23891 & ~n23898 ) | ( n23894 & ~n23898 ) ;
  assign n23900 = n19973 ^ n18375 ^ n9293 ;
  assign n23901 = n19704 ^ n3612 ^ n2002 ;
  assign n23902 = ( n3133 & n11686 ) | ( n3133 & ~n23901 ) | ( n11686 & ~n23901 ) ;
  assign n23903 = n14082 | n20624 ;
  assign n23904 = n23903 ^ n2304 ^ 1'b0 ;
  assign n23905 = n14809 ^ n11762 ^ n4723 ;
  assign n23906 = n23905 ^ n1300 ^ 1'b0 ;
  assign n23907 = n23904 & ~n23906 ;
  assign n23908 = ( n7796 & ~n8282 ) | ( n7796 & n14104 ) | ( ~n8282 & n14104 ) ;
  assign n23909 = ( ~n3692 & n10191 ) | ( ~n3692 & n23908 ) | ( n10191 & n23908 ) ;
  assign n23910 = ( n2175 & n8023 ) | ( n2175 & n23909 ) | ( n8023 & n23909 ) ;
  assign n23911 = n1064 | n11142 ;
  assign n23912 = n23910 | n23911 ;
  assign n23913 = ( n584 & n683 ) | ( n584 & n21364 ) | ( n683 & n21364 ) ;
  assign n23914 = n18014 & ~n18200 ;
  assign n23915 = n23914 ^ n11266 ^ 1'b0 ;
  assign n23916 = n23915 ^ n10568 ^ n9356 ;
  assign n23920 = n4419 ^ n3171 ^ 1'b0 ;
  assign n23921 = n8654 | n23920 ;
  assign n23922 = ( n5653 & ~n15366 ) | ( n5653 & n23921 ) | ( ~n15366 & n23921 ) ;
  assign n23917 = n6873 ^ n730 ^ n347 ;
  assign n23918 = n12324 ^ n7950 ^ 1'b0 ;
  assign n23919 = ~n23917 & n23918 ;
  assign n23923 = n23922 ^ n23919 ^ n14149 ;
  assign n23924 = ( n5794 & ~n6550 ) | ( n5794 & n11872 ) | ( ~n6550 & n11872 ) ;
  assign n23925 = n13558 ^ n7067 ^ n5871 ;
  assign n23927 = ( ~n3911 & n14704 ) | ( ~n3911 & n17953 ) | ( n14704 & n17953 ) ;
  assign n23926 = ~n6054 & n16386 ;
  assign n23928 = n23927 ^ n23926 ^ n10181 ;
  assign n23929 = n23928 ^ n19840 ^ 1'b0 ;
  assign n23930 = n7399 & n23929 ;
  assign n23931 = n15113 ^ n12816 ^ n11045 ;
  assign n23932 = n23931 ^ n12743 ^ n8125 ;
  assign n23933 = ( n369 & n9669 ) | ( n369 & ~n23932 ) | ( n9669 & ~n23932 ) ;
  assign n23934 = n14377 ^ n9337 ^ n7886 ;
  assign n23937 = n3230 & n17719 ;
  assign n23938 = n23937 ^ n14489 ^ 1'b0 ;
  assign n23939 = n23938 ^ n15635 ^ n10386 ;
  assign n23940 = n23939 ^ n13833 ^ 1'b0 ;
  assign n23935 = ( ~n1968 & n6915 ) | ( ~n1968 & n13189 ) | ( n6915 & n13189 ) ;
  assign n23936 = n8297 & n23935 ;
  assign n23941 = n23940 ^ n23936 ^ n21888 ;
  assign n23942 = n13534 ^ n10008 ^ n1776 ;
  assign n23943 = n17977 ^ n9632 ^ 1'b0 ;
  assign n23944 = ~n19375 & n23943 ;
  assign n23945 = ( n1904 & n4189 ) | ( n1904 & ~n9346 ) | ( n4189 & ~n9346 ) ;
  assign n23946 = n11467 ^ n3368 ^ 1'b0 ;
  assign n23947 = n19128 ^ n11545 ^ n4278 ;
  assign n23953 = ( ~n4934 & n5298 ) | ( ~n4934 & n6514 ) | ( n5298 & n6514 ) ;
  assign n23949 = n12369 ^ n11852 ^ n10089 ;
  assign n23950 = n23949 ^ n10065 ^ n7335 ;
  assign n23951 = n11032 ^ n7019 ^ 1'b0 ;
  assign n23952 = n23950 & n23951 ;
  assign n23948 = n22421 ^ n12605 ^ n1001 ;
  assign n23954 = n23953 ^ n23952 ^ n23948 ;
  assign n23955 = n10772 & ~n22648 ;
  assign n23956 = n1840 & n23955 ;
  assign n23957 = ~n893 & n5796 ;
  assign n23958 = ~n4930 & n23957 ;
  assign n23959 = n23958 ^ n16511 ^ 1'b0 ;
  assign n23960 = n14160 ^ n13699 ^ n787 ;
  assign n23961 = n23960 ^ n9821 ^ n5389 ;
  assign n23962 = ( ~n16858 & n17806 ) | ( ~n16858 & n23961 ) | ( n17806 & n23961 ) ;
  assign n23963 = ( ~n676 & n1432 ) | ( ~n676 & n19127 ) | ( n1432 & n19127 ) ;
  assign n23964 = n15629 ^ n8199 ^ 1'b0 ;
  assign n23965 = ( n9127 & ~n16959 ) | ( n9127 & n23721 ) | ( ~n16959 & n23721 ) ;
  assign n23966 = ( n729 & n14023 ) | ( n729 & ~n23965 ) | ( n14023 & ~n23965 ) ;
  assign n23967 = n17105 ^ n9033 ^ n8135 ;
  assign n23968 = ( n3334 & ~n6753 ) | ( n3334 & n23967 ) | ( ~n6753 & n23967 ) ;
  assign n23972 = n412 | n5901 ;
  assign n23973 = n23972 ^ n5668 ^ 1'b0 ;
  assign n23974 = n23973 ^ n6202 ^ x34 ;
  assign n23975 = n3814 & ~n23974 ;
  assign n23976 = n23975 ^ n10264 ^ n4645 ;
  assign n23969 = n23226 ^ n9721 ^ n1865 ;
  assign n23970 = ( ~n12800 & n15562 ) | ( ~n12800 & n23969 ) | ( n15562 & n23969 ) ;
  assign n23971 = n23970 ^ n17114 ^ n11829 ;
  assign n23977 = n23976 ^ n23971 ^ n2528 ;
  assign n23978 = ( n12723 & n23968 ) | ( n12723 & n23977 ) | ( n23968 & n23977 ) ;
  assign n23979 = n17814 ^ n5550 ^ n2631 ;
  assign n23980 = n23979 ^ n8218 ^ n6194 ;
  assign n23981 = n23980 ^ n19739 ^ n1657 ;
  assign n23982 = n23981 ^ n8006 ^ n2033 ;
  assign n23983 = n16196 & n19339 ;
  assign n23984 = ( n12485 & ~n13708 ) | ( n12485 & n23983 ) | ( ~n13708 & n23983 ) ;
  assign n23985 = ( n4381 & n5026 ) | ( n4381 & n11092 ) | ( n5026 & n11092 ) ;
  assign n23986 = n11254 ^ n8361 ^ x18 ;
  assign n23987 = n23986 ^ n1669 ^ 1'b0 ;
  assign n23988 = n3847 & n15838 ;
  assign n23989 = n15109 ^ n3051 ^ n2821 ;
  assign n23990 = n22803 ^ x5 ^ 1'b0 ;
  assign n23991 = ( n13744 & ~n17022 ) | ( n13744 & n21879 ) | ( ~n17022 & n21879 ) ;
  assign n23992 = ( n23989 & n23990 ) | ( n23989 & n23991 ) | ( n23990 & n23991 ) ;
  assign n23995 = n2957 | n14802 ;
  assign n23996 = n14229 | n23995 ;
  assign n23993 = x59 & ~n17499 ;
  assign n23994 = n14363 & n23993 ;
  assign n23997 = n23996 ^ n23994 ^ n6487 ;
  assign n23998 = n23997 ^ n20006 ^ 1'b0 ;
  assign n23999 = ( ~n2920 & n3428 ) | ( ~n2920 & n12694 ) | ( n3428 & n12694 ) ;
  assign n24000 = n14001 & n23999 ;
  assign n24001 = n24000 ^ n17675 ^ 1'b0 ;
  assign n24002 = ( n2635 & n19418 ) | ( n2635 & n24001 ) | ( n19418 & n24001 ) ;
  assign n24003 = n12146 ^ n250 ^ 1'b0 ;
  assign n24004 = ( n2461 & n19216 ) | ( n2461 & ~n24003 ) | ( n19216 & ~n24003 ) ;
  assign n24005 = n24004 ^ n19887 ^ n11965 ;
  assign n24006 = n22971 ^ n21801 ^ n13667 ;
  assign n24007 = ( n7575 & n9509 ) | ( n7575 & n10702 ) | ( n9509 & n10702 ) ;
  assign n24008 = ( ~n2891 & n4739 ) | ( ~n2891 & n15643 ) | ( n4739 & n15643 ) ;
  assign n24009 = n6840 ^ n4595 ^ n3986 ;
  assign n24010 = n6352 & n24009 ;
  assign n24011 = n24010 ^ n5549 ^ 1'b0 ;
  assign n24012 = n20239 ^ n6512 ^ 1'b0 ;
  assign n24013 = n503 & ~n24012 ;
  assign n24014 = ( n3652 & n8406 ) | ( n3652 & ~n16916 ) | ( n8406 & ~n16916 ) ;
  assign n24015 = n24014 ^ n12515 ^ 1'b0 ;
  assign n24016 = n12091 ^ n1251 ^ x101 ;
  assign n24017 = ( n17865 & n23791 ) | ( n17865 & n24016 ) | ( n23791 & n24016 ) ;
  assign n24018 = n9602 ^ n6386 ^ n4494 ;
  assign n24019 = ( n17019 & ~n20996 ) | ( n17019 & n24018 ) | ( ~n20996 & n24018 ) ;
  assign n24020 = n17914 ^ n13675 ^ n4878 ;
  assign n24021 = n18595 ^ n10946 ^ n2663 ;
  assign n24022 = n868 | n24021 ;
  assign n24024 = n4494 | n7373 ;
  assign n24023 = ( ~n3147 & n4222 ) | ( ~n3147 & n18507 ) | ( n4222 & n18507 ) ;
  assign n24025 = n24024 ^ n24023 ^ n12177 ;
  assign n24026 = n13471 ^ n6447 ^ n925 ;
  assign n24027 = n24026 ^ n18513 ^ 1'b0 ;
  assign n24028 = ( n4451 & n8528 ) | ( n4451 & ~n14878 ) | ( n8528 & ~n14878 ) ;
  assign n24029 = ( n7515 & n19382 ) | ( n7515 & ~n24028 ) | ( n19382 & ~n24028 ) ;
  assign n24030 = ( n3601 & n14996 ) | ( n3601 & ~n19134 ) | ( n14996 & ~n19134 ) ;
  assign n24031 = ( n16814 & n22913 ) | ( n16814 & ~n24030 ) | ( n22913 & ~n24030 ) ;
  assign n24035 = n5145 & ~n21018 ;
  assign n24036 = ~n15960 & n24035 ;
  assign n24033 = n12441 ^ n8313 ^ n3376 ;
  assign n24032 = ( n8839 & ~n12708 ) | ( n8839 & n18588 ) | ( ~n12708 & n18588 ) ;
  assign n24034 = n24033 ^ n24032 ^ n11274 ;
  assign n24037 = n24036 ^ n24034 ^ n13827 ;
  assign n24038 = n9845 & ~n10397 ;
  assign n24039 = ~n15302 & n24038 ;
  assign n24040 = ( n4701 & n19790 ) | ( n4701 & ~n24039 ) | ( n19790 & ~n24039 ) ;
  assign n24041 = n7040 & n8970 ;
  assign n24042 = n24041 ^ n2487 ^ 1'b0 ;
  assign n24043 = ( n1028 & ~n6417 ) | ( n1028 & n24042 ) | ( ~n6417 & n24042 ) ;
  assign n24044 = n10525 & ~n24043 ;
  assign n24045 = n4956 & n24044 ;
  assign n24046 = ( n2536 & ~n12620 ) | ( n2536 & n20251 ) | ( ~n12620 & n20251 ) ;
  assign n24049 = ( n11981 & ~n16688 ) | ( n11981 & n20064 ) | ( ~n16688 & n20064 ) ;
  assign n24047 = n8101 ^ n6777 ^ 1'b0 ;
  assign n24048 = n22312 & ~n24047 ;
  assign n24050 = n24049 ^ n24048 ^ n6553 ;
  assign n24051 = n7004 ^ n6560 ^ 1'b0 ;
  assign n24052 = ( n3020 & n9887 ) | ( n3020 & ~n24051 ) | ( n9887 & ~n24051 ) ;
  assign n24053 = ( ~n3119 & n21583 ) | ( ~n3119 & n24052 ) | ( n21583 & n24052 ) ;
  assign n24054 = n8688 ^ n3950 ^ 1'b0 ;
  assign n24055 = ( n3633 & ~n15517 ) | ( n3633 & n24054 ) | ( ~n15517 & n24054 ) ;
  assign n24056 = ( n4423 & n24053 ) | ( n4423 & ~n24055 ) | ( n24053 & ~n24055 ) ;
  assign n24057 = n3710 & ~n4109 ;
  assign n24058 = ~n4914 & n24057 ;
  assign n24059 = ( n2530 & n11850 ) | ( n2530 & ~n24058 ) | ( n11850 & ~n24058 ) ;
  assign n24060 = n24059 ^ n19641 ^ n6635 ;
  assign n24061 = n20419 ^ n12550 ^ n4890 ;
  assign n24062 = ~n7677 & n17022 ;
  assign n24063 = ~n6466 & n23659 ;
  assign n24064 = ~n3301 & n24063 ;
  assign n24065 = ( n406 & n5359 ) | ( n406 & n17046 ) | ( n5359 & n17046 ) ;
  assign n24066 = ( n9933 & ~n20224 ) | ( n9933 & n24065 ) | ( ~n20224 & n24065 ) ;
  assign n24067 = ~n23544 & n24066 ;
  assign n24068 = ~n9241 & n24067 ;
  assign n24069 = n21764 ^ n5964 ^ n5365 ;
  assign n24070 = n10628 & n10876 ;
  assign n24071 = ( n1026 & n24069 ) | ( n1026 & ~n24070 ) | ( n24069 & ~n24070 ) ;
  assign n24072 = ( n2507 & n4419 ) | ( n2507 & ~n17263 ) | ( n4419 & ~n17263 ) ;
  assign n24073 = n12223 ^ n6429 ^ x88 ;
  assign n24074 = ( ~n20076 & n24072 ) | ( ~n20076 & n24073 ) | ( n24072 & n24073 ) ;
  assign n24075 = ( n1742 & ~n5561 ) | ( n1742 & n24074 ) | ( ~n5561 & n24074 ) ;
  assign n24076 = ( ~n1788 & n1806 ) | ( ~n1788 & n4386 ) | ( n1806 & n4386 ) ;
  assign n24077 = ( ~n3650 & n12848 ) | ( ~n3650 & n24076 ) | ( n12848 & n24076 ) ;
  assign n24078 = n21813 ^ n21063 ^ n4764 ;
  assign n24080 = n10649 ^ n9834 ^ 1'b0 ;
  assign n24081 = n4724 | n24080 ;
  assign n24079 = n23755 ^ n7567 ^ 1'b0 ;
  assign n24082 = n24081 ^ n24079 ^ 1'b0 ;
  assign n24083 = n4488 ^ n3773 ^ 1'b0 ;
  assign n24084 = n24083 ^ n23021 ^ n3356 ;
  assign n24089 = n4842 | n12749 ;
  assign n24090 = n20797 & ~n24089 ;
  assign n24085 = n9491 ^ n5476 ^ n5379 ;
  assign n24086 = n24085 ^ n10633 ^ 1'b0 ;
  assign n24087 = ~n19061 & n24086 ;
  assign n24088 = ~n11528 & n24087 ;
  assign n24091 = n24090 ^ n24088 ^ 1'b0 ;
  assign n24092 = n8461 ^ n672 ^ 1'b0 ;
  assign n24093 = n24092 ^ n20438 ^ n12217 ;
  assign n24094 = n16892 ^ n7996 ^ n7886 ;
  assign n24095 = ( n2167 & n3070 ) | ( n2167 & n3564 ) | ( n3070 & n3564 ) ;
  assign n24096 = ( ~n3089 & n13040 ) | ( ~n3089 & n24095 ) | ( n13040 & n24095 ) ;
  assign n24097 = n24096 ^ n7564 ^ n3426 ;
  assign n24098 = n22024 ^ n17961 ^ n16842 ;
  assign n24099 = n162 | n4956 ;
  assign n24100 = ( n9362 & n15660 ) | ( n9362 & ~n17556 ) | ( n15660 & ~n17556 ) ;
  assign n24101 = n24100 ^ n22955 ^ n497 ;
  assign n24102 = ( n17804 & ~n21258 ) | ( n17804 & n24101 ) | ( ~n21258 & n24101 ) ;
  assign n24103 = n5248 ^ n4978 ^ n3179 ;
  assign n24104 = n6271 | n24103 ;
  assign n24105 = n20056 ^ n7024 ^ n3025 ;
  assign n24106 = ( x119 & n697 ) | ( x119 & ~n2326 ) | ( n697 & ~n2326 ) ;
  assign n24107 = ( n3879 & n10481 ) | ( n3879 & ~n24106 ) | ( n10481 & ~n24106 ) ;
  assign n24108 = n9531 & n24107 ;
  assign n24109 = ~n21866 & n24108 ;
  assign n24110 = n24109 ^ n21611 ^ n12835 ;
  assign n24113 = n20075 ^ n4474 ^ n1930 ;
  assign n24111 = n8932 & ~n14101 ;
  assign n24112 = n6664 & n24111 ;
  assign n24114 = n24113 ^ n24112 ^ n11033 ;
  assign n24115 = n18407 ^ n12800 ^ 1'b0 ;
  assign n24116 = n3488 & n7786 ;
  assign n24117 = ( n3700 & n24115 ) | ( n3700 & ~n24116 ) | ( n24115 & ~n24116 ) ;
  assign n24118 = n7976 & n14500 ;
  assign n24119 = n16776 & n24118 ;
  assign n24120 = ( ~n1631 & n17197 ) | ( ~n1631 & n24119 ) | ( n17197 & n24119 ) ;
  assign n24121 = ( n9443 & n9506 ) | ( n9443 & ~n20217 ) | ( n9506 & ~n20217 ) ;
  assign n24124 = n8775 ^ n5851 ^ n1045 ;
  assign n24123 = n19391 ^ n6411 ^ n3835 ;
  assign n24122 = n20564 ^ n7904 ^ n3173 ;
  assign n24125 = n24124 ^ n24123 ^ n24122 ;
  assign n24126 = n24125 ^ n20262 ^ n5340 ;
  assign n24127 = ~n5007 & n15690 ;
  assign n24129 = n14454 ^ n6713 ^ n2418 ;
  assign n24130 = n1940 | n24129 ;
  assign n24131 = n2353 & ~n24130 ;
  assign n24128 = n1257 & n16649 ;
  assign n24132 = n24131 ^ n24128 ^ 1'b0 ;
  assign n24133 = n24132 ^ n2603 ^ n2267 ;
  assign n24134 = n1188 & ~n22744 ;
  assign n24135 = ~n2820 & n24134 ;
  assign n24136 = n22971 ^ n7658 ^ 1'b0 ;
  assign n24137 = ( ~n753 & n2554 ) | ( ~n753 & n11768 ) | ( n2554 & n11768 ) ;
  assign n24138 = n9695 & n18039 ;
  assign n24139 = ~n24137 & n24138 ;
  assign n24140 = n24139 ^ n20764 ^ n7359 ;
  assign n24141 = n24140 ^ n19378 ^ 1'b0 ;
  assign n24142 = n21764 & n24141 ;
  assign n24151 = n2808 ^ n2708 ^ 1'b0 ;
  assign n24152 = ~n22978 & n24151 ;
  assign n24147 = n7772 ^ n5719 ^ n4220 ;
  assign n24148 = n20284 ^ n2372 ^ 1'b0 ;
  assign n24149 = n24147 & ~n24148 ;
  assign n24150 = n24149 ^ n10410 ^ n5641 ;
  assign n24153 = n24152 ^ n24150 ^ n10569 ;
  assign n24143 = ( n674 & ~n8300 ) | ( n674 & n18446 ) | ( ~n8300 & n18446 ) ;
  assign n24144 = ( n3171 & n11487 ) | ( n3171 & ~n24143 ) | ( n11487 & ~n24143 ) ;
  assign n24145 = n24144 ^ n12645 ^ n8930 ;
  assign n24146 = ( n5475 & n13439 ) | ( n5475 & ~n24145 ) | ( n13439 & ~n24145 ) ;
  assign n24154 = n24153 ^ n24146 ^ n8097 ;
  assign n24155 = n10472 ^ n2549 ^ n1480 ;
  assign n24156 = n15119 ^ n9957 ^ n8906 ;
  assign n24157 = ( n9862 & n15170 ) | ( n9862 & ~n20075 ) | ( n15170 & ~n20075 ) ;
  assign n24158 = ( n24155 & n24156 ) | ( n24155 & n24157 ) | ( n24156 & n24157 ) ;
  assign n24168 = ( ~n1284 & n1907 ) | ( ~n1284 & n11074 ) | ( n1907 & n11074 ) ;
  assign n24165 = n13375 ^ n11661 ^ n8627 ;
  assign n24166 = n3931 & n24165 ;
  assign n24159 = ( n1040 & n7551 ) | ( n1040 & ~n9043 ) | ( n7551 & ~n9043 ) ;
  assign n24160 = ( n6198 & ~n7461 ) | ( n6198 & n24159 ) | ( ~n7461 & n24159 ) ;
  assign n24161 = ( n408 & n1142 ) | ( n408 & n10335 ) | ( n1142 & n10335 ) ;
  assign n24162 = ( n18351 & n24160 ) | ( n18351 & ~n24161 ) | ( n24160 & ~n24161 ) ;
  assign n24163 = n24162 ^ n9208 ^ 1'b0 ;
  assign n24164 = n3135 & n24163 ;
  assign n24167 = n24166 ^ n24164 ^ n12036 ;
  assign n24169 = n24168 ^ n24167 ^ n14059 ;
  assign n24170 = n24169 ^ n10615 ^ n1105 ;
  assign n24171 = n13156 ^ n7096 ^ n7046 ;
  assign n24172 = n7233 ^ n3198 ^ 1'b0 ;
  assign n24173 = ( n12417 & ~n24171 ) | ( n12417 & n24172 ) | ( ~n24171 & n24172 ) ;
  assign n24174 = ( n10179 & ~n15281 ) | ( n10179 & n17544 ) | ( ~n15281 & n17544 ) ;
  assign n24175 = n24174 ^ n19213 ^ n14424 ;
  assign n24176 = n24175 ^ n13403 ^ n1588 ;
  assign n24177 = n6996 & n21813 ;
  assign n24178 = n24177 ^ n21665 ^ n17085 ;
  assign n24179 = ~n1704 & n6610 ;
  assign n24180 = n2320 & n24179 ;
  assign n24181 = n24180 ^ n17899 ^ n13010 ;
  assign n24182 = n20549 ^ n7303 ^ 1'b0 ;
  assign n24183 = n24181 | n24182 ;
  assign n24184 = n15801 ^ n15545 ^ n8646 ;
  assign n24185 = n16768 ^ n10438 ^ n4771 ;
  assign n24186 = n8465 & ~n11824 ;
  assign n24187 = ( n17899 & n24185 ) | ( n17899 & ~n24186 ) | ( n24185 & ~n24186 ) ;
  assign n24188 = ( n3276 & ~n24184 ) | ( n3276 & n24187 ) | ( ~n24184 & n24187 ) ;
  assign n24189 = ( n18934 & n24183 ) | ( n18934 & n24188 ) | ( n24183 & n24188 ) ;
  assign n24190 = n10029 ^ n5799 ^ n5092 ;
  assign n24191 = n442 & ~n24190 ;
  assign n24192 = ~n21787 & n24191 ;
  assign n24193 = n15874 ^ n10170 ^ n1262 ;
  assign n24194 = ~n3047 & n24193 ;
  assign n24198 = ( n414 & n19767 ) | ( n414 & ~n22021 ) | ( n19767 & ~n22021 ) ;
  assign n24195 = n323 & n12528 ;
  assign n24196 = n8414 & n24195 ;
  assign n24197 = n11948 | n24196 ;
  assign n24199 = n24198 ^ n24197 ^ 1'b0 ;
  assign n24200 = n7647 ^ n2532 ^ n1829 ;
  assign n24201 = n22002 ^ n1377 ^ 1'b0 ;
  assign n24202 = n12276 ^ n12229 ^ 1'b0 ;
  assign n24203 = n7469 ^ n3663 ^ 1'b0 ;
  assign n24204 = n24203 ^ n10327 ^ n2047 ;
  assign n24205 = ( n8144 & n15689 ) | ( n8144 & n24204 ) | ( n15689 & n24204 ) ;
  assign n24206 = n24205 ^ n16862 ^ n11185 ;
  assign n24207 = ( n178 & n872 ) | ( n178 & n8753 ) | ( n872 & n8753 ) ;
  assign n24208 = n19165 | n22301 ;
  assign n24209 = n12947 & ~n24208 ;
  assign n24210 = n1046 & n8342 ;
  assign n24211 = n24210 ^ n20061 ^ 1'b0 ;
  assign n24212 = ( n7602 & n24209 ) | ( n7602 & n24211 ) | ( n24209 & n24211 ) ;
  assign n24213 = ( n12818 & ~n14066 ) | ( n12818 & n24212 ) | ( ~n14066 & n24212 ) ;
  assign n24214 = ( n2119 & ~n4251 ) | ( n2119 & n7534 ) | ( ~n4251 & n7534 ) ;
  assign n24215 = n16879 & n24214 ;
  assign n24216 = n11990 & n24215 ;
  assign n24217 = n12318 ^ n11280 ^ 1'b0 ;
  assign n24218 = n6922 & ~n24217 ;
  assign n24219 = n13814 ^ n10570 ^ 1'b0 ;
  assign n24220 = n17302 ^ n10419 ^ n7943 ;
  assign n24223 = n462 & ~n15099 ;
  assign n24224 = n24223 ^ n10303 ^ 1'b0 ;
  assign n24221 = ~n6830 & n10217 ;
  assign n24222 = ~n1346 & n24221 ;
  assign n24225 = n24224 ^ n24222 ^ n19339 ;
  assign n24226 = n17788 & n19438 ;
  assign n24227 = n6520 & ~n15160 ;
  assign n24228 = n22370 & n24227 ;
  assign n24229 = ( n9734 & n19399 ) | ( n9734 & ~n24228 ) | ( n19399 & ~n24228 ) ;
  assign n24230 = ( n4292 & ~n5562 ) | ( n4292 & n11069 ) | ( ~n5562 & n11069 ) ;
  assign n24231 = n24196 ^ n2417 ^ n1281 ;
  assign n24232 = n17236 & ~n17465 ;
  assign n24233 = n14890 & n24232 ;
  assign n24234 = ( n8788 & ~n9017 ) | ( n8788 & n14250 ) | ( ~n9017 & n14250 ) ;
  assign n24235 = n8399 & ~n17603 ;
  assign n24236 = n24235 ^ n8841 ^ 1'b0 ;
  assign n24237 = n17573 & n24236 ;
  assign n24238 = n5855 & n24237 ;
  assign n24239 = ( n2721 & n23719 ) | ( n2721 & ~n24238 ) | ( n23719 & ~n24238 ) ;
  assign n24240 = ( n425 & n2906 ) | ( n425 & n15587 ) | ( n2906 & n15587 ) ;
  assign n24241 = n24240 ^ n18998 ^ n16603 ;
  assign n24247 = ( n1210 & n9347 ) | ( n1210 & n22783 ) | ( n9347 & n22783 ) ;
  assign n24243 = n4627 ^ n1886 ^ 1'b0 ;
  assign n24244 = n11189 ^ n3244 ^ n920 ;
  assign n24245 = ( n12484 & ~n24243 ) | ( n12484 & n24244 ) | ( ~n24243 & n24244 ) ;
  assign n24242 = ( n7196 & n8334 ) | ( n7196 & n18078 ) | ( n8334 & n18078 ) ;
  assign n24246 = n24245 ^ n24242 ^ 1'b0 ;
  assign n24248 = n24247 ^ n24246 ^ n4963 ;
  assign n24249 = n19252 ^ n8071 ^ n6417 ;
  assign n24250 = ( n5563 & ~n15277 ) | ( n5563 & n16644 ) | ( ~n15277 & n16644 ) ;
  assign n24251 = ( n12188 & n17220 ) | ( n12188 & ~n21059 ) | ( n17220 & ~n21059 ) ;
  assign n24252 = n14202 | n21177 ;
  assign n24253 = n8496 | n24252 ;
  assign n24257 = n11435 ^ n6220 ^ n1220 ;
  assign n24254 = n9008 ^ n7240 ^ n448 ;
  assign n24255 = ~n11806 & n12146 ;
  assign n24256 = n24254 & n24255 ;
  assign n24258 = n24257 ^ n24256 ^ n12698 ;
  assign n24259 = n3682 ^ n1470 ^ 1'b0 ;
  assign n24260 = n705 & n24259 ;
  assign n24261 = ( n8726 & n15928 ) | ( n8726 & n24260 ) | ( n15928 & n24260 ) ;
  assign n24262 = n18998 ^ n4444 ^ 1'b0 ;
  assign n24263 = n18682 ^ n18363 ^ n3872 ;
  assign n24264 = ( n10629 & n24262 ) | ( n10629 & n24263 ) | ( n24262 & n24263 ) ;
  assign n24265 = n15667 ^ n14021 ^ 1'b0 ;
  assign n24266 = ( n2294 & n5691 ) | ( n2294 & n15251 ) | ( n5691 & n15251 ) ;
  assign n24267 = n24266 ^ n6524 ^ n2699 ;
  assign n24268 = n24267 ^ n11490 ^ n11205 ;
  assign n24269 = n15273 ^ n4466 ^ 1'b0 ;
  assign n24270 = n9585 | n24269 ;
  assign n24271 = n24268 & n24270 ;
  assign n24272 = n20402 ^ n9439 ^ n3023 ;
  assign n24276 = n14623 ^ n8336 ^ n7195 ;
  assign n24275 = n18138 ^ n13504 ^ n1593 ;
  assign n24273 = n21488 ^ n2419 ^ 1'b0 ;
  assign n24274 = ~n11519 & n24273 ;
  assign n24277 = n24276 ^ n24275 ^ n24274 ;
  assign n24278 = ( n12360 & ~n24272 ) | ( n12360 & n24277 ) | ( ~n24272 & n24277 ) ;
  assign n24280 = ( n4951 & ~n5657 ) | ( n4951 & n13495 ) | ( ~n5657 & n13495 ) ;
  assign n24281 = n5856 ^ n5682 ^ n4269 ;
  assign n24282 = n24281 ^ n14281 ^ 1'b0 ;
  assign n24283 = n24280 & ~n24282 ;
  assign n24279 = ~n3315 & n5894 ;
  assign n24284 = n24283 ^ n24279 ^ 1'b0 ;
  assign n24285 = ( n2161 & n2609 ) | ( n2161 & n6885 ) | ( n2609 & n6885 ) ;
  assign n24286 = n12046 | n24285 ;
  assign n24287 = n24286 ^ n13809 ^ 1'b0 ;
  assign n24288 = n19468 ^ n18135 ^ 1'b0 ;
  assign n24289 = n24288 ^ n22677 ^ n11516 ;
  assign n24290 = ( n595 & n12728 ) | ( n595 & ~n15076 ) | ( n12728 & ~n15076 ) ;
  assign n24291 = ( n10089 & n21756 ) | ( n10089 & n24290 ) | ( n21756 & n24290 ) ;
  assign n24292 = ~n17310 & n24291 ;
  assign n24293 = n1305 & n3205 ;
  assign n24294 = n21894 & n24293 ;
  assign n24295 = n3249 ^ n243 ^ 1'b0 ;
  assign n24296 = ( ~n11173 & n24294 ) | ( ~n11173 & n24295 ) | ( n24294 & n24295 ) ;
  assign n24297 = ( n4390 & n4437 ) | ( n4390 & n4516 ) | ( n4437 & n4516 ) ;
  assign n24298 = ( n2606 & n13509 ) | ( n2606 & ~n24297 ) | ( n13509 & ~n24297 ) ;
  assign n24299 = n24298 ^ n11450 ^ 1'b0 ;
  assign n24300 = n23989 ^ n4831 ^ n1061 ;
  assign n24301 = ( n2531 & n9115 ) | ( n2531 & n24300 ) | ( n9115 & n24300 ) ;
  assign n24302 = n24301 ^ n20358 ^ n181 ;
  assign n24303 = n23492 ^ n19773 ^ 1'b0 ;
  assign n24304 = n14695 ^ n7235 ^ 1'b0 ;
  assign n24305 = ~n9215 & n24304 ;
  assign n24306 = n3585 ^ n2766 ^ n1830 ;
  assign n24307 = n24306 ^ n16177 ^ 1'b0 ;
  assign n24308 = x48 & ~n24307 ;
  assign n24309 = ( n8691 & n15487 ) | ( n8691 & ~n18766 ) | ( n15487 & ~n18766 ) ;
  assign n24310 = ~n3518 & n9261 ;
  assign n24311 = ( n2998 & n21567 ) | ( n2998 & n24310 ) | ( n21567 & n24310 ) ;
  assign n24315 = n19162 ^ n2123 ^ n774 ;
  assign n24313 = n13510 ^ n9256 ^ n4088 ;
  assign n24312 = n3683 | n6384 ;
  assign n24314 = n24313 ^ n24312 ^ 1'b0 ;
  assign n24316 = n24315 ^ n24314 ^ n10285 ;
  assign n24317 = ( n2255 & n13754 ) | ( n2255 & n24316 ) | ( n13754 & n24316 ) ;
  assign n24318 = ( ~n2464 & n7738 ) | ( ~n2464 & n13437 ) | ( n7738 & n13437 ) ;
  assign n24319 = ( n7036 & n23383 ) | ( n7036 & ~n24318 ) | ( n23383 & ~n24318 ) ;
  assign n24320 = ( ~n2666 & n18782 ) | ( ~n2666 & n24319 ) | ( n18782 & n24319 ) ;
  assign n24321 = n24320 ^ n1496 ^ 1'b0 ;
  assign n24322 = n9008 & n10553 ;
  assign n24323 = n24322 ^ n5676 ^ n956 ;
  assign n24324 = n24323 ^ n6030 ^ n5850 ;
  assign n24325 = n3188 & n19574 ;
  assign n24326 = n5814 ^ n3205 ^ 1'b0 ;
  assign n24327 = n1437 & ~n24326 ;
  assign n24328 = ( n9317 & n10622 ) | ( n9317 & n20088 ) | ( n10622 & n20088 ) ;
  assign n24329 = n13926 & n24328 ;
  assign n24330 = n24329 ^ n20838 ^ 1'b0 ;
  assign n24331 = n14985 | n20379 ;
  assign n24332 = n21129 ^ n18002 ^ 1'b0 ;
  assign n24333 = n18613 ^ n16758 ^ n11077 ;
  assign n24334 = n18452 ^ n5213 ^ 1'b0 ;
  assign n24335 = n24334 ^ n21778 ^ n3406 ;
  assign n24336 = n9846 ^ n6988 ^ n3895 ;
  assign n24337 = n2092 & ~n24336 ;
  assign n24338 = n9362 & n21647 ;
  assign n24339 = n24338 ^ n1789 ^ 1'b0 ;
  assign n24340 = n24339 ^ n12513 ^ n754 ;
  assign n24342 = n710 | n7534 ;
  assign n24341 = n14286 ^ n14196 ^ n1174 ;
  assign n24343 = n24342 ^ n24341 ^ n17157 ;
  assign n24344 = n7329 & ~n10104 ;
  assign n24345 = ( n2603 & n5886 ) | ( n2603 & ~n8285 ) | ( n5886 & ~n8285 ) ;
  assign n24346 = ( ~n7079 & n16408 ) | ( ~n7079 & n24345 ) | ( n16408 & n24345 ) ;
  assign n24347 = ( n2342 & ~n24344 ) | ( n2342 & n24346 ) | ( ~n24344 & n24346 ) ;
  assign n24350 = n7712 ^ n7698 ^ n2616 ;
  assign n24348 = n11547 ^ n10994 ^ 1'b0 ;
  assign n24349 = n8913 | n24348 ;
  assign n24351 = n24350 ^ n24349 ^ 1'b0 ;
  assign n24352 = n17844 ^ n2008 ^ n680 ;
  assign n24353 = n14480 & n24352 ;
  assign n24354 = n24353 ^ n16410 ^ 1'b0 ;
  assign n24355 = n24354 ^ n21214 ^ n16896 ;
  assign n24356 = n21095 ^ n8532 ^ n945 ;
  assign n24357 = ( n16578 & n21387 ) | ( n16578 & ~n21852 ) | ( n21387 & ~n21852 ) ;
  assign n24358 = ~n8413 & n12650 ;
  assign n24359 = n9336 & n24358 ;
  assign n24360 = n23529 ^ n16479 ^ n2859 ;
  assign n24361 = n24360 ^ n22388 ^ n7728 ;
  assign n24362 = n24361 ^ n14050 ^ 1'b0 ;
  assign n24363 = ~n12722 & n24362 ;
  assign n24364 = n4368 ^ n2989 ^ n2028 ;
  assign n24365 = n11855 ^ n3256 ^ n1268 ;
  assign n24366 = ( n5100 & ~n18037 ) | ( n5100 & n24365 ) | ( ~n18037 & n24365 ) ;
  assign n24367 = ( n6356 & ~n11902 ) | ( n6356 & n23764 ) | ( ~n11902 & n23764 ) ;
  assign n24368 = n24367 ^ n13334 ^ n8422 ;
  assign n24369 = n4586 & n12395 ;
  assign n24371 = n18190 ^ n11784 ^ n2561 ;
  assign n24370 = ~n5206 & n11989 ;
  assign n24372 = n24371 ^ n24370 ^ 1'b0 ;
  assign n24373 = ~n5122 & n24372 ;
  assign n24374 = ( n2083 & n3460 ) | ( n2083 & ~n4888 ) | ( n3460 & ~n4888 ) ;
  assign n24375 = ( n3046 & n17129 ) | ( n3046 & ~n24374 ) | ( n17129 & ~n24374 ) ;
  assign n24376 = n3879 | n5375 ;
  assign n24377 = n1004 & ~n24376 ;
  assign n24378 = n23335 ^ n19654 ^ n13083 ;
  assign n24379 = ( n13925 & n14422 ) | ( n13925 & ~n24378 ) | ( n14422 & ~n24378 ) ;
  assign n24380 = n24377 & n24379 ;
  assign n24381 = n21364 ^ n10099 ^ n6091 ;
  assign n24382 = ( n10170 & n11484 ) | ( n10170 & ~n24381 ) | ( n11484 & ~n24381 ) ;
  assign n24383 = n24382 ^ n5445 ^ n1934 ;
  assign n24384 = n9973 ^ n4708 ^ n3800 ;
  assign n24385 = n16217 ^ n15380 ^ n15019 ;
  assign n24386 = ( n4542 & ~n10843 ) | ( n4542 & n13785 ) | ( ~n10843 & n13785 ) ;
  assign n24387 = ( n6366 & n6450 ) | ( n6366 & ~n24386 ) | ( n6450 & ~n24386 ) ;
  assign n24388 = ( n254 & n1415 ) | ( n254 & ~n13126 ) | ( n1415 & ~n13126 ) ;
  assign n24389 = n24388 ^ n12390 ^ n214 ;
  assign n24390 = n22731 ^ n12461 ^ n5206 ;
  assign n24391 = ( ~n5935 & n24389 ) | ( ~n5935 & n24390 ) | ( n24389 & n24390 ) ;
  assign n24392 = n20795 ^ n1386 ^ 1'b0 ;
  assign n24393 = n5851 ^ n1034 ^ n846 ;
  assign n24394 = n24393 ^ n18790 ^ n7052 ;
  assign n24395 = n24394 ^ n16387 ^ n12470 ;
  assign n24396 = ~n8281 & n24395 ;
  assign n24397 = n13655 ^ n1343 ^ 1'b0 ;
  assign n24398 = ~n2593 & n24397 ;
  assign n24399 = ( x39 & n6610 ) | ( x39 & n7681 ) | ( n6610 & n7681 ) ;
  assign n24400 = n24399 ^ n10543 ^ 1'b0 ;
  assign n24401 = n24400 ^ n1410 ^ 1'b0 ;
  assign n24402 = n19186 ^ n18786 ^ n3759 ;
  assign n24403 = ( n4175 & ~n16638 ) | ( n4175 & n18440 ) | ( ~n16638 & n18440 ) ;
  assign n24404 = ( n3291 & n13803 ) | ( n3291 & n24403 ) | ( n13803 & n24403 ) ;
  assign n24405 = n19148 ^ n18579 ^ n1562 ;
  assign n24406 = ( n3472 & ~n6626 ) | ( n3472 & n19310 ) | ( ~n6626 & n19310 ) ;
  assign n24407 = n19407 ^ n18292 ^ n2515 ;
  assign n24408 = ( ~n1551 & n6814 ) | ( ~n1551 & n9058 ) | ( n6814 & n9058 ) ;
  assign n24409 = n24408 ^ n17670 ^ n12426 ;
  assign n24410 = n22373 | n24409 ;
  assign n24411 = n9502 ^ n9131 ^ 1'b0 ;
  assign n24412 = n24410 & n24411 ;
  assign n24415 = n1919 | n5467 ;
  assign n24413 = n18403 ^ n17966 ^ 1'b0 ;
  assign n24414 = n12959 & ~n24413 ;
  assign n24416 = n24415 ^ n24414 ^ n23242 ;
  assign n24417 = n10728 ^ n9104 ^ 1'b0 ;
  assign n24418 = n9164 ^ n3518 ^ n3315 ;
  assign n24419 = n24418 ^ n5316 ^ 1'b0 ;
  assign n24420 = n24419 ^ n15861 ^ 1'b0 ;
  assign n24421 = ( n13801 & n24417 ) | ( n13801 & ~n24420 ) | ( n24417 & ~n24420 ) ;
  assign n24422 = n5229 | n15354 ;
  assign n24423 = n10154 ^ n4599 ^ n2030 ;
  assign n24424 = n12230 & n22410 ;
  assign n24425 = n24423 & n24424 ;
  assign n24426 = n1930 & ~n24425 ;
  assign n24427 = n24426 ^ n6762 ^ 1'b0 ;
  assign n24428 = n7054 & n23891 ;
  assign n24429 = n24428 ^ n4535 ^ 1'b0 ;
  assign n24430 = ( n721 & n11992 ) | ( n721 & n12670 ) | ( n11992 & n12670 ) ;
  assign n24438 = ( ~n6186 & n14659 ) | ( ~n6186 & n20307 ) | ( n14659 & n20307 ) ;
  assign n24437 = n22557 ^ n8637 ^ n5337 ;
  assign n24439 = n24438 ^ n24437 ^ n989 ;
  assign n24435 = n8503 ^ n1249 ^ x47 ;
  assign n24431 = n140 & ~n1997 ;
  assign n24432 = n4278 & n24431 ;
  assign n24433 = n5828 | n24432 ;
  assign n24434 = n24433 ^ n21412 ^ 1'b0 ;
  assign n24436 = n24435 ^ n24434 ^ n16967 ;
  assign n24440 = n24439 ^ n24436 ^ n8795 ;
  assign n24441 = n14585 ^ n3026 ^ 1'b0 ;
  assign n24442 = n24441 ^ n13126 ^ n1174 ;
  assign n24443 = n1458 | n24442 ;
  assign n24444 = n16213 & ~n24443 ;
  assign n24445 = ( n9437 & n13143 ) | ( n9437 & ~n24444 ) | ( n13143 & ~n24444 ) ;
  assign n24446 = n11900 ^ n10155 ^ x93 ;
  assign n24447 = ( ~n7191 & n9779 ) | ( ~n7191 & n24446 ) | ( n9779 & n24446 ) ;
  assign n24448 = ( n3727 & n12137 ) | ( n3727 & ~n12674 ) | ( n12137 & ~n12674 ) ;
  assign n24449 = n7142 ^ n2405 ^ 1'b0 ;
  assign n24450 = ~n24448 & n24449 ;
  assign n24451 = n24450 ^ n20475 ^ n2651 ;
  assign n24459 = ( n1136 & n7381 ) | ( n1136 & n13775 ) | ( n7381 & n13775 ) ;
  assign n24458 = n6102 ^ x45 ^ 1'b0 ;
  assign n24456 = n18013 ^ n9941 ^ x72 ;
  assign n24457 = ( n15002 & ~n17061 ) | ( n15002 & n24456 ) | ( ~n17061 & n24456 ) ;
  assign n24460 = n24459 ^ n24458 ^ n24457 ;
  assign n24452 = n12402 ^ n7434 ^ n990 ;
  assign n24453 = n9183 & ~n24452 ;
  assign n24454 = ( n5018 & ~n11342 ) | ( n5018 & n24453 ) | ( ~n11342 & n24453 ) ;
  assign n24455 = n7940 | n24454 ;
  assign n24461 = n24460 ^ n24455 ^ 1'b0 ;
  assign n24462 = ( n5650 & n12229 ) | ( n5650 & n12925 ) | ( n12229 & n12925 ) ;
  assign n24463 = n4561 | n16360 ;
  assign n24464 = n24463 ^ n6279 ^ 1'b0 ;
  assign n24465 = ~n21505 & n24464 ;
  assign n24466 = ~n24462 & n24465 ;
  assign n24467 = n8465 ^ n3170 ^ 1'b0 ;
  assign n24468 = n526 | n24467 ;
  assign n24469 = n4973 ^ n2230 ^ n713 ;
  assign n24470 = n7113 ^ n6357 ^ n5271 ;
  assign n24471 = n24470 ^ n6616 ^ 1'b0 ;
  assign n24472 = n18696 ^ n15038 ^ n12715 ;
  assign n24473 = ( ~n1872 & n10331 ) | ( ~n1872 & n21028 ) | ( n10331 & n21028 ) ;
  assign n24474 = n21111 ^ n4624 ^ n2117 ;
  assign n24475 = n16386 ^ n12230 ^ n2933 ;
  assign n24476 = ( n6932 & n7865 ) | ( n6932 & ~n9887 ) | ( n7865 & ~n9887 ) ;
  assign n24477 = ( n7730 & n10283 ) | ( n7730 & n13801 ) | ( n10283 & n13801 ) ;
  assign n24478 = ( n1800 & n11077 ) | ( n1800 & n24477 ) | ( n11077 & n24477 ) ;
  assign n24479 = n24476 | n24478 ;
  assign n24480 = n24475 | n24479 ;
  assign n24481 = n24480 ^ n17149 ^ n13237 ;
  assign n24482 = ( n4640 & n12504 ) | ( n4640 & n14444 ) | ( n12504 & n14444 ) ;
  assign n24483 = n20034 & ~n22157 ;
  assign n24484 = ~n24482 & n24483 ;
  assign n24485 = n8068 ^ n4413 ^ x6 ;
  assign n24486 = n869 & n2993 ;
  assign n24487 = n24485 & n24486 ;
  assign n24488 = ( n2559 & ~n9616 ) | ( n2559 & n13678 ) | ( ~n9616 & n13678 ) ;
  assign n24489 = n6238 ^ n5355 ^ n4032 ;
  assign n24490 = n12495 & ~n24489 ;
  assign n24492 = n18209 ^ n4647 ^ n1790 ;
  assign n24491 = n17621 ^ n8591 ^ n6614 ;
  assign n24493 = n24492 ^ n24491 ^ n21978 ;
  assign n24494 = ( n5520 & n6643 ) | ( n5520 & n10546 ) | ( n6643 & n10546 ) ;
  assign n24495 = ( ~n19837 & n21822 ) | ( ~n19837 & n24494 ) | ( n21822 & n24494 ) ;
  assign n24496 = n14886 ^ n1854 ^ 1'b0 ;
  assign n24497 = ( ~n7442 & n8288 ) | ( ~n7442 & n12583 ) | ( n8288 & n12583 ) ;
  assign n24498 = n13101 & ~n24497 ;
  assign n24506 = ( n2235 & ~n6172 ) | ( n2235 & n17046 ) | ( ~n6172 & n17046 ) ;
  assign n24504 = ( n183 & n12367 ) | ( n183 & ~n22863 ) | ( n12367 & ~n22863 ) ;
  assign n24502 = n14098 ^ n6980 ^ n5828 ;
  assign n24503 = n24502 ^ n17123 ^ n16285 ;
  assign n24505 = n24504 ^ n24503 ^ n3324 ;
  assign n24499 = n4877 & n6829 ;
  assign n24500 = ~n1287 & n24499 ;
  assign n24501 = ( n9565 & n16280 ) | ( n9565 & ~n24500 ) | ( n16280 & ~n24500 ) ;
  assign n24507 = n24506 ^ n24505 ^ n24501 ;
  assign n24508 = n7476 ^ n5536 ^ n1110 ;
  assign n24509 = ( n6770 & n13981 ) | ( n6770 & ~n24508 ) | ( n13981 & ~n24508 ) ;
  assign n24511 = n7194 ^ n6245 ^ 1'b0 ;
  assign n24512 = ~n12996 & n24511 ;
  assign n24510 = n2131 ^ n421 ^ x86 ;
  assign n24513 = n24512 ^ n24510 ^ n1984 ;
  assign n24514 = n10952 ^ n8916 ^ 1'b0 ;
  assign n24515 = ( n1503 & n2478 ) | ( n1503 & n4073 ) | ( n2478 & n4073 ) ;
  assign n24516 = n24515 ^ n11237 ^ n729 ;
  assign n24517 = n3882 ^ n665 ^ x9 ;
  assign n24518 = n24517 ^ n22837 ^ n15582 ;
  assign n24519 = n8502 ^ n2709 ^ n240 ;
  assign n24520 = n24519 ^ n23723 ^ 1'b0 ;
  assign n24521 = n24055 & n24520 ;
  assign n24522 = n773 & n20809 ;
  assign n24523 = n3138 ^ n2496 ^ 1'b0 ;
  assign n24524 = ( n7034 & n19829 ) | ( n7034 & n24523 ) | ( n19829 & n24523 ) ;
  assign n24525 = n19873 ^ n18855 ^ n9605 ;
  assign n24526 = ( n1413 & n19439 ) | ( n1413 & ~n24525 ) | ( n19439 & ~n24525 ) ;
  assign n24529 = ( n6959 & n11736 ) | ( n6959 & n14235 ) | ( n11736 & n14235 ) ;
  assign n24528 = n7540 ^ n3173 ^ n1251 ;
  assign n24527 = ( n701 & n3943 ) | ( n701 & ~n8713 ) | ( n3943 & ~n8713 ) ;
  assign n24530 = n24529 ^ n24528 ^ n24527 ;
  assign n24531 = ( x89 & n2465 ) | ( x89 & n24530 ) | ( n2465 & n24530 ) ;
  assign n24532 = ( n3003 & n5885 ) | ( n3003 & n20654 ) | ( n5885 & n20654 ) ;
  assign n24533 = n13433 & ~n19492 ;
  assign n24534 = ( x59 & ~n4282 ) | ( x59 & n20351 ) | ( ~n4282 & n20351 ) ;
  assign n24535 = ~n16105 & n24534 ;
  assign n24536 = n5012 & n24535 ;
  assign n24537 = n23692 ^ n14157 ^ n2435 ;
  assign n24538 = ( n14884 & n24536 ) | ( n14884 & ~n24537 ) | ( n24536 & ~n24537 ) ;
  assign n24539 = ( n7998 & ~n8847 ) | ( n7998 & n18664 ) | ( ~n8847 & n18664 ) ;
  assign n24540 = n22823 ^ n14493 ^ 1'b0 ;
  assign n24541 = n24539 & ~n24540 ;
  assign n24542 = n16424 ^ n11417 ^ n10982 ;
  assign n24543 = ( n12456 & n21393 ) | ( n12456 & n24542 ) | ( n21393 & n24542 ) ;
  assign n24544 = n24543 ^ n23275 ^ n16729 ;
  assign n24548 = n4940 | n8282 ;
  assign n24545 = n19665 ^ n9544 ^ 1'b0 ;
  assign n24546 = ( ~n6225 & n7634 ) | ( ~n6225 & n24545 ) | ( n7634 & n24545 ) ;
  assign n24547 = n24546 ^ n16883 ^ n1484 ;
  assign n24549 = n24548 ^ n24547 ^ n9721 ;
  assign n24550 = n10221 & n10744 ;
  assign n24551 = n24550 ^ n6957 ^ 1'b0 ;
  assign n24552 = n24551 ^ n16782 ^ n6204 ;
  assign n24553 = n20142 ^ n13864 ^ n12583 ;
  assign n24554 = n24553 ^ n13172 ^ n12153 ;
  assign n24555 = n24554 ^ n20270 ^ n4073 ;
  assign n24556 = n12887 ^ n12724 ^ n10008 ;
  assign n24557 = n15728 ^ n3617 ^ 1'b0 ;
  assign n24558 = ( ~n995 & n11885 ) | ( ~n995 & n17204 ) | ( n11885 & n17204 ) ;
  assign n24559 = n8655 ^ n526 ^ 1'b0 ;
  assign n24560 = n24558 & n24559 ;
  assign n24561 = ( n15569 & n18270 ) | ( n15569 & n20775 ) | ( n18270 & n20775 ) ;
  assign n24562 = ( n428 & n2605 ) | ( n428 & ~n10091 ) | ( n2605 & ~n10091 ) ;
  assign n24563 = n24562 ^ n23307 ^ n9197 ;
  assign n24564 = n24349 ^ n1911 ^ 1'b0 ;
  assign n24565 = n11847 | n17527 ;
  assign n24566 = n2071 | n24565 ;
  assign n24567 = n24566 ^ n19421 ^ n17041 ;
  assign n24568 = ( n2011 & ~n2938 ) | ( n2011 & n13651 ) | ( ~n2938 & n13651 ) ;
  assign n24569 = n462 & n1820 ;
  assign n24570 = n24569 ^ n16443 ^ 1'b0 ;
  assign n24571 = ( ~n4160 & n20817 ) | ( ~n4160 & n24570 ) | ( n20817 & n24570 ) ;
  assign n24572 = ~n18323 & n24571 ;
  assign n24573 = n14992 ^ n668 ^ n527 ;
  assign n24574 = n3217 & ~n10738 ;
  assign n24575 = n24574 ^ n17140 ^ n2747 ;
  assign n24576 = n24575 ^ n20681 ^ n958 ;
  assign n24577 = n24576 ^ n4625 ^ 1'b0 ;
  assign n24578 = ( n5375 & ~n24573 ) | ( n5375 & n24577 ) | ( ~n24573 & n24577 ) ;
  assign n24579 = n20972 ^ n586 ^ 1'b0 ;
  assign n24580 = ( n12775 & n24113 ) | ( n12775 & n24579 ) | ( n24113 & n24579 ) ;
  assign n24581 = n18510 ^ n16686 ^ n8128 ;
  assign n24582 = n9912 & ~n24581 ;
  assign n24583 = ( n8297 & ~n14640 ) | ( n8297 & n24582 ) | ( ~n14640 & n24582 ) ;
  assign n24584 = ( n8414 & ~n10508 ) | ( n8414 & n24583 ) | ( ~n10508 & n24583 ) ;
  assign n24585 = n576 & n22768 ;
  assign n24586 = n5058 ^ n4838 ^ n3397 ;
  assign n24587 = ( ~x107 & n17379 ) | ( ~x107 & n24586 ) | ( n17379 & n24586 ) ;
  assign n24588 = n12728 ^ n7269 ^ n432 ;
  assign n24589 = n24588 ^ n22500 ^ n18327 ;
  assign n24590 = n24589 ^ n6571 ^ n3136 ;
  assign n24591 = ( ~n5293 & n11985 ) | ( ~n5293 & n19922 ) | ( n11985 & n19922 ) ;
  assign n24592 = ( n988 & n9783 ) | ( n988 & ~n24591 ) | ( n9783 & ~n24591 ) ;
  assign n24593 = n9761 ^ n6148 ^ x68 ;
  assign n24594 = ( n3040 & n10652 ) | ( n3040 & n24593 ) | ( n10652 & n24593 ) ;
  assign n24595 = n15796 ^ n3976 ^ 1'b0 ;
  assign n24596 = n3702 | n24595 ;
  assign n24597 = n1865 & n15701 ;
  assign n24598 = n24597 ^ n8365 ^ 1'b0 ;
  assign n24599 = n3050 & ~n24598 ;
  assign n24600 = n2835 & ~n9113 ;
  assign n24604 = n7956 & n10589 ;
  assign n24605 = n24604 ^ n7945 ^ 1'b0 ;
  assign n24601 = x69 & ~n9931 ;
  assign n24602 = n24601 ^ n3191 ^ 1'b0 ;
  assign n24603 = ( n3466 & n5550 ) | ( n3466 & ~n24602 ) | ( n5550 & ~n24602 ) ;
  assign n24606 = n24605 ^ n24603 ^ n20641 ;
  assign n24607 = ~n2039 & n9592 ;
  assign n24608 = n24607 ^ n17237 ^ 1'b0 ;
  assign n24609 = ( ~n1611 & n22265 ) | ( ~n1611 & n24608 ) | ( n22265 & n24608 ) ;
  assign n24610 = n7675 ^ n3400 ^ n2901 ;
  assign n24611 = n24610 ^ n16026 ^ 1'b0 ;
  assign n24612 = n6757 | n8742 ;
  assign n24613 = n24612 ^ n918 ^ 1'b0 ;
  assign n24614 = n12301 | n18828 ;
  assign n24615 = n24614 ^ n21282 ^ n9097 ;
  assign n24616 = n7377 | n24615 ;
  assign n24617 = n24613 | n24616 ;
  assign n24618 = n8573 & n22476 ;
  assign n24619 = n5724 & ~n8791 ;
  assign n24620 = n24619 ^ n11949 ^ 1'b0 ;
  assign n24621 = n16369 ^ n7092 ^ n6868 ;
  assign n24622 = ( n9205 & ~n9658 ) | ( n9205 & n24621 ) | ( ~n9658 & n24621 ) ;
  assign n24623 = n19018 ^ n8947 ^ n7981 ;
  assign n24624 = ( ~n8024 & n23444 ) | ( ~n8024 & n24623 ) | ( n23444 & n24623 ) ;
  assign n24632 = n2664 ^ n2608 ^ n2449 ;
  assign n24633 = n24632 ^ n5585 ^ n738 ;
  assign n24630 = n4326 | n12092 ;
  assign n24631 = n2727 | n24630 ;
  assign n24634 = n24633 ^ n24631 ^ n12049 ;
  assign n24627 = n12453 ^ n3170 ^ 1'b0 ;
  assign n24628 = n1636 & n24627 ;
  assign n24625 = n12318 ^ n10197 ^ n5036 ;
  assign n24626 = ( x59 & n1464 ) | ( x59 & ~n24625 ) | ( n1464 & ~n24625 ) ;
  assign n24629 = n24628 ^ n24626 ^ n20595 ;
  assign n24635 = n24634 ^ n24629 ^ n20725 ;
  assign n24636 = ( n896 & n6214 ) | ( n896 & ~n24635 ) | ( n6214 & ~n24635 ) ;
  assign n24637 = n2388 | n16721 ;
  assign n24638 = n3028 | n24637 ;
  assign n24639 = n5090 ^ n763 ^ 1'b0 ;
  assign n24640 = n4678 & ~n24639 ;
  assign n24641 = ~n19734 & n24640 ;
  assign n24642 = n24641 ^ n6340 ^ 1'b0 ;
  assign n24643 = ( n6999 & ~n16893 ) | ( n6999 & n19981 ) | ( ~n16893 & n19981 ) ;
  assign n24644 = n24643 ^ n4371 ^ 1'b0 ;
  assign n24645 = n17136 ^ n9756 ^ n4290 ;
  assign n24646 = n17774 ^ n14337 ^ 1'b0 ;
  assign n24647 = n24646 ^ n14638 ^ n4320 ;
  assign n24648 = n15272 ^ n13108 ^ n2444 ;
  assign n24649 = n24648 ^ n18408 ^ n855 ;
  assign n24650 = n8036 ^ n6590 ^ n6396 ;
  assign n24651 = n9732 | n19366 ;
  assign n24652 = ( n4253 & n24650 ) | ( n4253 & ~n24651 ) | ( n24650 & ~n24651 ) ;
  assign n24653 = n18074 ^ n17202 ^ n5800 ;
  assign n24654 = n5398 ^ n1386 ^ 1'b0 ;
  assign n24655 = ~n14076 & n24654 ;
  assign n24656 = n765 & ~n16085 ;
  assign n24657 = n24656 ^ n4975 ^ 1'b0 ;
  assign n24658 = ( n3458 & n12059 ) | ( n3458 & n14211 ) | ( n12059 & n14211 ) ;
  assign n24660 = n13448 ^ n10467 ^ n1777 ;
  assign n24659 = ( n2156 & ~n14989 ) | ( n2156 & n19574 ) | ( ~n14989 & n19574 ) ;
  assign n24661 = n24660 ^ n24659 ^ n2504 ;
  assign n24662 = n20972 ^ n14126 ^ 1'b0 ;
  assign n24663 = n1554 & ~n24662 ;
  assign n24664 = n24663 ^ n23224 ^ n12848 ;
  assign n24665 = n23831 ^ n13412 ^ n10532 ;
  assign n24666 = n24665 ^ n896 ^ 1'b0 ;
  assign n24674 = n20140 ^ n3973 ^ 1'b0 ;
  assign n24671 = ~x55 & n10593 ;
  assign n24672 = n24671 ^ n14787 ^ 1'b0 ;
  assign n24667 = n3122 | n8642 ;
  assign n24668 = n18857 & ~n24667 ;
  assign n24669 = n16473 | n24668 ;
  assign n24670 = n24669 ^ n7080 ^ 1'b0 ;
  assign n24673 = n24672 ^ n24670 ^ n20122 ;
  assign n24675 = n24674 ^ n24673 ^ n21686 ;
  assign n24676 = ( ~n15361 & n19326 ) | ( ~n15361 & n20610 ) | ( n19326 & n20610 ) ;
  assign n24677 = n7620 | n7668 ;
  assign n24678 = ( n10730 & n15895 ) | ( n10730 & n24677 ) | ( n15895 & n24677 ) ;
  assign n24679 = n800 & n11820 ;
  assign n24680 = n9542 ^ n5137 ^ 1'b0 ;
  assign n24681 = ~n2783 & n3276 ;
  assign n24682 = n24681 ^ n24389 ^ 1'b0 ;
  assign n24683 = ( n626 & n4290 ) | ( n626 & ~n18878 ) | ( n4290 & ~n18878 ) ;
  assign n24684 = ( ~n3108 & n20225 ) | ( ~n3108 & n24683 ) | ( n20225 & n24683 ) ;
  assign n24685 = ( n8785 & ~n14791 ) | ( n8785 & n17702 ) | ( ~n14791 & n17702 ) ;
  assign n24686 = n20459 & ~n24685 ;
  assign n24687 = ( x52 & ~n276 ) | ( x52 & n739 ) | ( ~n276 & n739 ) ;
  assign n24688 = n24687 ^ n2409 ^ 1'b0 ;
  assign n24689 = n19127 ^ n13754 ^ n12650 ;
  assign n24690 = n24689 ^ n19439 ^ n3564 ;
  assign n24691 = n2258 ^ n2164 ^ 1'b0 ;
  assign n24692 = n14800 & ~n24691 ;
  assign n24693 = n24319 ^ n17006 ^ n10884 ;
  assign n24694 = n5676 | n7164 ;
  assign n24695 = ( n1889 & ~n8256 ) | ( n1889 & n22561 ) | ( ~n8256 & n22561 ) ;
  assign n24696 = ( n5440 & n7324 ) | ( n5440 & ~n13220 ) | ( n7324 & ~n13220 ) ;
  assign n24697 = n2770 | n7312 ;
  assign n24698 = n3362 & n24697 ;
  assign n24699 = n24698 ^ n7074 ^ 1'b0 ;
  assign n24700 = ( n3814 & n8323 ) | ( n3814 & ~n24699 ) | ( n8323 & ~n24699 ) ;
  assign n24701 = ( n3643 & ~n10030 ) | ( n3643 & n24700 ) | ( ~n10030 & n24700 ) ;
  assign n24702 = n12996 ^ n3068 ^ n524 ;
  assign n24703 = n14966 ^ n14388 ^ n7807 ;
  assign n24704 = n24703 ^ n23198 ^ n9397 ;
  assign n24705 = ( n2090 & n15160 ) | ( n2090 & ~n24704 ) | ( n15160 & ~n24704 ) ;
  assign n24706 = ( n24701 & ~n24702 ) | ( n24701 & n24705 ) | ( ~n24702 & n24705 ) ;
  assign n24707 = n2068 & n18786 ;
  assign n24708 = n24707 ^ n7091 ^ 1'b0 ;
  assign n24709 = n24708 ^ n20986 ^ n14937 ;
  assign n24710 = n4543 ^ n2549 ^ 1'b0 ;
  assign n24711 = n18694 & n19627 ;
  assign n24712 = n24711 ^ n17819 ^ n12050 ;
  assign n24713 = ( n4162 & n8145 ) | ( n4162 & n24712 ) | ( n8145 & n24712 ) ;
  assign n24714 = ( ~n13114 & n24710 ) | ( ~n13114 & n24713 ) | ( n24710 & n24713 ) ;
  assign n24716 = n1038 ^ n611 ^ n458 ;
  assign n24717 = n24716 ^ n21140 ^ n7962 ;
  assign n24715 = ( n6977 & n15178 ) | ( n6977 & n23927 ) | ( n15178 & n23927 ) ;
  assign n24718 = n24717 ^ n24715 ^ n21874 ;
  assign n24719 = n24718 ^ n15575 ^ n6945 ;
  assign n24720 = ( ~n1721 & n12520 ) | ( ~n1721 & n23580 ) | ( n12520 & n23580 ) ;
  assign n24721 = n20179 ^ n18657 ^ n8545 ;
  assign n24722 = n14352 ^ n13800 ^ n1752 ;
  assign n24723 = ( ~n9750 & n15458 ) | ( ~n9750 & n19867 ) | ( n15458 & n19867 ) ;
  assign n24724 = ( ~n9430 & n13200 ) | ( ~n9430 & n14858 ) | ( n13200 & n14858 ) ;
  assign n24725 = ( n5687 & n12119 ) | ( n5687 & n24724 ) | ( n12119 & n24724 ) ;
  assign n24726 = n507 & n6800 ;
  assign n24729 = n12187 ^ n3219 ^ n563 ;
  assign n24727 = n287 & n17187 ;
  assign n24728 = ~n7721 & n24727 ;
  assign n24730 = n24729 ^ n24728 ^ n4948 ;
  assign n24731 = ~n2822 & n20957 ;
  assign n24732 = n24731 ^ n23013 ^ 1'b0 ;
  assign n24733 = ( n1610 & n5407 ) | ( n1610 & n24732 ) | ( n5407 & n24732 ) ;
  assign n24734 = n14402 ^ n4425 ^ 1'b0 ;
  assign n24735 = ~n24733 & n24734 ;
  assign n24736 = ( ~n11928 & n24730 ) | ( ~n11928 & n24735 ) | ( n24730 & n24735 ) ;
  assign n24737 = n22701 ^ n10193 ^ n8187 ;
  assign n24738 = n4203 ^ n2890 ^ n348 ;
  assign n24739 = n9734 ^ n8986 ^ n6894 ;
  assign n24740 = ( n12581 & n22607 ) | ( n12581 & n24739 ) | ( n22607 & n24739 ) ;
  assign n24741 = n10598 ^ n8932 ^ n8039 ;
  assign n24742 = n24741 ^ n9400 ^ 1'b0 ;
  assign n24743 = n23640 ^ n4627 ^ 1'b0 ;
  assign n24744 = n8146 & ~n24743 ;
  assign n24745 = n21768 ^ n21653 ^ n15385 ;
  assign n24746 = n6405 ^ x40 ^ 1'b0 ;
  assign n24747 = n2118 & n24746 ;
  assign n24748 = n24747 ^ n14051 ^ 1'b0 ;
  assign n24749 = n21921 ^ n19930 ^ n5134 ;
  assign n24750 = n14731 ^ n12554 ^ n5870 ;
  assign n24751 = ( n2086 & n7757 ) | ( n2086 & n14336 ) | ( n7757 & n14336 ) ;
  assign n24752 = n11026 & ~n21503 ;
  assign n24753 = ~x64 & n24752 ;
  assign n24754 = n17736 ^ n1384 ^ 1'b0 ;
  assign n24755 = n23862 & ~n24754 ;
  assign n24756 = n13154 | n17992 ;
  assign n24757 = n8821 ^ n8219 ^ 1'b0 ;
  assign n24758 = ( n1765 & n6761 ) | ( n1765 & ~n7609 ) | ( n6761 & ~n7609 ) ;
  assign n24759 = n24758 ^ n20818 ^ n19782 ;
  assign n24761 = n5532 ^ n2240 ^ 1'b0 ;
  assign n24762 = n15901 | n24761 ;
  assign n24760 = ( n14164 & n15319 ) | ( n14164 & n22790 ) | ( n15319 & n22790 ) ;
  assign n24763 = n24762 ^ n24760 ^ n7824 ;
  assign n24764 = n24763 ^ n23700 ^ n16578 ;
  assign n24765 = n14768 | n24313 ;
  assign n24766 = n18013 & ~n24765 ;
  assign n24767 = n24766 ^ n17601 ^ n11213 ;
  assign n24770 = n2461 | n14991 ;
  assign n24771 = n7445 | n24770 ;
  assign n24772 = n24771 ^ n15519 ^ n9120 ;
  assign n24768 = n11796 ^ n6377 ^ 1'b0 ;
  assign n24769 = n24768 ^ n20363 ^ n2892 ;
  assign n24773 = n24772 ^ n24769 ^ n7481 ;
  assign n24774 = n11635 ^ n4535 ^ n3905 ;
  assign n24775 = n19595 ^ n6870 ^ 1'b0 ;
  assign n24776 = ( n17174 & n24774 ) | ( n17174 & ~n24775 ) | ( n24774 & ~n24775 ) ;
  assign n24777 = ( ~n4399 & n6087 ) | ( ~n4399 & n8787 ) | ( n6087 & n8787 ) ;
  assign n24778 = n407 & n5093 ;
  assign n24779 = n24778 ^ n4304 ^ 1'b0 ;
  assign n24780 = ( n15873 & n19733 ) | ( n15873 & n24779 ) | ( n19733 & n24779 ) ;
  assign n24781 = ( n2849 & n20788 ) | ( n2849 & n24780 ) | ( n20788 & n24780 ) ;
  assign n24782 = n2464 & n3485 ;
  assign n24783 = n24782 ^ n6586 ^ 1'b0 ;
  assign n24784 = ( ~n11396 & n18335 ) | ( ~n11396 & n24783 ) | ( n18335 & n24783 ) ;
  assign n24785 = n10708 ^ n3382 ^ n1972 ;
  assign n24786 = n24785 ^ n23265 ^ n10462 ;
  assign n24787 = ( n3384 & ~n18370 ) | ( n3384 & n19236 ) | ( ~n18370 & n19236 ) ;
  assign n24788 = ( ~n3597 & n14342 ) | ( ~n3597 & n24787 ) | ( n14342 & n24787 ) ;
  assign n24789 = n24788 ^ n8576 ^ 1'b0 ;
  assign n24790 = n14313 | n24789 ;
  assign n24791 = n4299 ^ n3750 ^ 1'b0 ;
  assign n24792 = ( n4631 & n19685 ) | ( n4631 & n24791 ) | ( n19685 & n24791 ) ;
  assign n24793 = x105 & ~n6466 ;
  assign n24794 = n4278 & n24793 ;
  assign n24795 = n1659 & ~n3409 ;
  assign n24796 = ( n6499 & n24794 ) | ( n6499 & ~n24795 ) | ( n24794 & ~n24795 ) ;
  assign n24797 = n19282 ^ n8416 ^ 1'b0 ;
  assign n24798 = n834 & n24797 ;
  assign n24799 = ( n6773 & n17419 ) | ( n6773 & ~n24798 ) | ( n17419 & ~n24798 ) ;
  assign n24800 = ( n7294 & n8428 ) | ( n7294 & n10942 ) | ( n8428 & n10942 ) ;
  assign n24801 = n24800 ^ n10242 ^ 1'b0 ;
  assign n24802 = n19234 & n24801 ;
  assign n24803 = ( ~n10971 & n18416 ) | ( ~n10971 & n24802 ) | ( n18416 & n24802 ) ;
  assign n24804 = ( n11330 & n14751 ) | ( n11330 & ~n17071 ) | ( n14751 & ~n17071 ) ;
  assign n24805 = n22815 ^ n18973 ^ n6801 ;
  assign n24806 = n19725 & n21350 ;
  assign n24807 = n24806 ^ n12883 ^ 1'b0 ;
  assign n24808 = n1647 | n18633 ;
  assign n24809 = ( n14664 & ~n20475 ) | ( n14664 & n24808 ) | ( ~n20475 & n24808 ) ;
  assign n24810 = n7921 & ~n24809 ;
  assign n24811 = ~n9922 & n24810 ;
  assign n24812 = n16601 ^ n9690 ^ 1'b0 ;
  assign n24813 = ~n12544 & n24812 ;
  assign n24814 = ( ~n10788 & n11155 ) | ( ~n10788 & n17496 ) | ( n11155 & n17496 ) ;
  assign n24815 = ( n1344 & n2705 ) | ( n1344 & n4577 ) | ( n2705 & n4577 ) ;
  assign n24816 = n3264 & n9392 ;
  assign n24817 = n4135 | n7053 ;
  assign n24818 = x125 & ~n6113 ;
  assign n24819 = n24818 ^ n3467 ^ 1'b0 ;
  assign n24820 = ( n8276 & n13940 ) | ( n8276 & ~n24819 ) | ( n13940 & ~n24819 ) ;
  assign n24821 = n24820 ^ n22765 ^ n2093 ;
  assign n24822 = ( ~n24816 & n24817 ) | ( ~n24816 & n24821 ) | ( n24817 & n24821 ) ;
  assign n24823 = ( n2749 & ~n8820 ) | ( n2749 & n21339 ) | ( ~n8820 & n21339 ) ;
  assign n24824 = n22370 ^ n16926 ^ n3948 ;
  assign n24825 = n24824 ^ n19544 ^ n2559 ;
  assign n24826 = ( n8608 & n24823 ) | ( n8608 & n24825 ) | ( n24823 & n24825 ) ;
  assign n24827 = n6424 ^ n3057 ^ 1'b0 ;
  assign n24828 = n10760 | n24827 ;
  assign n24829 = n560 & ~n3659 ;
  assign n24830 = ~n2107 & n24829 ;
  assign n24831 = n24828 & n24830 ;
  assign n24832 = ( n6567 & ~n22521 ) | ( n6567 & n24831 ) | ( ~n22521 & n24831 ) ;
  assign n24833 = n4810 & n7335 ;
  assign n24834 = n24833 ^ n3968 ^ 1'b0 ;
  assign n24835 = n3700 & ~n6045 ;
  assign n24836 = n24835 ^ n7370 ^ 1'b0 ;
  assign n24837 = n4434 ^ n1117 ^ 1'b0 ;
  assign n24838 = ( n8640 & n11985 ) | ( n8640 & ~n24837 ) | ( n11985 & ~n24837 ) ;
  assign n24839 = ( n12994 & ~n22459 ) | ( n12994 & n24838 ) | ( ~n22459 & n24838 ) ;
  assign n24840 = ~n1178 & n19392 ;
  assign n24841 = ~n12666 & n24840 ;
  assign n24842 = n24841 ^ n14163 ^ n6366 ;
  assign n24843 = n12689 ^ n4653 ^ n593 ;
  assign n24844 = n24843 ^ n10333 ^ n9801 ;
  assign n24845 = n24844 ^ n19828 ^ n8823 ;
  assign n24846 = ~n7767 & n11227 ;
  assign n24847 = ~n13791 & n24846 ;
  assign n24849 = n14725 ^ n11990 ^ 1'b0 ;
  assign n24850 = ( n5411 & n15574 ) | ( n5411 & ~n24849 ) | ( n15574 & ~n24849 ) ;
  assign n24851 = n24850 ^ n14335 ^ n8057 ;
  assign n24852 = ( n4369 & n18675 ) | ( n4369 & n24851 ) | ( n18675 & n24851 ) ;
  assign n24853 = n24852 ^ n16685 ^ n8197 ;
  assign n24848 = ~n2677 & n8281 ;
  assign n24854 = n24853 ^ n24848 ^ 1'b0 ;
  assign n24855 = n24854 ^ n6020 ^ n5955 ;
  assign n24856 = n3567 ^ n543 ^ 1'b0 ;
  assign n24857 = n545 | n24856 ;
  assign n24858 = n4236 | n10667 ;
  assign n24859 = n24858 ^ n13917 ^ 1'b0 ;
  assign n24860 = ( n15898 & n16709 ) | ( n15898 & n18128 ) | ( n16709 & n18128 ) ;
  assign n24861 = ( n5980 & n10728 ) | ( n5980 & n24860 ) | ( n10728 & n24860 ) ;
  assign n24862 = ( n24857 & n24859 ) | ( n24857 & ~n24861 ) | ( n24859 & ~n24861 ) ;
  assign n24863 = ( n142 & n4006 ) | ( n142 & n23439 ) | ( n4006 & n23439 ) ;
  assign n24864 = ( n5317 & n11011 ) | ( n5317 & n16513 ) | ( n11011 & n16513 ) ;
  assign n24867 = ( n1123 & n3119 ) | ( n1123 & n13892 ) | ( n3119 & n13892 ) ;
  assign n24866 = ( ~n8329 & n11942 ) | ( ~n8329 & n12555 ) | ( n11942 & n12555 ) ;
  assign n24868 = n24867 ^ n24866 ^ n14997 ;
  assign n24869 = n24868 ^ n21789 ^ n7185 ;
  assign n24865 = n19226 ^ n5000 ^ x87 ;
  assign n24870 = n24869 ^ n24865 ^ n17728 ;
  assign n24871 = n6649 ^ n5041 ^ n3678 ;
  assign n24872 = n3651 & ~n14164 ;
  assign n24873 = n24871 & n24872 ;
  assign n24874 = n24729 ^ n23021 ^ n5464 ;
  assign n24875 = ( ~n23896 & n24242 ) | ( ~n23896 & n24874 ) | ( n24242 & n24874 ) ;
  assign n24876 = ( ~n7988 & n19707 ) | ( ~n7988 & n21765 ) | ( n19707 & n21765 ) ;
  assign n24877 = n8072 ^ n3197 ^ n1333 ;
  assign n24878 = n24877 ^ n8399 ^ n4860 ;
  assign n24879 = n20795 ^ n20415 ^ n8413 ;
  assign n24880 = n5399 ^ n2084 ^ 1'b0 ;
  assign n24881 = n3493 & n24880 ;
  assign n24882 = n13557 | n24881 ;
  assign n24883 = n5465 & ~n20540 ;
  assign n24884 = ( ~n14120 & n24882 ) | ( ~n14120 & n24883 ) | ( n24882 & n24883 ) ;
  assign n24885 = ( n1576 & n2506 ) | ( n1576 & ~n2579 ) | ( n2506 & ~n2579 ) ;
  assign n24886 = ( n1470 & ~n1912 ) | ( n1470 & n4909 ) | ( ~n1912 & n4909 ) ;
  assign n24887 = ( ~n6310 & n24885 ) | ( ~n6310 & n24886 ) | ( n24885 & n24886 ) ;
  assign n24894 = ( ~n10380 & n12098 ) | ( ~n10380 & n23444 ) | ( n12098 & n23444 ) ;
  assign n24895 = n24894 ^ n9959 ^ n1777 ;
  assign n24896 = n797 & ~n24895 ;
  assign n24897 = n24896 ^ n9787 ^ 1'b0 ;
  assign n24888 = n3970 ^ n3822 ^ n1379 ;
  assign n24889 = n24888 ^ n22356 ^ n18223 ;
  assign n24890 = n14047 ^ n742 ^ 1'b0 ;
  assign n24891 = n9395 & ~n12592 ;
  assign n24892 = ~n24890 & n24891 ;
  assign n24893 = ( n5784 & n24889 ) | ( n5784 & n24892 ) | ( n24889 & n24892 ) ;
  assign n24898 = n24897 ^ n24893 ^ n24079 ;
  assign n24899 = n14178 & n24685 ;
  assign n24900 = ( ~x3 & n14044 ) | ( ~x3 & n19727 ) | ( n14044 & n19727 ) ;
  assign n24901 = ( n9479 & n15648 ) | ( n9479 & ~n24900 ) | ( n15648 & ~n24900 ) ;
  assign n24902 = ( n10947 & ~n24899 ) | ( n10947 & n24901 ) | ( ~n24899 & n24901 ) ;
  assign n24903 = ( n1278 & n1972 ) | ( n1278 & ~n7305 ) | ( n1972 & ~n7305 ) ;
  assign n24904 = n10829 ^ n1357 ^ 1'b0 ;
  assign n24905 = ( n16332 & n24903 ) | ( n16332 & ~n24904 ) | ( n24903 & ~n24904 ) ;
  assign n24906 = ( ~n7269 & n14337 ) | ( ~n7269 & n14806 ) | ( n14337 & n14806 ) ;
  assign n24908 = n16679 ^ n6411 ^ n5264 ;
  assign n24909 = ~n6500 & n24908 ;
  assign n24907 = n1648 & ~n14746 ;
  assign n24910 = n24909 ^ n24907 ^ 1'b0 ;
  assign n24912 = ( ~n4383 & n7976 ) | ( ~n4383 & n13629 ) | ( n7976 & n13629 ) ;
  assign n24911 = n9312 & n23189 ;
  assign n24913 = n24912 ^ n24911 ^ 1'b0 ;
  assign n24914 = ( ~n9957 & n12366 ) | ( ~n9957 & n18197 ) | ( n12366 & n18197 ) ;
  assign n24915 = n24914 ^ n12885 ^ n1198 ;
  assign n24916 = n24915 ^ n3912 ^ 1'b0 ;
  assign n24917 = n14853 ^ n12553 ^ n5202 ;
  assign n24918 = n24917 ^ n1268 ^ 1'b0 ;
  assign n24919 = n24916 & n24918 ;
  assign n24920 = ( n850 & n10516 ) | ( n850 & ~n12720 ) | ( n10516 & ~n12720 ) ;
  assign n24921 = ( ~n1838 & n13493 ) | ( ~n1838 & n24920 ) | ( n13493 & n24920 ) ;
  assign n24922 = ( n3606 & n7163 ) | ( n3606 & ~n21801 ) | ( n7163 & ~n21801 ) ;
  assign n24923 = n13427 & n24922 ;
  assign n24924 = n14826 ^ n7439 ^ n6180 ;
  assign n24925 = ( ~n3064 & n8888 ) | ( ~n3064 & n24924 ) | ( n8888 & n24924 ) ;
  assign n24926 = ( ~n2552 & n10223 ) | ( ~n2552 & n10322 ) | ( n10223 & n10322 ) ;
  assign n24927 = n24926 ^ n17837 ^ n9865 ;
  assign n24930 = ( ~n3667 & n6785 ) | ( ~n3667 & n14040 ) | ( n6785 & n14040 ) ;
  assign n24931 = ( ~n7781 & n8592 ) | ( ~n7781 & n8797 ) | ( n8592 & n8797 ) ;
  assign n24932 = n304 & ~n24931 ;
  assign n24933 = ~n24930 & n24932 ;
  assign n24929 = n9961 ^ n3919 ^ n3865 ;
  assign n24928 = ( n12782 & ~n14450 ) | ( n12782 & n17230 ) | ( ~n14450 & n17230 ) ;
  assign n24934 = n24933 ^ n24929 ^ n24928 ;
  assign n24935 = ( n24925 & ~n24927 ) | ( n24925 & n24934 ) | ( ~n24927 & n24934 ) ;
  assign n24936 = n19569 & ~n23009 ;
  assign n24937 = ~n9757 & n24936 ;
  assign n24938 = ( x0 & n6299 ) | ( x0 & ~n24937 ) | ( n6299 & ~n24937 ) ;
  assign n24939 = ( n454 & n3215 ) | ( n454 & n19839 ) | ( n3215 & n19839 ) ;
  assign n24940 = ( ~n8072 & n11612 ) | ( ~n8072 & n24939 ) | ( n11612 & n24939 ) ;
  assign n24941 = ( n8178 & ~n24704 ) | ( n8178 & n24940 ) | ( ~n24704 & n24940 ) ;
  assign n24942 = ~n4723 & n6230 ;
  assign n24943 = n14307 ^ n2556 ^ n2079 ;
  assign n24944 = n6219 ^ n4356 ^ n2433 ;
  assign n24945 = ( n8106 & n24943 ) | ( n8106 & ~n24944 ) | ( n24943 & ~n24944 ) ;
  assign n24946 = ( n14978 & n24942 ) | ( n14978 & ~n24945 ) | ( n24942 & ~n24945 ) ;
  assign n24947 = n24946 ^ n15233 ^ n10894 ;
  assign n24948 = ( n3035 & ~n5283 ) | ( n3035 & n6280 ) | ( ~n5283 & n6280 ) ;
  assign n24949 = n18280 ^ n1990 ^ 1'b0 ;
  assign n24950 = n445 & n13404 ;
  assign n24951 = n21595 & n24950 ;
  assign n24952 = ( n5630 & n9225 ) | ( n5630 & ~n15042 ) | ( n9225 & ~n15042 ) ;
  assign n24953 = ( ~n9451 & n23856 ) | ( ~n9451 & n24952 ) | ( n23856 & n24952 ) ;
  assign n24954 = n18979 ^ n4934 ^ n3966 ;
  assign n24955 = ( ~n2427 & n12633 ) | ( ~n2427 & n24954 ) | ( n12633 & n24954 ) ;
  assign n24956 = ( n2513 & n2920 ) | ( n2513 & n11272 ) | ( n2920 & n11272 ) ;
  assign n24957 = n3451 ^ n344 ^ 1'b0 ;
  assign n24958 = n18905 & ~n24957 ;
  assign n24959 = ( n10629 & n24956 ) | ( n10629 & n24958 ) | ( n24956 & n24958 ) ;
  assign n24960 = ( x27 & ~n2472 ) | ( x27 & n6464 ) | ( ~n2472 & n6464 ) ;
  assign n24961 = ( n5392 & ~n12830 ) | ( n5392 & n24960 ) | ( ~n12830 & n24960 ) ;
  assign n24962 = n1821 & n24961 ;
  assign n24963 = n24962 ^ n23628 ^ n1618 ;
  assign n24964 = ~n4361 & n24963 ;
  assign n24965 = ( n7292 & ~n9375 ) | ( n7292 & n18106 ) | ( ~n9375 & n18106 ) ;
  assign n24966 = ( ~n12125 & n12232 ) | ( ~n12125 & n24965 ) | ( n12232 & n24965 ) ;
  assign n24967 = ( n3833 & n17527 ) | ( n3833 & n24966 ) | ( n17527 & n24966 ) ;
  assign n24968 = ( ~n6532 & n24964 ) | ( ~n6532 & n24967 ) | ( n24964 & n24967 ) ;
  assign n24970 = ( n2496 & n12216 ) | ( n2496 & ~n12437 ) | ( n12216 & ~n12437 ) ;
  assign n24969 = ~n2225 & n6238 ;
  assign n24971 = n24970 ^ n24969 ^ 1'b0 ;
  assign n24972 = ( ~n7417 & n14358 ) | ( ~n7417 & n17295 ) | ( n14358 & n17295 ) ;
  assign n24973 = n21940 ^ n14284 ^ 1'b0 ;
  assign n24974 = n15535 ^ n10893 ^ 1'b0 ;
  assign n24975 = ~n18424 & n24974 ;
  assign n24976 = n24975 ^ n636 ^ 1'b0 ;
  assign n24977 = n18348 & ~n24976 ;
  assign n24978 = ( n8060 & ~n18831 ) | ( n8060 & n20648 ) | ( ~n18831 & n20648 ) ;
  assign n24979 = n22845 ^ n22730 ^ n3823 ;
  assign n24980 = ( n6503 & n9814 ) | ( n6503 & ~n24979 ) | ( n9814 & ~n24979 ) ;
  assign n24981 = ~n15041 & n23193 ;
  assign n24982 = n17048 & ~n24981 ;
  assign n24983 = n23831 ^ n9699 ^ 1'b0 ;
  assign n24984 = n4612 & ~n24983 ;
  assign n24985 = n24984 ^ n20764 ^ n14325 ;
  assign n24986 = ~n21368 & n24985 ;
  assign n24987 = ( ~n3346 & n15281 ) | ( ~n3346 & n23273 ) | ( n15281 & n23273 ) ;
  assign n24988 = n24987 ^ n11209 ^ n1602 ;
  assign n24989 = n3191 & ~n7540 ;
  assign n24990 = n24989 ^ n10333 ^ 1'b0 ;
  assign n24991 = n12446 ^ n9771 ^ n8923 ;
  assign n24993 = n4697 ^ n1336 ^ n464 ;
  assign n24992 = n11662 ^ n10216 ^ 1'b0 ;
  assign n24994 = n24993 ^ n24992 ^ n13792 ;
  assign n24995 = n7979 ^ n3751 ^ 1'b0 ;
  assign n24996 = ( ~n1560 & n9828 ) | ( ~n1560 & n15071 ) | ( n9828 & n15071 ) ;
  assign n24998 = n1848 & n12750 ;
  assign n24999 = n24998 ^ n13646 ^ 1'b0 ;
  assign n24997 = n5956 | n10930 ;
  assign n25000 = n24999 ^ n24997 ^ 1'b0 ;
  assign n25001 = ( n12866 & n23812 ) | ( n12866 & ~n25000 ) | ( n23812 & ~n25000 ) ;
  assign n25002 = n11005 ^ n7226 ^ n5052 ;
  assign n25003 = n2268 | n6177 ;
  assign n25004 = ( n14652 & ~n21626 ) | ( n14652 & n25003 ) | ( ~n21626 & n25003 ) ;
  assign n25005 = n11971 ^ n228 ^ 1'b0 ;
  assign n25006 = n20858 & n25005 ;
  assign n25007 = n8053 & ~n17883 ;
  assign n25008 = n372 & n25007 ;
  assign n25009 = n19624 ^ n7078 ^ n3478 ;
  assign n25010 = n362 | n11137 ;
  assign n25011 = n25010 ^ n8057 ^ n1127 ;
  assign n25012 = ( n20322 & ~n22460 ) | ( n20322 & n25011 ) | ( ~n22460 & n25011 ) ;
  assign n25013 = n25012 ^ n16953 ^ n12453 ;
  assign n25014 = n5925 ^ n4311 ^ 1'b0 ;
  assign n25015 = n14630 | n25014 ;
  assign n25016 = n20325 & ~n25015 ;
  assign n25020 = ( ~n2389 & n5593 ) | ( ~n2389 & n10347 ) | ( n5593 & n10347 ) ;
  assign n25021 = n25020 ^ n16492 ^ n10000 ;
  assign n25017 = n16620 | n22228 ;
  assign n25018 = n25017 ^ n6940 ^ 1'b0 ;
  assign n25019 = n25018 ^ n11968 ^ n9534 ;
  assign n25022 = n25021 ^ n25019 ^ n6418 ;
  assign n25023 = ( n13650 & ~n19721 ) | ( n13650 & n25022 ) | ( ~n19721 & n25022 ) ;
  assign n25024 = ( n1565 & n3712 ) | ( n1565 & ~n21224 ) | ( n3712 & ~n21224 ) ;
  assign n25027 = n20163 ^ n15878 ^ n10466 ;
  assign n25025 = n1940 & n8069 ;
  assign n25026 = ( n2717 & n4513 ) | ( n2717 & n25025 ) | ( n4513 & n25025 ) ;
  assign n25028 = n25027 ^ n25026 ^ n5370 ;
  assign n25029 = n14002 ^ n9935 ^ n7272 ;
  assign n25030 = ~n21572 & n25029 ;
  assign n25032 = ( n1343 & n3009 ) | ( n1343 & ~n17305 ) | ( n3009 & ~n17305 ) ;
  assign n25033 = n2852 & n25032 ;
  assign n25034 = ~n9235 & n25033 ;
  assign n25031 = ~n8213 & n14964 ;
  assign n25035 = n25034 ^ n25031 ^ n7827 ;
  assign n25036 = n2182 & ~n9290 ;
  assign n25037 = ~n3713 & n21179 ;
  assign n25038 = ~n20385 & n25037 ;
  assign n25039 = n1798 | n10534 ;
  assign n25040 = ( n11181 & n14923 ) | ( n11181 & n25039 ) | ( n14923 & n25039 ) ;
  assign n25041 = n23953 ^ n15985 ^ n1570 ;
  assign n25042 = n25041 ^ n24156 ^ n16116 ;
  assign n25043 = n751 | n1478 ;
  assign n25044 = ( n3262 & ~n5753 ) | ( n3262 & n9707 ) | ( ~n5753 & n9707 ) ;
  assign n25045 = n5193 ^ n4323 ^ 1'b0 ;
  assign n25046 = n25045 ^ n10071 ^ n9116 ;
  assign n25047 = ( n10551 & n25044 ) | ( n10551 & n25046 ) | ( n25044 & n25046 ) ;
  assign n25048 = ( n18249 & ~n25043 ) | ( n18249 & n25047 ) | ( ~n25043 & n25047 ) ;
  assign n25052 = n9806 ^ n9646 ^ n1059 ;
  assign n25050 = n5993 ^ n4780 ^ x69 ;
  assign n25051 = n25050 ^ n8338 ^ n477 ;
  assign n25049 = n9228 ^ n1713 ^ n631 ;
  assign n25053 = n25052 ^ n25051 ^ n25049 ;
  assign n25054 = n1840 | n8988 ;
  assign n25055 = n25054 ^ n1632 ^ 1'b0 ;
  assign n25056 = n25055 ^ n16603 ^ n8311 ;
  assign n25057 = n25056 ^ n19526 ^ n14957 ;
  assign n25058 = n19266 & ~n25057 ;
  assign n25059 = n17865 ^ n13795 ^ n13787 ;
  assign n25060 = n25059 ^ n11984 ^ n11064 ;
  assign n25061 = n17504 ^ n15531 ^ n12609 ;
  assign n25062 = n25061 ^ n5122 ^ 1'b0 ;
  assign n25063 = n1822 & ~n25062 ;
  assign n25064 = ( n4799 & ~n11470 ) | ( n4799 & n18676 ) | ( ~n11470 & n18676 ) ;
  assign n25065 = n18698 ^ n12275 ^ 1'b0 ;
  assign n25066 = n7963 & ~n25065 ;
  assign n25067 = ( ~x98 & n25064 ) | ( ~x98 & n25066 ) | ( n25064 & n25066 ) ;
  assign n25068 = ( n6493 & n7673 ) | ( n6493 & ~n7807 ) | ( n7673 & ~n7807 ) ;
  assign n25069 = n25068 ^ n12120 ^ 1'b0 ;
  assign n25070 = n25067 | n25069 ;
  assign n25071 = n14152 ^ n9155 ^ n3406 ;
  assign n25072 = n11411 ^ n4780 ^ x88 ;
  assign n25073 = n18786 ^ n18103 ^ n2265 ;
  assign n25074 = ( n3683 & n14504 ) | ( n3683 & ~n15214 ) | ( n14504 & ~n15214 ) ;
  assign n25075 = n25074 ^ n15668 ^ n1232 ;
  assign n25076 = ( n9351 & n25073 ) | ( n9351 & ~n25075 ) | ( n25073 & ~n25075 ) ;
  assign n25077 = n21619 ^ n16270 ^ n7302 ;
  assign n25078 = n7960 ^ n4948 ^ 1'b0 ;
  assign n25079 = ( n5650 & n10315 ) | ( n5650 & ~n24410 ) | ( n10315 & ~n24410 ) ;
  assign n25080 = ( ~n25077 & n25078 ) | ( ~n25077 & n25079 ) | ( n25078 & n25079 ) ;
  assign n25081 = n25080 ^ n19587 ^ n8027 ;
  assign n25082 = n23530 ^ n21563 ^ 1'b0 ;
  assign n25083 = ( n3485 & ~n13680 ) | ( n3485 & n16944 ) | ( ~n13680 & n16944 ) ;
  assign n25084 = n25083 ^ n10940 ^ 1'b0 ;
  assign n25085 = n25082 | n25084 ;
  assign n25086 = n10541 ^ n9675 ^ 1'b0 ;
  assign n25087 = n5584 ^ n4817 ^ n816 ;
  assign n25088 = n25087 ^ n23219 ^ n11811 ;
  assign n25089 = ( ~x100 & n12957 ) | ( ~x100 & n24374 ) | ( n12957 & n24374 ) ;
  assign n25090 = ( n159 & ~n1780 ) | ( n159 & n11742 ) | ( ~n1780 & n11742 ) ;
  assign n25091 = n25090 ^ n17742 ^ n10839 ;
  assign n25092 = n25091 ^ n22610 ^ n12744 ;
  assign n25097 = n12260 ^ n3447 ^ 1'b0 ;
  assign n25098 = n7040 & ~n25097 ;
  assign n25093 = n19531 ^ n12333 ^ n1119 ;
  assign n25094 = n1059 | n9560 ;
  assign n25095 = n3365 | n25094 ;
  assign n25096 = ( n11444 & n25093 ) | ( n11444 & n25095 ) | ( n25093 & n25095 ) ;
  assign n25099 = n25098 ^ n25096 ^ n13097 ;
  assign n25100 = n14864 ^ n7608 ^ n5531 ;
  assign n25101 = n25100 ^ n11515 ^ n8111 ;
  assign n25102 = n16035 ^ n6717 ^ 1'b0 ;
  assign n25103 = n16840 ^ n16747 ^ n1145 ;
  assign n25104 = n5340 ^ n5019 ^ 1'b0 ;
  assign n25105 = n14638 ^ n1645 ^ n859 ;
  assign n25106 = ( n596 & n25104 ) | ( n596 & n25105 ) | ( n25104 & n25105 ) ;
  assign n25107 = ( n7529 & n17631 ) | ( n7529 & n22901 ) | ( n17631 & n22901 ) ;
  assign n25108 = ( n11732 & n25106 ) | ( n11732 & n25107 ) | ( n25106 & n25107 ) ;
  assign n25109 = ( n6092 & n15695 ) | ( n6092 & ~n19312 ) | ( n15695 & ~n19312 ) ;
  assign n25110 = n25109 ^ n7389 ^ n7278 ;
  assign n25112 = n18348 ^ n11707 ^ n2374 ;
  assign n25111 = ( n3276 & ~n12850 ) | ( n3276 & n17452 ) | ( ~n12850 & n17452 ) ;
  assign n25113 = n25112 ^ n25111 ^ n17372 ;
  assign n25116 = ( n1829 & n8627 ) | ( n1829 & ~n22411 ) | ( n8627 & ~n22411 ) ;
  assign n25114 = n3540 & n16644 ;
  assign n25115 = n4696 & n25114 ;
  assign n25117 = n25116 ^ n25115 ^ n9579 ;
  assign n25118 = n25117 ^ n16559 ^ n1081 ;
  assign n25119 = ~n355 & n22238 ;
  assign n25120 = n25119 ^ n15907 ^ 1'b0 ;
  assign n25124 = ( ~n2182 & n5704 ) | ( ~n2182 & n6649 ) | ( n5704 & n6649 ) ;
  assign n25123 = n1036 | n1862 ;
  assign n25125 = n25124 ^ n25123 ^ 1'b0 ;
  assign n25126 = n6901 | n25125 ;
  assign n25127 = n1258 | n25126 ;
  assign n25121 = n4558 & ~n10925 ;
  assign n25122 = ~n18387 & n25121 ;
  assign n25128 = n25127 ^ n25122 ^ n19465 ;
  assign n25129 = ( n2902 & n18741 ) | ( n2902 & n19226 ) | ( n18741 & n19226 ) ;
  assign n25130 = ( n3929 & n13256 ) | ( n3929 & ~n25129 ) | ( n13256 & ~n25129 ) ;
  assign n25131 = ( n154 & n4560 ) | ( n154 & ~n13783 ) | ( n4560 & ~n13783 ) ;
  assign n25132 = n2457 & ~n2906 ;
  assign n25133 = n25132 ^ n16688 ^ n12936 ;
  assign n25134 = n25133 ^ n15348 ^ n12354 ;
  assign n25135 = n19749 ^ n14445 ^ n342 ;
  assign n25136 = n25135 ^ n20859 ^ n14808 ;
  assign n25137 = n18443 ^ n6514 ^ n3787 ;
  assign n25138 = ( ~n5192 & n8330 ) | ( ~n5192 & n25137 ) | ( n8330 & n25137 ) ;
  assign n25139 = n24732 ^ n19749 ^ n6696 ;
  assign n25140 = n13216 ^ n3263 ^ 1'b0 ;
  assign n25141 = ( ~n25138 & n25139 ) | ( ~n25138 & n25140 ) | ( n25139 & n25140 ) ;
  assign n25142 = n18782 ^ n11745 ^ n8129 ;
  assign n25143 = n8283 & ~n15572 ;
  assign n25144 = ~n5733 & n25143 ;
  assign n25145 = n1296 | n6356 ;
  assign n25146 = n6809 ^ n887 ^ 1'b0 ;
  assign n25147 = ~n14009 & n25146 ;
  assign n25148 = ( n13329 & n19997 ) | ( n13329 & n25147 ) | ( n19997 & n25147 ) ;
  assign n25149 = ( n404 & ~n9400 ) | ( n404 & n17955 ) | ( ~n9400 & n17955 ) ;
  assign n25150 = ( n8484 & ~n11440 ) | ( n8484 & n25149 ) | ( ~n11440 & n25149 ) ;
  assign n25151 = ( n14639 & n24409 ) | ( n14639 & n25150 ) | ( n24409 & n25150 ) ;
  assign n25152 = n19225 ^ n8843 ^ 1'b0 ;
  assign n25153 = ( n4053 & n9167 ) | ( n4053 & n13761 ) | ( n9167 & n13761 ) ;
  assign n25154 = n11656 & n25153 ;
  assign n25155 = n17333 ^ n6953 ^ n6231 ;
  assign n25156 = n20016 ^ n12232 ^ 1'b0 ;
  assign n25157 = n18360 ^ x58 ^ 1'b0 ;
  assign n25158 = ~n9938 & n20726 ;
  assign n25159 = ( n689 & n15167 ) | ( n689 & n16620 ) | ( n15167 & n16620 ) ;
  assign n25160 = n19154 ^ n6865 ^ n3387 ;
  assign n25161 = ( n11152 & n11707 ) | ( n11152 & ~n25160 ) | ( n11707 & ~n25160 ) ;
  assign n25162 = n25161 ^ n5081 ^ 1'b0 ;
  assign n25163 = n7198 & n25162 ;
  assign n25164 = ~n6275 & n25163 ;
  assign n25165 = ( n1865 & n15265 ) | ( n1865 & ~n25059 ) | ( n15265 & ~n25059 ) ;
  assign n25166 = n24480 ^ n12551 ^ 1'b0 ;
  assign n25167 = n423 & n23523 ;
  assign n25168 = n25167 ^ n16961 ^ 1'b0 ;
  assign n25169 = n25168 ^ n14445 ^ n559 ;
  assign n25170 = n7840 & ~n12541 ;
  assign n25171 = ( ~n842 & n5281 ) | ( ~n842 & n10126 ) | ( n5281 & n10126 ) ;
  assign n25172 = n10103 | n12816 ;
  assign n25173 = n25171 & ~n25172 ;
  assign n25174 = n25173 ^ n7940 ^ n2719 ;
  assign n25175 = ( ~n3688 & n22621 ) | ( ~n3688 & n25174 ) | ( n22621 & n25174 ) ;
  assign n25176 = n7266 & n19774 ;
  assign n25177 = n25176 ^ n18205 ^ n4691 ;
  assign n25178 = ( ~n567 & n4513 ) | ( ~n567 & n9563 ) | ( n4513 & n9563 ) ;
  assign n25179 = n17447 ^ n11956 ^ n7904 ;
  assign n25180 = n25179 ^ n1496 ^ x123 ;
  assign n25181 = ~n11307 & n25180 ;
  assign n25182 = ~n10090 & n25181 ;
  assign n25183 = ( n9840 & n25178 ) | ( n9840 & n25182 ) | ( n25178 & n25182 ) ;
  assign n25186 = n3543 ^ n3191 ^ n523 ;
  assign n25184 = n22826 ^ n12595 ^ n10701 ;
  assign n25185 = ( n5271 & n19453 ) | ( n5271 & ~n25184 ) | ( n19453 & ~n25184 ) ;
  assign n25187 = n25186 ^ n25185 ^ n23881 ;
  assign n25188 = n21077 ^ n11258 ^ 1'b0 ;
  assign n25189 = ( ~n1251 & n6380 ) | ( ~n1251 & n10382 ) | ( n6380 & n10382 ) ;
  assign n25190 = n25189 ^ n20201 ^ n2783 ;
  assign n25191 = n10540 ^ n3628 ^ 1'b0 ;
  assign n25192 = n16863 & n25191 ;
  assign n25193 = n18446 ^ n10299 ^ n3624 ;
  assign n25194 = ( n17781 & n23390 ) | ( n17781 & ~n25193 ) | ( n23390 & ~n25193 ) ;
  assign n25195 = ( n1235 & n12333 ) | ( n1235 & n19073 ) | ( n12333 & n19073 ) ;
  assign n25200 = n199 | n12313 ;
  assign n25201 = n25200 ^ n11113 ^ 1'b0 ;
  assign n25196 = n18633 | n21682 ;
  assign n25197 = ( ~n1100 & n6593 ) | ( ~n1100 & n25196 ) | ( n6593 & n25196 ) ;
  assign n25198 = n25197 ^ n17581 ^ n11466 ;
  assign n25199 = ( ~n1395 & n8461 ) | ( ~n1395 & n25198 ) | ( n8461 & n25198 ) ;
  assign n25202 = n25201 ^ n25199 ^ n14021 ;
  assign n25203 = n13537 ^ n12565 ^ n10058 ;
  assign n25204 = n25203 ^ n18501 ^ n12711 ;
  assign n25205 = n24733 ^ n17766 ^ n5298 ;
  assign n25206 = n7468 & ~n19192 ;
  assign n25207 = ~n16295 & n25206 ;
  assign n25213 = ( n2519 & n13919 ) | ( n2519 & ~n20511 ) | ( n13919 & ~n20511 ) ;
  assign n25209 = ~n1179 & n12594 ;
  assign n25210 = ~n15103 & n25209 ;
  assign n25208 = ~n1670 & n4190 ;
  assign n25211 = n25210 ^ n25208 ^ 1'b0 ;
  assign n25212 = ~n23084 & n25211 ;
  assign n25214 = n25213 ^ n25212 ^ 1'b0 ;
  assign n25215 = ( n2622 & n2766 ) | ( n2622 & ~n11107 ) | ( n2766 & ~n11107 ) ;
  assign n25216 = n13617 ^ n10546 ^ n2776 ;
  assign n25217 = ( n3821 & n25215 ) | ( n3821 & ~n25216 ) | ( n25215 & ~n25216 ) ;
  assign n25218 = n25217 ^ n14642 ^ n9719 ;
  assign n25219 = n3334 ^ n2468 ^ n1971 ;
  assign n25220 = n25219 ^ n24001 ^ n14202 ;
  assign n25221 = n4848 ^ n4006 ^ n2448 ;
  assign n25222 = n25221 ^ n13085 ^ n10784 ;
  assign n25223 = n24399 & n25222 ;
  assign n25224 = ( n14738 & n22860 ) | ( n14738 & n25223 ) | ( n22860 & n25223 ) ;
  assign n25225 = n25224 ^ n21659 ^ n202 ;
  assign n25226 = ( n859 & n1582 ) | ( n859 & n7057 ) | ( n1582 & n7057 ) ;
  assign n25227 = n25226 ^ n21854 ^ n5502 ;
  assign n25228 = n19355 ^ n11490 ^ n305 ;
  assign n25229 = n25228 ^ n24825 ^ n13278 ;
  assign n25230 = n1982 & ~n12059 ;
  assign n25231 = ~n4090 & n25230 ;
  assign n25232 = ( n15022 & n20509 ) | ( n15022 & ~n25231 ) | ( n20509 & ~n25231 ) ;
  assign n25233 = ~n10310 & n12088 ;
  assign n25234 = n18799 ^ n9510 ^ n1406 ;
  assign n25235 = ( n6886 & n12632 ) | ( n6886 & n16405 ) | ( n12632 & n16405 ) ;
  assign n25236 = n25235 ^ n5104 ^ n2034 ;
  assign n25237 = n689 & n17825 ;
  assign n25238 = ( ~n17696 & n22810 ) | ( ~n17696 & n25237 ) | ( n22810 & n25237 ) ;
  assign n25239 = ( n2149 & ~n6200 ) | ( n2149 & n19090 ) | ( ~n6200 & n19090 ) ;
  assign n25240 = n144 & n19562 ;
  assign n25241 = ~n25239 & n25240 ;
  assign n25248 = ( ~x91 & x93 ) | ( ~x91 & n1752 ) | ( x93 & n1752 ) ;
  assign n25244 = ( n1550 & n4169 ) | ( n1550 & n19574 ) | ( n4169 & n19574 ) ;
  assign n25245 = ( ~n391 & n10030 ) | ( ~n391 & n25244 ) | ( n10030 & n25244 ) ;
  assign n25242 = ~n545 & n19818 ;
  assign n25243 = n25242 ^ n12305 ^ 1'b0 ;
  assign n25246 = n25245 ^ n25243 ^ n3080 ;
  assign n25247 = n25246 ^ n14499 ^ n7670 ;
  assign n25249 = n25248 ^ n25247 ^ n1008 ;
  assign n25250 = ( ~n16284 & n25241 ) | ( ~n16284 & n25249 ) | ( n25241 & n25249 ) ;
  assign n25251 = n18934 ^ n4445 ^ n3937 ;
  assign n25252 = ~n17536 & n25251 ;
  assign n25253 = n25252 ^ n21222 ^ 1'b0 ;
  assign n25254 = ( n1435 & n8815 ) | ( n1435 & ~n16888 ) | ( n8815 & ~n16888 ) ;
  assign n25255 = ( n2348 & n11638 ) | ( n2348 & n12557 ) | ( n11638 & n12557 ) ;
  assign n25256 = n25255 ^ n1462 ^ 1'b0 ;
  assign n25257 = n25254 | n25256 ;
  assign n25258 = n22274 ^ n11345 ^ n1755 ;
  assign n25259 = n25258 ^ n23228 ^ n10963 ;
  assign n25260 = ( n11967 & n13098 ) | ( n11967 & n16361 ) | ( n13098 & n16361 ) ;
  assign n25261 = ( n1940 & n16742 ) | ( n1940 & ~n25260 ) | ( n16742 & ~n25260 ) ;
  assign n25262 = n23981 ^ n21778 ^ n15715 ;
  assign n25263 = n7985 ^ n1241 ^ 1'b0 ;
  assign n25264 = n3062 & ~n25263 ;
  assign n25265 = ( n9257 & ~n20018 ) | ( n9257 & n25264 ) | ( ~n20018 & n25264 ) ;
  assign n25266 = n14367 ^ n3920 ^ n3302 ;
  assign n25267 = n25265 & n25266 ;
  assign n25268 = ~n5400 & n23569 ;
  assign n25269 = ( n3392 & n25246 ) | ( n3392 & ~n25268 ) | ( n25246 & ~n25268 ) ;
  assign n25270 = n25269 ^ n18209 ^ n1574 ;
  assign n25271 = ( ~n2142 & n25267 ) | ( ~n2142 & n25270 ) | ( n25267 & n25270 ) ;
  assign n25272 = n19707 ^ n5479 ^ n2549 ;
  assign n25273 = n25272 ^ n14441 ^ n4321 ;
  assign n25274 = ( n1712 & n8569 ) | ( n1712 & n25273 ) | ( n8569 & n25273 ) ;
  assign n25275 = n16415 ^ n7248 ^ n3654 ;
  assign n25276 = ( n5356 & n8287 ) | ( n5356 & ~n25275 ) | ( n8287 & ~n25275 ) ;
  assign n25277 = ( ~n419 & n5019 ) | ( ~n419 & n25276 ) | ( n5019 & n25276 ) ;
  assign n25278 = ~n7350 & n25277 ;
  assign n25279 = ~n8186 & n25278 ;
  assign n25280 = ~n495 & n6800 ;
  assign n25281 = n25280 ^ n19796 ^ 1'b0 ;
  assign n25282 = n17121 & ~n22913 ;
  assign n25283 = n19531 ^ n16209 ^ n2395 ;
  assign n25284 = ( ~n4150 & n6253 ) | ( ~n4150 & n25283 ) | ( n6253 & n25283 ) ;
  assign n25285 = n18680 ^ n7426 ^ n3263 ;
  assign n25286 = ( n10703 & ~n20414 ) | ( n10703 & n25285 ) | ( ~n20414 & n25285 ) ;
  assign n25287 = ( n11597 & n14686 ) | ( n11597 & ~n25286 ) | ( n14686 & ~n25286 ) ;
  assign n25288 = ( n4361 & ~n6635 ) | ( n4361 & n6686 ) | ( ~n6635 & n6686 ) ;
  assign n25289 = n25288 ^ n2493 ^ 1'b0 ;
  assign n25290 = n15316 ^ n13523 ^ n11687 ;
  assign n25291 = ~n6923 & n7870 ;
  assign n25292 = n18117 ^ n16601 ^ n2630 ;
  assign n25293 = ( ~n8428 & n15386 ) | ( ~n8428 & n25292 ) | ( n15386 & n25292 ) ;
  assign n25294 = n23930 & ~n25293 ;
  assign n25295 = n25294 ^ n16386 ^ 1'b0 ;
  assign n25296 = ~n19160 & n20887 ;
  assign n25297 = n19822 ^ n6792 ^ n3224 ;
  assign n25298 = n8307 & n25297 ;
  assign n25299 = ( n10012 & n19258 ) | ( n10012 & ~n25298 ) | ( n19258 & ~n25298 ) ;
  assign n25300 = ( n7323 & ~n18184 ) | ( n7323 & n18293 ) | ( ~n18184 & n18293 ) ;
  assign n25301 = n22965 ^ n19391 ^ n11263 ;
  assign n25302 = ( n1156 & ~n2655 ) | ( n1156 & n22937 ) | ( ~n2655 & n22937 ) ;
  assign n25303 = ~n10889 & n18525 ;
  assign n25304 = ~n25302 & n25303 ;
  assign n25305 = ( n15997 & n17121 ) | ( n15997 & n18075 ) | ( n17121 & n18075 ) ;
  assign n25306 = n8751 ^ x62 ^ 1'b0 ;
  assign n25307 = n11736 | n25306 ;
  assign n25308 = ( n7482 & n25305 ) | ( n7482 & n25307 ) | ( n25305 & n25307 ) ;
  assign n25309 = ( ~n5360 & n15687 ) | ( ~n5360 & n23153 ) | ( n15687 & n23153 ) ;
  assign n25312 = n2987 | n7972 ;
  assign n25313 = n25312 ^ n9674 ^ 1'b0 ;
  assign n25310 = ( ~x74 & n4413 ) | ( ~x74 & n4665 ) | ( n4413 & n4665 ) ;
  assign n25311 = n25310 ^ n14305 ^ n6265 ;
  assign n25314 = n25313 ^ n25311 ^ n9618 ;
  assign n25315 = n13102 ^ n9968 ^ n2985 ;
  assign n25316 = ( n7465 & ~n10089 ) | ( n7465 & n25315 ) | ( ~n10089 & n25315 ) ;
  assign n25317 = n25316 ^ n20605 ^ n4532 ;
  assign n25318 = n9783 ^ n3971 ^ 1'b0 ;
  assign n25319 = n10295 & n25318 ;
  assign n25320 = n17285 ^ n7440 ^ 1'b0 ;
  assign n25321 = n2022 & ~n25320 ;
  assign n25322 = n25321 ^ n17499 ^ n11501 ;
  assign n25323 = ~n2142 & n8244 ;
  assign n25324 = n25323 ^ n4128 ^ 1'b0 ;
  assign n25325 = n12961 ^ n5674 ^ 1'b0 ;
  assign n25326 = n9708 & ~n25325 ;
  assign n25327 = ( n10652 & ~n11155 ) | ( n10652 & n11440 ) | ( ~n11155 & n11440 ) ;
  assign n25328 = n12553 ^ n1731 ^ 1'b0 ;
  assign n25329 = n25328 ^ n10939 ^ n6643 ;
  assign n25330 = n25327 | n25329 ;
  assign n25331 = ( ~n198 & n2769 ) | ( ~n198 & n23771 ) | ( n2769 & n23771 ) ;
  assign n25332 = n2139 ^ n1586 ^ n906 ;
  assign n25333 = ~n1732 & n18800 ;
  assign n25334 = n25333 ^ n593 ^ 1'b0 ;
  assign n25335 = n21410 ^ n14445 ^ n14009 ;
  assign n25336 = n6848 & ~n22634 ;
  assign n25337 = ~n25335 & n25336 ;
  assign n25338 = n9955 & n24826 ;
  assign n25339 = ~n11236 & n25338 ;
  assign n25341 = n2978 & n10579 ;
  assign n25342 = ~n5260 & n25341 ;
  assign n25343 = n14335 ^ n2381 ^ n2015 ;
  assign n25344 = ( ~n1940 & n25342 ) | ( ~n1940 & n25343 ) | ( n25342 & n25343 ) ;
  assign n25340 = ( n669 & n4533 ) | ( n669 & n22022 ) | ( n4533 & n22022 ) ;
  assign n25345 = n25344 ^ n25340 ^ n23655 ;
  assign n25348 = n11002 ^ n9198 ^ n1504 ;
  assign n25346 = n7436 ^ n6650 ^ 1'b0 ;
  assign n25347 = n18680 | n25346 ;
  assign n25349 = n25348 ^ n25347 ^ n25080 ;
  assign n25350 = n11056 & n24052 ;
  assign n25351 = n25350 ^ n12017 ^ n9799 ;
  assign n25352 = n18097 ^ n4969 ^ 1'b0 ;
  assign n25353 = n25352 ^ n23542 ^ n8294 ;
  assign n25354 = n763 & n10130 ;
  assign n25355 = ( n5362 & n10818 ) | ( n5362 & ~n12198 ) | ( n10818 & ~n12198 ) ;
  assign n25356 = n25355 ^ n18405 ^ n5060 ;
  assign n25357 = n25356 ^ n7108 ^ 1'b0 ;
  assign n25358 = n11701 | n25357 ;
  assign n25361 = n5769 & ~n16105 ;
  assign n25362 = n25361 ^ n7928 ^ 1'b0 ;
  assign n25363 = ( n725 & n11641 ) | ( n725 & ~n13067 ) | ( n11641 & ~n13067 ) ;
  assign n25364 = ( n9208 & n25362 ) | ( n9208 & ~n25363 ) | ( n25362 & ~n25363 ) ;
  assign n25359 = ( n7996 & n9783 ) | ( n7996 & n20720 ) | ( n9783 & n20720 ) ;
  assign n25360 = n3919 & ~n25359 ;
  assign n25365 = n25364 ^ n25360 ^ 1'b0 ;
  assign n25366 = n11760 ^ n11246 ^ n4608 ;
  assign n25367 = n24419 ^ n17405 ^ n15978 ;
  assign n25368 = ( ~n7744 & n25366 ) | ( ~n7744 & n25367 ) | ( n25366 & n25367 ) ;
  assign n25369 = n23128 ^ n16384 ^ n12198 ;
  assign n25370 = n13045 ^ n3012 ^ 1'b0 ;
  assign n25371 = ( n392 & n2453 ) | ( n392 & ~n25370 ) | ( n2453 & ~n25370 ) ;
  assign n25372 = n25371 ^ n19937 ^ n19739 ;
  assign n25373 = ~n6560 & n8158 ;
  assign n25374 = ( n4896 & n6310 ) | ( n4896 & ~n25373 ) | ( n6310 & ~n25373 ) ;
  assign n25375 = n25374 ^ n9383 ^ n2703 ;
  assign n25376 = n9987 ^ n8875 ^ 1'b0 ;
  assign n25377 = n5618 & n25376 ;
  assign n25378 = n25377 ^ n4816 ^ 1'b0 ;
  assign n25379 = n7426 & n23159 ;
  assign n25381 = n22930 ^ n1740 ^ n220 ;
  assign n25380 = n1844 & n22742 ;
  assign n25382 = n25381 ^ n25380 ^ 1'b0 ;
  assign n25383 = n18740 ^ n12963 ^ n5804 ;
  assign n25384 = n1708 & n14412 ;
  assign n25385 = n25384 ^ n254 ^ 1'b0 ;
  assign n25386 = n7053 | n20756 ;
  assign n25387 = n13859 & ~n25386 ;
  assign n25388 = ( n4870 & ~n7574 ) | ( n4870 & n9522 ) | ( ~n7574 & n9522 ) ;
  assign n25389 = n10036 ^ n7245 ^ n1581 ;
  assign n25390 = n25389 ^ n22912 ^ n15981 ;
  assign n25391 = n25390 ^ n13019 ^ n12534 ;
  assign n25392 = n7938 & n18413 ;
  assign n25393 = n25392 ^ n11609 ^ 1'b0 ;
  assign n25394 = n4240 ^ n3863 ^ 1'b0 ;
  assign n25395 = ( n3665 & ~n25393 ) | ( n3665 & n25394 ) | ( ~n25393 & n25394 ) ;
  assign n25397 = n8385 ^ n6597 ^ n2427 ;
  assign n25396 = n4663 | n11853 ;
  assign n25398 = n25397 ^ n25396 ^ 1'b0 ;
  assign n25399 = ( n1069 & ~n16168 ) | ( n1069 & n25398 ) | ( ~n16168 & n25398 ) ;
  assign n25400 = n25399 ^ n10008 ^ n6020 ;
  assign n25403 = n6249 ^ n5911 ^ n3236 ;
  assign n25404 = ~n9861 & n25403 ;
  assign n25405 = ( n11852 & ~n16823 ) | ( n11852 & n25404 ) | ( ~n16823 & n25404 ) ;
  assign n25401 = ~n2472 & n24042 ;
  assign n25402 = n25401 ^ n187 ^ 1'b0 ;
  assign n25406 = n25405 ^ n25402 ^ n2070 ;
  assign n25407 = ( x116 & n4627 ) | ( x116 & ~n20918 ) | ( n4627 & ~n20918 ) ;
  assign n25408 = n23128 ^ n14594 ^ 1'b0 ;
  assign n25409 = n2756 | n4629 ;
  assign n25410 = n25409 ^ n8732 ^ 1'b0 ;
  assign n25411 = n25410 ^ n17911 ^ n9186 ;
  assign n25412 = n14300 & n25411 ;
  assign n25413 = ( n10888 & ~n12192 ) | ( n10888 & n25412 ) | ( ~n12192 & n25412 ) ;
  assign n25414 = n6659 ^ n5794 ^ 1'b0 ;
  assign n25415 = n11827 & ~n25414 ;
  assign n25416 = ( n11850 & ~n17364 ) | ( n11850 & n25415 ) | ( ~n17364 & n25415 ) ;
  assign n25417 = ( n7876 & ~n17212 ) | ( n7876 & n18626 ) | ( ~n17212 & n18626 ) ;
  assign n25418 = ( n24491 & n25416 ) | ( n24491 & n25417 ) | ( n25416 & n25417 ) ;
  assign n25419 = n7454 ^ n6150 ^ n4139 ;
  assign n25420 = n25419 ^ n9693 ^ 1'b0 ;
  assign n25421 = ~n13473 & n19249 ;
  assign n25422 = n25421 ^ n23521 ^ 1'b0 ;
  assign n25423 = n13312 ^ n4777 ^ n4362 ;
  assign n25424 = n25423 ^ n20977 ^ n342 ;
  assign n25425 = ( n11699 & n20620 ) | ( n11699 & ~n23835 ) | ( n20620 & ~n23835 ) ;
  assign n25426 = ( ~n340 & n13808 ) | ( ~n340 & n25425 ) | ( n13808 & n25425 ) ;
  assign n25427 = ( n918 & n8194 ) | ( n918 & n14087 ) | ( n8194 & n14087 ) ;
  assign n25428 = n25427 ^ n8283 ^ n1573 ;
  assign n25429 = ( n8474 & n22332 ) | ( n8474 & ~n25428 ) | ( n22332 & ~n25428 ) ;
  assign n25430 = ~n6982 & n7396 ;
  assign n25431 = ~n25429 & n25430 ;
  assign n25432 = n25431 ^ n19733 ^ n14271 ;
  assign n25433 = n20560 ^ n3433 ^ n3045 ;
  assign n25434 = n25433 ^ n5752 ^ n831 ;
  assign n25435 = n1597 | n4013 ;
  assign n25436 = ( n1147 & n14222 ) | ( n1147 & n19857 ) | ( n14222 & n19857 ) ;
  assign n25437 = n25435 | n25436 ;
  assign n25438 = ( n1909 & n3200 ) | ( n1909 & n4309 ) | ( n3200 & n4309 ) ;
  assign n25442 = ~n6019 & n14908 ;
  assign n25443 = n25442 ^ n10708 ^ 1'b0 ;
  assign n25439 = n13015 ^ n11416 ^ n4150 ;
  assign n25440 = n25147 ^ n11290 ^ 1'b0 ;
  assign n25441 = n25439 & ~n25440 ;
  assign n25444 = n25443 ^ n25441 ^ 1'b0 ;
  assign n25445 = n14693 ^ n5583 ^ 1'b0 ;
  assign n25447 = n1876 ^ n620 ^ n562 ;
  assign n25446 = n5826 & ~n23050 ;
  assign n25448 = n25447 ^ n25446 ^ 1'b0 ;
  assign n25449 = n18164 | n18744 ;
  assign n25450 = ( n10496 & n15168 ) | ( n10496 & n18044 ) | ( n15168 & n18044 ) ;
  assign n25451 = ~n5529 & n17821 ;
  assign n25452 = ~n2465 & n25451 ;
  assign n25453 = n25452 ^ n6463 ^ 1'b0 ;
  assign n25454 = n2900 | n3339 ;
  assign n25455 = n25454 ^ n11618 ^ n3046 ;
  assign n25456 = ( n17252 & n19277 ) | ( n17252 & ~n25203 ) | ( n19277 & ~n25203 ) ;
  assign n25457 = n1057 & ~n2639 ;
  assign n25458 = n25457 ^ n3219 ^ 1'b0 ;
  assign n25459 = ~n1564 & n25458 ;
  assign n25460 = n17695 & n25459 ;
  assign n25461 = n6506 & ~n6685 ;
  assign n25462 = n15816 & n25461 ;
  assign n25463 = n10295 ^ n6143 ^ n3899 ;
  assign n25464 = n5948 ^ n5012 ^ 1'b0 ;
  assign n25465 = ( n4139 & n15264 ) | ( n4139 & ~n25464 ) | ( n15264 & ~n25464 ) ;
  assign n25466 = ( n6841 & n6949 ) | ( n6841 & n25465 ) | ( n6949 & n25465 ) ;
  assign n25467 = ( n5816 & n7592 ) | ( n5816 & ~n23060 ) | ( n7592 & ~n23060 ) ;
  assign n25468 = ( n1886 & n3022 ) | ( n1886 & ~n16814 ) | ( n3022 & ~n16814 ) ;
  assign n25469 = ( n19853 & n22347 ) | ( n19853 & n25468 ) | ( n22347 & n25468 ) ;
  assign n25470 = n25469 ^ n22405 ^ n4762 ;
  assign n25471 = ( n2780 & n3851 ) | ( n2780 & ~n5608 ) | ( n3851 & ~n5608 ) ;
  assign n25472 = ( n2927 & n6689 ) | ( n2927 & ~n25471 ) | ( n6689 & ~n25471 ) ;
  assign n25473 = n22472 ^ n9835 ^ n5937 ;
  assign n25474 = ~n396 & n11458 ;
  assign n25475 = ~n2247 & n25474 ;
  assign n25477 = n23756 ^ n15451 ^ n7883 ;
  assign n25476 = n13197 ^ n2064 ^ n513 ;
  assign n25478 = n25477 ^ n25476 ^ n7531 ;
  assign n25479 = ( n2452 & n13074 ) | ( n2452 & ~n20261 ) | ( n13074 & ~n20261 ) ;
  assign n25483 = ( n1444 & n6397 ) | ( n1444 & ~n10305 ) | ( n6397 & ~n10305 ) ;
  assign n25480 = ~n9168 & n15391 ;
  assign n25481 = n25480 ^ n19787 ^ 1'b0 ;
  assign n25482 = ( n12439 & n16026 ) | ( n12439 & n25481 ) | ( n16026 & n25481 ) ;
  assign n25484 = n25483 ^ n25482 ^ n611 ;
  assign n25485 = ( n15365 & n25479 ) | ( n15365 & n25484 ) | ( n25479 & n25484 ) ;
  assign n25486 = n17621 ^ n8533 ^ 1'b0 ;
  assign n25487 = n1170 | n9413 ;
  assign n25488 = ( n5611 & ~n16859 ) | ( n5611 & n25487 ) | ( ~n16859 & n25487 ) ;
  assign n25489 = ~n6303 & n25488 ;
  assign n25490 = ( n12299 & n25486 ) | ( n12299 & ~n25489 ) | ( n25486 & ~n25489 ) ;
  assign n25491 = ( n1456 & n6507 ) | ( n1456 & ~n15180 ) | ( n6507 & ~n15180 ) ;
  assign n25492 = ( ~n7411 & n12152 ) | ( ~n7411 & n21355 ) | ( n12152 & n21355 ) ;
  assign n25493 = ( n826 & n9707 ) | ( n826 & n19757 ) | ( n9707 & n19757 ) ;
  assign n25494 = ( n15450 & n25492 ) | ( n15450 & n25493 ) | ( n25492 & n25493 ) ;
  assign n25495 = n25494 ^ n10328 ^ 1'b0 ;
  assign n25496 = n25495 ^ n16203 ^ n2799 ;
  assign n25497 = n25496 ^ n17391 ^ n12458 ;
  assign n25500 = ( ~n3126 & n16642 ) | ( ~n3126 & n19216 ) | ( n16642 & n19216 ) ;
  assign n25498 = n11476 ^ n3526 ^ 1'b0 ;
  assign n25499 = ~n20726 & n25498 ;
  assign n25501 = n25500 ^ n25499 ^ n18723 ;
  assign n25502 = n24984 ^ n19700 ^ n13007 ;
  assign n25503 = n24530 ^ n6956 ^ 1'b0 ;
  assign n25504 = n18740 & n25503 ;
  assign n25505 = n23069 ^ n7655 ^ n1109 ;
  assign n25506 = ( n299 & n20510 ) | ( n299 & n25505 ) | ( n20510 & n25505 ) ;
  assign n25507 = n25506 ^ n21751 ^ n4660 ;
  assign n25513 = n18212 ^ n14039 ^ n13385 ;
  assign n25514 = ( n495 & n15898 ) | ( n495 & ~n25513 ) | ( n15898 & ~n25513 ) ;
  assign n25508 = ( n15113 & ~n16367 ) | ( n15113 & n16831 ) | ( ~n16367 & n16831 ) ;
  assign n25509 = n25508 ^ n21396 ^ n1738 ;
  assign n25510 = ( n5475 & n9461 ) | ( n5475 & ~n25509 ) | ( n9461 & ~n25509 ) ;
  assign n25511 = ( n9219 & n20776 ) | ( n9219 & ~n25510 ) | ( n20776 & ~n25510 ) ;
  assign n25512 = ( n4281 & ~n14654 ) | ( n4281 & n25511 ) | ( ~n14654 & n25511 ) ;
  assign n25515 = n25514 ^ n25512 ^ n16360 ;
  assign n25516 = n11543 ^ n9771 ^ n896 ;
  assign n25517 = n25516 ^ n9745 ^ n3467 ;
  assign n25518 = ~n9719 & n23310 ;
  assign n25519 = ( n11290 & n12353 ) | ( n11290 & ~n25518 ) | ( n12353 & ~n25518 ) ;
  assign n25520 = n25519 ^ n13374 ^ n2862 ;
  assign n25521 = ( n2473 & n12993 ) | ( n2473 & n22779 ) | ( n12993 & n22779 ) ;
  assign n25522 = n17191 | n24453 ;
  assign n25523 = n25522 ^ n10071 ^ 1'b0 ;
  assign n25524 = ~n4659 & n6964 ;
  assign n25525 = n5818 & n25524 ;
  assign n25526 = ( n20813 & ~n21037 ) | ( n20813 & n25525 ) | ( ~n21037 & n25525 ) ;
  assign n25527 = n12919 ^ n707 ^ 1'b0 ;
  assign n25528 = n25527 ^ n22392 ^ n19276 ;
  assign n25529 = n25528 ^ n12289 ^ n10097 ;
  assign n25530 = ( ~n736 & n6978 ) | ( ~n736 & n11284 ) | ( n6978 & n11284 ) ;
  assign n25531 = ( n4654 & n5697 ) | ( n4654 & ~n17157 ) | ( n5697 & ~n17157 ) ;
  assign n25532 = n25531 ^ n10977 ^ 1'b0 ;
  assign n25533 = n25530 & n25532 ;
  assign n25534 = n25533 ^ n4985 ^ 1'b0 ;
  assign n25535 = ( ~n22126 & n25529 ) | ( ~n22126 & n25534 ) | ( n25529 & n25534 ) ;
  assign n25536 = n6655 & n15832 ;
  assign n25537 = n5268 ^ n4925 ^ 1'b0 ;
  assign n25538 = n5774 | n25537 ;
  assign n25539 = n25538 ^ n20956 ^ n668 ;
  assign n25540 = n11069 ^ n7261 ^ 1'b0 ;
  assign n25541 = n25539 & ~n25540 ;
  assign n25542 = ( ~n14149 & n17742 ) | ( ~n14149 & n25541 ) | ( n17742 & n25541 ) ;
  assign n25546 = n24685 ^ n1653 ^ 1'b0 ;
  assign n25543 = n10646 ^ n10154 ^ n5922 ;
  assign n25544 = ( ~n1912 & n5752 ) | ( ~n1912 & n25543 ) | ( n5752 & n25543 ) ;
  assign n25545 = ( n7124 & n16025 ) | ( n7124 & n25544 ) | ( n16025 & n25544 ) ;
  assign n25547 = n25546 ^ n25545 ^ n11969 ;
  assign n25548 = ( n3430 & n6157 ) | ( n3430 & n16645 ) | ( n6157 & n16645 ) ;
  assign n25549 = n1850 ^ n1653 ^ 1'b0 ;
  assign n25550 = n14539 ^ n12544 ^ n486 ;
  assign n25551 = ( n18358 & ~n25549 ) | ( n18358 & n25550 ) | ( ~n25549 & n25550 ) ;
  assign n25552 = ( ~x2 & n5392 ) | ( ~x2 & n9417 ) | ( n5392 & n9417 ) ;
  assign n25553 = n4281 & n4823 ;
  assign n25554 = n1114 & n25553 ;
  assign n25555 = ( n8969 & n21182 ) | ( n8969 & ~n22705 ) | ( n21182 & ~n22705 ) ;
  assign n25556 = ( ~n7034 & n15750 ) | ( ~n7034 & n25555 ) | ( n15750 & n25555 ) ;
  assign n25557 = ( ~n890 & n10108 ) | ( ~n890 & n25556 ) | ( n10108 & n25556 ) ;
  assign n25558 = n14212 ^ n3852 ^ 1'b0 ;
  assign n25559 = ( n4404 & ~n5210 ) | ( n4404 & n25558 ) | ( ~n5210 & n25558 ) ;
  assign n25560 = ( n451 & ~n1040 ) | ( n451 & n25559 ) | ( ~n1040 & n25559 ) ;
  assign n25561 = n24551 ^ n18633 ^ n16813 ;
  assign n25562 = n13135 & n25189 ;
  assign n25563 = n25562 ^ n16229 ^ 1'b0 ;
  assign n25564 = n13756 & ~n18108 ;
  assign n25565 = n17855 ^ n8513 ^ n1160 ;
  assign n25566 = n21264 ^ n12620 ^ n11098 ;
  assign n25567 = ( n3118 & n19850 ) | ( n3118 & ~n25566 ) | ( n19850 & ~n25566 ) ;
  assign n25568 = ( ~n946 & n1865 ) | ( ~n946 & n21831 ) | ( n1865 & n21831 ) ;
  assign n25569 = n10120 ^ n6827 ^ n4764 ;
  assign n25570 = n25569 ^ n10262 ^ n677 ;
  assign n25571 = n25570 ^ n10720 ^ n7175 ;
  assign n25574 = ( n3423 & n3516 ) | ( n3423 & n15385 ) | ( n3516 & n15385 ) ;
  assign n25572 = n4764 ^ n3135 ^ n215 ;
  assign n25573 = ~n22144 & n25572 ;
  assign n25575 = n25574 ^ n25573 ^ 1'b0 ;
  assign n25576 = n4299 | n25575 ;
  assign n25577 = n4096 & ~n25576 ;
  assign n25578 = ( n4452 & ~n8524 ) | ( n4452 & n18149 ) | ( ~n8524 & n18149 ) ;
  assign n25579 = ( n8741 & ~n17731 ) | ( n8741 & n22264 ) | ( ~n17731 & n22264 ) ;
  assign n25580 = ( n1861 & ~n7229 ) | ( n1861 & n25579 ) | ( ~n7229 & n25579 ) ;
  assign n25581 = n6295 | n25580 ;
  assign n25582 = n25578 | n25581 ;
  assign n25584 = n15358 ^ n12462 ^ n7121 ;
  assign n25583 = ~n337 & n15450 ;
  assign n25585 = n25584 ^ n25583 ^ 1'b0 ;
  assign n25588 = ( n10013 & ~n10312 ) | ( n10013 & n13232 ) | ( ~n10312 & n13232 ) ;
  assign n25586 = ( ~n1325 & n2851 ) | ( ~n1325 & n5399 ) | ( n2851 & n5399 ) ;
  assign n25587 = n25586 ^ n15673 ^ n13275 ;
  assign n25589 = n25588 ^ n25587 ^ 1'b0 ;
  assign n25590 = n17105 ^ n13983 ^ n2012 ;
  assign n25591 = n25590 ^ n5023 ^ 1'b0 ;
  assign n25592 = ( n348 & n2643 ) | ( n348 & n14937 ) | ( n2643 & n14937 ) ;
  assign n25593 = n20605 | n25592 ;
  assign n25594 = n2425 | n25593 ;
  assign n25595 = n12959 ^ n9244 ^ n1481 ;
  assign n25596 = n25595 ^ n20595 ^ n18694 ;
  assign n25597 = n9080 ^ n3931 ^ 1'b0 ;
  assign n25598 = ~n5471 & n25597 ;
  assign n25599 = ( n9167 & n16357 ) | ( n9167 & n25598 ) | ( n16357 & n25598 ) ;
  assign n25600 = n17962 ^ n17834 ^ 1'b0 ;
  assign n25601 = ~n10472 & n16875 ;
  assign n25602 = n6476 & n9974 ;
  assign n25603 = ~n15369 & n25602 ;
  assign n25606 = n20952 ^ n10001 ^ n7191 ;
  assign n25604 = n793 | n14496 ;
  assign n25605 = n1351 & ~n25604 ;
  assign n25607 = n25606 ^ n25605 ^ 1'b0 ;
  assign n25608 = n6371 ^ n4522 ^ 1'b0 ;
  assign n25609 = n4107 & n25608 ;
  assign n25610 = n25609 ^ n8515 ^ n6662 ;
  assign n25611 = n25610 ^ n24415 ^ n2909 ;
  assign n25612 = n25611 ^ n6481 ^ 1'b0 ;
  assign n25613 = ~n15616 & n25612 ;
  assign n25614 = n25613 ^ n10330 ^ n7804 ;
  assign n25615 = ( n7098 & n13407 ) | ( n7098 & ~n21821 ) | ( n13407 & ~n21821 ) ;
  assign n25616 = ( n4865 & n7733 ) | ( n4865 & n25615 ) | ( n7733 & n25615 ) ;
  assign n25617 = ( n10210 & n15128 ) | ( n10210 & ~n15403 ) | ( n15128 & ~n15403 ) ;
  assign n25618 = n19940 ^ n7559 ^ n6527 ;
  assign n25619 = ( ~n24419 & n25617 ) | ( ~n24419 & n25618 ) | ( n25617 & n25618 ) ;
  assign n25620 = ( ~n3973 & n24168 ) | ( ~n3973 & n25619 ) | ( n24168 & n25619 ) ;
  assign n25621 = n17681 ^ n17361 ^ n5003 ;
  assign n25622 = ~n20882 & n25621 ;
  assign n25623 = n2823 | n9360 ;
  assign n25624 = n25623 ^ n13556 ^ n13383 ;
  assign n25625 = ~n19408 & n19547 ;
  assign n25626 = n15016 & n25625 ;
  assign n25627 = n9826 ^ n1960 ^ 1'b0 ;
  assign n25628 = n16271 & ~n25627 ;
  assign n25630 = n12502 ^ n2027 ^ n1749 ;
  assign n25629 = n9611 ^ n2712 ^ n1158 ;
  assign n25631 = n25630 ^ n25629 ^ n1928 ;
  assign n25632 = n10464 ^ n10065 ^ 1'b0 ;
  assign n25633 = x76 & ~n7313 ;
  assign n25634 = n25633 ^ n13074 ^ 1'b0 ;
  assign n25635 = ( ~n7948 & n9912 ) | ( ~n7948 & n15770 ) | ( n9912 & n15770 ) ;
  assign n25636 = ( ~n4097 & n25634 ) | ( ~n4097 & n25635 ) | ( n25634 & n25635 ) ;
  assign n25637 = n3217 ^ n736 ^ n731 ;
  assign n25638 = ( n17802 & n19241 ) | ( n17802 & ~n25637 ) | ( n19241 & ~n25637 ) ;
  assign n25639 = n22673 ^ n15431 ^ 1'b0 ;
  assign n25640 = n25538 ^ n20964 ^ n2776 ;
  assign n25641 = n25640 ^ n22557 ^ n4791 ;
  assign n25642 = n25641 ^ n24072 ^ n7689 ;
  assign n25643 = n25315 ^ n11858 ^ 1'b0 ;
  assign n25644 = n7405 ^ n6244 ^ n3319 ;
  assign n25645 = n25644 ^ n6812 ^ n945 ;
  assign n25646 = n13147 & ~n25645 ;
  assign n25647 = n2678 & ~n25646 ;
  assign n25648 = n25647 ^ n14759 ^ 1'b0 ;
  assign n25649 = n144 & n4104 ;
  assign n25650 = n25649 ^ n13499 ^ 1'b0 ;
  assign n25651 = n21421 ^ n13307 ^ n3034 ;
  assign n25652 = ( ~n5803 & n25650 ) | ( ~n5803 & n25651 ) | ( n25650 & n25651 ) ;
  assign n25653 = n15419 & n25652 ;
  assign n25654 = n25653 ^ n12483 ^ 1'b0 ;
  assign n25655 = n25654 ^ n17848 ^ n15063 ;
  assign n25656 = n24456 ^ n20265 ^ n9546 ;
  assign n25657 = ( n5548 & n6442 ) | ( n5548 & n21083 ) | ( n6442 & n21083 ) ;
  assign n25658 = ~n21072 & n25657 ;
  assign n25659 = ( ~n2565 & n11361 ) | ( ~n2565 & n13275 ) | ( n11361 & n13275 ) ;
  assign n25660 = ( ~n6098 & n14161 ) | ( ~n6098 & n25659 ) | ( n14161 & n25659 ) ;
  assign n25661 = n9237 ^ n8004 ^ 1'b0 ;
  assign n25662 = n14481 | n25661 ;
  assign n25663 = n6423 & ~n25662 ;
  assign n25664 = n16927 | n25663 ;
  assign n25666 = n1420 & n1751 ;
  assign n25667 = ~n16565 & n25666 ;
  assign n25665 = ~n7309 & n10112 ;
  assign n25668 = n25667 ^ n25665 ^ n15045 ;
  assign n25669 = n12754 ^ n9652 ^ n8832 ;
  assign n25670 = n12221 ^ n9897 ^ n9743 ;
  assign n25671 = n25670 ^ n11327 ^ n10623 ;
  assign n25672 = ( ~n11813 & n17862 ) | ( ~n11813 & n20534 ) | ( n17862 & n20534 ) ;
  assign n25673 = n25672 ^ n16340 ^ n5619 ;
  assign n25679 = ( n12094 & n12295 ) | ( n12094 & ~n13945 ) | ( n12295 & ~n13945 ) ;
  assign n25675 = n16435 ^ n5882 ^ n653 ;
  assign n25676 = ( n9469 & n10181 ) | ( n9469 & ~n25675 ) | ( n10181 & ~n25675 ) ;
  assign n25674 = n2396 | n10847 ;
  assign n25677 = n25676 ^ n25674 ^ n20744 ;
  assign n25678 = ( n3106 & ~n7129 ) | ( n3106 & n25677 ) | ( ~n7129 & n25677 ) ;
  assign n25680 = n25679 ^ n25678 ^ 1'b0 ;
  assign n25683 = n20368 ^ n8050 ^ n1942 ;
  assign n25684 = n25683 ^ n14656 ^ n12748 ;
  assign n25685 = ( n5408 & ~n11830 ) | ( n5408 & n25684 ) | ( ~n11830 & n25684 ) ;
  assign n25681 = n1209 & n3745 ;
  assign n25682 = n2776 & ~n25681 ;
  assign n25686 = n25685 ^ n25682 ^ 1'b0 ;
  assign n25688 = n10957 ^ n7590 ^ n337 ;
  assign n25687 = n8601 | n21132 ;
  assign n25689 = n25688 ^ n25687 ^ 1'b0 ;
  assign n25690 = n25689 ^ n4315 ^ 1'b0 ;
  assign n25691 = n16636 & n25690 ;
  assign n25696 = ( n153 & n21142 ) | ( n153 & ~n21787 ) | ( n21142 & ~n21787 ) ;
  assign n25692 = n23367 ^ n7840 ^ n2045 ;
  assign n25693 = ( n10699 & ~n12953 ) | ( n10699 & n25692 ) | ( ~n12953 & n25692 ) ;
  assign n25694 = n25693 ^ n13897 ^ n10207 ;
  assign n25695 = n2873 & ~n25694 ;
  assign n25697 = n25696 ^ n25695 ^ 1'b0 ;
  assign n25698 = n8172 & n25697 ;
  assign n25699 = ( n6378 & n6792 ) | ( n6378 & n9940 ) | ( n6792 & n9940 ) ;
  assign n25700 = n25699 ^ n20818 ^ n13976 ;
  assign n25701 = ( n5410 & ~n11761 ) | ( n5410 & n12949 ) | ( ~n11761 & n12949 ) ;
  assign n25702 = n20419 ^ n6743 ^ n4445 ;
  assign n25703 = n17242 ^ n9459 ^ 1'b0 ;
  assign n25704 = n4508 & n25703 ;
  assign n25705 = ( n14250 & n20864 ) | ( n14250 & ~n25704 ) | ( n20864 & ~n25704 ) ;
  assign n25706 = n19307 ^ n9434 ^ 1'b0 ;
  assign n25707 = n15128 & n25706 ;
  assign n25708 = n3165 & n18175 ;
  assign n25709 = ~n25707 & n25708 ;
  assign n25710 = ( ~n7726 & n10657 ) | ( ~n7726 & n19636 ) | ( n10657 & n19636 ) ;
  assign n25711 = n2546 & n2608 ;
  assign n25712 = ~n25710 & n25711 ;
  assign n25713 = ( ~n18388 & n18595 ) | ( ~n18388 & n25712 ) | ( n18595 & n25712 ) ;
  assign n25714 = ( ~n766 & n8249 ) | ( ~n766 & n11663 ) | ( n8249 & n11663 ) ;
  assign n25715 = ( n8144 & n25713 ) | ( n8144 & ~n25714 ) | ( n25713 & ~n25714 ) ;
  assign n25716 = ( n213 & n4629 ) | ( n213 & n14105 ) | ( n4629 & n14105 ) ;
  assign n25717 = n24730 ^ n3590 ^ 1'b0 ;
  assign n25718 = ~n8721 & n25717 ;
  assign n25719 = ( ~n832 & n21901 ) | ( ~n832 & n25718 ) | ( n21901 & n25718 ) ;
  assign n25720 = n15281 ^ n8665 ^ n7935 ;
  assign n25721 = n18483 ^ n10704 ^ 1'b0 ;
  assign n25722 = n3058 | n5951 ;
  assign n25723 = n25722 ^ n17862 ^ n1661 ;
  assign n25724 = ( n25720 & ~n25721 ) | ( n25720 & n25723 ) | ( ~n25721 & n25723 ) ;
  assign n25725 = n6844 & ~n6984 ;
  assign n25726 = n25725 ^ n21307 ^ 1'b0 ;
  assign n25727 = ( n4788 & n5193 ) | ( n4788 & ~n6357 ) | ( n5193 & ~n6357 ) ;
  assign n25728 = n1167 & n25727 ;
  assign n25729 = n25728 ^ n15559 ^ 1'b0 ;
  assign n25730 = n8212 ^ n6022 ^ 1'b0 ;
  assign n25731 = ( n2242 & n6945 ) | ( n2242 & ~n17961 ) | ( n6945 & ~n17961 ) ;
  assign n25732 = n25435 ^ n15197 ^ n7795 ;
  assign n25733 = n25732 ^ n24536 ^ n3309 ;
  assign n25734 = ( n13307 & n23575 ) | ( n13307 & n25733 ) | ( n23575 & n25733 ) ;
  assign n25735 = n10646 ^ n8092 ^ n7427 ;
  assign n25736 = ( n1483 & n1545 ) | ( n1483 & n25735 ) | ( n1545 & n25735 ) ;
  assign n25737 = n25736 ^ n22554 ^ n4321 ;
  assign n25738 = n14833 ^ n5636 ^ 1'b0 ;
  assign n25739 = ~n4143 & n16754 ;
  assign n25740 = n4834 | n24766 ;
  assign n25741 = n25739 & ~n25740 ;
  assign n25742 = n15817 ^ n1479 ^ 1'b0 ;
  assign n25743 = n20264 & ~n25742 ;
  assign n25744 = n948 | n19152 ;
  assign n25745 = n25744 ^ n8350 ^ 1'b0 ;
  assign n25746 = n14595 ^ n9611 ^ n3616 ;
  assign n25747 = n16814 ^ n10735 ^ n3004 ;
  assign n25748 = ( ~n6323 & n12055 ) | ( ~n6323 & n25747 ) | ( n12055 & n25747 ) ;
  assign n25749 = n25748 ^ n20258 ^ n11606 ;
  assign n25750 = n25749 ^ n473 ^ n442 ;
  assign n25751 = n12121 ^ n8230 ^ 1'b0 ;
  assign n25752 = ( n12734 & n23756 ) | ( n12734 & n25751 ) | ( n23756 & n25751 ) ;
  assign n25753 = ( n2493 & ~n18805 ) | ( n2493 & n25707 ) | ( ~n18805 & n25707 ) ;
  assign n25754 = n16436 ^ n15115 ^ n10310 ;
  assign n25755 = n7380 ^ n603 ^ 1'b0 ;
  assign n25756 = n13326 & n25755 ;
  assign n25757 = n25756 ^ n19008 ^ n9097 ;
  assign n25758 = ( n18314 & n25754 ) | ( n18314 & ~n25757 ) | ( n25754 & ~n25757 ) ;
  assign n25759 = n5379 & ~n9011 ;
  assign n25760 = n9011 & n25759 ;
  assign n25761 = n25760 ^ n19323 ^ n2247 ;
  assign n25762 = n25761 ^ n1152 ^ n362 ;
  assign n25763 = n9036 ^ n5774 ^ n3882 ;
  assign n25764 = n6984 | n25056 ;
  assign n25765 = n25763 | n25764 ;
  assign n25766 = ( n3896 & ~n4246 ) | ( n3896 & n21751 ) | ( ~n4246 & n21751 ) ;
  assign n25767 = n25766 ^ n3814 ^ 1'b0 ;
  assign n25768 = ~n18297 & n25767 ;
  assign n25769 = ( ~n5571 & n7149 ) | ( ~n5571 & n12697 ) | ( n7149 & n12697 ) ;
  assign n25770 = ( ~n4088 & n5958 ) | ( ~n4088 & n22554 ) | ( n5958 & n22554 ) ;
  assign n25771 = ( ~n9482 & n12666 ) | ( ~n9482 & n13709 ) | ( n12666 & n13709 ) ;
  assign n25772 = n22489 ^ n5990 ^ 1'b0 ;
  assign n25773 = ~n19901 & n25772 ;
  assign n25774 = ( ~n3460 & n3854 ) | ( ~n3460 & n11764 ) | ( n3854 & n11764 ) ;
  assign n25775 = ( n5753 & n25773 ) | ( n5753 & n25774 ) | ( n25773 & n25774 ) ;
  assign n25776 = n23524 ^ n21924 ^ 1'b0 ;
  assign n25777 = n2967 & ~n4080 ;
  assign n25778 = n25777 ^ n21139 ^ n21079 ;
  assign n25779 = n21669 ^ n15852 ^ 1'b0 ;
  assign n25780 = ~n18600 & n25779 ;
  assign n25781 = n25780 ^ n21579 ^ n9056 ;
  assign n25782 = ( ~n18128 & n21059 ) | ( ~n18128 & n25781 ) | ( n21059 & n25781 ) ;
  assign n25783 = n2688 ^ n1784 ^ n784 ;
  assign n25784 = ( ~n9075 & n19382 ) | ( ~n9075 & n25783 ) | ( n19382 & n25783 ) ;
  assign n25785 = n18495 ^ n2154 ^ 1'b0 ;
  assign n25786 = n25784 & n25785 ;
  assign n25787 = n7292 ^ n6082 ^ 1'b0 ;
  assign n25788 = n25786 & n25787 ;
  assign n25789 = n11439 | n13606 ;
  assign n25790 = ( n1441 & ~n7633 ) | ( n1441 & n9686 ) | ( ~n7633 & n9686 ) ;
  assign n25791 = n25789 & ~n25790 ;
  assign n25792 = n4810 & n5036 ;
  assign n25793 = n25792 ^ n5063 ^ 1'b0 ;
  assign n25794 = n25793 ^ n5058 ^ 1'b0 ;
  assign n25795 = ( n19449 & ~n19869 ) | ( n19449 & n25794 ) | ( ~n19869 & n25794 ) ;
  assign n25796 = n25795 ^ n3441 ^ n3087 ;
  assign n25797 = ~n7818 & n15759 ;
  assign n25798 = ~n21462 & n25797 ;
  assign n25799 = n25798 ^ n12149 ^ n173 ;
  assign n25800 = n23821 ^ n5519 ^ 1'b0 ;
  assign n25801 = n17170 ^ n7212 ^ n7006 ;
  assign n25802 = ( ~n10768 & n18928 ) | ( ~n10768 & n19556 ) | ( n18928 & n19556 ) ;
  assign n25803 = n5459 | n25802 ;
  assign n25804 = n25803 ^ n22723 ^ 1'b0 ;
  assign n25805 = n16436 ^ n16327 ^ n7465 ;
  assign n25806 = ( ~n1573 & n11951 ) | ( ~n1573 & n25423 ) | ( n11951 & n25423 ) ;
  assign n25807 = n12621 & ~n25806 ;
  assign n25808 = ~n5308 & n7152 ;
  assign n25809 = n11236 ^ n865 ^ 1'b0 ;
  assign n25810 = ~n22002 & n25809 ;
  assign n25811 = n25810 ^ n12808 ^ n4846 ;
  assign n25812 = ( ~n5836 & n25808 ) | ( ~n5836 & n25811 ) | ( n25808 & n25811 ) ;
  assign n25813 = n16163 ^ n14896 ^ n11508 ;
  assign n25814 = ( ~n939 & n24314 ) | ( ~n939 & n25813 ) | ( n24314 & n25813 ) ;
  assign n25815 = n25814 ^ n23979 ^ n8932 ;
  assign n25816 = n7016 ^ n4271 ^ n3328 ;
  assign n25817 = ( x97 & ~n3195 ) | ( x97 & n8044 ) | ( ~n3195 & n8044 ) ;
  assign n25818 = ( n7198 & n12856 ) | ( n7198 & ~n25817 ) | ( n12856 & ~n25817 ) ;
  assign n25819 = ( n7798 & n18506 ) | ( n7798 & ~n25818 ) | ( n18506 & ~n25818 ) ;
  assign n25820 = n25819 ^ n23262 ^ n11628 ;
  assign n25821 = ( n6465 & n17524 ) | ( n6465 & ~n25820 ) | ( n17524 & ~n25820 ) ;
  assign n25822 = n25410 ^ n5410 ^ n2998 ;
  assign n25823 = n25822 ^ n19129 ^ 1'b0 ;
  assign n25824 = n3004 & ~n25823 ;
  assign n25825 = ( n1108 & n5881 ) | ( n1108 & ~n22519 ) | ( n5881 & ~n22519 ) ;
  assign n25826 = n3054 & ~n25825 ;
  assign n25827 = n2695 & n25826 ;
  assign n25828 = ~n2316 & n6668 ;
  assign n25829 = n3968 & n25828 ;
  assign n25830 = n25829 ^ n2062 ^ n1731 ;
  assign n25831 = n3585 ^ n2965 ^ n2270 ;
  assign n25832 = ( n14284 & n15182 ) | ( n14284 & n25831 ) | ( n15182 & n25831 ) ;
  assign n25833 = n3228 & ~n7366 ;
  assign n25834 = n6668 ^ n6608 ^ n3928 ;
  assign n25838 = n7345 ^ n6977 ^ n2323 ;
  assign n25837 = ( n1695 & n4817 ) | ( n1695 & n12115 ) | ( n4817 & n12115 ) ;
  assign n25835 = ( n1414 & ~n9989 ) | ( n1414 & n20507 ) | ( ~n9989 & n20507 ) ;
  assign n25836 = n25835 ^ n8716 ^ n6325 ;
  assign n25839 = n25838 ^ n25837 ^ n25836 ;
  assign n25840 = n4955 & ~n22436 ;
  assign n25841 = n25839 & n25840 ;
  assign n25842 = ( n12123 & n25834 ) | ( n12123 & n25841 ) | ( n25834 & n25841 ) ;
  assign n25843 = ( ~n1657 & n1725 ) | ( ~n1657 & n1775 ) | ( n1725 & n1775 ) ;
  assign n25844 = ( n12521 & n12888 ) | ( n12521 & ~n16263 ) | ( n12888 & ~n16263 ) ;
  assign n25845 = ~n6817 & n9192 ;
  assign n25846 = ~n4574 & n25845 ;
  assign n25847 = n8209 ^ n4414 ^ 1'b0 ;
  assign n25848 = ~n3703 & n25847 ;
  assign n25849 = n25846 | n25848 ;
  assign n25850 = ~n3668 & n9762 ;
  assign n25851 = n25850 ^ n21649 ^ 1'b0 ;
  assign n25852 = n5666 & ~n16701 ;
  assign n25853 = n25852 ^ n10800 ^ 1'b0 ;
  assign n25854 = ~n3545 & n3640 ;
  assign n25855 = ( ~n8731 & n19590 ) | ( ~n8731 & n25854 ) | ( n19590 & n25854 ) ;
  assign n25856 = n6446 & n13751 ;
  assign n25857 = n25856 ^ n20419 ^ 1'b0 ;
  assign n25858 = n25857 ^ n12468 ^ 1'b0 ;
  assign n25859 = n22455 ^ n3583 ^ n1799 ;
  assign n25860 = n25362 ^ n22557 ^ 1'b0 ;
  assign n25861 = ( n5719 & n16241 ) | ( n5719 & n17401 ) | ( n16241 & n17401 ) ;
  assign n25862 = n12679 ^ n10351 ^ n3657 ;
  assign n25863 = ( n406 & n4465 ) | ( n406 & n6513 ) | ( n4465 & n6513 ) ;
  assign n25864 = ( ~n24106 & n24772 ) | ( ~n24106 & n25863 ) | ( n24772 & n25863 ) ;
  assign n25865 = n2153 & n8774 ;
  assign n25866 = ~n4606 & n25865 ;
  assign n25868 = n19276 ^ n9274 ^ n4190 ;
  assign n25867 = n25505 ^ n22151 ^ n16754 ;
  assign n25869 = n25868 ^ n25867 ^ n8801 ;
  assign n25870 = n23835 ^ n12698 ^ n725 ;
  assign n25871 = ( n4732 & n11709 ) | ( n4732 & ~n19702 ) | ( n11709 & ~n19702 ) ;
  assign n25872 = n25871 ^ n11984 ^ 1'b0 ;
  assign n25873 = n25870 | n25872 ;
  assign n25874 = n25869 & ~n25873 ;
  assign n25875 = ( n270 & ~n10632 ) | ( n270 & n10983 ) | ( ~n10632 & n10983 ) ;
  assign n25876 = n25875 ^ n18888 ^ n2981 ;
  assign n25877 = n18877 ^ n16949 ^ n7911 ;
  assign n25878 = ( n3114 & ~n25876 ) | ( n3114 & n25877 ) | ( ~n25876 & n25877 ) ;
  assign n25879 = ( n4539 & n13321 ) | ( n4539 & ~n25878 ) | ( n13321 & ~n25878 ) ;
  assign n25880 = ( n2504 & ~n14187 ) | ( n2504 & n19275 ) | ( ~n14187 & n19275 ) ;
  assign n25881 = n8034 | n23808 ;
  assign n25882 = n13005 | n23629 ;
  assign n25883 = ( n3031 & n13371 ) | ( n3031 & n25882 ) | ( n13371 & n25882 ) ;
  assign n25884 = n4524 ^ n3965 ^ n1560 ;
  assign n25885 = ( n6728 & n22029 ) | ( n6728 & n25884 ) | ( n22029 & n25884 ) ;
  assign n25891 = n20624 ^ n4975 ^ n4973 ;
  assign n25892 = n25891 ^ n21164 ^ n1032 ;
  assign n25889 = n18833 ^ n5911 ^ n5077 ;
  assign n25887 = n25795 ^ n4889 ^ 1'b0 ;
  assign n25888 = n1780 & ~n25887 ;
  assign n25886 = n8513 ^ n4729 ^ n1434 ;
  assign n25890 = n25889 ^ n25888 ^ n25886 ;
  assign n25893 = n25892 ^ n25890 ^ n15803 ;
  assign n25894 = n16760 ^ n10771 ^ n3982 ;
  assign n25895 = n23483 ^ n11669 ^ n6613 ;
  assign n25896 = n25895 ^ n10242 ^ n5921 ;
  assign n25897 = ( n2609 & n4532 ) | ( n2609 & n5680 ) | ( n4532 & n5680 ) ;
  assign n25898 = n25897 ^ n11718 ^ n5809 ;
  assign n25899 = ( n8724 & n12600 ) | ( n8724 & n25898 ) | ( n12600 & n25898 ) ;
  assign n25900 = ( ~n3102 & n12115 ) | ( ~n3102 & n14584 ) | ( n12115 & n14584 ) ;
  assign n25901 = n5356 | n19598 ;
  assign n25902 = n22923 & ~n25901 ;
  assign n25903 = ( n3430 & n15652 ) | ( n3430 & n25902 ) | ( n15652 & n25902 ) ;
  assign n25904 = n25903 ^ n15258 ^ n6822 ;
  assign n25906 = ( n5065 & n7284 ) | ( n5065 & n11611 ) | ( n7284 & n11611 ) ;
  assign n25905 = n19463 ^ n14131 ^ 1'b0 ;
  assign n25907 = n25906 ^ n25905 ^ n3297 ;
  assign n25909 = n24425 ^ n15850 ^ n10404 ;
  assign n25908 = n6218 ^ n2434 ^ n841 ;
  assign n25910 = n25909 ^ n25908 ^ n4326 ;
  assign n25911 = n9161 ^ n6073 ^ n1617 ;
  assign n25912 = n25911 ^ n16609 ^ n7726 ;
  assign n25913 = n23326 ^ n21754 ^ n14734 ;
  assign n25914 = n9110 ^ n4930 ^ n429 ;
  assign n25915 = ( n11247 & ~n14807 ) | ( n11247 & n25914 ) | ( ~n14807 & n25914 ) ;
  assign n25916 = ~n1854 & n24913 ;
  assign n25917 = ~n25258 & n25916 ;
  assign n25918 = n10465 ^ n9790 ^ 1'b0 ;
  assign n25919 = n1304 & ~n5287 ;
  assign n25920 = n25919 ^ n3082 ^ 1'b0 ;
  assign n25921 = n25920 ^ n20322 ^ 1'b0 ;
  assign n25922 = ~n4948 & n25921 ;
  assign n25923 = n14545 ^ n9447 ^ n4165 ;
  assign n25924 = n24072 & n25923 ;
  assign n25925 = n23148 ^ n16926 ^ n8684 ;
  assign n25926 = ( n25922 & n25924 ) | ( n25922 & ~n25925 ) | ( n25924 & ~n25925 ) ;
  assign n25927 = ( n10381 & n16796 ) | ( n10381 & n25926 ) | ( n16796 & n25926 ) ;
  assign n25930 = ( n1076 & n12036 ) | ( n1076 & n21334 ) | ( n12036 & n21334 ) ;
  assign n25928 = n7168 | n8701 ;
  assign n25929 = n25928 ^ n22124 ^ n10583 ;
  assign n25931 = n25930 ^ n25929 ^ n3823 ;
  assign n25932 = ( n15319 & ~n15956 ) | ( n15319 & n25931 ) | ( ~n15956 & n25931 ) ;
  assign n25933 = n948 | n8696 ;
  assign n25934 = n22546 ^ n4831 ^ n668 ;
  assign n25935 = ( ~n5684 & n25933 ) | ( ~n5684 & n25934 ) | ( n25933 & n25934 ) ;
  assign n25936 = n2225 & ~n11566 ;
  assign n25937 = n25936 ^ n24157 ^ 1'b0 ;
  assign n25938 = n21389 ^ n11177 ^ 1'b0 ;
  assign n25943 = ( n1582 & n15898 ) | ( n1582 & ~n18346 ) | ( n15898 & ~n18346 ) ;
  assign n25940 = n8000 & n14352 ;
  assign n25941 = n25940 ^ n9551 ^ 1'b0 ;
  assign n25942 = ( ~n306 & n17653 ) | ( ~n306 & n25941 ) | ( n17653 & n25941 ) ;
  assign n25939 = n8624 | n16047 ;
  assign n25944 = n25943 ^ n25942 ^ n25939 ;
  assign n25945 = n15351 ^ n8027 ^ n3873 ;
  assign n25946 = n20863 ^ n18306 ^ n16209 ;
  assign n25947 = ( n12076 & ~n13183 ) | ( n12076 & n25946 ) | ( ~n13183 & n25946 ) ;
  assign n25948 = ( ~n20958 & n25945 ) | ( ~n20958 & n25947 ) | ( n25945 & n25947 ) ;
  assign n25949 = ( n2524 & ~n10907 ) | ( n2524 & n23879 ) | ( ~n10907 & n23879 ) ;
  assign n25950 = n24754 ^ n21255 ^ n20585 ;
  assign n25951 = n15614 ^ n14262 ^ n11720 ;
  assign n25952 = ( n15587 & n25371 ) | ( n15587 & ~n25951 ) | ( n25371 & ~n25951 ) ;
  assign n25953 = ( n6536 & ~n25217 ) | ( n6536 & n25514 ) | ( ~n25217 & n25514 ) ;
  assign n25954 = n13194 ^ n6281 ^ x84 ;
  assign n25955 = n22331 & ~n25954 ;
  assign n25956 = n21092 ^ n16906 ^ 1'b0 ;
  assign n25957 = ~n9670 & n25956 ;
  assign n25958 = n14877 ^ n5668 ^ n4472 ;
  assign n25959 = n4388 & n25958 ;
  assign n25961 = n17802 ^ n8337 ^ 1'b0 ;
  assign n25960 = n24103 ^ n20186 ^ n8639 ;
  assign n25962 = n25961 ^ n25960 ^ n7496 ;
  assign n25963 = ~n9807 & n14985 ;
  assign n25964 = n23088 ^ n5956 ^ n2480 ;
  assign n25965 = n16747 ^ n10580 ^ 1'b0 ;
  assign n25966 = n11577 & ~n25965 ;
  assign n25967 = n25966 ^ n2202 ^ 1'b0 ;
  assign n25968 = n2764 | n25967 ;
  assign n25969 = n3994 | n25968 ;
  assign n25970 = n22603 ^ n7958 ^ n3273 ;
  assign n25971 = ( n3686 & n7727 ) | ( n3686 & ~n7885 ) | ( n7727 & ~n7885 ) ;
  assign n25972 = n9904 & ~n25971 ;
  assign n25973 = n25972 ^ n24767 ^ 1'b0 ;
  assign n25974 = ~n7507 & n19694 ;
  assign n25975 = n25974 ^ n4045 ^ 1'b0 ;
  assign n25976 = ( n10618 & n10686 ) | ( n10618 & n25975 ) | ( n10686 & n25975 ) ;
  assign n25977 = ( x58 & ~n1006 ) | ( x58 & n3614 ) | ( ~n1006 & n3614 ) ;
  assign n25978 = n7065 ^ n5975 ^ n4895 ;
  assign n25979 = ~n3035 & n9987 ;
  assign n25980 = n25979 ^ n1657 ^ 1'b0 ;
  assign n25981 = ( ~n1691 & n17390 ) | ( ~n1691 & n25980 ) | ( n17390 & n25980 ) ;
  assign n25982 = n12026 ^ n3561 ^ n1588 ;
  assign n25983 = ( n1749 & n24095 ) | ( n1749 & n25982 ) | ( n24095 & n25982 ) ;
  assign n25985 = n2948 ^ n2653 ^ 1'b0 ;
  assign n25984 = n1675 | n17438 ;
  assign n25986 = n25985 ^ n25984 ^ n25696 ;
  assign n25987 = ~n1049 & n3559 ;
  assign n25988 = n25987 ^ n17532 ^ 1'b0 ;
  assign n25989 = n25988 ^ n8986 ^ n6446 ;
  assign n25990 = ~n25983 & n25989 ;
  assign n25991 = n25990 ^ n2437 ^ 1'b0 ;
  assign n25992 = n22140 | n22940 ;
  assign n25993 = n5932 | n25992 ;
  assign n25994 = n8306 & n25993 ;
  assign n25995 = ~n4167 & n25994 ;
  assign n26003 = ( n239 & ~n18817 ) | ( n239 & n21495 ) | ( ~n18817 & n21495 ) ;
  assign n26001 = n19639 ^ n18192 ^ n5272 ;
  assign n25998 = n1462 & ~n24222 ;
  assign n25999 = ~n10762 & n25998 ;
  assign n25996 = ( n412 & ~n799 ) | ( n412 & n1264 ) | ( ~n799 & n1264 ) ;
  assign n25997 = ( n5954 & n13870 ) | ( n5954 & n25996 ) | ( n13870 & n25996 ) ;
  assign n26000 = n25999 ^ n25997 ^ n22723 ;
  assign n26002 = n26001 ^ n26000 ^ n17779 ;
  assign n26004 = n26003 ^ n26002 ^ n8364 ;
  assign n26005 = ( n3882 & n21136 ) | ( n3882 & ~n21260 ) | ( n21136 & ~n21260 ) ;
  assign n26006 = ( n9271 & ~n16664 ) | ( n9271 & n23786 ) | ( ~n16664 & n23786 ) ;
  assign n26007 = ( ~n763 & n4598 ) | ( ~n763 & n22512 ) | ( n4598 & n22512 ) ;
  assign n26013 = n8350 ^ n5928 ^ 1'b0 ;
  assign n26014 = ~n7328 & n26013 ;
  assign n26009 = n18222 ^ n4581 ^ n1732 ;
  assign n26008 = ( n857 & ~n14154 ) | ( n857 & n16066 ) | ( ~n14154 & n16066 ) ;
  assign n26010 = n26009 ^ n26008 ^ n5546 ;
  assign n26011 = n2095 | n26010 ;
  assign n26012 = ( ~n9656 & n18032 ) | ( ~n9656 & n26011 ) | ( n18032 & n26011 ) ;
  assign n26015 = n26014 ^ n26012 ^ n21348 ;
  assign n26016 = ( n1317 & n1422 ) | ( n1317 & n15214 ) | ( n1422 & n15214 ) ;
  assign n26017 = n26016 ^ n18163 ^ 1'b0 ;
  assign n26018 = n5998 | n26017 ;
  assign n26019 = n26018 ^ n16150 ^ 1'b0 ;
  assign n26020 = n5221 & n10790 ;
  assign n26021 = ~n14171 & n26020 ;
  assign n26022 = ~n4883 & n19861 ;
  assign n26023 = n26022 ^ n14100 ^ 1'b0 ;
  assign n26024 = n24674 & ~n26023 ;
  assign n26026 = n6985 ^ n4939 ^ x30 ;
  assign n26025 = n18082 ^ n13918 ^ n3867 ;
  assign n26027 = n26026 ^ n26025 ^ n20150 ;
  assign n26028 = ( n4065 & n4202 ) | ( n4065 & ~n11971 ) | ( n4202 & ~n11971 ) ;
  assign n26029 = n26028 ^ n25869 ^ n23725 ;
  assign n26030 = ( n12553 & n17091 ) | ( n12553 & ~n24205 ) | ( n17091 & ~n24205 ) ;
  assign n26031 = n862 & ~n8302 ;
  assign n26032 = n26031 ^ n9045 ^ 1'b0 ;
  assign n26033 = ( ~n9608 & n19797 ) | ( ~n9608 & n25640 ) | ( n19797 & n25640 ) ;
  assign n26034 = ( n5932 & n26032 ) | ( n5932 & n26033 ) | ( n26032 & n26033 ) ;
  assign n26035 = ( n761 & n9216 ) | ( n761 & ~n10782 ) | ( n9216 & ~n10782 ) ;
  assign n26037 = n16352 ^ n1244 ^ 1'b0 ;
  assign n26036 = ( n8679 & ~n14000 ) | ( n8679 & n16393 ) | ( ~n14000 & n16393 ) ;
  assign n26038 = n26037 ^ n26036 ^ n14056 ;
  assign n26039 = ( ~x26 & n9683 ) | ( ~x26 & n21301 ) | ( n9683 & n21301 ) ;
  assign n26040 = n26039 ^ n14026 ^ n1731 ;
  assign n26041 = n4563 & n26040 ;
  assign n26042 = n26041 ^ n11511 ^ 1'b0 ;
  assign n26043 = ( n5132 & ~n11757 ) | ( n5132 & n17116 ) | ( ~n11757 & n17116 ) ;
  assign n26044 = n12187 & n26043 ;
  assign n26045 = n16483 ^ n14079 ^ n3344 ;
  assign n26046 = ( n211 & ~n1354 ) | ( n211 & n13365 ) | ( ~n1354 & n13365 ) ;
  assign n26047 = ~n4804 & n26046 ;
  assign n26048 = ( ~n6382 & n6597 ) | ( ~n6382 & n26047 ) | ( n6597 & n26047 ) ;
  assign n26049 = n26048 ^ n12473 ^ n1174 ;
  assign n26050 = n26049 ^ n9584 ^ n5232 ;
  assign n26051 = n2760 | n14905 ;
  assign n26052 = n496 | n26051 ;
  assign n26053 = ( n18751 & ~n20287 ) | ( n18751 & n26052 ) | ( ~n20287 & n26052 ) ;
  assign n26054 = ( n26045 & n26050 ) | ( n26045 & n26053 ) | ( n26050 & n26053 ) ;
  assign n26055 = ( n2888 & n3789 ) | ( n2888 & n4499 ) | ( n3789 & n4499 ) ;
  assign n26056 = ( n1419 & n4091 ) | ( n1419 & n26055 ) | ( n4091 & n26055 ) ;
  assign n26057 = ( n1416 & n12216 ) | ( n1416 & ~n25837 ) | ( n12216 & ~n25837 ) ;
  assign n26058 = n26057 ^ n15879 ^ n12032 ;
  assign n26059 = n16047 ^ n4700 ^ 1'b0 ;
  assign n26060 = n26058 & n26059 ;
  assign n26061 = n24026 ^ n15726 ^ n2489 ;
  assign n26062 = n26061 ^ n4680 ^ n434 ;
  assign n26063 = ( ~n26056 & n26060 ) | ( ~n26056 & n26062 ) | ( n26060 & n26062 ) ;
  assign n26064 = n15793 ^ n1662 ^ n1298 ;
  assign n26065 = n16791 ^ n3373 ^ n1388 ;
  assign n26067 = ( n2797 & n13442 ) | ( n2797 & ~n18048 ) | ( n13442 & ~n18048 ) ;
  assign n26066 = ( n2846 & ~n6094 ) | ( n2846 & n13156 ) | ( ~n6094 & n13156 ) ;
  assign n26068 = n26067 ^ n26066 ^ n2207 ;
  assign n26069 = n23965 ^ n21055 ^ n1210 ;
  assign n26070 = x5 | n9981 ;
  assign n26071 = n26070 ^ n20122 ^ 1'b0 ;
  assign n26072 = n22349 ^ n21591 ^ 1'b0 ;
  assign n26073 = ( n18072 & ~n26071 ) | ( n18072 & n26072 ) | ( ~n26071 & n26072 ) ;
  assign n26075 = n10446 ^ n7130 ^ n170 ;
  assign n26074 = n862 & n12195 ;
  assign n26076 = n26075 ^ n26074 ^ 1'b0 ;
  assign n26077 = ( n4630 & ~n12833 ) | ( n4630 & n21339 ) | ( ~n12833 & n21339 ) ;
  assign n26078 = ( n1941 & n3530 ) | ( n1941 & n10875 ) | ( n3530 & n10875 ) ;
  assign n26079 = ~n4162 & n26078 ;
  assign n26080 = ( ~n7207 & n15140 ) | ( ~n7207 & n20171 ) | ( n15140 & n20171 ) ;
  assign n26081 = n9557 & ~n19609 ;
  assign n26082 = n4227 | n20834 ;
  assign n26083 = ( ~n18292 & n26081 ) | ( ~n18292 & n26082 ) | ( n26081 & n26082 ) ;
  assign n26084 = n19577 ^ n17309 ^ n9098 ;
  assign n26085 = n26084 ^ n22178 ^ n19208 ;
  assign n26087 = ( n1022 & ~n4698 ) | ( n1022 & n24491 ) | ( ~n4698 & n24491 ) ;
  assign n26086 = n16513 ^ n10706 ^ n4194 ;
  assign n26088 = n26087 ^ n26086 ^ n20352 ;
  assign n26089 = n3038 & ~n17141 ;
  assign n26090 = n26089 ^ n4269 ^ 1'b0 ;
  assign n26091 = n26090 ^ n23511 ^ n298 ;
  assign n26092 = n20446 ^ n15498 ^ n15340 ;
  assign n26093 = n14379 ^ n7139 ^ 1'b0 ;
  assign n26094 = n26092 | n26093 ;
  assign n26095 = n18719 ^ n16233 ^ 1'b0 ;
  assign n26096 = ~n474 & n13831 ;
  assign n26097 = n26096 ^ n10534 ^ 1'b0 ;
  assign n26098 = ( n3467 & n7190 ) | ( n3467 & n10892 ) | ( n7190 & n10892 ) ;
  assign n26099 = ( ~n2054 & n16066 ) | ( ~n2054 & n26098 ) | ( n16066 & n26098 ) ;
  assign n26100 = n1711 & ~n2363 ;
  assign n26101 = n7317 & ~n26100 ;
  assign n26102 = ( n813 & n3301 ) | ( n813 & ~n16248 ) | ( n3301 & ~n16248 ) ;
  assign n26103 = ( n9262 & n14017 ) | ( n9262 & ~n15137 ) | ( n14017 & ~n15137 ) ;
  assign n26104 = ( ~n26101 & n26102 ) | ( ~n26101 & n26103 ) | ( n26102 & n26103 ) ;
  assign n26105 = n6901 ^ n4363 ^ 1'b0 ;
  assign n26106 = ( n5351 & n18168 ) | ( n5351 & n26105 ) | ( n18168 & n26105 ) ;
  assign n26107 = ( n5611 & n16837 ) | ( n5611 & n26106 ) | ( n16837 & n26106 ) ;
  assign n26108 = ~n6766 & n9835 ;
  assign n26109 = n26108 ^ n19356 ^ n17574 ;
  assign n26110 = n26109 ^ n5257 ^ 1'b0 ;
  assign n26111 = n6513 ^ n186 ^ 1'b0 ;
  assign n26112 = n20822 ^ n16467 ^ n11704 ;
  assign n26113 = ( ~n21631 & n26111 ) | ( ~n21631 & n26112 ) | ( n26111 & n26112 ) ;
  assign n26114 = n26113 ^ n12082 ^ n7261 ;
  assign n26117 = n5672 ^ n3176 ^ 1'b0 ;
  assign n26118 = n6179 | n26117 ;
  assign n26119 = n26118 ^ n12068 ^ n6034 ;
  assign n26120 = n26119 ^ n8687 ^ n5047 ;
  assign n26115 = ~n8386 & n19178 ;
  assign n26116 = ( n5813 & n13853 ) | ( n5813 & ~n26115 ) | ( n13853 & ~n26115 ) ;
  assign n26121 = n26120 ^ n26116 ^ n19155 ;
  assign n26122 = ~n3045 & n18722 ;
  assign n26123 = ( n3637 & n5962 ) | ( n3637 & n7132 ) | ( n5962 & n7132 ) ;
  assign n26124 = n26123 ^ n3189 ^ 1'b0 ;
  assign n26125 = n26124 ^ n8064 ^ n4032 ;
  assign n26126 = n14836 ^ n3137 ^ n1559 ;
  assign n26127 = n9605 ^ n5477 ^ 1'b0 ;
  assign n26128 = n26126 & ~n26127 ;
  assign n26129 = ( ~n14021 & n15969 ) | ( ~n14021 & n22166 ) | ( n15969 & n22166 ) ;
  assign n26130 = n26129 ^ n24767 ^ 1'b0 ;
  assign n26131 = ~n16666 & n26130 ;
  assign n26132 = ( ~n1457 & n13532 ) | ( ~n1457 & n25211 ) | ( n13532 & n25211 ) ;
  assign n26133 = ( n4876 & n22222 ) | ( n4876 & ~n26132 ) | ( n22222 & ~n26132 ) ;
  assign n26134 = n17446 ^ n17271 ^ n13391 ;
  assign n26135 = ( n7924 & n16168 ) | ( n7924 & ~n26134 ) | ( n16168 & ~n26134 ) ;
  assign n26136 = n22792 ^ n14158 ^ 1'b0 ;
  assign n26137 = n25373 ^ n21677 ^ 1'b0 ;
  assign n26138 = n14286 ^ n4181 ^ 1'b0 ;
  assign n26139 = n26138 ^ n20754 ^ n16909 ;
  assign n26140 = n26139 ^ n14420 ^ n12679 ;
  assign n26141 = n18324 ^ n9384 ^ 1'b0 ;
  assign n26142 = n26141 ^ n22370 ^ n7071 ;
  assign n26143 = n12816 ^ n6765 ^ n185 ;
  assign n26144 = n26143 ^ n6624 ^ 1'b0 ;
  assign n26145 = n18914 ^ n8063 ^ n7378 ;
  assign n26146 = ( ~n3810 & n7646 ) | ( ~n3810 & n14354 ) | ( n7646 & n14354 ) ;
  assign n26147 = n18373 ^ n5211 ^ 1'b0 ;
  assign n26148 = n26147 ^ n8502 ^ n2997 ;
  assign n26149 = ( n4681 & ~n9534 ) | ( n4681 & n26148 ) | ( ~n9534 & n26148 ) ;
  assign n26150 = ( n9864 & n13374 ) | ( n9864 & n26149 ) | ( n13374 & n26149 ) ;
  assign n26151 = n23514 ^ n7769 ^ n4285 ;
  assign n26152 = ( n9665 & ~n14736 ) | ( n9665 & n23791 ) | ( ~n14736 & n23791 ) ;
  assign n26153 = ~n14943 & n22001 ;
  assign n26154 = ( x44 & n3752 ) | ( x44 & n26153 ) | ( n3752 & n26153 ) ;
  assign n26155 = n9851 ^ n2412 ^ 1'b0 ;
  assign n26156 = n26155 ^ n25943 ^ n19464 ;
  assign n26157 = ~n24207 & n26156 ;
  assign n26158 = n26157 ^ n1954 ^ 1'b0 ;
  assign n26159 = n20625 ^ n19243 ^ n5551 ;
  assign n26160 = n11421 & n26159 ;
  assign n26161 = ~n4127 & n26160 ;
  assign n26162 = ( n2601 & n8500 ) | ( n2601 & ~n22087 ) | ( n8500 & ~n22087 ) ;
  assign n26163 = ( n5702 & n6015 ) | ( n5702 & n11480 ) | ( n6015 & n11480 ) ;
  assign n26164 = n21312 ^ n20993 ^ n4162 ;
  assign n26165 = n11087 | n26164 ;
  assign n26166 = ( n26162 & ~n26163 ) | ( n26162 & n26165 ) | ( ~n26163 & n26165 ) ;
  assign n26167 = n7675 | n10030 ;
  assign n26168 = n18962 & ~n26167 ;
  assign n26169 = ( n1425 & n11174 ) | ( n1425 & n26168 ) | ( n11174 & n26168 ) ;
  assign n26170 = n26169 ^ n20615 ^ n6261 ;
  assign n26171 = ( n11661 & n19432 ) | ( n11661 & ~n26170 ) | ( n19432 & ~n26170 ) ;
  assign n26172 = n26171 ^ n15084 ^ n3555 ;
  assign n26173 = n20267 ^ n18719 ^ n8982 ;
  assign n26174 = ( n17696 & n19134 ) | ( n17696 & n26173 ) | ( n19134 & n26173 ) ;
  assign n26175 = ( n13146 & n18416 ) | ( n13146 & ~n22144 ) | ( n18416 & ~n22144 ) ;
  assign n26176 = ( n3370 & n25531 ) | ( n3370 & ~n26175 ) | ( n25531 & ~n26175 ) ;
  assign n26177 = n22621 ^ n9597 ^ n829 ;
  assign n26179 = n15436 ^ n14972 ^ 1'b0 ;
  assign n26180 = n18826 & n26179 ;
  assign n26178 = ( n10687 & ~n12118 ) | ( n10687 & n23915 ) | ( ~n12118 & n23915 ) ;
  assign n26181 = n26180 ^ n26178 ^ n7106 ;
  assign n26182 = ~n8749 & n25316 ;
  assign n26183 = n24059 & n26182 ;
  assign n26184 = n15521 ^ n6262 ^ n5165 ;
  assign n26185 = ~n7427 & n26184 ;
  assign n26186 = n5256 & n26185 ;
  assign n26187 = n26186 ^ n23958 ^ n5671 ;
  assign n26188 = n16051 ^ n10621 ^ n6210 ;
  assign n26189 = ( n2336 & ~n6867 ) | ( n2336 & n18058 ) | ( ~n6867 & n18058 ) ;
  assign n26190 = n8431 ^ n4871 ^ 1'b0 ;
  assign n26191 = ( n14039 & n26189 ) | ( n14039 & ~n26190 ) | ( n26189 & ~n26190 ) ;
  assign n26192 = ( x65 & n5666 ) | ( x65 & n12237 ) | ( n5666 & n12237 ) ;
  assign n26193 = n26192 ^ n20434 ^ n7536 ;
  assign n26194 = n25011 ^ n19199 ^ n3814 ;
  assign n26195 = ( ~n11720 & n13791 ) | ( ~n11720 & n26194 ) | ( n13791 & n26194 ) ;
  assign n26196 = n21270 ^ n19060 ^ n8053 ;
  assign n26197 = n26196 ^ n10115 ^ n9436 ;
  assign n26198 = n3591 & ~n26197 ;
  assign n26199 = n18323 & n26198 ;
  assign n26200 = n465 & ~n15326 ;
  assign n26201 = ~n23023 & n26200 ;
  assign n26202 = n13723 ^ n8175 ^ n4841 ;
  assign n26203 = n3192 ^ n2615 ^ n1142 ;
  assign n26204 = ( ~n11948 & n26202 ) | ( ~n11948 & n26203 ) | ( n26202 & n26203 ) ;
  assign n26205 = n2556 & n15353 ;
  assign n26206 = n7691 ^ n4802 ^ 1'b0 ;
  assign n26207 = ( ~n2024 & n4386 ) | ( ~n2024 & n11631 ) | ( n4386 & n11631 ) ;
  assign n26208 = n3814 | n12966 ;
  assign n26209 = ( ~n26206 & n26207 ) | ( ~n26206 & n26208 ) | ( n26207 & n26208 ) ;
  assign n26210 = n8873 ^ n8235 ^ x67 ;
  assign n26211 = n26210 ^ n15275 ^ n13407 ;
  assign n26212 = ( ~n21338 & n21521 ) | ( ~n21338 & n26211 ) | ( n21521 & n26211 ) ;
  assign n26213 = n10417 ^ n557 ^ n344 ;
  assign n26214 = n26213 ^ n9400 ^ n5412 ;
  assign n26215 = ( ~n1970 & n4898 ) | ( ~n1970 & n14249 ) | ( n4898 & n14249 ) ;
  assign n26216 = n26215 ^ n12042 ^ 1'b0 ;
  assign n26217 = n16358 ^ n10610 ^ 1'b0 ;
  assign n26218 = ( n4901 & ~n8377 ) | ( n4901 & n26217 ) | ( ~n8377 & n26217 ) ;
  assign n26219 = ( n11430 & ~n26216 ) | ( n11430 & n26218 ) | ( ~n26216 & n26218 ) ;
  assign n26220 = n22875 ^ n11909 ^ n917 ;
  assign n26221 = ( n7486 & n11145 ) | ( n7486 & n12488 ) | ( n11145 & n12488 ) ;
  assign n26222 = n26221 ^ n12272 ^ 1'b0 ;
  assign n26223 = n26220 & ~n26222 ;
  assign n26224 = n22741 ^ n8014 ^ 1'b0 ;
  assign n26225 = n2622 & n26224 ;
  assign n26226 = ( ~n3423 & n7041 ) | ( ~n3423 & n26225 ) | ( n7041 & n26225 ) ;
  assign n26227 = ~n2389 & n26226 ;
  assign n26228 = n6653 & ~n22588 ;
  assign n26229 = n26228 ^ n13437 ^ n376 ;
  assign n26230 = ( n11852 & n17286 ) | ( n11852 & n19394 ) | ( n17286 & n19394 ) ;
  assign n26231 = n15866 ^ n13744 ^ n575 ;
  assign n26232 = ( n10296 & n13751 ) | ( n10296 & ~n26231 ) | ( n13751 & ~n26231 ) ;
  assign n26233 = ( n5029 & ~n12018 ) | ( n5029 & n15784 ) | ( ~n12018 & n15784 ) ;
  assign n26234 = ( n3258 & n19256 ) | ( n3258 & n26233 ) | ( n19256 & n26233 ) ;
  assign n26235 = ( n1528 & n4424 ) | ( n1528 & ~n4485 ) | ( n4424 & ~n4485 ) ;
  assign n26236 = ( n21405 & n24281 ) | ( n21405 & n26235 ) | ( n24281 & n26235 ) ;
  assign n26237 = ( n988 & ~n19968 ) | ( n988 & n26236 ) | ( ~n19968 & n26236 ) ;
  assign n26238 = n26237 ^ n25665 ^ n7089 ;
  assign n26239 = n21632 ^ n15052 ^ n12033 ;
  assign n26240 = ( n3178 & n8431 ) | ( n3178 & n19788 ) | ( n8431 & n19788 ) ;
  assign n26241 = n26240 ^ n529 ^ 1'b0 ;
  assign n26242 = n9455 & n10670 ;
  assign n26243 = n18398 ^ n7349 ^ n5148 ;
  assign n26244 = n26243 ^ n10869 ^ n4550 ;
  assign n26245 = n26244 ^ n10112 ^ n841 ;
  assign n26246 = n13789 ^ n5471 ^ n5406 ;
  assign n26247 = ( n4650 & n8000 ) | ( n4650 & n11306 ) | ( n8000 & n11306 ) ;
  assign n26248 = ( ~n2995 & n21022 ) | ( ~n2995 & n26247 ) | ( n21022 & n26247 ) ;
  assign n26250 = n1058 & ~n14548 ;
  assign n26251 = n26250 ^ n10763 ^ 1'b0 ;
  assign n26249 = n12267 ^ n1505 ^ x46 ;
  assign n26252 = n26251 ^ n26249 ^ n5247 ;
  assign n26253 = ( n8743 & n16820 ) | ( n8743 & n23291 ) | ( n16820 & n23291 ) ;
  assign n26254 = n6152 ^ n1560 ^ n879 ;
  assign n26255 = ( n18769 & n18821 ) | ( n18769 & n26254 ) | ( n18821 & n26254 ) ;
  assign n26256 = n26255 ^ n18407 ^ n16424 ;
  assign n26257 = ( n1717 & n6084 ) | ( n1717 & ~n6275 ) | ( n6084 & ~n6275 ) ;
  assign n26258 = n26257 ^ n9005 ^ 1'b0 ;
  assign n26259 = ~n6154 & n26258 ;
  assign n26260 = n26259 ^ n14157 ^ 1'b0 ;
  assign n26261 = n9884 & n26260 ;
  assign n26262 = n8333 ^ n3581 ^ 1'b0 ;
  assign n26263 = n20587 ^ n4791 ^ x53 ;
  assign n26264 = ( ~n9279 & n26262 ) | ( ~n9279 & n26263 ) | ( n26262 & n26263 ) ;
  assign n26265 = n17012 ^ n8990 ^ n4504 ;
  assign n26266 = n3056 & ~n26265 ;
  assign n26267 = ( n4646 & n11990 ) | ( n4646 & n22281 ) | ( n11990 & n22281 ) ;
  assign n26268 = n24410 ^ n18801 ^ n16055 ;
  assign n26272 = ( n7239 & n8573 ) | ( n7239 & ~n18365 ) | ( n8573 & ~n18365 ) ;
  assign n26269 = ( n4155 & n4200 ) | ( n4155 & n18732 ) | ( n4200 & n18732 ) ;
  assign n26270 = ~n25056 & n26269 ;
  assign n26271 = n6798 & n26270 ;
  assign n26273 = n26272 ^ n26271 ^ n11900 ;
  assign n26274 = ( n3605 & ~n4972 ) | ( n3605 & n8983 ) | ( ~n4972 & n8983 ) ;
  assign n26275 = ~n512 & n14623 ;
  assign n26276 = n619 ^ n171 ^ 1'b0 ;
  assign n26277 = n26276 ^ n6389 ^ n3400 ;
  assign n26278 = n26277 ^ n9247 ^ 1'b0 ;
  assign n26279 = n3735 & n11457 ;
  assign n26280 = ~n15531 & n26279 ;
  assign n26281 = n379 | n7111 ;
  assign n26282 = ( ~n5984 & n15704 ) | ( ~n5984 & n17551 ) | ( n15704 & n17551 ) ;
  assign n26283 = n18031 ^ n9556 ^ n4044 ;
  assign n26284 = ( ~n580 & n3904 ) | ( ~n580 & n11055 ) | ( n3904 & n11055 ) ;
  assign n26285 = ( n12091 & ~n25211 ) | ( n12091 & n26284 ) | ( ~n25211 & n26284 ) ;
  assign n26286 = n24965 ^ n22695 ^ n2960 ;
  assign n26287 = ( ~n1012 & n7287 ) | ( ~n1012 & n26286 ) | ( n7287 & n26286 ) ;
  assign n26288 = n25342 ^ n7916 ^ n159 ;
  assign n26289 = ( ~n582 & n26287 ) | ( ~n582 & n26288 ) | ( n26287 & n26288 ) ;
  assign n26290 = n10888 ^ n9349 ^ n2602 ;
  assign n26291 = ( n3784 & n14984 ) | ( n3784 & ~n26290 ) | ( n14984 & ~n26290 ) ;
  assign n26292 = ( n1262 & n7895 ) | ( n1262 & n26291 ) | ( n7895 & n26291 ) ;
  assign n26293 = ( ~n4597 & n10179 ) | ( ~n4597 & n17137 ) | ( n10179 & n17137 ) ;
  assign n26294 = ( n14920 & n17677 ) | ( n14920 & n26293 ) | ( n17677 & n26293 ) ;
  assign n26295 = ( ~n14791 & n19984 ) | ( ~n14791 & n26294 ) | ( n19984 & n26294 ) ;
  assign n26296 = n17197 & ~n17532 ;
  assign n26297 = ~n20862 & n26296 ;
  assign n26298 = ( ~n4104 & n5831 ) | ( ~n4104 & n8806 ) | ( n5831 & n8806 ) ;
  assign n26299 = n26298 ^ n10644 ^ n5538 ;
  assign n26300 = ~n4682 & n9524 ;
  assign n26301 = n26299 & n26300 ;
  assign n26302 = ( n3093 & n5183 ) | ( n3093 & n23138 ) | ( n5183 & n23138 ) ;
  assign n26303 = ( n1395 & n12842 ) | ( n1395 & ~n12868 ) | ( n12842 & ~n12868 ) ;
  assign n26304 = n8817 ^ n7113 ^ n3787 ;
  assign n26305 = n26304 ^ n3091 ^ 1'b0 ;
  assign n26306 = n7156 & n7532 ;
  assign n26307 = n5736 & ~n9846 ;
  assign n26308 = n26306 & n26307 ;
  assign n26309 = n26308 ^ n17015 ^ n14993 ;
  assign n26310 = ( n10986 & n17115 ) | ( n10986 & n26309 ) | ( n17115 & n26309 ) ;
  assign n26311 = ( n2055 & n26305 ) | ( n2055 & ~n26310 ) | ( n26305 & ~n26310 ) ;
  assign n26312 = n17473 ^ n9100 ^ 1'b0 ;
  assign n26313 = n15276 & n26312 ;
  assign n26314 = ( ~n3863 & n22165 ) | ( ~n3863 & n26313 ) | ( n22165 & n26313 ) ;
  assign n26315 = n14539 ^ n9616 ^ 1'b0 ;
  assign n26316 = n667 & n16356 ;
  assign n26317 = n14677 & n26316 ;
  assign n26318 = n26317 ^ n18719 ^ 1'b0 ;
  assign n26319 = n985 | n26318 ;
  assign n26320 = n6834 & n20956 ;
  assign n26321 = n26320 ^ n10889 ^ 1'b0 ;
  assign n26322 = ( n743 & ~n1561 ) | ( n743 & n3472 ) | ( ~n1561 & n3472 ) ;
  assign n26323 = ( ~n20681 & n24928 ) | ( ~n20681 & n26322 ) | ( n24928 & n26322 ) ;
  assign n26324 = n1645 & n2808 ;
  assign n26325 = ( n1600 & n24323 ) | ( n1600 & n25316 ) | ( n24323 & n25316 ) ;
  assign n26326 = n19896 & ~n26325 ;
  assign n26327 = ~n3754 & n12852 ;
  assign n26328 = ~n2540 & n26327 ;
  assign n26329 = n26328 ^ n4085 ^ 1'b0 ;
  assign n26330 = n26329 ^ n24341 ^ n21059 ;
  assign n26331 = n15671 ^ n7682 ^ n1695 ;
  assign n26332 = ( n2654 & ~n20379 ) | ( n2654 & n26331 ) | ( ~n20379 & n26331 ) ;
  assign n26333 = ( n3972 & n15488 ) | ( n3972 & n22149 ) | ( n15488 & n22149 ) ;
  assign n26339 = n17243 ^ n11638 ^ n8441 ;
  assign n26337 = n21245 ^ n12372 ^ 1'b0 ;
  assign n26338 = ~n6422 & n26337 ;
  assign n26335 = ( n3868 & ~n7329 ) | ( n3868 & n14056 ) | ( ~n7329 & n14056 ) ;
  assign n26336 = ( x25 & ~n26207 ) | ( x25 & n26335 ) | ( ~n26207 & n26335 ) ;
  assign n26340 = n26339 ^ n26338 ^ n26336 ;
  assign n26334 = n3324 & n21484 ;
  assign n26341 = n26340 ^ n26334 ^ 1'b0 ;
  assign n26342 = ~n4658 & n15854 ;
  assign n26343 = ~n21523 & n26342 ;
  assign n26344 = n9346 ^ n376 ^ 1'b0 ;
  assign n26345 = n6172 & ~n26344 ;
  assign n26346 = n26345 ^ n16478 ^ n6341 ;
  assign n26347 = ( n3370 & n3379 ) | ( n3370 & n13264 ) | ( n3379 & n13264 ) ;
  assign n26348 = ( n5994 & ~n18673 ) | ( n5994 & n24123 ) | ( ~n18673 & n24123 ) ;
  assign n26349 = n21327 ^ n16466 ^ 1'b0 ;
  assign n26350 = n26348 | n26349 ;
  assign n26351 = ( ~n9846 & n26347 ) | ( ~n9846 & n26350 ) | ( n26347 & n26350 ) ;
  assign n26352 = n18354 ^ n13371 ^ 1'b0 ;
  assign n26353 = ( n4630 & ~n5074 ) | ( n4630 & n25667 ) | ( ~n5074 & n25667 ) ;
  assign n26354 = n24987 & ~n26353 ;
  assign n26355 = ~n5121 & n26354 ;
  assign n26356 = n14723 ^ n9816 ^ 1'b0 ;
  assign n26357 = n19863 | n26356 ;
  assign n26358 = ( ~n675 & n3508 ) | ( ~n675 & n21019 ) | ( n3508 & n21019 ) ;
  assign n26359 = ( n4441 & n6150 ) | ( n4441 & ~n26358 ) | ( n6150 & ~n26358 ) ;
  assign n26360 = ( n5701 & n14669 ) | ( n5701 & ~n16898 ) | ( n14669 & ~n16898 ) ;
  assign n26361 = n8641 ^ n6087 ^ n4965 ;
  assign n26362 = n26361 ^ n15148 ^ x23 ;
  assign n26363 = n26362 ^ n16939 ^ 1'b0 ;
  assign n26364 = n8404 & n9731 ;
  assign n26365 = n26364 ^ n10957 ^ 1'b0 ;
  assign n26366 = ( n17998 & n23775 ) | ( n17998 & ~n26365 ) | ( n23775 & ~n26365 ) ;
  assign n26367 = ( n976 & ~n6470 ) | ( n976 & n21634 ) | ( ~n6470 & n21634 ) ;
  assign n26368 = n21690 ^ n11276 ^ n4088 ;
  assign n26369 = ( n1428 & ~n2521 ) | ( n1428 & n4573 ) | ( ~n2521 & n4573 ) ;
  assign n26370 = n15638 & n26369 ;
  assign n26371 = n17458 & ~n25544 ;
  assign n26372 = n26370 & n26371 ;
  assign n26373 = ( n2378 & n2766 ) | ( n2378 & ~n2774 ) | ( n2766 & ~n2774 ) ;
  assign n26374 = ( n578 & ~n17716 ) | ( n578 & n26373 ) | ( ~n17716 & n26373 ) ;
  assign n26375 = n23847 ^ n18304 ^ n16553 ;
  assign n26376 = n21809 ^ n19029 ^ n5950 ;
  assign n26377 = ( n873 & n5578 ) | ( n873 & n22028 ) | ( n5578 & n22028 ) ;
  assign n26378 = ( n1456 & ~n16067 ) | ( n1456 & n26377 ) | ( ~n16067 & n26377 ) ;
  assign n26379 = ( n9754 & n14851 ) | ( n9754 & ~n15545 ) | ( n14851 & ~n15545 ) ;
  assign n26380 = n8603 ^ n4879 ^ 1'b0 ;
  assign n26381 = ~n6329 & n26380 ;
  assign n26382 = ( ~n4612 & n17010 ) | ( ~n4612 & n26381 ) | ( n17010 & n26381 ) ;
  assign n26383 = ( ~n5990 & n17236 ) | ( ~n5990 & n26382 ) | ( n17236 & n26382 ) ;
  assign n26384 = n26383 ^ n22821 ^ n16341 ;
  assign n26385 = ~n9308 & n22537 ;
  assign n26386 = ~n19109 & n26385 ;
  assign n26387 = n10458 ^ n9622 ^ n7351 ;
  assign n26391 = n7716 ^ n7164 ^ n3458 ;
  assign n26392 = ( n4848 & n17071 ) | ( n4848 & n26391 ) | ( n17071 & n26391 ) ;
  assign n26394 = n7426 & n8325 ;
  assign n26393 = n394 & ~n4087 ;
  assign n26395 = n26394 ^ n26393 ^ 1'b0 ;
  assign n26396 = n26395 ^ n19062 ^ n4376 ;
  assign n26397 = ( n2392 & ~n26392 ) | ( n2392 & n26396 ) | ( ~n26392 & n26396 ) ;
  assign n26388 = n6214 ^ n154 ^ x11 ;
  assign n26389 = n19316 ^ n13582 ^ n477 ;
  assign n26390 = ( n951 & n26388 ) | ( n951 & n26389 ) | ( n26388 & n26389 ) ;
  assign n26398 = n26397 ^ n26390 ^ n8383 ;
  assign n26399 = n6733 | n23796 ;
  assign n26400 = n26399 ^ n18072 ^ n14584 ;
  assign n26401 = n11577 & n14154 ;
  assign n26402 = n26401 ^ n13870 ^ 1'b0 ;
  assign n26403 = ( n275 & ~n2034 ) | ( n275 & n15174 ) | ( ~n2034 & n15174 ) ;
  assign n26404 = n26403 ^ n25546 ^ n10124 ;
  assign n26405 = n14570 ^ n12567 ^ n1428 ;
  assign n26406 = n26404 & n26405 ;
  assign n26407 = ( n24341 & n26402 ) | ( n24341 & ~n26406 ) | ( n26402 & ~n26406 ) ;
  assign n26408 = n19518 ^ n3415 ^ 1'b0 ;
  assign n26409 = n15924 | n26408 ;
  assign n26410 = ( ~n8131 & n24798 ) | ( ~n8131 & n26409 ) | ( n24798 & n26409 ) ;
  assign n26411 = ( ~n646 & n2233 ) | ( ~n646 & n5795 ) | ( n2233 & n5795 ) ;
  assign n26412 = ( ~n2599 & n6299 ) | ( ~n2599 & n26411 ) | ( n6299 & n26411 ) ;
  assign n26413 = ( n20080 & ~n25045 ) | ( n20080 & n26412 ) | ( ~n25045 & n26412 ) ;
  assign n26414 = n5565 ^ n3048 ^ 1'b0 ;
  assign n26415 = n26414 ^ n14324 ^ 1'b0 ;
  assign n26416 = n23488 ^ n1903 ^ n1269 ;
  assign n26417 = ( n2920 & ~n12979 ) | ( n2920 & n15425 ) | ( ~n12979 & n15425 ) ;
  assign n26418 = ( ~n3485 & n11648 ) | ( ~n3485 & n20876 ) | ( n11648 & n20876 ) ;
  assign n26419 = ( n14851 & n26417 ) | ( n14851 & n26418 ) | ( n26417 & n26418 ) ;
  assign n26420 = n7145 ^ n6709 ^ n5598 ;
  assign n26421 = n26420 ^ n15115 ^ n1121 ;
  assign n26425 = n1841 | n7645 ;
  assign n26426 = n26425 ^ n16467 ^ n9359 ;
  assign n26427 = ( ~n18541 & n25051 ) | ( ~n18541 & n26426 ) | ( n25051 & n26426 ) ;
  assign n26423 = ( ~n4828 & n20415 ) | ( ~n4828 & n23655 ) | ( n20415 & n23655 ) ;
  assign n26422 = ( n3028 & n6592 ) | ( n3028 & ~n8709 ) | ( n6592 & ~n8709 ) ;
  assign n26424 = n26423 ^ n26422 ^ n25020 ;
  assign n26428 = n26427 ^ n26424 ^ n8214 ;
  assign n26429 = ~n366 & n25329 ;
  assign n26430 = n409 & n10942 ;
  assign n26431 = n26430 ^ n2124 ^ 1'b0 ;
  assign n26432 = n4972 | n9069 ;
  assign n26433 = n9368 | n26432 ;
  assign n26434 = n18170 ^ n3707 ^ 1'b0 ;
  assign n26435 = n26433 & n26434 ;
  assign n26436 = n6385 ^ n2346 ^ n302 ;
  assign n26437 = n26436 ^ n22565 ^ 1'b0 ;
  assign n26438 = n18424 ^ n12866 ^ n10490 ;
  assign n26439 = ( n1428 & n17184 ) | ( n1428 & ~n26438 ) | ( n17184 & ~n26438 ) ;
  assign n26440 = n9328 ^ n1712 ^ n834 ;
  assign n26441 = n5656 & n26440 ;
  assign n26442 = n14905 & n26441 ;
  assign n26443 = n26442 ^ n9479 ^ 1'b0 ;
  assign n26444 = ~n18581 & n26443 ;
  assign n26445 = n26444 ^ n2515 ^ 1'b0 ;
  assign n26451 = n3136 ^ n2438 ^ n350 ;
  assign n26449 = n2304 & ~n15472 ;
  assign n26450 = n7373 & n26449 ;
  assign n26446 = ( n6884 & ~n7138 ) | ( n6884 & n16898 ) | ( ~n7138 & n16898 ) ;
  assign n26447 = ~n3991 & n26446 ;
  assign n26448 = n12284 & n26447 ;
  assign n26452 = n26451 ^ n26450 ^ n26448 ;
  assign n26453 = ( n770 & n6006 ) | ( n770 & ~n15738 ) | ( n6006 & ~n15738 ) ;
  assign n26454 = n24613 ^ n19749 ^ n7034 ;
  assign n26455 = n26454 ^ n15702 ^ n13874 ;
  assign n26456 = ~n2132 & n11768 ;
  assign n26457 = n26456 ^ n1625 ^ 1'b0 ;
  assign n26458 = n26457 ^ n19377 ^ n4890 ;
  assign n26459 = ~n11857 & n21988 ;
  assign n26460 = n2430 | n9568 ;
  assign n26461 = n10727 ^ n6030 ^ 1'b0 ;
  assign n26462 = n26460 & ~n26461 ;
  assign n26463 = n731 ^ n546 ^ x61 ;
  assign n26464 = n26463 ^ n8008 ^ 1'b0 ;
  assign n26465 = ~n10916 & n15907 ;
  assign n26466 = ( n460 & ~n3951 ) | ( n460 & n22001 ) | ( ~n3951 & n22001 ) ;
  assign n26467 = n24420 ^ n16993 ^ n2755 ;
  assign n26468 = ( n25307 & n26466 ) | ( n25307 & n26467 ) | ( n26466 & n26467 ) ;
  assign n26469 = ~n7283 & n23687 ;
  assign n26470 = n26469 ^ n7300 ^ n7184 ;
  assign n26471 = ( n4292 & n18612 ) | ( n4292 & ~n22073 ) | ( n18612 & ~n22073 ) ;
  assign n26472 = n6191 ^ n1780 ^ 1'b0 ;
  assign n26473 = n6956 ^ n1672 ^ n172 ;
  assign n26474 = ( n12929 & ~n18855 ) | ( n12929 & n26473 ) | ( ~n18855 & n26473 ) ;
  assign n26475 = ( n172 & ~n26472 ) | ( n172 & n26474 ) | ( ~n26472 & n26474 ) ;
  assign n26476 = n26475 ^ n10651 ^ n10352 ;
  assign n26480 = ( n8368 & n8985 ) | ( n8368 & n9027 ) | ( n8985 & n9027 ) ;
  assign n26481 = n26480 ^ n25733 ^ n8020 ;
  assign n26477 = n8984 ^ n6836 ^ n5155 ;
  assign n26478 = n12435 ^ n11726 ^ 1'b0 ;
  assign n26479 = ~n26477 & n26478 ;
  assign n26482 = n26481 ^ n26479 ^ n6691 ;
  assign n26483 = n6220 ^ n5843 ^ n257 ;
  assign n26484 = ~n15174 & n26483 ;
  assign n26485 = ( ~n9799 & n22414 ) | ( ~n9799 & n26484 ) | ( n22414 & n26484 ) ;
  assign n26486 = n11592 ^ n7988 ^ 1'b0 ;
  assign n26487 = n20066 & n26486 ;
  assign n26488 = n13673 ^ n9280 ^ n2279 ;
  assign n26489 = n26488 ^ n19024 ^ n15364 ;
  assign n26490 = n4760 ^ n1674 ^ 1'b0 ;
  assign n26491 = ( n2291 & ~n9775 ) | ( n2291 & n26490 ) | ( ~n9775 & n26490 ) ;
  assign n26492 = n26491 ^ n17526 ^ n6379 ;
  assign n26493 = n12740 ^ n10829 ^ n8947 ;
  assign n26494 = ( n256 & ~n7421 ) | ( n256 & n14524 ) | ( ~n7421 & n14524 ) ;
  assign n26495 = n8365 ^ n368 ^ 1'b0 ;
  assign n26496 = n26494 & n26495 ;
  assign n26497 = ( ~n183 & n3605 ) | ( ~n183 & n26496 ) | ( n3605 & n26496 ) ;
  assign n26498 = ( n6455 & ~n24702 ) | ( n6455 & n26497 ) | ( ~n24702 & n26497 ) ;
  assign n26499 = n11373 | n26498 ;
  assign n26500 = n20194 ^ n18068 ^ 1'b0 ;
  assign n26501 = n10096 & ~n26500 ;
  assign n26502 = n26501 ^ n17398 ^ n6720 ;
  assign n26503 = n20200 ^ n11605 ^ n7514 ;
  assign n26504 = ( n5744 & n12030 ) | ( n5744 & ~n14759 ) | ( n12030 & ~n14759 ) ;
  assign n26505 = ( n23398 & n23833 ) | ( n23398 & ~n26504 ) | ( n23833 & ~n26504 ) ;
  assign n26506 = n19426 | n19774 ;
  assign n26507 = n924 | n14174 ;
  assign n26508 = n13445 ^ n12199 ^ n1112 ;
  assign n26509 = n5903 & ~n26508 ;
  assign n26510 = ( ~n3785 & n14235 ) | ( ~n3785 & n26509 ) | ( n14235 & n26509 ) ;
  assign n26511 = ( n9067 & n12242 ) | ( n9067 & n25838 ) | ( n12242 & n25838 ) ;
  assign n26512 = n3469 | n22054 ;
  assign n26513 = n19457 | n26512 ;
  assign n26514 = n26513 ^ n13507 ^ n9822 ;
  assign n26515 = ~n257 & n13748 ;
  assign n26516 = n15226 & n26515 ;
  assign n26517 = n26516 ^ n21018 ^ 1'b0 ;
  assign n26518 = ( n4070 & n12529 ) | ( n4070 & ~n14795 ) | ( n12529 & ~n14795 ) ;
  assign n26519 = ( ~n2129 & n3714 ) | ( ~n2129 & n23881 ) | ( n3714 & n23881 ) ;
  assign n26520 = n17332 ^ n11577 ^ n4752 ;
  assign n26521 = n15059 & n18446 ;
  assign n26522 = n26521 ^ n17028 ^ 1'b0 ;
  assign n26523 = n26522 ^ n20530 ^ n4295 ;
  assign n26524 = n20188 ^ n2906 ^ 1'b0 ;
  assign n26525 = n14734 ^ n11152 ^ n4766 ;
  assign n26526 = n26525 ^ n14285 ^ n2242 ;
  assign n26529 = ~n4131 & n19888 ;
  assign n26530 = n23569 & n26529 ;
  assign n26531 = n24916 | n26530 ;
  assign n26527 = n22783 ^ n16297 ^ n4309 ;
  assign n26528 = ( n5943 & n14556 ) | ( n5943 & ~n26527 ) | ( n14556 & ~n26527 ) ;
  assign n26532 = n26531 ^ n26528 ^ n8239 ;
  assign n26533 = n17474 ^ n3748 ^ 1'b0 ;
  assign n26534 = ( ~n7119 & n9212 ) | ( ~n7119 & n19238 ) | ( n9212 & n19238 ) ;
  assign n26535 = n26534 ^ n20401 ^ n16587 ;
  assign n26536 = ( n21589 & n26533 ) | ( n21589 & ~n26535 ) | ( n26533 & ~n26535 ) ;
  assign n26539 = n10295 ^ n3912 ^ n3615 ;
  assign n26540 = ( ~n1456 & n17024 ) | ( ~n1456 & n26539 ) | ( n17024 & n26539 ) ;
  assign n26538 = ( n5264 & n7590 ) | ( n5264 & ~n17682 ) | ( n7590 & ~n17682 ) ;
  assign n26537 = n24036 ^ n9235 ^ n2215 ;
  assign n26541 = n26540 ^ n26538 ^ n26537 ;
  assign n26542 = ( n1436 & ~n6676 ) | ( n1436 & n13506 ) | ( ~n6676 & n13506 ) ;
  assign n26543 = n8058 ^ n4368 ^ 1'b0 ;
  assign n26544 = n20148 ^ n17094 ^ n865 ;
  assign n26545 = ( n917 & n26543 ) | ( n917 & n26544 ) | ( n26543 & n26544 ) ;
  assign n26546 = n25264 ^ n17947 ^ x98 ;
  assign n26547 = n26546 ^ n13138 ^ n4626 ;
  assign n26548 = n26547 ^ n6934 ^ n3458 ;
  assign n26549 = n20017 ^ n7528 ^ n3079 ;
  assign n26550 = n1115 | n15060 ;
  assign n26551 = n26550 ^ n4088 ^ 1'b0 ;
  assign n26552 = n3547 & n22498 ;
  assign n26553 = n25068 ^ n13582 ^ 1'b0 ;
  assign n26554 = ( n18884 & n26009 ) | ( n18884 & ~n26553 ) | ( n26009 & ~n26553 ) ;
  assign n26555 = ( x19 & ~n2788 ) | ( x19 & n5253 ) | ( ~n2788 & n5253 ) ;
  assign n26561 = n8242 ^ n3013 ^ 1'b0 ;
  assign n26556 = n14187 ^ n8803 ^ n3897 ;
  assign n26557 = ( n356 & n9649 ) | ( n356 & ~n18853 ) | ( n9649 & ~n18853 ) ;
  assign n26558 = ( ~n23968 & n26556 ) | ( ~n23968 & n26557 ) | ( n26556 & n26557 ) ;
  assign n26559 = ( n12524 & n18006 ) | ( n12524 & ~n18634 ) | ( n18006 & ~n18634 ) ;
  assign n26560 = n26558 & ~n26559 ;
  assign n26562 = n26561 ^ n26560 ^ n9341 ;
  assign n26563 = n12023 ^ n10191 ^ n2788 ;
  assign n26564 = ( n14235 & n19803 ) | ( n14235 & ~n26563 ) | ( n19803 & ~n26563 ) ;
  assign n26565 = ( n2912 & n10644 ) | ( n2912 & n26564 ) | ( n10644 & n26564 ) ;
  assign n26566 = ( n17297 & n21076 ) | ( n17297 & ~n26565 ) | ( n21076 & ~n26565 ) ;
  assign n26567 = n21517 ^ n3063 ^ 1'b0 ;
  assign n26568 = n3253 | n5738 ;
  assign n26569 = n12000 & ~n26568 ;
  assign n26570 = ( n22144 & n24732 ) | ( n22144 & ~n26569 ) | ( n24732 & ~n26569 ) ;
  assign n26573 = ~n4350 & n8479 ;
  assign n26574 = ( n2529 & n14610 ) | ( n2529 & ~n26573 ) | ( n14610 & ~n26573 ) ;
  assign n26571 = n20072 ^ n14325 ^ n5808 ;
  assign n26572 = n9309 & n26571 ;
  assign n26575 = n26574 ^ n26572 ^ 1'b0 ;
  assign n26576 = n26575 ^ n4495 ^ n1265 ;
  assign n26577 = n8236 ^ n2764 ^ n647 ;
  assign n26578 = n26577 ^ n19088 ^ n13022 ;
  assign n26581 = n15356 ^ n13189 ^ n1551 ;
  assign n26579 = ( n1872 & n4252 ) | ( n1872 & n5507 ) | ( n4252 & n5507 ) ;
  assign n26580 = n26579 ^ n20067 ^ n18435 ;
  assign n26582 = n26581 ^ n26580 ^ n12683 ;
  assign n26588 = n9072 ^ n8247 ^ n566 ;
  assign n26585 = n14451 ^ n3652 ^ n529 ;
  assign n26583 = n6945 & n14412 ;
  assign n26584 = n26583 ^ n16619 ^ 1'b0 ;
  assign n26586 = n26585 ^ n26584 ^ 1'b0 ;
  assign n26587 = n2369 & ~n26586 ;
  assign n26589 = n26588 ^ n26587 ^ n7410 ;
  assign n26590 = ( n17693 & ~n19142 ) | ( n17693 & n22512 ) | ( ~n19142 & n22512 ) ;
  assign n26591 = n13453 ^ n2745 ^ 1'b0 ;
  assign n26592 = n6722 & ~n26591 ;
  assign n26593 = n26592 ^ n10565 ^ n7404 ;
  assign n26594 = ( n9947 & n26590 ) | ( n9947 & n26593 ) | ( n26590 & n26593 ) ;
  assign n26595 = ( n4068 & n6015 ) | ( n4068 & ~n14966 ) | ( n6015 & ~n14966 ) ;
  assign n26596 = ( n6439 & ~n11019 ) | ( n6439 & n26595 ) | ( ~n11019 & n26595 ) ;
  assign n26597 = n22816 ^ n22204 ^ n18509 ;
  assign n26598 = ( n2262 & n8691 ) | ( n2262 & ~n16321 ) | ( n8691 & ~n16321 ) ;
  assign n26599 = n8193 & n26598 ;
  assign n26600 = n26597 & n26599 ;
  assign n26601 = ~n1456 & n23554 ;
  assign n26602 = ~n11421 & n26601 ;
  assign n26603 = n13750 | n26602 ;
  assign n26604 = n25292 & ~n26603 ;
  assign n26605 = n10493 ^ n3190 ^ n818 ;
  assign n26606 = n4737 & n8613 ;
  assign n26607 = n25138 ^ n24316 ^ n8352 ;
  assign n26608 = n21083 ^ n11219 ^ n3092 ;
  assign n26609 = n15799 ^ n5399 ^ n4468 ;
  assign n26610 = ( n3633 & ~n4560 ) | ( n3633 & n26609 ) | ( ~n4560 & n26609 ) ;
  assign n26611 = ( n8861 & ~n26608 ) | ( n8861 & n26610 ) | ( ~n26608 & n26610 ) ;
  assign n26613 = ( n3017 & n3248 ) | ( n3017 & n6503 ) | ( n3248 & n6503 ) ;
  assign n26612 = n11662 ^ n4231 ^ n2871 ;
  assign n26614 = n26613 ^ n26612 ^ n11115 ;
  assign n26615 = n17888 ^ n4720 ^ 1'b0 ;
  assign n26616 = ~n8445 & n26615 ;
  assign n26617 = n26616 ^ n15780 ^ n3283 ;
  assign n26618 = ( n1142 & n8342 ) | ( n1142 & ~n13495 ) | ( n8342 & ~n13495 ) ;
  assign n26619 = n12353 ^ n11879 ^ 1'b0 ;
  assign n26620 = n1189 | n26619 ;
  assign n26621 = ( n329 & n19700 ) | ( n329 & n26620 ) | ( n19700 & n26620 ) ;
  assign n26622 = ~n26306 & n26621 ;
  assign n26624 = n6527 ^ n2929 ^ n2115 ;
  assign n26623 = n1243 & ~n14076 ;
  assign n26625 = n26624 ^ n26623 ^ 1'b0 ;
  assign n26626 = n26625 ^ n19677 ^ 1'b0 ;
  assign n26627 = ( n5700 & n5828 ) | ( n5700 & n26626 ) | ( n5828 & n26626 ) ;
  assign n26628 = n17231 & ~n22634 ;
  assign n26630 = n18290 ^ n4058 ^ 1'b0 ;
  assign n26631 = n1657 & ~n26630 ;
  assign n26629 = n7044 ^ n4204 ^ 1'b0 ;
  assign n26632 = n26631 ^ n26629 ^ n12011 ;
  assign n26633 = ( ~n5549 & n7873 ) | ( ~n5549 & n22275 ) | ( n7873 & n22275 ) ;
  assign n26634 = ( ~n349 & n424 ) | ( ~n349 & n26633 ) | ( n424 & n26633 ) ;
  assign n26635 = n3526 & ~n21112 ;
  assign n26636 = n26635 ^ n7120 ^ 1'b0 ;
  assign n26637 = n26636 ^ n16180 ^ n11884 ;
  assign n26638 = n2957 & n6914 ;
  assign n26639 = n11364 ^ n8441 ^ n3840 ;
  assign n26640 = n2560 ^ x15 ^ 1'b0 ;
  assign n26641 = n26639 | n26640 ;
  assign n26642 = n16635 ^ n6634 ^ 1'b0 ;
  assign n26643 = n26642 ^ n23478 ^ n3426 ;
  assign n26644 = ( ~n20049 & n23428 ) | ( ~n20049 & n26643 ) | ( n23428 & n26643 ) ;
  assign n26645 = ~n1926 & n14932 ;
  assign n26646 = n248 & n1554 ;
  assign n26647 = ~n18291 & n26646 ;
  assign n26648 = ( n3090 & ~n26645 ) | ( n3090 & n26647 ) | ( ~n26645 & n26647 ) ;
  assign n26649 = n1105 | n25173 ;
  assign n26650 = n1699 | n6192 ;
  assign n26651 = n26650 ^ n20366 ^ 1'b0 ;
  assign n26652 = ( n13577 & n15164 ) | ( n13577 & ~n26651 ) | ( n15164 & ~n26651 ) ;
  assign n26653 = n26652 ^ n16839 ^ 1'b0 ;
  assign n26654 = ( n11671 & n14814 ) | ( n11671 & ~n17944 ) | ( n14814 & ~n17944 ) ;
  assign n26655 = n26654 ^ n15850 ^ 1'b0 ;
  assign n26656 = n26655 ^ n10923 ^ n2813 ;
  assign n26657 = ~n23717 & n26656 ;
  assign n26658 = n14498 ^ n12187 ^ n529 ;
  assign n26659 = ~n20164 & n26658 ;
  assign n26660 = n19437 & n26659 ;
  assign n26661 = x107 & ~n26459 ;
  assign n26662 = ~n18005 & n26661 ;
  assign n26663 = n18346 ^ n9916 ^ n6183 ;
  assign n26664 = n26663 ^ n22588 ^ n19994 ;
  assign n26667 = ( n2029 & ~n2107 ) | ( n2029 & n8383 ) | ( ~n2107 & n8383 ) ;
  assign n26665 = n6124 & n10935 ;
  assign n26666 = n26665 ^ n12274 ^ 1'b0 ;
  assign n26668 = n26667 ^ n26666 ^ n15262 ;
  assign n26669 = n26668 ^ n2858 ^ n1893 ;
  assign n26670 = n23045 ^ n16704 ^ n2683 ;
  assign n26671 = n26670 ^ n25046 ^ n1867 ;
  assign n26672 = n919 & n7117 ;
  assign n26673 = n13615 ^ n9905 ^ n5043 ;
  assign n26674 = n1243 & n10124 ;
  assign n26675 = ~n3149 & n26674 ;
  assign n26676 = ( n3822 & n7101 ) | ( n3822 & n7771 ) | ( n7101 & n7771 ) ;
  assign n26677 = n26676 ^ n12240 ^ 1'b0 ;
  assign n26678 = n18587 ^ n7943 ^ 1'b0 ;
  assign n26679 = n5526 | n26678 ;
  assign n26680 = ( n3144 & n6078 ) | ( n3144 & ~n26679 ) | ( n6078 & ~n26679 ) ;
  assign n26681 = n10658 & ~n26680 ;
  assign n26682 = ( n5551 & n8311 ) | ( n5551 & ~n26681 ) | ( n8311 & ~n26681 ) ;
  assign n26683 = n12058 ^ n5895 ^ n3847 ;
  assign n26684 = n26683 ^ n17720 ^ 1'b0 ;
  assign n26685 = n2749 ^ n1871 ^ n936 ;
  assign n26686 = ( n10655 & n22269 ) | ( n10655 & n26685 ) | ( n22269 & n26685 ) ;
  assign n26687 = n22126 ^ n16212 ^ 1'b0 ;
  assign n26688 = n20683 ^ n4388 ^ n4315 ;
  assign n26689 = ( n12945 & n18669 ) | ( n12945 & n24685 ) | ( n18669 & n24685 ) ;
  assign n26690 = n26689 ^ n16206 ^ n1638 ;
  assign n26691 = ( n26687 & n26688 ) | ( n26687 & ~n26690 ) | ( n26688 & ~n26690 ) ;
  assign n26692 = n22984 ^ n20194 ^ 1'b0 ;
  assign n26693 = n5282 & ~n26692 ;
  assign n26694 = n26693 ^ n6665 ^ n4513 ;
  assign n26695 = n20636 ^ n14894 ^ n7498 ;
  assign n26696 = ~n5508 & n9317 ;
  assign n26697 = n26695 & n26696 ;
  assign n26698 = n19532 ^ n15257 ^ n8791 ;
  assign n26699 = ( ~n5468 & n18031 ) | ( ~n5468 & n23348 ) | ( n18031 & n23348 ) ;
  assign n26700 = ( ~n10250 & n26698 ) | ( ~n10250 & n26699 ) | ( n26698 & n26699 ) ;
  assign n26701 = n20506 ^ n11077 ^ 1'b0 ;
  assign n26702 = n14254 ^ n11342 ^ n4587 ;
  assign n26703 = n18350 ^ n1903 ^ 1'b0 ;
  assign n26704 = n19189 | n26703 ;
  assign n26705 = n8249 ^ n2244 ^ 1'b0 ;
  assign n26706 = n951 | n26705 ;
  assign n26707 = ( ~n18460 & n19999 ) | ( ~n18460 & n26706 ) | ( n19999 & n26706 ) ;
  assign n26711 = n9255 ^ n4252 ^ 1'b0 ;
  assign n26708 = n17389 ^ n1072 ^ n520 ;
  assign n26709 = n15886 & ~n26708 ;
  assign n26710 = n10990 & n26709 ;
  assign n26712 = n26711 ^ n26710 ^ n18468 ;
  assign n26713 = n21745 ^ n17591 ^ n12031 ;
  assign n26714 = n8308 | n26713 ;
  assign n26715 = n26714 ^ n26313 ^ 1'b0 ;
  assign n26716 = n20757 ^ n18854 ^ 1'b0 ;
  assign n26717 = n18270 | n26716 ;
  assign n26718 = n8834 ^ n4925 ^ n2623 ;
  assign n26719 = ( x36 & n9062 ) | ( x36 & ~n11103 ) | ( n9062 & ~n11103 ) ;
  assign n26720 = ( n3863 & ~n26718 ) | ( n3863 & n26719 ) | ( ~n26718 & n26719 ) ;
  assign n26721 = n3867 & n6657 ;
  assign n26722 = ( n1354 & ~n5816 ) | ( n1354 & n26721 ) | ( ~n5816 & n26721 ) ;
  assign n26723 = ( n16790 & ~n18159 ) | ( n16790 & n19455 ) | ( ~n18159 & n19455 ) ;
  assign n26724 = n15026 ^ n11108 ^ n3277 ;
  assign n26725 = ( ~n195 & n3807 ) | ( ~n195 & n26724 ) | ( n3807 & n26724 ) ;
  assign n26729 = n6948 & ~n12605 ;
  assign n26726 = n4680 & n9405 ;
  assign n26727 = n22803 & n26726 ;
  assign n26728 = ( ~n4809 & n8797 ) | ( ~n4809 & n26727 ) | ( n8797 & n26727 ) ;
  assign n26730 = n26729 ^ n26728 ^ n1339 ;
  assign n26731 = n2124 ^ n377 ^ n268 ;
  assign n26732 = ( n6471 & n11565 ) | ( n6471 & ~n12795 ) | ( n11565 & ~n12795 ) ;
  assign n26733 = n26732 ^ n5384 ^ n1691 ;
  assign n26734 = n26733 ^ n1828 ^ n1286 ;
  assign n26735 = ( n11584 & n26731 ) | ( n11584 & ~n26734 ) | ( n26731 & ~n26734 ) ;
  assign n26736 = ( n3010 & ~n3215 ) | ( n3010 & n3726 ) | ( ~n3215 & n3726 ) ;
  assign n26737 = n4855 & ~n26736 ;
  assign n26738 = n7145 ^ n2479 ^ 1'b0 ;
  assign n26739 = n16012 & ~n24139 ;
  assign n26740 = n26739 ^ n1780 ^ 1'b0 ;
  assign n26741 = n18321 & ~n26740 ;
  assign n26742 = n26741 ^ n16195 ^ 1'b0 ;
  assign n26743 = ( n2066 & n3077 ) | ( n2066 & ~n6471 ) | ( n3077 & ~n6471 ) ;
  assign n26744 = ( n8672 & n18921 ) | ( n8672 & ~n26743 ) | ( n18921 & ~n26743 ) ;
  assign n26745 = n16875 ^ n6407 ^ n5546 ;
  assign n26746 = n6478 ^ n4376 ^ 1'b0 ;
  assign n26747 = n1161 & n26746 ;
  assign n26748 = ( n2456 & n2619 ) | ( n2456 & n7769 ) | ( n2619 & n7769 ) ;
  assign n26749 = ( n1119 & ~n26747 ) | ( n1119 & n26748 ) | ( ~n26747 & n26748 ) ;
  assign n26750 = n17913 ^ n4048 ^ 1'b0 ;
  assign n26751 = ~n2639 & n26750 ;
  assign n26752 = n26751 ^ n26025 ^ n7218 ;
  assign n26753 = n9383 ^ n8524 ^ n2918 ;
  assign n26754 = ( ~n6325 & n9106 ) | ( ~n6325 & n26411 ) | ( n9106 & n26411 ) ;
  assign n26755 = ( n9855 & n26753 ) | ( n9855 & ~n26754 ) | ( n26753 & ~n26754 ) ;
  assign n26757 = n3747 & ~n6869 ;
  assign n26758 = n26757 ^ n16100 ^ n3671 ;
  assign n26756 = n10686 ^ n6547 ^ n4997 ;
  assign n26759 = n26758 ^ n26756 ^ n25574 ;
  assign n26760 = ( ~n2202 & n5720 ) | ( ~n2202 & n11894 ) | ( n5720 & n11894 ) ;
  assign n26761 = n13803 | n26760 ;
  assign n26762 = n2846 & ~n26761 ;
  assign n26763 = ( n12593 & ~n20937 ) | ( n12593 & n26762 ) | ( ~n20937 & n26762 ) ;
  assign n26764 = n5627 & n25897 ;
  assign n26765 = ~n20688 & n26764 ;
  assign n26766 = n5154 ^ n2614 ^ n880 ;
  assign n26767 = n22023 ^ n12488 ^ n11232 ;
  assign n26768 = n19408 ^ n18296 ^ n2391 ;
  assign n26769 = n4076 & n4480 ;
  assign n26770 = n26769 ^ n2249 ^ 1'b0 ;
  assign n26771 = ( n2770 & n9648 ) | ( n2770 & n26770 ) | ( n9648 & n26770 ) ;
  assign n26772 = n14834 ^ n10122 ^ 1'b0 ;
  assign n26773 = n5192 & n26772 ;
  assign n26774 = n26773 ^ n25914 ^ n22334 ;
  assign n26775 = n7153 | n9865 ;
  assign n26776 = n26775 ^ n6734 ^ 1'b0 ;
  assign n26777 = ( n10878 & n11022 ) | ( n10878 & ~n26776 ) | ( n11022 & ~n26776 ) ;
  assign n26778 = n26777 ^ n14712 ^ n629 ;
  assign n26779 = ( n17558 & n25525 ) | ( n17558 & n26778 ) | ( n25525 & n26778 ) ;
  assign n26780 = ( n1392 & n2859 ) | ( n1392 & n8308 ) | ( n2859 & n8308 ) ;
  assign n26781 = n4704 & ~n21370 ;
  assign n26782 = ~n18635 & n24450 ;
  assign n26783 = n26782 ^ n25247 ^ 1'b0 ;
  assign n26784 = ( ~n8868 & n26781 ) | ( ~n8868 & n26783 ) | ( n26781 & n26783 ) ;
  assign n26785 = n26784 ^ n25405 ^ n15981 ;
  assign n26786 = n20484 ^ n17670 ^ n4779 ;
  assign n26787 = n26786 ^ n17985 ^ 1'b0 ;
  assign n26788 = n15107 | n26787 ;
  assign n26789 = n1744 & ~n9736 ;
  assign n26790 = n18355 ^ n3111 ^ n599 ;
  assign n26791 = ( n11651 & ~n21464 ) | ( n11651 & n26790 ) | ( ~n21464 & n26790 ) ;
  assign n26792 = n26348 ^ n12723 ^ n10966 ;
  assign n26793 = n26792 ^ n18749 ^ n10769 ;
  assign n26794 = ( n4409 & n5164 ) | ( n4409 & n8779 ) | ( n5164 & n8779 ) ;
  assign n26795 = n10595 ^ n5920 ^ n5250 ;
  assign n26796 = n26795 ^ n6820 ^ 1'b0 ;
  assign n26797 = n4661 ^ n3087 ^ n1523 ;
  assign n26798 = ( n3237 & ~n15675 ) | ( n3237 & n26797 ) | ( ~n15675 & n26797 ) ;
  assign n26799 = n8799 | n26798 ;
  assign n26800 = n26799 ^ n13846 ^ n3953 ;
  assign n26801 = ( n16747 & n20875 ) | ( n16747 & ~n25080 ) | ( n20875 & ~n25080 ) ;
  assign n26804 = ( n3985 & n8078 ) | ( n3985 & ~n22767 ) | ( n8078 & ~n22767 ) ;
  assign n26805 = ( n8898 & n14571 ) | ( n8898 & n26804 ) | ( n14571 & n26804 ) ;
  assign n26802 = ~n7589 & n20288 ;
  assign n26803 = n3696 & n26802 ;
  assign n26806 = n26805 ^ n26803 ^ n25129 ;
  assign n26807 = ( n7392 & n9249 ) | ( n7392 & ~n13327 ) | ( n9249 & ~n13327 ) ;
  assign n26808 = n26807 ^ n20843 ^ n10623 ;
  assign n26809 = n14630 ^ n5065 ^ 1'b0 ;
  assign n26810 = n26808 & ~n26809 ;
  assign n26811 = n6015 | n11034 ;
  assign n26812 = n8368 & ~n26811 ;
  assign n26813 = ~n26207 & n26812 ;
  assign n26814 = n10971 & n19019 ;
  assign n26815 = n26814 ^ n9732 ^ 1'b0 ;
  assign n26816 = n19438 ^ n4685 ^ 1'b0 ;
  assign n26817 = n26815 & n26816 ;
  assign n26818 = ( ~n392 & n2085 ) | ( ~n392 & n5391 ) | ( n2085 & n5391 ) ;
  assign n26819 = n26818 ^ n18636 ^ n15572 ;
  assign n26820 = n2944 ^ n1660 ^ 1'b0 ;
  assign n26821 = n8575 & ~n26820 ;
  assign n26822 = ( ~n15578 & n25355 ) | ( ~n15578 & n26821 ) | ( n25355 & n26821 ) ;
  assign n26823 = n26822 ^ n9666 ^ 1'b0 ;
  assign n26824 = n1621 ^ n1072 ^ n677 ;
  assign n26825 = n26824 ^ n25193 ^ n24912 ;
  assign n26826 = n26825 ^ n15890 ^ n15218 ;
  assign n26827 = n21698 ^ n21453 ^ n338 ;
  assign n26828 = n26827 ^ n6470 ^ 1'b0 ;
  assign n26829 = n4294 | n26828 ;
  assign n26830 = n22770 ^ n18167 ^ 1'b0 ;
  assign n26831 = n26830 ^ n4102 ^ 1'b0 ;
  assign n26832 = ~n26829 & n26831 ;
  assign n26833 = ( ~n14239 & n26535 ) | ( ~n14239 & n26832 ) | ( n26535 & n26832 ) ;
  assign n26834 = n17528 ^ n16098 ^ n15801 ;
  assign n26835 = ( ~n2426 & n4992 ) | ( ~n2426 & n14169 ) | ( n4992 & n14169 ) ;
  assign n26836 = ~n13355 & n26835 ;
  assign n26837 = ~n7814 & n26836 ;
  assign n26838 = n737 | n11528 ;
  assign n26839 = n1046 & ~n5126 ;
  assign n26840 = n26839 ^ n3026 ^ 1'b0 ;
  assign n26841 = n26840 ^ n6987 ^ n5979 ;
  assign n26842 = ( n837 & n1972 ) | ( n837 & n6579 ) | ( n1972 & n6579 ) ;
  assign n26844 = ( ~n386 & n2446 ) | ( ~n386 & n3367 ) | ( n2446 & n3367 ) ;
  assign n26843 = n2069 & ~n13704 ;
  assign n26845 = n26844 ^ n26843 ^ n13373 ;
  assign n26846 = n12119 ^ n4251 ^ 1'b0 ;
  assign n26847 = n22670 ^ n4021 ^ n1159 ;
  assign n26848 = n5147 | n14285 ;
  assign n26849 = n9167 & ~n26848 ;
  assign n26850 = ( n3442 & n26847 ) | ( n3442 & ~n26849 ) | ( n26847 & ~n26849 ) ;
  assign n26851 = ( n1711 & ~n4320 ) | ( n1711 & n11440 ) | ( ~n4320 & n11440 ) ;
  assign n26852 = ( ~n9762 & n10483 ) | ( ~n9762 & n26851 ) | ( n10483 & n26851 ) ;
  assign n26853 = n20167 ^ n5393 ^ 1'b0 ;
  assign n26854 = ~n12245 & n26853 ;
  assign n26855 = ( n436 & ~n6989 ) | ( n436 & n13867 ) | ( ~n6989 & n13867 ) ;
  assign n26856 = n17395 | n26855 ;
  assign n26857 = n26856 ^ n7162 ^ 1'b0 ;
  assign n26858 = n14434 ^ n7856 ^ n5126 ;
  assign n26859 = n26858 ^ n2607 ^ 1'b0 ;
  assign n26860 = ( n4024 & ~n9111 ) | ( n4024 & n11569 ) | ( ~n9111 & n11569 ) ;
  assign n26861 = ( ~n9509 & n23003 ) | ( ~n9509 & n26860 ) | ( n23003 & n26860 ) ;
  assign n26862 = n12168 ^ n2845 ^ 1'b0 ;
  assign n26863 = ( n7241 & n7367 ) | ( n7241 & ~n8234 ) | ( n7367 & ~n8234 ) ;
  assign n26864 = n26863 ^ n11845 ^ n9018 ;
  assign n26865 = n13022 | n26864 ;
  assign n26866 = ( n11661 & n16501 ) | ( n11661 & ~n26865 ) | ( n16501 & ~n26865 ) ;
  assign n26867 = n2561 & n7556 ;
  assign n26868 = ( n3447 & ~n7382 ) | ( n3447 & n26867 ) | ( ~n7382 & n26867 ) ;
  assign n26869 = n18358 ^ n8316 ^ 1'b0 ;
  assign n26870 = ~n8256 & n15980 ;
  assign n26871 = ~n7788 & n26870 ;
  assign n26872 = ( n7671 & n10633 ) | ( n7671 & ~n18002 ) | ( n10633 & ~n18002 ) ;
  assign n26873 = ( n2377 & ~n2970 ) | ( n2377 & n3626 ) | ( ~n2970 & n3626 ) ;
  assign n26874 = n26873 ^ n7405 ^ n5131 ;
  assign n26875 = n26874 ^ n21447 ^ 1'b0 ;
  assign n26876 = n713 & n22892 ;
  assign n26877 = ~n15524 & n26876 ;
  assign n26878 = n26877 ^ n22441 ^ n3878 ;
  assign n26879 = n25029 ^ n7462 ^ n6256 ;
  assign n26880 = n17187 ^ n16358 ^ 1'b0 ;
  assign n26881 = n452 | n4896 ;
  assign n26882 = ( n19995 & n25817 ) | ( n19995 & n26881 ) | ( n25817 & n26881 ) ;
  assign n26883 = n916 | n5428 ;
  assign n26884 = n1971 | n26883 ;
  assign n26885 = ( n13538 & ~n18400 ) | ( n13538 & n20445 ) | ( ~n18400 & n20445 ) ;
  assign n26886 = n26885 ^ n18754 ^ n15368 ;
  assign n26887 = n26886 ^ n21452 ^ 1'b0 ;
  assign n26888 = n9345 & n26887 ;
  assign n26889 = n171 & ~n7075 ;
  assign n26890 = ( n2235 & n5796 ) | ( n2235 & ~n20598 ) | ( n5796 & ~n20598 ) ;
  assign n26891 = ( ~n1158 & n20386 ) | ( ~n1158 & n26890 ) | ( n20386 & n26890 ) ;
  assign n26892 = ( n2368 & n4711 ) | ( n2368 & n6186 ) | ( n4711 & n6186 ) ;
  assign n26893 = n25447 ^ n17818 ^ n8568 ;
  assign n26894 = n9475 ^ n5411 ^ n3542 ;
  assign n26895 = n26894 ^ n10228 ^ 1'b0 ;
  assign n26896 = n12033 | n26895 ;
  assign n26897 = n21142 ^ n19093 ^ n2956 ;
  assign n26898 = n12942 ^ n11158 ^ n1048 ;
  assign n26899 = ( ~n8296 & n9813 ) | ( ~n8296 & n26898 ) | ( n9813 & n26898 ) ;
  assign n26900 = ~n26897 & n26899 ;
  assign n26901 = n26900 ^ n17961 ^ 1'b0 ;
  assign n26902 = n14107 ^ n7117 ^ n5384 ;
  assign n26903 = ( n21563 & n23215 ) | ( n21563 & ~n26902 ) | ( n23215 & ~n26902 ) ;
  assign n26904 = n26903 ^ n13655 ^ n12354 ;
  assign n26905 = n1110 & ~n24342 ;
  assign n26906 = ~n3427 & n26905 ;
  assign n26909 = ( n18617 & n19236 ) | ( n18617 & n26751 ) | ( n19236 & n26751 ) ;
  assign n26907 = ~n3989 & n14591 ;
  assign n26908 = n26907 ^ n1588 ^ 1'b0 ;
  assign n26910 = n26909 ^ n26908 ^ n6712 ;
  assign n26911 = ( n11880 & n26906 ) | ( n11880 & n26910 ) | ( n26906 & n26910 ) ;
  assign n26912 = n4792 ^ n2118 ^ n212 ;
  assign n26913 = ( n14066 & ~n17646 ) | ( n14066 & n26912 ) | ( ~n17646 & n26912 ) ;
  assign n26914 = ( n535 & n18280 ) | ( n535 & ~n26913 ) | ( n18280 & ~n26913 ) ;
  assign n26915 = n26914 ^ n3901 ^ 1'b0 ;
  assign n26916 = n21716 ^ n8850 ^ n1920 ;
  assign n26917 = n19106 & n26916 ;
  assign n26918 = ( ~n8153 & n18075 ) | ( ~n8153 & n26917 ) | ( n18075 & n26917 ) ;
  assign n26919 = n10099 & n17621 ;
  assign n26920 = n23358 ^ n11462 ^ n8074 ;
  assign n26921 = ( n13067 & ~n13359 ) | ( n13067 & n26920 ) | ( ~n13359 & n26920 ) ;
  assign n26922 = ( ~n3754 & n4565 ) | ( ~n3754 & n9232 ) | ( n4565 & n9232 ) ;
  assign n26923 = ( n19665 & n20736 ) | ( n19665 & n26922 ) | ( n20736 & n26922 ) ;
  assign n26924 = ~n12408 & n25550 ;
  assign n26925 = ( n16459 & n26923 ) | ( n16459 & n26924 ) | ( n26923 & n26924 ) ;
  assign n26926 = n22140 ^ n13188 ^ n11715 ;
  assign n26927 = n19311 | n26458 ;
  assign n26928 = n24631 | n26927 ;
  assign n26929 = ( n5231 & n9560 ) | ( n5231 & n19835 ) | ( n9560 & n19835 ) ;
  assign n26930 = n9008 & ~n26929 ;
  assign n26931 = n26930 ^ n6823 ^ n2477 ;
  assign n26932 = ( n14883 & n16154 ) | ( n14883 & n20173 ) | ( n16154 & n20173 ) ;
  assign n26933 = n11416 ^ n11117 ^ n2923 ;
  assign n26934 = ( n564 & n1614 ) | ( n564 & n26933 ) | ( n1614 & n26933 ) ;
  assign n26935 = n10535 ^ n8297 ^ n154 ;
  assign n26938 = ( n4089 & ~n7352 ) | ( n4089 & n12853 ) | ( ~n7352 & n12853 ) ;
  assign n26936 = n7232 & ~n8174 ;
  assign n26937 = n23367 & ~n26936 ;
  assign n26939 = n26938 ^ n26937 ^ n21157 ;
  assign n26940 = ( ~n855 & n13814 ) | ( ~n855 & n20028 ) | ( n13814 & n20028 ) ;
  assign n26941 = ( n3918 & n24965 ) | ( n3918 & n26940 ) | ( n24965 & n26940 ) ;
  assign n26942 = ( n6961 & ~n21675 ) | ( n6961 & n24457 ) | ( ~n21675 & n24457 ) ;
  assign n26943 = n5271 ^ n4900 ^ n435 ;
  assign n26944 = n26943 ^ n6150 ^ 1'b0 ;
  assign n26945 = ~n9991 & n26944 ;
  assign n26946 = n26945 ^ n7442 ^ 1'b0 ;
  assign n26947 = n26946 ^ n23031 ^ n10840 ;
  assign n26948 = n12403 ^ n3158 ^ 1'b0 ;
  assign n26949 = n7821 | n26948 ;
  assign n26950 = n26949 ^ n26108 ^ n22251 ;
  assign n26951 = ( ~n5134 & n11409 ) | ( ~n5134 & n26369 ) | ( n11409 & n26369 ) ;
  assign n26952 = ( ~n16599 & n17142 ) | ( ~n16599 & n18595 ) | ( n17142 & n18595 ) ;
  assign n26953 = n23663 ^ n8731 ^ n4547 ;
  assign n26954 = n4949 | n17238 ;
  assign n26955 = n9854 | n26954 ;
  assign n26956 = n26955 ^ n6361 ^ n1946 ;
  assign n26957 = n659 | n3801 ;
  assign n26958 = n26957 ^ n4742 ^ 1'b0 ;
  assign n26959 = n22005 ^ n17157 ^ n15842 ;
  assign n26960 = n7187 ^ n5520 ^ n1652 ;
  assign n26961 = ( n2797 & n17069 ) | ( n2797 & n17965 ) | ( n17069 & n17965 ) ;
  assign n26962 = ( n1664 & n18324 ) | ( n1664 & ~n26961 ) | ( n18324 & ~n26961 ) ;
  assign n26963 = ~n5667 & n15615 ;
  assign n26964 = ( n17085 & n19298 ) | ( n17085 & ~n26963 ) | ( n19298 & ~n26963 ) ;
  assign n26965 = ( ~x125 & n8742 ) | ( ~x125 & n26964 ) | ( n8742 & n26964 ) ;
  assign n26966 = n8742 ^ n8570 ^ n5498 ;
  assign n26967 = ( n1741 & n5439 ) | ( n1741 & ~n11617 ) | ( n5439 & ~n11617 ) ;
  assign n26968 = ( n352 & n14264 ) | ( n352 & n19243 ) | ( n14264 & n19243 ) ;
  assign n26969 = ( n9887 & n15625 ) | ( n9887 & n26968 ) | ( n15625 & n26968 ) ;
  assign n26970 = ( n7535 & n26967 ) | ( n7535 & ~n26969 ) | ( n26967 & ~n26969 ) ;
  assign n26971 = ( n11491 & n21636 ) | ( n11491 & ~n26970 ) | ( n21636 & ~n26970 ) ;
  assign n26972 = n4975 | n10403 ;
  assign n26973 = n26972 ^ n7086 ^ 1'b0 ;
  assign n26974 = n26973 ^ n25174 ^ n9807 ;
  assign n26975 = n5273 | n16041 ;
  assign n26976 = n26975 ^ n13123 ^ 1'b0 ;
  assign n26977 = n16954 ^ n14422 ^ n3812 ;
  assign n26978 = ( ~n6545 & n14100 ) | ( ~n6545 & n26977 ) | ( n14100 & n26977 ) ;
  assign n26979 = n26978 ^ n11998 ^ 1'b0 ;
  assign n26980 = ~n18152 & n26979 ;
  assign n26981 = ( n10653 & n19178 ) | ( n10653 & ~n22196 ) | ( n19178 & ~n22196 ) ;
  assign n26982 = n24457 ^ n17291 ^ 1'b0 ;
  assign n26983 = n26982 ^ n17591 ^ n4840 ;
  assign n26984 = n5345 & n14332 ;
  assign n26985 = n18296 & n26984 ;
  assign n26986 = n13424 & ~n26985 ;
  assign n26987 = n21784 & n26986 ;
  assign n26988 = n3622 & ~n26987 ;
  assign n26989 = n26988 ^ n21545 ^ n12364 ;
  assign n26990 = ~n10022 & n20729 ;
  assign n26991 = n26990 ^ n3339 ^ 1'b0 ;
  assign n26992 = ( ~n5618 & n17238 ) | ( ~n5618 & n26991 ) | ( n17238 & n26991 ) ;
  assign n26993 = n7953 & ~n11206 ;
  assign n26994 = ~n14114 & n26993 ;
  assign n26995 = x46 & n3422 ;
  assign n26996 = ( ~n25525 & n26994 ) | ( ~n25525 & n26995 ) | ( n26994 & n26995 ) ;
  assign n26997 = n25180 ^ n19199 ^ n8211 ;
  assign n26998 = n26997 ^ n22286 ^ 1'b0 ;
  assign n26999 = n15022 ^ n14097 ^ 1'b0 ;
  assign n27000 = n9077 & ~n26999 ;
  assign n27001 = n6985 ^ n5310 ^ n2480 ;
  assign n27002 = n21261 ^ n16196 ^ 1'b0 ;
  assign n27003 = n27001 & ~n27002 ;
  assign n27004 = n13605 & n27003 ;
  assign n27005 = n27004 ^ n8451 ^ 1'b0 ;
  assign n27006 = ( n10215 & ~n14277 ) | ( n10215 & n20054 ) | ( ~n14277 & n20054 ) ;
  assign n27008 = ( n914 & n2381 ) | ( n914 & n7518 ) | ( n2381 & n7518 ) ;
  assign n27007 = ( ~n1231 & n9125 ) | ( ~n1231 & n15483 ) | ( n9125 & n15483 ) ;
  assign n27009 = n27008 ^ n27007 ^ n26052 ;
  assign n27010 = ( n10192 & n12177 ) | ( n10192 & n17651 ) | ( n12177 & n17651 ) ;
  assign n27011 = ( n12961 & n25890 ) | ( n12961 & ~n27010 ) | ( n25890 & ~n27010 ) ;
  assign n27012 = n2502 & ~n26165 ;
  assign n27013 = ( n7837 & n8155 ) | ( n7837 & n12439 ) | ( n8155 & n12439 ) ;
  assign n27014 = ( n6143 & ~n6412 ) | ( n6143 & n27013 ) | ( ~n6412 & n27013 ) ;
  assign n27015 = n26797 ^ n13216 ^ n6072 ;
  assign n27016 = n747 & n25437 ;
  assign n27017 = n9831 & n27016 ;
  assign n27018 = n8568 ^ n1025 ^ 1'b0 ;
  assign n27019 = ~n3800 & n27018 ;
  assign n27020 = n27019 ^ n26658 ^ 1'b0 ;
  assign n27021 = n6158 ^ n5623 ^ n2033 ;
  assign n27022 = ( n2009 & n12492 ) | ( n2009 & ~n27021 ) | ( n12492 & ~n27021 ) ;
  assign n27027 = n8167 ^ n1903 ^ 1'b0 ;
  assign n27028 = ~n1359 & n27027 ;
  assign n27025 = ( n6939 & ~n7102 ) | ( n6939 & n14332 ) | ( ~n7102 & n14332 ) ;
  assign n27026 = ( n765 & n5207 ) | ( n765 & n27025 ) | ( n5207 & n27025 ) ;
  assign n27023 = n1463 & n5047 ;
  assign n27024 = n4700 & n27023 ;
  assign n27029 = n27028 ^ n27026 ^ n27024 ;
  assign n27030 = n2105 & n15660 ;
  assign n27031 = n5194 ^ n1927 ^ x73 ;
  assign n27032 = ( n3646 & n6465 ) | ( n3646 & n13141 ) | ( n6465 & n13141 ) ;
  assign n27033 = ( n13329 & n17123 ) | ( n13329 & ~n27032 ) | ( n17123 & ~n27032 ) ;
  assign n27034 = ( ~n1994 & n6429 ) | ( ~n1994 & n21031 ) | ( n6429 & n21031 ) ;
  assign n27035 = n10145 & n25773 ;
  assign n27036 = n27035 ^ n7336 ^ 1'b0 ;
  assign n27037 = n6671 & ~n27036 ;
  assign n27038 = ( n430 & ~n5261 ) | ( n430 & n27037 ) | ( ~n5261 & n27037 ) ;
  assign n27039 = ( n1150 & n2868 ) | ( n1150 & ~n20676 ) | ( n2868 & ~n20676 ) ;
  assign n27043 = n8171 ^ n5425 ^ 1'b0 ;
  assign n27040 = ( ~n2395 & n11439 ) | ( ~n2395 & n12466 ) | ( n11439 & n12466 ) ;
  assign n27041 = n27040 ^ n22312 ^ n16107 ;
  assign n27042 = n22913 | n27041 ;
  assign n27044 = n27043 ^ n27042 ^ 1'b0 ;
  assign n27047 = n2602 & n8497 ;
  assign n27048 = ~n21126 & n27047 ;
  assign n27045 = n19656 ^ n17382 ^ n14954 ;
  assign n27046 = n27045 ^ n19870 ^ n15924 ;
  assign n27049 = n27048 ^ n27046 ^ n612 ;
  assign n27050 = n3221 & ~n12805 ;
  assign n27051 = n11928 ^ n2494 ^ 1'b0 ;
  assign n27052 = n6550 | n27051 ;
  assign n27053 = ( n19238 & ~n27050 ) | ( n19238 & n27052 ) | ( ~n27050 & n27052 ) ;
  assign n27054 = n21139 ^ n8076 ^ n727 ;
  assign n27055 = n24408 & n27054 ;
  assign n27056 = n8392 | n27055 ;
  assign n27057 = n27056 ^ n8389 ^ 1'b0 ;
  assign n27058 = ( n1888 & n9131 ) | ( n1888 & ~n27057 ) | ( n9131 & ~n27057 ) ;
  assign n27059 = n12976 ^ n12411 ^ n3277 ;
  assign n27060 = n11150 & ~n13384 ;
  assign n27061 = ~n14731 & n27060 ;
  assign n27062 = ( n21410 & n22490 ) | ( n21410 & n27061 ) | ( n22490 & n27061 ) ;
  assign n27063 = ( n4573 & n7369 ) | ( n4573 & n7788 ) | ( n7369 & n7788 ) ;
  assign n27064 = n27063 ^ n19333 ^ n15144 ;
  assign n27065 = ( n14205 & ~n21227 ) | ( n14205 & n27064 ) | ( ~n21227 & n27064 ) ;
  assign n27066 = ( n15228 & n16443 ) | ( n15228 & n27065 ) | ( n16443 & n27065 ) ;
  assign n27067 = n22648 ^ n21916 ^ n18221 ;
  assign n27068 = ~n1927 & n3648 ;
  assign n27069 = n27068 ^ n8098 ^ 1'b0 ;
  assign n27070 = n13560 ^ n12139 ^ 1'b0 ;
  assign n27071 = ~n12462 & n27070 ;
  assign n27072 = ( ~n2322 & n19258 ) | ( ~n2322 & n27071 ) | ( n19258 & n27071 ) ;
  assign n27073 = ~n1388 & n3101 ;
  assign n27074 = ( ~n1783 & n4104 ) | ( ~n1783 & n27073 ) | ( n4104 & n27073 ) ;
  assign n27075 = ( n15136 & n20838 ) | ( n15136 & n27074 ) | ( n20838 & n27074 ) ;
  assign n27076 = n24288 ^ n17252 ^ n299 ;
  assign n27078 = ( n6475 & n8810 ) | ( n6475 & ~n10404 ) | ( n8810 & ~n10404 ) ;
  assign n27077 = ( n1232 & n5632 ) | ( n1232 & ~n15247 ) | ( n5632 & ~n15247 ) ;
  assign n27079 = n27078 ^ n27077 ^ 1'b0 ;
  assign n27080 = ~n7192 & n27079 ;
  assign n27081 = n27080 ^ n13872 ^ n9032 ;
  assign n27082 = n27081 ^ n16691 ^ n1562 ;
  assign n27083 = n8476 ^ n1213 ^ x17 ;
  assign n27084 = ( n5006 & n9981 ) | ( n5006 & ~n27083 ) | ( n9981 & ~n27083 ) ;
  assign n27086 = ( n3495 & n7959 ) | ( n3495 & ~n20983 ) | ( n7959 & ~n20983 ) ;
  assign n27085 = ~n1084 & n4885 ;
  assign n27087 = n27086 ^ n27085 ^ n7692 ;
  assign n27088 = n23673 ^ n15600 ^ n3224 ;
  assign n27089 = ( ~n16843 & n27087 ) | ( ~n16843 & n27088 ) | ( n27087 & n27088 ) ;
  assign n27090 = ~n2214 & n4674 ;
  assign n27091 = n27090 ^ n13382 ^ n6223 ;
  assign n27094 = n19515 ^ n4536 ^ n423 ;
  assign n27092 = n16330 ^ n2466 ^ n644 ;
  assign n27093 = n5607 & n27092 ;
  assign n27095 = n27094 ^ n27093 ^ 1'b0 ;
  assign n27096 = ( ~n12660 & n22792 ) | ( ~n12660 & n26711 ) | ( n22792 & n26711 ) ;
  assign n27097 = n26790 ^ n6261 ^ 1'b0 ;
  assign n27098 = n13090 ^ n5701 ^ n2698 ;
  assign n27099 = x114 & ~n15159 ;
  assign n27103 = n6895 & ~n8528 ;
  assign n27100 = ( n2123 & n8279 ) | ( n2123 & n12883 ) | ( n8279 & n12883 ) ;
  assign n27101 = n14840 ^ n9086 ^ 1'b0 ;
  assign n27102 = n27100 & ~n27101 ;
  assign n27104 = n27103 ^ n27102 ^ n2856 ;
  assign n27105 = ( n21787 & n27099 ) | ( n21787 & n27104 ) | ( n27099 & n27104 ) ;
  assign n27106 = ( n6655 & n6770 ) | ( n6655 & ~n10888 ) | ( n6770 & ~n10888 ) ;
  assign n27107 = n11182 ^ n3012 ^ 1'b0 ;
  assign n27108 = ( n20963 & n27106 ) | ( n20963 & n27107 ) | ( n27106 & n27107 ) ;
  assign n27109 = ( n14761 & n15751 ) | ( n14761 & n23685 ) | ( n15751 & n23685 ) ;
  assign n27110 = x48 & ~n14438 ;
  assign n27111 = n27110 ^ n16374 ^ 1'b0 ;
  assign n27112 = n201 & n9974 ;
  assign n27113 = n23752 ^ n10008 ^ 1'b0 ;
  assign n27114 = ~n19790 & n25399 ;
  assign n27115 = n22871 ^ n15818 ^ n2351 ;
  assign n27116 = n148 & ~n8122 ;
  assign n27117 = n27116 ^ n9366 ^ 1'b0 ;
  assign n27118 = n7315 & ~n27117 ;
  assign n27119 = n27118 ^ n10189 ^ n1799 ;
  assign n27120 = ( n2082 & n15852 ) | ( n2082 & n25876 ) | ( n15852 & n25876 ) ;
  assign n27121 = ( n3507 & n14026 ) | ( n3507 & ~n19869 ) | ( n14026 & ~n19869 ) ;
  assign n27122 = ( n3103 & ~n25182 ) | ( n3103 & n27121 ) | ( ~n25182 & n27121 ) ;
  assign n27123 = n4216 & ~n13978 ;
  assign n27124 = n27123 ^ n19016 ^ 1'b0 ;
  assign n27125 = ( n3147 & ~n24886 ) | ( n3147 & n27124 ) | ( ~n24886 & n27124 ) ;
  assign n27126 = ~n9800 & n19660 ;
  assign n27127 = n27126 ^ n8821 ^ 1'b0 ;
  assign n27128 = n6679 & n27127 ;
  assign n27129 = n7065 | n27128 ;
  assign n27130 = ~n12077 & n27129 ;
  assign n27131 = n27130 ^ n4425 ^ 1'b0 ;
  assign n27132 = ( n1581 & ~n2008 ) | ( n1581 & n6380 ) | ( ~n2008 & n6380 ) ;
  assign n27133 = n24776 ^ n22196 ^ 1'b0 ;
  assign n27134 = n27132 & ~n27133 ;
  assign n27135 = ( n4373 & ~n5279 ) | ( n4373 & n10210 ) | ( ~n5279 & n10210 ) ;
  assign n27136 = n9618 ^ n5200 ^ n1055 ;
  assign n27137 = n15295 & ~n27136 ;
  assign n27138 = ( n26844 & ~n27135 ) | ( n26844 & n27137 ) | ( ~n27135 & n27137 ) ;
  assign n27139 = n23326 ^ n3350 ^ n1005 ;
  assign n27140 = ( n2049 & ~n2964 ) | ( n2049 & n27139 ) | ( ~n2964 & n27139 ) ;
  assign n27141 = n17943 ^ n8653 ^ n8503 ;
  assign n27142 = n27141 ^ n10441 ^ n6948 ;
  assign n27143 = n24774 ^ n7530 ^ 1'b0 ;
  assign n27144 = ( n7072 & ~n23375 ) | ( n7072 & n27143 ) | ( ~n23375 & n27143 ) ;
  assign n27145 = n26106 ^ n18839 ^ 1'b0 ;
  assign n27146 = n22584 & ~n27145 ;
  assign n27147 = ~n25554 & n27146 ;
  assign n27148 = n26818 & n27147 ;
  assign n27149 = n22628 ^ n3228 ^ 1'b0 ;
  assign n27150 = n21108 & ~n27149 ;
  assign n27151 = n27150 ^ n25966 ^ n13367 ;
  assign n27152 = ( n11604 & n13054 ) | ( n11604 & n22124 ) | ( n13054 & n22124 ) ;
  assign n27153 = n27152 ^ n16979 ^ n7271 ;
  assign n27156 = ( ~n1025 & n8937 ) | ( ~n1025 & n13380 ) | ( n8937 & n13380 ) ;
  assign n27157 = n27156 ^ n3281 ^ n2112 ;
  assign n27154 = ~n7534 & n12911 ;
  assign n27155 = n27154 ^ n17263 ^ 1'b0 ;
  assign n27158 = n27157 ^ n27155 ^ n6260 ;
  assign n27159 = n12023 ^ n8820 ^ n4708 ;
  assign n27160 = n7944 ^ n4880 ^ n4507 ;
  assign n27161 = n27160 ^ n18451 ^ n13317 ;
  assign n27162 = n1731 & ~n15814 ;
  assign n27163 = n27154 ^ n24400 ^ 1'b0 ;
  assign n27164 = n11711 & n21591 ;
  assign n27165 = n27164 ^ n25471 ^ 1'b0 ;
  assign n27166 = ( n1050 & n5162 ) | ( n1050 & ~n26647 ) | ( n5162 & ~n26647 ) ;
  assign n27167 = ( ~n2335 & n4066 ) | ( ~n2335 & n21258 ) | ( n4066 & n21258 ) ;
  assign n27168 = n5284 ^ n4945 ^ 1'b0 ;
  assign n27169 = n14958 ^ n12222 ^ n4076 ;
  assign n27170 = ( ~n27167 & n27168 ) | ( ~n27167 & n27169 ) | ( n27168 & n27169 ) ;
  assign n27173 = ( ~n6443 & n16397 ) | ( ~n6443 & n18672 ) | ( n16397 & n18672 ) ;
  assign n27171 = n18072 ^ n13049 ^ n12318 ;
  assign n27172 = n27171 ^ n13321 ^ n2616 ;
  assign n27174 = n27173 ^ n27172 ^ n7323 ;
  assign n27175 = n18370 ^ n6762 ^ 1'b0 ;
  assign n27176 = ~n4689 & n27175 ;
  assign n27177 = n14770 & n27176 ;
  assign n27178 = ( n2754 & n26262 ) | ( n2754 & n27177 ) | ( n26262 & n27177 ) ;
  assign n27179 = ( n10231 & n14007 ) | ( n10231 & n16849 ) | ( n14007 & n16849 ) ;
  assign n27180 = ( n6441 & n9402 ) | ( n6441 & ~n27179 ) | ( n9402 & ~n27179 ) ;
  assign n27181 = n27160 ^ n10989 ^ n1419 ;
  assign n27182 = n27181 ^ n26899 ^ n8398 ;
  assign n27183 = ( n6983 & n8469 ) | ( n6983 & n23693 ) | ( n8469 & n23693 ) ;
  assign n27184 = n9947 & n16888 ;
  assign n27185 = n9276 ^ n7889 ^ n1282 ;
  assign n27186 = ( n12528 & n16420 ) | ( n12528 & ~n27185 ) | ( n16420 & ~n27185 ) ;
  assign n27191 = ( n2542 & n16123 ) | ( n2542 & n19872 ) | ( n16123 & n19872 ) ;
  assign n27192 = ( n3555 & n15753 ) | ( n3555 & ~n21208 ) | ( n15753 & ~n21208 ) ;
  assign n27193 = ( n2643 & n27191 ) | ( n2643 & n27192 ) | ( n27191 & n27192 ) ;
  assign n27189 = ( n3911 & n8411 ) | ( n3911 & n13171 ) | ( n8411 & n13171 ) ;
  assign n27187 = ~n3246 & n5155 ;
  assign n27188 = ~n24417 & n27187 ;
  assign n27190 = n27189 ^ n27188 ^ n16954 ;
  assign n27194 = n27193 ^ n27190 ^ n2666 ;
  assign n27195 = n7574 | n9496 ;
  assign n27196 = n1287 | n27195 ;
  assign n27197 = n19364 | n27196 ;
  assign n27198 = n10653 ^ n4872 ^ 1'b0 ;
  assign n27199 = n11096 & ~n27198 ;
  assign n27200 = ( n5678 & n23614 ) | ( n5678 & ~n27199 ) | ( n23614 & ~n27199 ) ;
  assign n27201 = ( ~n2979 & n3045 ) | ( ~n2979 & n13795 ) | ( n3045 & n13795 ) ;
  assign n27202 = ( n5632 & n12475 ) | ( n5632 & n27201 ) | ( n12475 & n27201 ) ;
  assign n27203 = ( n14913 & n16656 ) | ( n14913 & n27202 ) | ( n16656 & n27202 ) ;
  assign n27204 = n4502 ^ n1474 ^ 1'b0 ;
  assign n27205 = n27204 ^ n20741 ^ 1'b0 ;
  assign n27206 = n9503 & n27205 ;
  assign n27207 = ~n917 & n27206 ;
  assign n27208 = n27207 ^ n3236 ^ 1'b0 ;
  assign n27209 = n14680 ^ n5200 ^ 1'b0 ;
  assign n27210 = ( n707 & n12277 ) | ( n707 & ~n15578 ) | ( n12277 & ~n15578 ) ;
  assign n27211 = ( n691 & ~n1022 ) | ( n691 & n3120 ) | ( ~n1022 & n3120 ) ;
  assign n27212 = n15301 ^ n10472 ^ n3995 ;
  assign n27213 = n26511 ^ n20066 ^ 1'b0 ;
  assign n27214 = n20351 & ~n27213 ;
  assign n27215 = ( n16538 & n27212 ) | ( n16538 & n27214 ) | ( n27212 & n27214 ) ;
  assign n27220 = ( ~n3802 & n5494 ) | ( ~n3802 & n8026 ) | ( n5494 & n8026 ) ;
  assign n27221 = ( n14192 & n22512 ) | ( n14192 & n27220 ) | ( n22512 & n27220 ) ;
  assign n27216 = n9235 ^ n516 ^ 1'b0 ;
  assign n27217 = ( n6616 & ~n8319 ) | ( n6616 & n12554 ) | ( ~n8319 & n12554 ) ;
  assign n27218 = n5164 & n27217 ;
  assign n27219 = ~n27216 & n27218 ;
  assign n27222 = n27221 ^ n27219 ^ n6323 ;
  assign n27223 = ( n386 & n3205 ) | ( n386 & n3331 ) | ( n3205 & n3331 ) ;
  assign n27224 = n27223 ^ n23529 ^ n17995 ;
  assign n27227 = n10193 ^ n1193 ^ 1'b0 ;
  assign n27228 = ~n10646 & n27227 ;
  assign n27225 = n8804 ^ n6877 ^ n2566 ;
  assign n27226 = ( n17911 & n20260 ) | ( n17911 & ~n27225 ) | ( n20260 & ~n27225 ) ;
  assign n27229 = n27228 ^ n27226 ^ n16076 ;
  assign n27230 = n22039 ^ n770 ^ 1'b0 ;
  assign n27231 = n20475 | n27230 ;
  assign n27232 = n15650 ^ n7021 ^ 1'b0 ;
  assign n27233 = n4708 & n27232 ;
  assign n27234 = n10190 ^ n6459 ^ n2455 ;
  assign n27235 = ( n9546 & n16499 ) | ( n9546 & n27234 ) | ( n16499 & n27234 ) ;
  assign n27236 = n27235 ^ n25427 ^ n243 ;
  assign n27237 = n25604 ^ n7124 ^ n6949 ;
  assign n27238 = ( n390 & ~n6006 ) | ( n390 & n27237 ) | ( ~n6006 & n27237 ) ;
  assign n27239 = ( n9306 & n11893 ) | ( n9306 & ~n23665 ) | ( n11893 & ~n23665 ) ;
  assign n27240 = n27239 ^ n25122 ^ n2723 ;
  assign n27241 = ( n3460 & n13044 ) | ( n3460 & n17524 ) | ( n13044 & n17524 ) ;
  assign n27242 = n25137 ^ n13209 ^ n9957 ;
  assign n27243 = n17759 ^ n15639 ^ n12894 ;
  assign n27244 = n296 & ~n3251 ;
  assign n27245 = ( n6851 & n8188 ) | ( n6851 & n17244 ) | ( n8188 & n17244 ) ;
  assign n27246 = n143 | n27245 ;
  assign n27247 = n27244 & ~n27246 ;
  assign n27248 = n20416 ^ n20224 ^ n2342 ;
  assign n27249 = ( x70 & n656 ) | ( x70 & n8856 ) | ( n656 & n8856 ) ;
  assign n27250 = n26985 ^ n12947 ^ n10197 ;
  assign n27251 = ( n7072 & n17574 ) | ( n7072 & n27250 ) | ( n17574 & n27250 ) ;
  assign n27252 = ~n10149 & n11770 ;
  assign n27253 = n8541 | n15286 ;
  assign n27254 = ( n10664 & ~n14406 ) | ( n10664 & n27253 ) | ( ~n14406 & n27253 ) ;
  assign n27255 = ( n6265 & ~n10927 ) | ( n6265 & n12359 ) | ( ~n10927 & n12359 ) ;
  assign n27256 = n27255 ^ n26111 ^ n7842 ;
  assign n27257 = ( n729 & ~n1825 ) | ( n729 & n5583 ) | ( ~n1825 & n5583 ) ;
  assign n27258 = ( n6822 & ~n17491 ) | ( n6822 & n27257 ) | ( ~n17491 & n27257 ) ;
  assign n27259 = n27258 ^ n16877 ^ 1'b0 ;
  assign n27260 = n18252 & ~n27259 ;
  assign n27261 = n19790 ^ n16139 ^ n2337 ;
  assign n27262 = n12199 | n27261 ;
  assign n27263 = ~n7053 & n11671 ;
  assign n27264 = ( n1926 & n14680 ) | ( n1926 & n27263 ) | ( n14680 & n27263 ) ;
  assign n27265 = n26100 ^ n15213 ^ n616 ;
  assign n27266 = n7261 & ~n11963 ;
  assign n27267 = n27266 ^ n25960 ^ n14492 ;
  assign n27268 = n25559 ^ n15825 ^ n1010 ;
  assign n27269 = n27268 ^ n23493 ^ n9917 ;
  assign n27270 = ( n4587 & n9010 ) | ( n4587 & ~n10333 ) | ( n9010 & ~n10333 ) ;
  assign n27271 = n4532 ^ n4075 ^ n2008 ;
  assign n27272 = n27271 ^ n5042 ^ n3233 ;
  assign n27280 = n22182 ^ n4150 ^ n2387 ;
  assign n27273 = ( ~n563 & n5551 ) | ( ~n563 & n20615 ) | ( n5551 & n20615 ) ;
  assign n27274 = ( n3972 & n14459 ) | ( n3972 & ~n27273 ) | ( n14459 & ~n27273 ) ;
  assign n27275 = n15997 & ~n27274 ;
  assign n27276 = n23317 & ~n27275 ;
  assign n27277 = ~n9528 & n27276 ;
  assign n27278 = n27277 ^ n17928 ^ n8127 ;
  assign n27279 = n21304 | n27278 ;
  assign n27281 = n27280 ^ n27279 ^ n3017 ;
  assign n27284 = ( ~n925 & n20509 ) | ( ~n925 & n22909 ) | ( n20509 & n22909 ) ;
  assign n27285 = ( ~n16979 & n19466 ) | ( ~n16979 & n27284 ) | ( n19466 & n27284 ) ;
  assign n27282 = ( n4166 & n12372 ) | ( n4166 & ~n22029 ) | ( n12372 & ~n22029 ) ;
  assign n27283 = n1104 & ~n27282 ;
  assign n27286 = n27285 ^ n27283 ^ 1'b0 ;
  assign n27287 = n16039 ^ n13981 ^ 1'b0 ;
  assign n27288 = n24316 ^ n20113 ^ n1876 ;
  assign n27289 = ( n6754 & ~n7103 ) | ( n6754 & n12031 ) | ( ~n7103 & n12031 ) ;
  assign n27290 = n3227 | n11775 ;
  assign n27291 = n9219 & ~n27290 ;
  assign n27292 = n27291 ^ n3059 ^ n1009 ;
  assign n27293 = n12998 | n27292 ;
  assign n27294 = n19926 | n27293 ;
  assign n27295 = n27263 | n27294 ;
  assign n27296 = n14644 ^ n14302 ^ n6499 ;
  assign n27297 = ( n20284 & n22290 ) | ( n20284 & ~n27296 ) | ( n22290 & ~n27296 ) ;
  assign n27298 = ( n8511 & n13596 ) | ( n8511 & n20361 ) | ( n13596 & n20361 ) ;
  assign n27299 = n21372 ^ n1797 ^ 1'b0 ;
  assign n27300 = n5486 & ~n27299 ;
  assign n27301 = n426 & ~n1244 ;
  assign n27302 = ( n3901 & n4793 ) | ( n3901 & ~n10066 ) | ( n4793 & ~n10066 ) ;
  assign n27303 = n27302 ^ n25458 ^ 1'b0 ;
  assign n27304 = ( ~n962 & n10001 ) | ( ~n962 & n10864 ) | ( n10001 & n10864 ) ;
  assign n27305 = ( n11760 & ~n13468 ) | ( n11760 & n14006 ) | ( ~n13468 & n14006 ) ;
  assign n27306 = ( n3001 & ~n20994 ) | ( n3001 & n27305 ) | ( ~n20994 & n27305 ) ;
  assign n27307 = ( ~n670 & n4478 ) | ( ~n670 & n6535 ) | ( n4478 & n6535 ) ;
  assign n27308 = n27307 ^ n22200 ^ n4866 ;
  assign n27309 = ( n7369 & n23458 ) | ( n7369 & ~n27308 ) | ( n23458 & ~n27308 ) ;
  assign n27310 = n16560 ^ n6340 ^ 1'b0 ;
  assign n27314 = ( n11441 & n17408 ) | ( n11441 & n19587 ) | ( n17408 & n19587 ) ;
  assign n27311 = n6628 | n17508 ;
  assign n27312 = n27311 ^ n8722 ^ n3339 ;
  assign n27313 = ~n6745 & n27312 ;
  assign n27315 = n27314 ^ n27313 ^ n14677 ;
  assign n27316 = n15226 ^ n8594 ^ n2926 ;
  assign n27317 = n25025 ^ n3372 ^ n3279 ;
  assign n27318 = ( n4696 & ~n6728 ) | ( n4696 & n27317 ) | ( ~n6728 & n27317 ) ;
  assign n27319 = n2769 | n27318 ;
  assign n27320 = n6565 ^ n6008 ^ 1'b0 ;
  assign n27322 = n7414 ^ n5630 ^ n3728 ;
  assign n27321 = n14144 ^ n11429 ^ n4489 ;
  assign n27323 = n27322 ^ n27321 ^ n11936 ;
  assign n27324 = ~n6469 & n18112 ;
  assign n27325 = ~n27323 & n27324 ;
  assign n27326 = n14414 ^ n4666 ^ n1232 ;
  assign n27327 = n15651 ^ n14913 ^ n8983 ;
  assign n27328 = ( n8165 & n27326 ) | ( n8165 & ~n27327 ) | ( n27326 & ~n27327 ) ;
  assign n27332 = ( n2544 & n11594 ) | ( n2544 & ~n13415 ) | ( n11594 & ~n13415 ) ;
  assign n27333 = ( n265 & n2182 ) | ( n265 & ~n27332 ) | ( n2182 & ~n27332 ) ;
  assign n27334 = n27333 ^ n17153 ^ 1'b0 ;
  assign n27329 = n10464 ^ n6901 ^ 1'b0 ;
  assign n27330 = n17537 | n27329 ;
  assign n27331 = n27330 ^ n16804 ^ n7083 ;
  assign n27335 = n27334 ^ n27331 ^ n10572 ;
  assign n27336 = ~n8826 & n13741 ;
  assign n27337 = ~n4154 & n27336 ;
  assign n27338 = ( n22085 & ~n24069 ) | ( n22085 & n27337 ) | ( ~n24069 & n27337 ) ;
  assign n27339 = ( n1655 & n14805 ) | ( n1655 & n23891 ) | ( n14805 & n23891 ) ;
  assign n27340 = ( ~n2860 & n11985 ) | ( ~n2860 & n20630 ) | ( n11985 & n20630 ) ;
  assign n27341 = ( n1210 & ~n14010 ) | ( n1210 & n20419 ) | ( ~n14010 & n20419 ) ;
  assign n27342 = n27341 ^ n3923 ^ 1'b0 ;
  assign n27343 = n2402 & n27342 ;
  assign n27344 = ( ~n5858 & n20690 ) | ( ~n5858 & n27343 ) | ( n20690 & n27343 ) ;
  assign n27345 = ( n1014 & ~n2186 ) | ( n1014 & n15818 ) | ( ~n2186 & n15818 ) ;
  assign n27346 = n27345 ^ n13017 ^ n9268 ;
  assign n27347 = ( ~n9080 & n18682 ) | ( ~n9080 & n19018 ) | ( n18682 & n19018 ) ;
  assign n27348 = n10512 ^ n9067 ^ n1305 ;
  assign n27349 = n27348 ^ n3613 ^ 1'b0 ;
  assign n27350 = n27347 & n27349 ;
  assign n27351 = ~n7007 & n15653 ;
  assign n27352 = n27351 ^ n19010 ^ 1'b0 ;
  assign n27353 = n7102 & n13365 ;
  assign n27354 = n27353 ^ n6270 ^ 1'b0 ;
  assign n27355 = n22056 ^ n11394 ^ n8192 ;
  assign n27356 = n27355 ^ n2322 ^ 1'b0 ;
  assign n27357 = n27354 | n27356 ;
  assign n27358 = n20610 ^ n15065 ^ n14913 ;
  assign n27359 = n6285 ^ n2872 ^ 1'b0 ;
  assign n27360 = n2882 | n27359 ;
  assign n27361 = n27360 ^ n19109 ^ n1417 ;
  assign n27362 = n27361 ^ n11925 ^ n10869 ;
  assign n27369 = ( n805 & n8457 ) | ( n805 & n13040 ) | ( n8457 & n13040 ) ;
  assign n27370 = n27369 ^ n23124 ^ n15860 ;
  assign n27371 = ( n11136 & ~n23109 ) | ( n11136 & n27370 ) | ( ~n23109 & n27370 ) ;
  assign n27367 = ( n489 & n4403 ) | ( n489 & ~n11301 ) | ( n4403 & ~n11301 ) ;
  assign n27368 = ( n6297 & n21470 ) | ( n6297 & ~n27367 ) | ( n21470 & ~n27367 ) ;
  assign n27363 = n8947 ^ n5658 ^ 1'b0 ;
  assign n27364 = x27 & n27363 ;
  assign n27365 = ( n8854 & n9454 ) | ( n8854 & n13754 ) | ( n9454 & n13754 ) ;
  assign n27366 = n27364 & ~n27365 ;
  assign n27372 = n27371 ^ n27368 ^ n27366 ;
  assign n27373 = n12705 ^ n11538 ^ n1777 ;
  assign n27374 = ( n11006 & n15507 ) | ( n11006 & n27373 ) | ( n15507 & n27373 ) ;
  assign n27375 = n27374 ^ n23939 ^ n2569 ;
  assign n27376 = n24539 ^ n943 ^ n868 ;
  assign n27377 = ( n22758 & ~n27375 ) | ( n22758 & n27376 ) | ( ~n27375 & n27376 ) ;
  assign n27378 = n3375 | n5968 ;
  assign n27379 = n27378 ^ n9893 ^ 1'b0 ;
  assign n27380 = n27379 ^ n7825 ^ 1'b0 ;
  assign n27381 = n2962 & ~n27380 ;
  assign n27382 = ( n422 & n2803 ) | ( n422 & ~n16363 ) | ( n2803 & ~n16363 ) ;
  assign n27383 = n27382 ^ n3238 ^ n3023 ;
  assign n27384 = ( n2138 & ~n27381 ) | ( n2138 & n27383 ) | ( ~n27381 & n27383 ) ;
  assign n27385 = n10572 | n22344 ;
  assign n27386 = ~n19403 & n24699 ;
  assign n27387 = n20131 ^ n7487 ^ 1'b0 ;
  assign n27388 = n27386 & n27387 ;
  assign n27389 = n12312 ^ n6338 ^ n6319 ;
  assign n27390 = n20070 & ~n24711 ;
  assign n27391 = n27390 ^ n1425 ^ 1'b0 ;
  assign n27392 = n27391 ^ n26735 ^ 1'b0 ;
  assign n27393 = n27389 & n27392 ;
  assign n27394 = n13147 ^ n11307 ^ n3221 ;
  assign n27395 = n18495 ^ n5331 ^ 1'b0 ;
  assign n27396 = ( ~n5161 & n10079 ) | ( ~n5161 & n14808 ) | ( n10079 & n14808 ) ;
  assign n27397 = n6999 ^ n851 ^ 1'b0 ;
  assign n27398 = ( n2904 & n6369 ) | ( n2904 & n27397 ) | ( n6369 & n27397 ) ;
  assign n27399 = n18058 ^ n7850 ^ n5828 ;
  assign n27400 = n2589 & n3345 ;
  assign n27401 = n8028 ^ n4558 ^ 1'b0 ;
  assign n27402 = n27400 & n27401 ;
  assign n27403 = ~n7125 & n9065 ;
  assign n27404 = ~n27402 & n27403 ;
  assign n27405 = n4593 ^ n2210 ^ n331 ;
  assign n27406 = n4989 ^ n4822 ^ 1'b0 ;
  assign n27407 = ~n27405 & n27406 ;
  assign n27408 = n23288 ^ n22007 ^ 1'b0 ;
  assign n27409 = ~n3989 & n10109 ;
  assign n27410 = ( n3024 & n26753 ) | ( n3024 & n27409 ) | ( n26753 & n27409 ) ;
  assign n27411 = ( ~n4321 & n5367 ) | ( ~n4321 & n13131 ) | ( n5367 & n13131 ) ;
  assign n27412 = ( ~n4191 & n4525 ) | ( ~n4191 & n5431 ) | ( n4525 & n5431 ) ;
  assign n27413 = n27412 ^ n18897 ^ 1'b0 ;
  assign n27414 = ( n7592 & n10010 ) | ( n7592 & n27413 ) | ( n10010 & n27413 ) ;
  assign n27415 = n7443 | n10013 ;
  assign n27416 = n5257 ^ n4217 ^ n450 ;
  assign n27417 = ( n1445 & ~n18526 ) | ( n1445 & n27416 ) | ( ~n18526 & n27416 ) ;
  assign n27418 = n2594 & n27417 ;
  assign n27419 = n27418 ^ n14911 ^ 1'b0 ;
  assign n27420 = n27419 ^ n13445 ^ n7959 ;
  assign n27421 = ( ~n5979 & n8155 ) | ( ~n5979 & n11751 ) | ( n8155 & n11751 ) ;
  assign n27422 = n27421 ^ n15756 ^ n8310 ;
  assign n27423 = n27422 ^ n7125 ^ n6772 ;
  assign n27424 = n25160 ^ n1985 ^ 1'b0 ;
  assign n27425 = n1159 & n27424 ;
  assign n27426 = ( n495 & ~n4300 ) | ( n495 & n15614 ) | ( ~n4300 & n15614 ) ;
  assign n27427 = n8719 & ~n27426 ;
  assign n27428 = n27427 ^ n12795 ^ 1'b0 ;
  assign n27429 = n8302 ^ n3844 ^ 1'b0 ;
  assign n27430 = n27429 ^ n17886 ^ 1'b0 ;
  assign n27432 = ( n164 & n1065 ) | ( n164 & ~n7258 ) | ( n1065 & ~n7258 ) ;
  assign n27431 = ( ~n3243 & n22036 ) | ( ~n3243 & n26912 ) | ( n22036 & n26912 ) ;
  assign n27433 = n27432 ^ n27431 ^ n25061 ;
  assign n27434 = n21746 ^ n7883 ^ n3254 ;
  assign n27435 = ( n14761 & n17074 ) | ( n14761 & ~n27434 ) | ( n17074 & ~n27434 ) ;
  assign n27436 = n6967 ^ n6175 ^ x34 ;
  assign n27437 = ( ~n9652 & n21412 ) | ( ~n9652 & n27436 ) | ( n21412 & n27436 ) ;
  assign n27438 = ( n5873 & n9122 ) | ( n5873 & n14421 ) | ( n9122 & n14421 ) ;
  assign n27439 = x60 | n27438 ;
  assign n27441 = n21114 ^ n1983 ^ 1'b0 ;
  assign n27440 = ( n5825 & ~n19818 ) | ( n5825 & n24107 ) | ( ~n19818 & n24107 ) ;
  assign n27442 = n27441 ^ n27440 ^ n10934 ;
  assign n27443 = n27442 ^ n6314 ^ n4310 ;
  assign n27444 = ( ~n3304 & n16135 ) | ( ~n3304 & n21327 ) | ( n16135 & n21327 ) ;
  assign n27445 = n7465 & n12668 ;
  assign n27446 = n27444 & n27445 ;
  assign n27451 = n8825 & n9840 ;
  assign n27448 = n2789 & n7575 ;
  assign n27449 = ~n9531 & n27448 ;
  assign n27447 = n21396 ^ n20177 ^ n5674 ;
  assign n27450 = n27449 ^ n27447 ^ n2885 ;
  assign n27452 = n27451 ^ n27450 ^ n3976 ;
  assign n27453 = n27452 ^ n23770 ^ n5381 ;
  assign n27454 = ( ~n26105 & n27446 ) | ( ~n26105 & n27453 ) | ( n27446 & n27453 ) ;
  assign n27455 = n7897 ^ n6553 ^ n2840 ;
  assign n27456 = ( ~n1495 & n8006 ) | ( ~n1495 & n27455 ) | ( n8006 & n27455 ) ;
  assign n27457 = n5912 & ~n13433 ;
  assign n27458 = ( n5645 & n16158 ) | ( n5645 & ~n19986 ) | ( n16158 & ~n19986 ) ;
  assign n27459 = n5959 ^ n5896 ^ 1'b0 ;
  assign n27460 = n1104 & n27459 ;
  assign n27461 = ~n2502 & n27460 ;
  assign n27462 = n27461 ^ n25727 ^ 1'b0 ;
  assign n27463 = ( ~n488 & n26290 ) | ( ~n488 & n27462 ) | ( n26290 & n27462 ) ;
  assign n27464 = ~n2379 & n27463 ;
  assign n27465 = ( n2254 & ~n19842 ) | ( n2254 & n22489 ) | ( ~n19842 & n22489 ) ;
  assign n27466 = ( n2925 & ~n18737 ) | ( n2925 & n27465 ) | ( ~n18737 & n27465 ) ;
  assign n27467 = ( ~n27458 & n27464 ) | ( ~n27458 & n27466 ) | ( n27464 & n27466 ) ;
  assign n27468 = ( n3142 & ~n13713 ) | ( n3142 & n16803 ) | ( ~n13713 & n16803 ) ;
  assign n27469 = n27468 ^ n13187 ^ n6315 ;
  assign n27470 = ( x9 & n1150 ) | ( x9 & ~n21410 ) | ( n1150 & ~n21410 ) ;
  assign n27471 = ~n7295 & n8407 ;
  assign n27472 = n9027 ^ n2360 ^ 1'b0 ;
  assign n27473 = ~n3463 & n27472 ;
  assign n27474 = ~n12364 & n27248 ;
  assign n27475 = n27474 ^ n23231 ^ 1'b0 ;
  assign n27477 = ( ~n2542 & n17263 ) | ( ~n2542 & n24960 ) | ( n17263 & n24960 ) ;
  assign n27476 = n4167 & ~n25683 ;
  assign n27478 = n27477 ^ n27476 ^ n24583 ;
  assign n27479 = n27478 ^ n21770 ^ n3081 ;
  assign n27480 = n7187 ^ n1781 ^ 1'b0 ;
  assign n27481 = ( n4697 & ~n13232 ) | ( n4697 & n27480 ) | ( ~n13232 & n27480 ) ;
  assign n27485 = n14395 ^ n6337 ^ n3593 ;
  assign n27483 = ( n759 & n3161 ) | ( n759 & ~n15756 ) | ( n3161 & ~n15756 ) ;
  assign n27482 = ~n3634 & n12752 ;
  assign n27484 = n27483 ^ n27482 ^ 1'b0 ;
  assign n27486 = n27485 ^ n27484 ^ n25251 ;
  assign n27487 = n1649 & n2211 ;
  assign n27488 = ~n4752 & n27487 ;
  assign n27489 = n23291 ^ n14593 ^ n6928 ;
  assign n27490 = n27489 ^ n15042 ^ n13033 ;
  assign n27491 = n2295 ^ n1484 ^ 1'b0 ;
  assign n27492 = ( ~n9125 & n15140 ) | ( ~n9125 & n27491 ) | ( n15140 & n27491 ) ;
  assign n27493 = n9271 ^ n9186 ^ 1'b0 ;
  assign n27494 = n27492 & ~n27493 ;
  assign n27495 = ( ~n10062 & n26469 ) | ( ~n10062 & n27494 ) | ( n26469 & n27494 ) ;
  assign n27496 = ( n14201 & ~n27490 ) | ( n14201 & n27495 ) | ( ~n27490 & n27495 ) ;
  assign n27497 = ( n17131 & n27488 ) | ( n17131 & ~n27496 ) | ( n27488 & ~n27496 ) ;
  assign n27498 = n4372 ^ n2257 ^ n1410 ;
  assign n27499 = n27498 ^ n15843 ^ n2262 ;
  assign n27502 = n12856 ^ n4756 ^ n2499 ;
  assign n27500 = ( n6108 & ~n10109 ) | ( n6108 & n14913 ) | ( ~n10109 & n14913 ) ;
  assign n27501 = n27500 ^ n23896 ^ n740 ;
  assign n27503 = n27502 ^ n27501 ^ n11682 ;
  assign n27504 = n3999 & n9430 ;
  assign n27505 = n27504 ^ n3993 ^ 1'b0 ;
  assign n27506 = n27505 ^ n21282 ^ n7688 ;
  assign n27508 = n13511 ^ n4698 ^ n4610 ;
  assign n27507 = ( n3936 & n7042 ) | ( n3936 & n24386 ) | ( n7042 & n24386 ) ;
  assign n27509 = n27508 ^ n27507 ^ 1'b0 ;
  assign n27510 = ~n26143 & n27509 ;
  assign n27511 = ( ~x51 & n10399 ) | ( ~x51 & n17417 ) | ( n10399 & n17417 ) ;
  assign n27512 = n13435 ^ n4143 ^ 1'b0 ;
  assign n27513 = n27511 & ~n27512 ;
  assign n27514 = ( n6681 & n14591 ) | ( n6681 & n18833 ) | ( n14591 & n18833 ) ;
  assign n27515 = n4580 ^ n3891 ^ x61 ;
  assign n27516 = n17311 | n27515 ;
  assign n27517 = n1071 | n25756 ;
  assign n27518 = x94 & ~n27517 ;
  assign n27519 = n3986 | n8375 ;
  assign n27520 = n1949 & ~n27519 ;
  assign n27521 = n2753 & n8309 ;
  assign n27522 = n8844 & n27521 ;
  assign n27523 = ( n1104 & n13628 ) | ( n1104 & n27522 ) | ( n13628 & n27522 ) ;
  assign n27524 = ( n12148 & n27520 ) | ( n12148 & n27523 ) | ( n27520 & n27523 ) ;
  assign n27525 = ( ~n4915 & n9026 ) | ( ~n4915 & n15805 ) | ( n9026 & n15805 ) ;
  assign n27526 = ( ~n762 & n3033 ) | ( ~n762 & n23308 ) | ( n3033 & n23308 ) ;
  assign n27527 = n6127 & n18749 ;
  assign n27528 = ~n23345 & n27527 ;
  assign n27529 = ~n2343 & n6593 ;
  assign n27530 = n3192 & n24107 ;
  assign n27531 = n27529 & n27530 ;
  assign n27532 = n21628 ^ n21626 ^ 1'b0 ;
  assign n27533 = n3270 | n27532 ;
  assign n27534 = n6655 ^ n3697 ^ n1269 ;
  assign n27535 = ~n16082 & n27534 ;
  assign n27536 = ~n10342 & n27535 ;
  assign n27537 = n27536 ^ n11606 ^ n1242 ;
  assign n27538 = ~n13089 & n27537 ;
  assign n27539 = ( n356 & ~n26045 ) | ( n356 & n27538 ) | ( ~n26045 & n27538 ) ;
  assign n27541 = n14965 ^ n1765 ^ 1'b0 ;
  assign n27542 = ( n5581 & n20166 ) | ( n5581 & ~n27541 ) | ( n20166 & ~n27541 ) ;
  assign n27540 = n6590 ^ n2673 ^ n613 ;
  assign n27543 = n27542 ^ n27540 ^ 1'b0 ;
  assign n27544 = ( n8592 & ~n10372 ) | ( n8592 & n20585 ) | ( ~n10372 & n20585 ) ;
  assign n27545 = n20034 ^ n14589 ^ n2268 ;
  assign n27546 = n3913 | n16281 ;
  assign n27547 = n27546 ^ n13424 ^ 1'b0 ;
  assign n27548 = ( n1275 & ~n3633 ) | ( n1275 & n19972 ) | ( ~n3633 & n19972 ) ;
  assign n27549 = ( n6350 & n27547 ) | ( n6350 & ~n27548 ) | ( n27547 & ~n27548 ) ;
  assign n27550 = n19901 ^ n16870 ^ n5643 ;
  assign n27551 = ( n204 & n19034 ) | ( n204 & n22668 ) | ( n19034 & n22668 ) ;
  assign n27552 = n13639 | n27551 ;
  assign n27553 = n10105 & ~n27552 ;
  assign n27554 = n21177 ^ n2625 ^ 1'b0 ;
  assign n27555 = n7094 | n27554 ;
  assign n27556 = n20014 & ~n27555 ;
  assign n27557 = n178 | n3557 ;
  assign n27558 = n27557 ^ n1564 ^ 1'b0 ;
  assign n27559 = n5052 | n15954 ;
  assign n27560 = n27559 ^ n783 ^ 1'b0 ;
  assign n27561 = n27560 ^ n11803 ^ n3192 ;
  assign n27562 = n15905 ^ n14964 ^ 1'b0 ;
  assign n27563 = n9579 ^ n3543 ^ 1'b0 ;
  assign n27564 = n24889 ^ n21535 ^ 1'b0 ;
  assign n27565 = ( n24437 & n27563 ) | ( n24437 & ~n27564 ) | ( n27563 & ~n27564 ) ;
  assign n27566 = n27565 ^ n26924 ^ n23986 ;
  assign n27567 = ( ~n3933 & n9302 ) | ( ~n3933 & n24583 ) | ( n9302 & n24583 ) ;
  assign n27568 = ( n7096 & n8976 ) | ( n7096 & ~n27567 ) | ( n8976 & ~n27567 ) ;
  assign n27569 = n27568 ^ n18352 ^ n2501 ;
  assign n27570 = n22476 ^ n7692 ^ n889 ;
  assign n27571 = n6868 & n18853 ;
  assign n27572 = n21403 & n27571 ;
  assign n27573 = n16327 ^ n16096 ^ 1'b0 ;
  assign n27574 = n20362 ^ n17309 ^ 1'b0 ;
  assign n27575 = n2576 & ~n27574 ;
  assign n27576 = n14087 ^ n11439 ^ n5211 ;
  assign n27582 = n15609 ^ n5984 ^ n1087 ;
  assign n27581 = n23535 ^ n2269 ^ n149 ;
  assign n27577 = n6464 ^ n6393 ^ n2377 ;
  assign n27578 = ( n8184 & n17677 ) | ( n8184 & n27577 ) | ( n17677 & n27577 ) ;
  assign n27579 = ~n14516 & n27578 ;
  assign n27580 = n22510 & n27579 ;
  assign n27583 = n27582 ^ n27581 ^ n27580 ;
  assign n27584 = ( ~n2459 & n4652 ) | ( ~n2459 & n25966 ) | ( n4652 & n25966 ) ;
  assign n27585 = ( n9119 & n10057 ) | ( n9119 & ~n14019 ) | ( n10057 & ~n14019 ) ;
  assign n27586 = ( n7668 & ~n17047 ) | ( n7668 & n27585 ) | ( ~n17047 & n27585 ) ;
  assign n27587 = ( n4677 & ~n21853 ) | ( n4677 & n25484 ) | ( ~n21853 & n25484 ) ;
  assign n27588 = n18390 ^ n16988 ^ n2690 ;
  assign n27590 = n12768 | n22437 ;
  assign n27591 = n27590 ^ n5856 ^ 1'b0 ;
  assign n27592 = n27591 ^ n23470 ^ n7936 ;
  assign n27589 = ( ~n989 & n10703 ) | ( ~n989 & n11077 ) | ( n10703 & n11077 ) ;
  assign n27593 = n27592 ^ n27589 ^ n25713 ;
  assign n27594 = ~n191 & n6839 ;
  assign n27595 = ~n7939 & n27594 ;
  assign n27596 = n10698 | n27595 ;
  assign n27597 = n13150 & ~n27596 ;
  assign n27598 = ( ~n14022 & n21408 ) | ( ~n14022 & n21560 ) | ( n21408 & n21560 ) ;
  assign n27599 = ( n6987 & n13704 ) | ( n6987 & ~n20473 ) | ( n13704 & ~n20473 ) ;
  assign n27600 = ( n359 & n19962 ) | ( n359 & ~n27599 ) | ( n19962 & ~n27599 ) ;
  assign n27601 = n14719 & ~n23840 ;
  assign n27602 = n27601 ^ n17577 ^ 1'b0 ;
  assign n27603 = n27602 ^ n13435 ^ n3445 ;
  assign n27604 = n6652 ^ n1275 ^ 1'b0 ;
  assign n27605 = n4364 & n27604 ;
  assign n27606 = ( ~n276 & n4556 ) | ( ~n276 & n27605 ) | ( n4556 & n27605 ) ;
  assign n27607 = ( n780 & n16196 ) | ( n780 & ~n19195 ) | ( n16196 & ~n19195 ) ;
  assign n27608 = n20711 ^ n14906 ^ n12470 ;
  assign n27609 = n27608 ^ n16459 ^ n5581 ;
  assign n27610 = n20579 ^ n17199 ^ 1'b0 ;
  assign n27611 = ~n15385 & n27610 ;
  assign n27612 = n27611 ^ n12217 ^ n2122 ;
  assign n27613 = n8345 ^ n2761 ^ n312 ;
  assign n27614 = ( ~n141 & n10195 ) | ( ~n141 & n27613 ) | ( n10195 & n27613 ) ;
  assign n27615 = n27614 ^ n22694 ^ x105 ;
  assign n27616 = n27615 ^ n11022 ^ n7776 ;
  assign n27617 = n27616 ^ n14884 ^ n299 ;
  assign n27618 = n15157 & ~n18202 ;
  assign n27619 = ~n22609 & n27618 ;
  assign n27620 = n762 & n4055 ;
  assign n27621 = n2417 & n27620 ;
  assign n27622 = n27621 ^ n15952 ^ 1'b0 ;
  assign n27623 = n21708 & n27622 ;
  assign n27624 = n19866 & ~n20511 ;
  assign n27625 = n27624 ^ n9728 ^ 1'b0 ;
  assign n27626 = ( n17764 & n22976 ) | ( n17764 & n27625 ) | ( n22976 & n27625 ) ;
  assign n27627 = n19162 ^ n17061 ^ n212 ;
  assign n27628 = n27627 ^ n18399 ^ n1257 ;
  assign n27629 = ( n1645 & n18050 ) | ( n1645 & n27628 ) | ( n18050 & n27628 ) ;
  assign n27630 = n645 & n2272 ;
  assign n27631 = n5458 | n27630 ;
  assign n27632 = n27631 ^ n20692 ^ n875 ;
  assign n27633 = ( n1091 & ~n1272 ) | ( n1091 & n27050 ) | ( ~n1272 & n27050 ) ;
  assign n27634 = n27633 ^ n21940 ^ n17108 ;
  assign n27635 = ( ~n3621 & n7077 ) | ( ~n3621 & n11005 ) | ( n7077 & n11005 ) ;
  assign n27636 = n5218 | n27635 ;
  assign n27637 = n23719 ^ n20481 ^ n5586 ;
  assign n27638 = n15818 | n18020 ;
  assign n27639 = ( n2773 & n2842 ) | ( n2773 & n6215 ) | ( n2842 & n6215 ) ;
  assign n27640 = ( n7693 & n14414 ) | ( n7693 & ~n27639 ) | ( n14414 & ~n27639 ) ;
  assign n27641 = n2972 & n23928 ;
  assign n27642 = n27640 & n27641 ;
  assign n27644 = n9568 ^ n5373 ^ 1'b0 ;
  assign n27645 = n963 & ~n27644 ;
  assign n27643 = ( n208 & n1770 ) | ( n208 & ~n21880 ) | ( n1770 & ~n21880 ) ;
  assign n27646 = n27645 ^ n27643 ^ n14875 ;
  assign n27647 = ( n18561 & n20991 ) | ( n18561 & ~n25756 ) | ( n20991 & ~n25756 ) ;
  assign n27652 = ~n5841 & n6863 ;
  assign n27653 = n20082 & n27652 ;
  assign n27648 = n678 & ~n14126 ;
  assign n27649 = n27648 ^ n1031 ^ 1'b0 ;
  assign n27650 = ( n5319 & ~n13199 ) | ( n5319 & n27649 ) | ( ~n13199 & n27649 ) ;
  assign n27651 = n2517 & n27650 ;
  assign n27654 = n27653 ^ n27651 ^ 1'b0 ;
  assign n27655 = ( n5167 & ~n27647 ) | ( n5167 & n27654 ) | ( ~n27647 & n27654 ) ;
  assign n27656 = n27655 ^ n1380 ^ 1'b0 ;
  assign n27657 = n27656 ^ n15616 ^ n14645 ;
  assign n27658 = n27135 ^ n5914 ^ 1'b0 ;
  assign n27659 = ~n133 & n8491 ;
  assign n27660 = ( n6343 & n27658 ) | ( n6343 & n27659 ) | ( n27658 & n27659 ) ;
  assign n27661 = n5108 ^ n5045 ^ 1'b0 ;
  assign n27662 = n24310 & n27661 ;
  assign n27663 = n27662 ^ n20372 ^ n7230 ;
  assign n27664 = n15517 ^ n5350 ^ n5030 ;
  assign n27665 = ( n4997 & n12524 ) | ( n4997 & n27664 ) | ( n12524 & n27664 ) ;
  assign n27666 = n3959 & ~n12290 ;
  assign n27667 = n27666 ^ n1735 ^ 1'b0 ;
  assign n27668 = n11745 & n14392 ;
  assign n27669 = n27667 & n27668 ;
  assign n27670 = ( n9043 & n16079 ) | ( n9043 & n27669 ) | ( n16079 & n27669 ) ;
  assign n27671 = n21114 ^ n16991 ^ 1'b0 ;
  assign n27672 = n19683 | n27671 ;
  assign n27673 = n2209 & n27672 ;
  assign n27674 = ( n10706 & n18934 ) | ( n10706 & n20179 ) | ( n18934 & n20179 ) ;
  assign n27675 = ( ~n7744 & n22111 ) | ( ~n7744 & n27674 ) | ( n22111 & n27674 ) ;
  assign n27676 = n18490 ^ n15582 ^ n3986 ;
  assign n27677 = n27676 ^ n15882 ^ n9725 ;
  assign n27678 = ( ~n2203 & n9258 ) | ( ~n2203 & n16507 ) | ( n9258 & n16507 ) ;
  assign n27679 = n21625 ^ n2799 ^ 1'b0 ;
  assign n27680 = n27679 ^ n15897 ^ n8547 ;
  assign n27681 = n26873 ^ n12679 ^ n4782 ;
  assign n27682 = ( ~n20380 & n26186 ) | ( ~n20380 & n27681 ) | ( n26186 & n27681 ) ;
  assign n27683 = ( n6637 & n7506 ) | ( n6637 & ~n9349 ) | ( n7506 & ~n9349 ) ;
  assign n27684 = n4448 & ~n27683 ;
  assign n27685 = n27684 ^ n13950 ^ 1'b0 ;
  assign n27686 = n21208 ^ n4890 ^ n4831 ;
  assign n27687 = ( n8950 & ~n27685 ) | ( n8950 & n27686 ) | ( ~n27685 & n27686 ) ;
  assign n27688 = n13943 ^ n6338 ^ n865 ;
  assign n27691 = ( n5340 & ~n5994 ) | ( n5340 & n23057 ) | ( ~n5994 & n23057 ) ;
  assign n27689 = ~n9506 & n11746 ;
  assign n27690 = n27689 ^ n25617 ^ n1998 ;
  assign n27692 = n27691 ^ n27690 ^ 1'b0 ;
  assign n27693 = n873 & n2948 ;
  assign n27694 = n27693 ^ n10198 ^ 1'b0 ;
  assign n27695 = ~n1592 & n23595 ;
  assign n27696 = n17828 ^ n8701 ^ 1'b0 ;
  assign n27697 = n20419 ^ n17219 ^ n2064 ;
  assign n27698 = n19903 ^ n10900 ^ n7918 ;
  assign n27699 = n4890 ^ n1285 ^ 1'b0 ;
  assign n27700 = ~n347 & n27699 ;
  assign n27701 = n27700 ^ n20625 ^ n13371 ;
  assign n27702 = n23447 ^ n4269 ^ 1'b0 ;
  assign n27703 = n4731 | n27702 ;
  assign n27704 = n27703 ^ n21895 ^ n8589 ;
  assign n27705 = n6351 & ~n23921 ;
  assign n27706 = ( n2212 & n4574 ) | ( n2212 & ~n27705 ) | ( n4574 & ~n27705 ) ;
  assign n27707 = n27706 ^ n16917 ^ n464 ;
  assign n27708 = n7386 ^ n5411 ^ 1'b0 ;
  assign n27709 = n15792 | n27708 ;
  assign n27710 = ( n2445 & n12740 ) | ( n2445 & ~n27709 ) | ( n12740 & ~n27709 ) ;
  assign n27711 = n4070 & ~n17224 ;
  assign n27712 = n27711 ^ n24697 ^ 1'b0 ;
  assign n27713 = ( ~n3924 & n20557 ) | ( ~n3924 & n27712 ) | ( n20557 & n27712 ) ;
  assign n27714 = n10457 | n18708 ;
  assign n27715 = n27713 & ~n27714 ;
  assign n27716 = ( n6755 & ~n7531 ) | ( n6755 & n9092 ) | ( ~n7531 & n9092 ) ;
  assign n27717 = ( n149 & n12208 ) | ( n149 & n27716 ) | ( n12208 & n27716 ) ;
  assign n27718 = n27717 ^ n12588 ^ 1'b0 ;
  assign n27719 = ~n27715 & n27718 ;
  assign n27720 = n13351 & ~n15316 ;
  assign n27721 = ~n26973 & n27720 ;
  assign n27722 = n27721 ^ n7976 ^ 1'b0 ;
  assign n27723 = n20015 ^ n4767 ^ 1'b0 ;
  assign n27724 = ( ~n3350 & n8762 ) | ( ~n3350 & n10012 ) | ( n8762 & n10012 ) ;
  assign n27725 = ( ~n14869 & n14880 ) | ( ~n14869 & n27724 ) | ( n14880 & n27724 ) ;
  assign n27726 = n26040 ^ n18236 ^ n9127 ;
  assign n27727 = n12337 ^ n8823 ^ n7021 ;
  assign n27728 = ( n1227 & n6180 ) | ( n1227 & ~n21453 ) | ( n6180 & ~n21453 ) ;
  assign n27729 = n27728 ^ n10618 ^ n1825 ;
  assign n27730 = n14957 ^ n12063 ^ n7469 ;
  assign n27731 = ( ~n11958 & n27729 ) | ( ~n11958 & n27730 ) | ( n27729 & n27730 ) ;
  assign n27732 = n20325 ^ n3841 ^ 1'b0 ;
  assign n27733 = n13025 ^ n1675 ^ 1'b0 ;
  assign n27734 = ~n19985 & n27733 ;
  assign n27735 = ( n4691 & ~n12640 ) | ( n4691 & n27734 ) | ( ~n12640 & n27734 ) ;
  assign n27736 = ( ~n22871 & n27732 ) | ( ~n22871 & n27735 ) | ( n27732 & n27735 ) ;
  assign n27737 = n2909 ^ n582 ^ 1'b0 ;
  assign n27738 = ~n27522 & n27737 ;
  assign n27739 = n27738 ^ n5869 ^ n5749 ;
  assign n27740 = n22923 ^ n19407 ^ n18529 ;
  assign n27741 = ( n9722 & n12106 ) | ( n9722 & ~n21096 ) | ( n12106 & ~n21096 ) ;
  assign n27742 = n7442 | n10845 ;
  assign n27743 = n19984 | n27742 ;
  assign n27744 = ( n27268 & n27741 ) | ( n27268 & n27743 ) | ( n27741 & n27743 ) ;
  assign n27745 = n7055 & n26257 ;
  assign n27746 = ~n27744 & n27745 ;
  assign n27747 = ( n2011 & ~n5600 ) | ( n2011 & n15481 ) | ( ~n5600 & n15481 ) ;
  assign n27748 = n4765 ^ n2236 ^ 1'b0 ;
  assign n27749 = ~n27747 & n27748 ;
  assign n27750 = ( n9139 & n18997 ) | ( n9139 & ~n26016 ) | ( n18997 & ~n26016 ) ;
  assign n27751 = ( n8467 & n13790 ) | ( n8467 & ~n20965 ) | ( n13790 & ~n20965 ) ;
  assign n27752 = n10106 ^ n9088 ^ n3845 ;
  assign n27753 = ( n15846 & ~n17423 ) | ( n15846 & n20105 ) | ( ~n17423 & n20105 ) ;
  assign n27754 = n22557 ^ n1228 ^ 1'b0 ;
  assign n27755 = n3805 & n27754 ;
  assign n27756 = ( ~n6367 & n11881 ) | ( ~n6367 & n27755 ) | ( n11881 & n27755 ) ;
  assign n27757 = n5836 | n27756 ;
  assign n27758 = ~n27753 & n27757 ;
  assign n27759 = n10833 ^ n7614 ^ 1'b0 ;
  assign n27760 = n26138 & n27759 ;
  assign n27761 = ( ~n4232 & n9537 ) | ( ~n4232 & n27760 ) | ( n9537 & n27760 ) ;
  assign n27764 = ( n1781 & ~n4508 ) | ( n1781 & n8431 ) | ( ~n4508 & n8431 ) ;
  assign n27765 = ( ~n15446 & n19311 ) | ( ~n15446 & n27764 ) | ( n19311 & n27764 ) ;
  assign n27762 = n4334 & ~n19717 ;
  assign n27763 = ~n26835 & n27762 ;
  assign n27766 = n27765 ^ n27763 ^ n19319 ;
  assign n27767 = n2815 ^ n1726 ^ 1'b0 ;
  assign n27768 = ( ~n1401 & n26075 ) | ( ~n1401 & n27767 ) | ( n26075 & n27767 ) ;
  assign n27769 = n27768 ^ n8068 ^ 1'b0 ;
  assign n27770 = n27766 | n27769 ;
  assign n27771 = n7493 ^ n6114 ^ n527 ;
  assign n27772 = n7089 & n27771 ;
  assign n27773 = n19142 ^ n13995 ^ 1'b0 ;
  assign n27774 = n1282 & n27773 ;
  assign n27775 = ~n1825 & n15764 ;
  assign n27776 = n21542 | n27775 ;
  assign n27777 = ( n5375 & n10250 ) | ( n5375 & n27776 ) | ( n10250 & n27776 ) ;
  assign n27778 = n17616 ^ n17405 ^ n16478 ;
  assign n27779 = ( ~n393 & n4559 ) | ( ~n393 & n22770 ) | ( n4559 & n22770 ) ;
  assign n27780 = n27779 ^ n11883 ^ n3186 ;
  assign n27781 = n1342 & ~n1451 ;
  assign n27782 = n20153 & n27781 ;
  assign n27783 = n817 ^ n516 ^ 1'b0 ;
  assign n27784 = n4962 & n27783 ;
  assign n27785 = n27784 ^ n25808 ^ n8072 ;
  assign n27786 = ( n27221 & n27782 ) | ( n27221 & n27785 ) | ( n27782 & n27785 ) ;
  assign n27787 = ( ~n2711 & n6169 ) | ( ~n2711 & n23896 ) | ( n6169 & n23896 ) ;
  assign n27788 = ( n5246 & n7323 ) | ( n5246 & ~n7469 ) | ( n7323 & ~n7469 ) ;
  assign n27789 = ( ~n16057 & n27787 ) | ( ~n16057 & n27788 ) | ( n27787 & n27788 ) ;
  assign n27790 = n10899 ^ n6149 ^ n2742 ;
  assign n27791 = ( n4374 & n9154 ) | ( n4374 & ~n13875 ) | ( n9154 & ~n13875 ) ;
  assign n27792 = ( n4114 & n7863 ) | ( n4114 & n27791 ) | ( n7863 & n27791 ) ;
  assign n27793 = ( n16754 & n27790 ) | ( n16754 & n27792 ) | ( n27790 & n27792 ) ;
  assign n27794 = n1615 & n13103 ;
  assign n27795 = n27794 ^ n25933 ^ 1'b0 ;
  assign n27796 = ( n19719 & n23489 ) | ( n19719 & n27795 ) | ( n23489 & n27795 ) ;
  assign n27797 = ~n611 & n21214 ;
  assign n27798 = n27797 ^ n20897 ^ 1'b0 ;
  assign n27799 = n14411 ^ n7206 ^ 1'b0 ;
  assign n27800 = n12120 & n27799 ;
  assign n27801 = ( ~n6391 & n18448 ) | ( ~n6391 & n20192 ) | ( n18448 & n20192 ) ;
  assign n27802 = ( ~n4965 & n10952 ) | ( ~n4965 & n13504 ) | ( n10952 & n13504 ) ;
  assign n27803 = ( ~n6370 & n16896 ) | ( ~n6370 & n27802 ) | ( n16896 & n27802 ) ;
  assign n27804 = n26460 ^ n7832 ^ n2060 ;
  assign n27805 = n356 & ~n5382 ;
  assign n27806 = ~n4090 & n27805 ;
  assign n27807 = n27806 ^ n20446 ^ n7829 ;
  assign n27808 = n24999 ^ n16660 ^ n9328 ;
  assign n27809 = n27808 ^ n22674 ^ n19853 ;
  assign n27810 = n4896 ^ n1051 ^ 1'b0 ;
  assign n27811 = ( n457 & ~n11762 ) | ( n457 & n27810 ) | ( ~n11762 & n27810 ) ;
  assign n27812 = ( n16420 & n17448 ) | ( n16420 & ~n27811 ) | ( n17448 & ~n27811 ) ;
  assign n27813 = ( ~n4024 & n7439 ) | ( ~n4024 & n22659 ) | ( n7439 & n22659 ) ;
  assign n27814 = ( n7932 & n20285 ) | ( n7932 & n27813 ) | ( n20285 & n27813 ) ;
  assign n27821 = n12846 ^ n9445 ^ n2596 ;
  assign n27822 = n27821 ^ n9526 ^ n3241 ;
  assign n27820 = ~n12334 & n24712 ;
  assign n27823 = n27822 ^ n27820 ^ n6169 ;
  assign n27815 = n11394 ^ n209 ^ x19 ;
  assign n27816 = n27815 ^ n17515 ^ n15175 ;
  assign n27817 = n16942 ^ n11290 ^ n1957 ;
  assign n27818 = n27817 ^ n26390 ^ n18864 ;
  assign n27819 = ( n4339 & n27816 ) | ( n4339 & ~n27818 ) | ( n27816 & ~n27818 ) ;
  assign n27824 = n27823 ^ n27819 ^ n6525 ;
  assign n27825 = n18323 ^ n11472 ^ 1'b0 ;
  assign n27826 = ~n8484 & n27825 ;
  assign n27827 = n23967 ^ n14386 ^ 1'b0 ;
  assign n27828 = n22790 & n27827 ;
  assign n27832 = n13212 ^ n13031 ^ n10062 ;
  assign n27829 = n2084 ^ n1215 ^ 1'b0 ;
  assign n27830 = n24871 ^ n10554 ^ n4165 ;
  assign n27831 = ( n6480 & ~n27829 ) | ( n6480 & n27830 ) | ( ~n27829 & n27830 ) ;
  assign n27833 = n27832 ^ n27831 ^ n9861 ;
  assign n27834 = n12331 ^ n969 ^ 1'b0 ;
  assign n27836 = ( n3257 & n8249 ) | ( n3257 & n12945 ) | ( n8249 & n12945 ) ;
  assign n27835 = n4874 | n6204 ;
  assign n27837 = n27836 ^ n27835 ^ 1'b0 ;
  assign n27838 = n27837 ^ n26109 ^ n7969 ;
  assign n27839 = n18045 ^ n11428 ^ 1'b0 ;
  assign n27840 = n9225 ^ n7063 ^ 1'b0 ;
  assign n27841 = n3594 & ~n27840 ;
  assign n27842 = n27841 ^ n2254 ^ 1'b0 ;
  assign n27843 = ( n10162 & n26683 ) | ( n10162 & ~n27842 ) | ( n26683 & ~n27842 ) ;
  assign n27844 = n10372 & ~n14609 ;
  assign n27845 = ~n1030 & n27844 ;
  assign n27846 = ( ~n4864 & n17082 ) | ( ~n4864 & n25246 ) | ( n17082 & n25246 ) ;
  assign n27847 = n8305 ^ n3909 ^ n2874 ;
  assign n27848 = ~n208 & n9439 ;
  assign n27849 = n4890 & n27848 ;
  assign n27850 = n27849 ^ n577 ^ 1'b0 ;
  assign n27851 = n6981 & n7670 ;
  assign n27852 = n13618 ^ n12687 ^ n4579 ;
  assign n27853 = ( ~n3291 & n13519 ) | ( ~n3291 & n27852 ) | ( n13519 & n27852 ) ;
  assign n27854 = n9328 ^ n6021 ^ 1'b0 ;
  assign n27855 = ( n2191 & ~n5350 ) | ( n2191 & n15691 ) | ( ~n5350 & n15691 ) ;
  assign n27857 = n22439 ^ n3954 ^ 1'b0 ;
  assign n27858 = ( ~n14235 & n22137 ) | ( ~n14235 & n27857 ) | ( n22137 & n27857 ) ;
  assign n27856 = n19642 | n20551 ;
  assign n27859 = n27858 ^ n27856 ^ 1'b0 ;
  assign n27860 = ( n6065 & n7675 ) | ( n6065 & n19001 ) | ( n7675 & n19001 ) ;
  assign n27861 = ( n16134 & n26748 ) | ( n16134 & n27860 ) | ( n26748 & n27860 ) ;
  assign n27862 = n27861 ^ n22151 ^ n19657 ;
  assign n27863 = ( n260 & n298 ) | ( n260 & ~n740 ) | ( n298 & ~n740 ) ;
  assign n27864 = n27863 ^ n5291 ^ n449 ;
  assign n27865 = n26475 ^ n7957 ^ 1'b0 ;
  assign n27866 = n1762 & n27865 ;
  assign n27867 = ~n23994 & n27866 ;
  assign n27868 = ~n598 & n18976 ;
  assign n27869 = ~n12255 & n27868 ;
  assign n27870 = n27869 ^ n25019 ^ n8008 ;
  assign n27871 = n18715 ^ n8799 ^ n4703 ;
  assign n27872 = n22122 ^ n7029 ^ n3464 ;
  assign n27873 = ( ~n3360 & n21960 ) | ( ~n3360 & n22997 ) | ( n21960 & n22997 ) ;
  assign n27874 = ( n5051 & n6554 ) | ( n5051 & ~n6986 ) | ( n6554 & ~n6986 ) ;
  assign n27875 = n6972 & n13755 ;
  assign n27876 = n27874 & n27875 ;
  assign n27877 = n11398 ^ n3052 ^ 1'b0 ;
  assign n27878 = n20712 & ~n27877 ;
  assign n27879 = n2764 & n25763 ;
  assign n27880 = n16200 ^ n1435 ^ 1'b0 ;
  assign n27881 = n1826 & n27880 ;
  assign n27882 = ( n10235 & ~n27879 ) | ( n10235 & n27881 ) | ( ~n27879 & n27881 ) ;
  assign n27883 = ( n7894 & n15269 ) | ( n7894 & ~n18048 ) | ( n15269 & ~n18048 ) ;
  assign n27884 = n15067 ^ n14254 ^ n4216 ;
  assign n27885 = n27884 ^ n20420 ^ 1'b0 ;
  assign n27886 = ~n27883 & n27885 ;
  assign n27887 = ( n19325 & n20189 ) | ( n19325 & n27886 ) | ( n20189 & n27886 ) ;
  assign n27888 = n23891 ^ n16715 ^ n196 ;
  assign n27889 = n7451 ^ n4076 ^ 1'b0 ;
  assign n27890 = ( n4299 & n10307 ) | ( n4299 & n27889 ) | ( n10307 & n27889 ) ;
  assign n27891 = ( n16842 & ~n17772 ) | ( n16842 & n26244 ) | ( ~n17772 & n26244 ) ;
  assign n27892 = n17474 ^ n16449 ^ 1'b0 ;
  assign n27893 = ~n177 & n6075 ;
  assign n27894 = n27893 ^ n16017 ^ 1'b0 ;
  assign n27895 = n27894 ^ n18293 ^ n14539 ;
  assign n27896 = n5474 ^ n319 ^ 1'b0 ;
  assign n27897 = n27895 & n27896 ;
  assign n27898 = ( n8791 & ~n27892 ) | ( n8791 & n27897 ) | ( ~n27892 & n27897 ) ;
  assign n27899 = ( n5453 & ~n6567 ) | ( n5453 & n13763 ) | ( ~n6567 & n13763 ) ;
  assign n27900 = n4669 & ~n4956 ;
  assign n27901 = n27900 ^ n12022 ^ n7242 ;
  assign n27902 = n27901 ^ n19916 ^ n4835 ;
  assign n27903 = ( ~n19074 & n19800 ) | ( ~n19074 & n23648 ) | ( n19800 & n23648 ) ;
  assign n27904 = ~n22548 & n27903 ;
  assign n27905 = n27904 ^ n17733 ^ 1'b0 ;
  assign n27906 = n2874 | n5828 ;
  assign n27907 = n27906 ^ n22121 ^ 1'b0 ;
  assign n27908 = ( ~n8926 & n16906 ) | ( ~n8926 & n26258 ) | ( n16906 & n26258 ) ;
  assign n27909 = n2447 & ~n19084 ;
  assign n27910 = n5380 & n27909 ;
  assign n27911 = n27910 ^ n12007 ^ n1938 ;
  assign n27912 = n8568 ^ n2686 ^ n828 ;
  assign n27913 = n27912 ^ n22839 ^ n1976 ;
  assign n27914 = ( n8435 & ~n18390 ) | ( n8435 & n27913 ) | ( ~n18390 & n27913 ) ;
  assign n27915 = ( n12782 & ~n20365 ) | ( n12782 & n26017 ) | ( ~n20365 & n26017 ) ;
  assign n27916 = ( n140 & ~n5695 ) | ( n140 & n11826 ) | ( ~n5695 & n11826 ) ;
  assign n27917 = n27916 ^ n13573 ^ n5049 ;
  assign n27918 = n20322 ^ n18637 ^ n3241 ;
  assign n27919 = ( ~n4371 & n16672 ) | ( ~n4371 & n19736 ) | ( n16672 & n19736 ) ;
  assign n27920 = ( n7588 & n8879 ) | ( n7588 & n10981 ) | ( n8879 & n10981 ) ;
  assign n27921 = n27920 ^ n25437 ^ 1'b0 ;
  assign n27922 = n27919 & n27921 ;
  assign n27923 = n13897 ^ n1166 ^ 1'b0 ;
  assign n27924 = n21003 ^ n18892 ^ 1'b0 ;
  assign n27925 = n23330 & n27924 ;
  assign n27926 = ( n18203 & n20456 ) | ( n18203 & n27925 ) | ( n20456 & n27925 ) ;
  assign n27927 = n14565 ^ n8510 ^ n1237 ;
  assign n27928 = n11951 | n14166 ;
  assign n27929 = ( n9939 & n27927 ) | ( n9939 & n27928 ) | ( n27927 & n27928 ) ;
  assign n27930 = n4543 & ~n14264 ;
  assign n27931 = n27930 ^ n7281 ^ 1'b0 ;
  assign n27932 = ( n8418 & n23485 ) | ( n8418 & n27931 ) | ( n23485 & n27931 ) ;
  assign n27933 = ( n2841 & n16595 ) | ( n2841 & ~n21433 ) | ( n16595 & ~n21433 ) ;
  assign n27934 = n26525 ^ n25247 ^ 1'b0 ;
  assign n27935 = n4506 & n18194 ;
  assign n27936 = n22948 ^ n3588 ^ 1'b0 ;
  assign n27937 = n15892 | n27936 ;
  assign n27938 = n4511 ^ n4386 ^ 1'b0 ;
  assign n27939 = n27938 ^ n13775 ^ n5965 ;
  assign n27940 = n26000 ^ n9503 ^ n3108 ;
  assign n27941 = ( n3820 & n9151 ) | ( n3820 & n14859 ) | ( n9151 & n14859 ) ;
  assign n27942 = ~n4214 & n22971 ;
  assign n27943 = ~n25011 & n27942 ;
  assign n27944 = ( ~n4473 & n27941 ) | ( ~n4473 & n27943 ) | ( n27941 & n27943 ) ;
  assign n27945 = ( n5229 & n5706 ) | ( n5229 & ~n14891 ) | ( n5706 & ~n14891 ) ;
  assign n27946 = n4167 ^ n1066 ^ 1'b0 ;
  assign n27947 = ~n309 & n27946 ;
  assign n27948 = n27947 ^ n10643 ^ n236 ;
  assign n27949 = ( n5870 & ~n22347 ) | ( n5870 & n27948 ) | ( ~n22347 & n27948 ) ;
  assign n27950 = n5040 ^ n3140 ^ 1'b0 ;
  assign n27951 = n21745 & ~n27950 ;
  assign n27952 = ( n20930 & ~n27819 ) | ( n20930 & n27951 ) | ( ~n27819 & n27951 ) ;
  assign n27953 = n16088 | n18177 ;
  assign n27954 = n14784 & ~n27953 ;
  assign n27955 = n18698 ^ n12827 ^ n5732 ;
  assign n27956 = n8929 ^ n8300 ^ 1'b0 ;
  assign n27957 = ~n27955 & n27956 ;
  assign n27958 = n7531 ^ n4213 ^ n1328 ;
  assign n27959 = n16446 & ~n27958 ;
  assign n27960 = n9721 ^ n3405 ^ 1'b0 ;
  assign n27961 = n27959 & n27960 ;
  assign n27962 = n27961 ^ n7184 ^ 1'b0 ;
  assign n27963 = ( n4485 & n8087 ) | ( n4485 & ~n9437 ) | ( n8087 & ~n9437 ) ;
  assign n27964 = n27963 ^ n8900 ^ 1'b0 ;
  assign n27966 = n3745 | n10071 ;
  assign n27967 = n27966 ^ n17208 ^ 1'b0 ;
  assign n27965 = n14988 ^ n8146 ^ n1134 ;
  assign n27968 = n27967 ^ n27965 ^ n16176 ;
  assign n27969 = n26165 ^ n24554 ^ n18324 ;
  assign n27970 = ( ~n2230 & n11717 ) | ( ~n2230 & n26581 ) | ( n11717 & n26581 ) ;
  assign n27971 = ~n427 & n27970 ;
  assign n27972 = ( n4022 & ~n10265 ) | ( n4022 & n27971 ) | ( ~n10265 & n27971 ) ;
  assign n27973 = n18686 ^ n18273 ^ n10996 ;
  assign n27974 = n15043 & ~n27973 ;
  assign n27975 = n18091 | n24181 ;
  assign n27976 = n27975 ^ n634 ^ 1'b0 ;
  assign n27978 = n18718 ^ n8656 ^ 1'b0 ;
  assign n27979 = n4461 | n27978 ;
  assign n27980 = n27979 ^ n23997 ^ n10334 ;
  assign n27977 = n14368 & ~n18706 ;
  assign n27981 = n27980 ^ n27977 ^ 1'b0 ;
  assign n27983 = ( ~n3608 & n7964 ) | ( ~n3608 & n16883 ) | ( n7964 & n16883 ) ;
  assign n27982 = n20461 ^ n13814 ^ n2696 ;
  assign n27984 = n27983 ^ n27982 ^ n23221 ;
  assign n27985 = ~n5450 & n27280 ;
  assign n27986 = n27985 ^ n1041 ^ 1'b0 ;
  assign n27987 = ( n5196 & n6877 ) | ( n5196 & ~n27986 ) | ( n6877 & ~n27986 ) ;
  assign n27988 = n16071 ^ n4857 ^ n3909 ;
  assign n27989 = ( n22442 & n27987 ) | ( n22442 & n27988 ) | ( n27987 & n27988 ) ;
  assign n27990 = ~n9018 & n11675 ;
  assign n27991 = ~n10009 & n27990 ;
  assign n27992 = n15349 ^ n5574 ^ n1047 ;
  assign n27993 = ( n13032 & ~n27991 ) | ( n13032 & n27992 ) | ( ~n27991 & n27992 ) ;
  assign n27994 = n18232 ^ n13088 ^ n3996 ;
  assign n27995 = ( ~n15850 & n27253 ) | ( ~n15850 & n27994 ) | ( n27253 & n27994 ) ;
  assign n27996 = n21056 ^ n15428 ^ n4560 ;
  assign n27997 = n7473 ^ n4272 ^ 1'b0 ;
  assign n27998 = ~n26778 & n27997 ;
  assign n27999 = n12087 ^ n10719 ^ n5224 ;
  assign n28000 = ( n3967 & ~n14997 ) | ( n3967 & n27999 ) | ( ~n14997 & n27999 ) ;
  assign n28002 = ( ~n3680 & n5795 ) | ( ~n3680 & n11650 ) | ( n5795 & n11650 ) ;
  assign n28003 = ( n3891 & n18311 ) | ( n3891 & n28002 ) | ( n18311 & n28002 ) ;
  assign n28001 = n9421 ^ n7641 ^ n3737 ;
  assign n28004 = n28003 ^ n28001 ^ n27402 ;
  assign n28005 = n24930 ^ n8261 ^ n4583 ;
  assign n28006 = n27239 ^ n19590 ^ 1'b0 ;
  assign n28007 = n5482 ^ n2933 ^ n512 ;
  assign n28008 = ( ~n1657 & n25464 ) | ( ~n1657 & n28007 ) | ( n25464 & n28007 ) ;
  assign n28009 = ( n2341 & ~n3820 ) | ( n2341 & n4041 ) | ( ~n3820 & n4041 ) ;
  assign n28010 = ~n7431 & n22479 ;
  assign n28011 = n28009 & n28010 ;
  assign n28012 = ( ~n20356 & n28008 ) | ( ~n20356 & n28011 ) | ( n28008 & n28011 ) ;
  assign n28013 = n20415 ^ n10235 ^ n4941 ;
  assign n28014 = n28013 ^ n10764 ^ n7052 ;
  assign n28015 = n4538 | n10089 ;
  assign n28016 = n11369 & ~n28015 ;
  assign n28017 = n2617 & n24504 ;
  assign n28018 = n15449 ^ n11685 ^ n8592 ;
  assign n28019 = ( n160 & ~n275 ) | ( n160 & n5555 ) | ( ~n275 & n5555 ) ;
  assign n28020 = ( n13138 & n28018 ) | ( n13138 & n28019 ) | ( n28018 & n28019 ) ;
  assign n28021 = ~n15636 & n22378 ;
  assign n28022 = n28021 ^ n26488 ^ n21397 ;
  assign n28023 = ( ~n12550 & n15654 ) | ( ~n12550 & n28022 ) | ( n15654 & n28022 ) ;
  assign n28024 = n20792 ^ n2481 ^ x107 ;
  assign n28025 = ( ~n15258 & n27578 ) | ( ~n15258 & n28024 ) | ( n27578 & n28024 ) ;
  assign n28026 = ( n5221 & n5796 ) | ( n5221 & n13066 ) | ( n5796 & n13066 ) ;
  assign n28027 = n19217 ^ n17336 ^ n17264 ;
  assign n28028 = ( n12061 & n27347 ) | ( n12061 & n28027 ) | ( n27347 & n28027 ) ;
  assign n28029 = ( ~n1191 & n3067 ) | ( ~n1191 & n17446 ) | ( n3067 & n17446 ) ;
  assign n28030 = ~n4601 & n5386 ;
  assign n28031 = ~n19517 & n28030 ;
  assign n28032 = n2810 ^ n543 ^ 1'b0 ;
  assign n28033 = n22121 | n28032 ;
  assign n28034 = ( n333 & n17574 ) | ( n333 & n28033 ) | ( n17574 & n28033 ) ;
  assign n28035 = n15892 ^ n10048 ^ n3600 ;
  assign n28036 = ( ~n3717 & n28034 ) | ( ~n3717 & n28035 ) | ( n28034 & n28035 ) ;
  assign n28037 = ( n9531 & n17444 ) | ( n9531 & n28036 ) | ( n17444 & n28036 ) ;
  assign n28038 = n6279 & ~n6424 ;
  assign n28039 = n28037 & n28038 ;
  assign n28040 = n10252 ^ n3756 ^ n832 ;
  assign n28041 = ( n325 & n14047 ) | ( n325 & n28040 ) | ( n14047 & n28040 ) ;
  assign n28042 = n22920 ^ n20874 ^ 1'b0 ;
  assign n28048 = n2100 | n21567 ;
  assign n28049 = n28048 ^ n12287 ^ 1'b0 ;
  assign n28043 = ~n2039 & n5797 ;
  assign n28044 = n3285 & n28043 ;
  assign n28045 = ( n387 & ~n15717 ) | ( n387 & n28044 ) | ( ~n15717 & n28044 ) ;
  assign n28046 = n9209 | n28045 ;
  assign n28047 = n14548 & ~n28046 ;
  assign n28050 = n28049 ^ n28047 ^ n8352 ;
  assign n28051 = n12945 ^ n3074 ^ x82 ;
  assign n28052 = ( n4701 & n15575 ) | ( n4701 & n28051 ) | ( n15575 & n28051 ) ;
  assign n28053 = ( n279 & n7359 ) | ( n279 & n19580 ) | ( n7359 & n19580 ) ;
  assign n28054 = n5909 ^ n4926 ^ n2262 ;
  assign n28055 = n713 ^ n334 ^ 1'b0 ;
  assign n28056 = n28054 & ~n28055 ;
  assign n28058 = ( n6665 & n19190 ) | ( n6665 & ~n19865 ) | ( n19190 & ~n19865 ) ;
  assign n28057 = n15876 | n26161 ;
  assign n28059 = n28058 ^ n28057 ^ 1'b0 ;
  assign n28060 = n21756 ^ n14347 ^ n7028 ;
  assign n28061 = n28060 ^ n26933 ^ n11052 ;
  assign n28062 = n510 & n18153 ;
  assign n28063 = ( n3166 & n10182 ) | ( n3166 & n23054 ) | ( n10182 & n23054 ) ;
  assign n28064 = n7705 ^ n6775 ^ n331 ;
  assign n28065 = n17118 ^ n15299 ^ 1'b0 ;
  assign n28066 = n28065 ^ n24116 ^ n6372 ;
  assign n28067 = ~n20985 & n28066 ;
  assign n28068 = n21584 ^ n14830 ^ n12620 ;
  assign n28069 = n19092 ^ n6006 ^ n370 ;
  assign n28070 = n28069 ^ n18504 ^ 1'b0 ;
  assign n28071 = ~n21996 & n28070 ;
  assign n28072 = n2425 | n8321 ;
  assign n28073 = n16200 ^ n3578 ^ 1'b0 ;
  assign n28074 = n28072 & n28073 ;
  assign n28076 = n13305 ^ n11010 ^ n9922 ;
  assign n28075 = ( n2654 & n5743 ) | ( n2654 & n8536 ) | ( n5743 & n8536 ) ;
  assign n28077 = n28076 ^ n28075 ^ n4499 ;
  assign n28078 = ~n8810 & n14171 ;
  assign n28079 = ( ~x23 & n3719 ) | ( ~x23 & n28078 ) | ( n3719 & n28078 ) ;
  assign n28080 = x48 & ~n7868 ;
  assign n28081 = n28080 ^ n4022 ^ 1'b0 ;
  assign n28082 = n23745 ^ n14539 ^ n886 ;
  assign n28083 = ( n1994 & n7338 ) | ( n1994 & n28082 ) | ( n7338 & n28082 ) ;
  assign n28084 = n13469 & ~n28083 ;
  assign n28085 = ( ~n28079 & n28081 ) | ( ~n28079 & n28084 ) | ( n28081 & n28084 ) ;
  assign n28086 = n6267 ^ n3535 ^ n1610 ;
  assign n28087 = ( n5115 & n10234 ) | ( n5115 & n28086 ) | ( n10234 & n28086 ) ;
  assign n28090 = n12211 & ~n15069 ;
  assign n28088 = n18925 ^ n3905 ^ 1'b0 ;
  assign n28089 = ~n4014 & n28088 ;
  assign n28091 = n28090 ^ n28089 ^ n999 ;
  assign n28094 = n12185 ^ n7249 ^ n6794 ;
  assign n28095 = n28094 ^ n14821 ^ n3077 ;
  assign n28092 = n350 & ~n6194 ;
  assign n28093 = n28092 ^ n25546 ^ n6072 ;
  assign n28096 = n28095 ^ n28093 ^ n27442 ;
  assign n28097 = n22705 ^ n14609 ^ n13220 ;
  assign n28098 = ( ~n23219 & n23326 ) | ( ~n23219 & n28097 ) | ( n23326 & n28097 ) ;
  assign n28099 = n28098 ^ n25098 ^ n5980 ;
  assign n28100 = n25427 | n28099 ;
  assign n28101 = ~n3445 & n23158 ;
  assign n28102 = ( n287 & ~n20696 ) | ( n287 & n28101 ) | ( ~n20696 & n28101 ) ;
  assign n28103 = ~n609 & n3387 ;
  assign n28104 = n28103 ^ n25878 ^ 1'b0 ;
  assign n28105 = ~n8450 & n27333 ;
  assign n28106 = ~n15149 & n28105 ;
  assign n28108 = ( n8399 & n17149 ) | ( n8399 & ~n18682 ) | ( n17149 & ~n18682 ) ;
  assign n28109 = ( ~n10528 & n19598 ) | ( ~n10528 & n28108 ) | ( n19598 & n28108 ) ;
  assign n28107 = n15376 | n22848 ;
  assign n28110 = n28109 ^ n28107 ^ 1'b0 ;
  assign n28111 = n17995 & ~n27307 ;
  assign n28112 = ~n1017 & n28111 ;
  assign n28113 = ( n1400 & n10740 ) | ( n1400 & ~n28112 ) | ( n10740 & ~n28112 ) ;
  assign n28114 = n10614 ^ n9243 ^ n5635 ;
  assign n28115 = n28114 ^ n8653 ^ n3273 ;
  assign n28116 = n3967 & n14242 ;
  assign n28117 = n28116 ^ n8564 ^ 1'b0 ;
  assign n28118 = ~n15948 & n28117 ;
  assign n28119 = ( n2011 & ~n10371 ) | ( n2011 & n24441 ) | ( ~n10371 & n24441 ) ;
  assign n28120 = n28119 ^ n5451 ^ 1'b0 ;
  assign n28122 = n1559 ^ n1362 ^ 1'b0 ;
  assign n28121 = n17107 ^ n16552 ^ n5333 ;
  assign n28123 = n28122 ^ n28121 ^ n2631 ;
  assign n28124 = ( n10352 & n28120 ) | ( n10352 & n28123 ) | ( n28120 & n28123 ) ;
  assign n28125 = n10324 ^ n2910 ^ 1'b0 ;
  assign n28126 = ( ~n4056 & n7159 ) | ( ~n4056 & n28125 ) | ( n7159 & n28125 ) ;
  assign n28127 = ~n5320 & n25248 ;
  assign n28128 = n18680 & n28127 ;
  assign n28129 = ( ~n3821 & n5250 ) | ( ~n3821 & n28128 ) | ( n5250 & n28128 ) ;
  assign n28130 = ( n9341 & ~n16046 ) | ( n9341 & n28129 ) | ( ~n16046 & n28129 ) ;
  assign n28131 = n24157 ^ n512 ^ 1'b0 ;
  assign n28133 = ~n3913 & n15274 ;
  assign n28134 = n28133 ^ n4452 ^ 1'b0 ;
  assign n28132 = n7760 & ~n7968 ;
  assign n28135 = n28134 ^ n28132 ^ n8424 ;
  assign n28136 = n17946 & ~n28135 ;
  assign n28137 = n28136 ^ n12137 ^ 1'b0 ;
  assign n28138 = n7793 ^ n2654 ^ 1'b0 ;
  assign n28139 = n2433 & n28138 ;
  assign n28140 = ( n6771 & n21506 ) | ( n6771 & n28139 ) | ( n21506 & n28139 ) ;
  assign n28141 = n28140 ^ n6361 ^ n4536 ;
  assign n28142 = n22701 ^ n14747 ^ n9640 ;
  assign n28144 = ( n4035 & ~n5902 ) | ( n4035 & n19598 ) | ( ~n5902 & n19598 ) ;
  assign n28145 = n28144 ^ n11678 ^ n2523 ;
  assign n28143 = n18903 ^ n7244 ^ n2930 ;
  assign n28146 = n28145 ^ n28143 ^ n18128 ;
  assign n28147 = n10987 ^ n9292 ^ 1'b0 ;
  assign n28148 = n28147 ^ n24809 ^ n1309 ;
  assign n28149 = ( n6427 & ~n6469 ) | ( n6427 & n18612 ) | ( ~n6469 & n18612 ) ;
  assign n28152 = ( ~n7426 & n9781 ) | ( ~n7426 & n10747 ) | ( n9781 & n10747 ) ;
  assign n28150 = n1020 & n1086 ;
  assign n28151 = n9209 & n28150 ;
  assign n28153 = n28152 ^ n28151 ^ n11589 ;
  assign n28154 = ( n5565 & ~n7068 ) | ( n5565 & n23663 ) | ( ~n7068 & n23663 ) ;
  assign n28155 = n388 | n8643 ;
  assign n28156 = n3090 & n12858 ;
  assign n28157 = n28156 ^ n8724 ^ 1'b0 ;
  assign n28158 = ( ~n2727 & n19486 ) | ( ~n2727 & n21647 ) | ( n19486 & n21647 ) ;
  assign n28159 = n10292 & ~n28158 ;
  assign n28160 = n18800 ^ n7588 ^ n1472 ;
  assign n28161 = n16180 | n20964 ;
  assign n28162 = n28160 | n28161 ;
  assign n28163 = n21380 ^ n10790 ^ n1322 ;
  assign n28168 = ( n4587 & n10958 ) | ( n4587 & ~n12529 ) | ( n10958 & ~n12529 ) ;
  assign n28167 = n20681 ^ n16325 ^ n476 ;
  assign n28164 = n7744 ^ n4891 ^ n1664 ;
  assign n28165 = n28164 ^ n15897 ^ 1'b0 ;
  assign n28166 = n9828 & n28165 ;
  assign n28169 = n28168 ^ n28167 ^ n28166 ;
  assign n28170 = ( n27767 & n28163 ) | ( n27767 & n28169 ) | ( n28163 & n28169 ) ;
  assign n28171 = n10485 ^ n6462 ^ 1'b0 ;
  assign n28172 = ~n15223 & n28171 ;
  assign n28173 = n28172 ^ n25665 ^ n2023 ;
  assign n28174 = ( ~n8626 & n18832 ) | ( ~n8626 & n28173 ) | ( n18832 & n28173 ) ;
  assign n28175 = n21180 ^ n20681 ^ n10126 ;
  assign n28176 = ( n14089 & n17273 ) | ( n14089 & ~n22628 ) | ( n17273 & ~n22628 ) ;
  assign n28177 = n28176 ^ n23671 ^ n5212 ;
  assign n28178 = ( ~n2766 & n13448 ) | ( ~n2766 & n17020 ) | ( n13448 & n17020 ) ;
  assign n28179 = ( n2293 & ~n8941 ) | ( n2293 & n12961 ) | ( ~n8941 & n12961 ) ;
  assign n28182 = n20268 ^ n14493 ^ n6670 ;
  assign n28180 = n25371 ^ n7465 ^ n6161 ;
  assign n28181 = n6424 | n28180 ;
  assign n28183 = n28182 ^ n28181 ^ 1'b0 ;
  assign n28184 = n23174 ^ n5357 ^ 1'b0 ;
  assign n28185 = n28183 & n28184 ;
  assign n28186 = n14802 | n19472 ;
  assign n28187 = n28186 ^ n10729 ^ 1'b0 ;
  assign n28188 = n815 & ~n16934 ;
  assign n28189 = ~n13857 & n28188 ;
  assign n28192 = n139 & ~n699 ;
  assign n28191 = n11372 & n16325 ;
  assign n28193 = n28192 ^ n28191 ^ 1'b0 ;
  assign n28190 = n19252 ^ n14959 ^ n4712 ;
  assign n28194 = n28193 ^ n28190 ^ 1'b0 ;
  assign n28195 = n24244 ^ n11775 ^ n8601 ;
  assign n28196 = n28195 ^ n8038 ^ n3499 ;
  assign n28197 = ( n1862 & ~n10744 ) | ( n1862 & n13249 ) | ( ~n10744 & n13249 ) ;
  assign n28198 = n11359 ^ n3555 ^ n2160 ;
  assign n28199 = n28198 ^ n5127 ^ 1'b0 ;
  assign n28200 = n16820 & ~n28199 ;
  assign n28201 = ( n11895 & n13482 ) | ( n11895 & ~n28200 ) | ( n13482 & ~n28200 ) ;
  assign n28205 = n25307 ^ n6157 ^ n6006 ;
  assign n28202 = n17199 ^ n349 ^ 1'b0 ;
  assign n28203 = ( x95 & ~n733 ) | ( x95 & n28202 ) | ( ~n733 & n28202 ) ;
  assign n28204 = ( n23630 & ~n26028 ) | ( n23630 & n28203 ) | ( ~n26028 & n28203 ) ;
  assign n28206 = n28205 ^ n28204 ^ 1'b0 ;
  assign n28207 = n23330 ^ n8703 ^ n7876 ;
  assign n28208 = n28207 ^ n25674 ^ n18945 ;
  assign n28209 = n2279 & ~n12452 ;
  assign n28210 = n28209 ^ n15040 ^ 1'b0 ;
  assign n28211 = n2087 | n2947 ;
  assign n28212 = n1245 | n28211 ;
  assign n28213 = n17199 & ~n28212 ;
  assign n28214 = n25727 ^ n6080 ^ n5298 ;
  assign n28215 = n15834 ^ n15772 ^ n11358 ;
  assign n28216 = n28215 ^ n25067 ^ n13924 ;
  assign n28217 = n28216 ^ n13153 ^ 1'b0 ;
  assign n28218 = ( n1922 & n6262 ) | ( n1922 & n10079 ) | ( n6262 & n10079 ) ;
  assign n28219 = n19981 ^ n7793 ^ 1'b0 ;
  assign n28220 = n15121 | n28219 ;
  assign n28221 = ( n10866 & n28218 ) | ( n10866 & n28220 ) | ( n28218 & n28220 ) ;
  assign n28222 = ( n16347 & n17594 ) | ( n16347 & n20589 ) | ( n17594 & n20589 ) ;
  assign n28223 = ~n1320 & n28222 ;
  assign n28224 = ( n7719 & n8300 ) | ( n7719 & n28223 ) | ( n8300 & n28223 ) ;
  assign n28226 = n5383 & n6707 ;
  assign n28225 = n25093 ^ n21567 ^ n12743 ;
  assign n28227 = n28226 ^ n28225 ^ n5839 ;
  assign n28228 = n28227 ^ n21640 ^ n20560 ;
  assign n28229 = ( n1961 & n2877 ) | ( n1961 & n26299 ) | ( n2877 & n26299 ) ;
  assign n28230 = ( n4434 & ~n10986 ) | ( n4434 & n28229 ) | ( ~n10986 & n28229 ) ;
  assign n28231 = n26208 ^ n20662 ^ 1'b0 ;
  assign n28232 = n1419 & n28231 ;
  assign n28233 = n15097 ^ n4832 ^ n1327 ;
  assign n28234 = n24795 ^ n17557 ^ n9488 ;
  assign n28235 = ( n2964 & ~n7469 ) | ( n2964 & n13947 ) | ( ~n7469 & n13947 ) ;
  assign n28236 = n2378 ^ n2327 ^ n1146 ;
  assign n28240 = n7893 ^ n5583 ^ 1'b0 ;
  assign n28241 = ~n4058 & n28240 ;
  assign n28238 = ( n603 & ~n6739 ) | ( n603 & n17576 ) | ( ~n6739 & n17576 ) ;
  assign n28237 = n20579 ^ n12584 ^ n8559 ;
  assign n28239 = n28238 ^ n28237 ^ n11056 ;
  assign n28242 = n28241 ^ n28239 ^ n15091 ;
  assign n28243 = ~n9781 & n13422 ;
  assign n28244 = n18280 ^ n12143 ^ n3340 ;
  assign n28245 = n17807 ^ n16186 ^ 1'b0 ;
  assign n28246 = n21942 ^ n7187 ^ n6845 ;
  assign n28247 = ( n7457 & n9938 ) | ( n7457 & ~n28246 ) | ( n9938 & ~n28246 ) ;
  assign n28248 = ( n10664 & ~n26383 ) | ( n10664 & n28247 ) | ( ~n26383 & n28247 ) ;
  assign n28249 = n28248 ^ n7171 ^ n1103 ;
  assign n28250 = n28249 ^ n14779 ^ 1'b0 ;
  assign n28251 = ~n28245 & n28250 ;
  assign n28252 = n14945 ^ n9935 ^ n6769 ;
  assign n28253 = n4294 | n21355 ;
  assign n28254 = n16066 | n28253 ;
  assign n28255 = ( n9351 & ~n28252 ) | ( n9351 & n28254 ) | ( ~n28252 & n28254 ) ;
  assign n28256 = ( n3492 & ~n18297 ) | ( n3492 & n19232 ) | ( ~n18297 & n19232 ) ;
  assign n28257 = n28256 ^ n15844 ^ n10247 ;
  assign n28258 = ( n14468 & n23470 ) | ( n14468 & ~n28257 ) | ( n23470 & ~n28257 ) ;
  assign n28259 = n17828 & ~n18256 ;
  assign n28261 = ( n11663 & n12780 ) | ( n11663 & n14498 ) | ( n12780 & n14498 ) ;
  assign n28260 = ( ~n11230 & n11874 ) | ( ~n11230 & n17622 ) | ( n11874 & n17622 ) ;
  assign n28262 = n28261 ^ n28260 ^ n771 ;
  assign n28263 = n17302 & n25489 ;
  assign n28264 = ( n1807 & n27522 ) | ( n1807 & n28263 ) | ( n27522 & n28263 ) ;
  assign n28265 = n22525 ^ n18447 ^ 1'b0 ;
  assign n28266 = n27782 | n28265 ;
  assign n28267 = n20348 ^ n1102 ^ 1'b0 ;
  assign n28268 = x62 & n28267 ;
  assign n28269 = n23852 ^ n12508 ^ n4566 ;
  assign n28270 = ( n25857 & n28268 ) | ( n25857 & n28269 ) | ( n28268 & n28269 ) ;
  assign n28272 = n21525 ^ n7886 ^ 1'b0 ;
  assign n28273 = n19526 & n28272 ;
  assign n28271 = n21619 ^ n20838 ^ n5491 ;
  assign n28274 = n28273 ^ n28271 ^ n2329 ;
  assign n28275 = n17537 ^ n5354 ^ n3603 ;
  assign n28276 = ( n18814 & n19248 ) | ( n18814 & n28275 ) | ( n19248 & n28275 ) ;
  assign n28277 = n6965 & ~n8016 ;
  assign n28278 = n11933 ^ n6924 ^ n4796 ;
  assign n28279 = n3704 ^ n3215 ^ n1884 ;
  assign n28280 = ( n5020 & n28278 ) | ( n5020 & n28279 ) | ( n28278 & n28279 ) ;
  assign n28281 = ( n27317 & ~n28277 ) | ( n27317 & n28280 ) | ( ~n28277 & n28280 ) ;
  assign n28282 = n21600 ^ n4883 ^ n1961 ;
  assign n28283 = ( n16870 & ~n18776 ) | ( n16870 & n25786 ) | ( ~n18776 & n25786 ) ;
  assign n28284 = n24144 ^ n19773 ^ 1'b0 ;
  assign n28285 = n4444 & n28284 ;
  assign n28287 = ( n6117 & n9333 ) | ( n6117 & ~n14520 ) | ( n9333 & ~n14520 ) ;
  assign n28286 = n17139 ^ n6329 ^ n4202 ;
  assign n28288 = n28287 ^ n28286 ^ n15231 ;
  assign n28289 = n28285 & ~n28288 ;
  assign n28290 = n14077 ^ n4964 ^ 1'b0 ;
  assign n28291 = n3620 | n28290 ;
  assign n28292 = n28291 ^ n24345 ^ n2719 ;
  assign n28293 = n11466 ^ n7422 ^ n6322 ;
  assign n28294 = n2788 & n28293 ;
  assign n28295 = n25572 ^ n23097 ^ n9863 ;
  assign n28296 = n6194 ^ n3036 ^ 1'b0 ;
  assign n28297 = n13994 & n28296 ;
  assign n28298 = n28295 & n28297 ;
  assign n28299 = n10645 ^ n8393 ^ n5079 ;
  assign n28300 = n28299 ^ n4958 ^ n4680 ;
  assign n28301 = ( n8339 & n14891 ) | ( n8339 & ~n28300 ) | ( n14891 & ~n28300 ) ;
  assign n28302 = n22302 ^ n10241 ^ 1'b0 ;
  assign n28303 = n28302 ^ n26987 ^ n4546 ;
  assign n28304 = ( ~n7278 & n9117 ) | ( ~n7278 & n9968 ) | ( n9117 & n9968 ) ;
  assign n28305 = n24980 ^ n8207 ^ 1'b0 ;
  assign n28306 = n28304 & ~n28305 ;
  assign n28307 = n28306 ^ n9271 ^ n1348 ;
  assign n28308 = ( n1606 & n14266 ) | ( n1606 & n21800 ) | ( n14266 & n21800 ) ;
  assign n28309 = ( ~n17265 & n17546 ) | ( ~n17265 & n28308 ) | ( n17546 & n28308 ) ;
  assign n28310 = ( n4171 & ~n15519 ) | ( n4171 & n28309 ) | ( ~n15519 & n28309 ) ;
  assign n28311 = n28310 ^ n15984 ^ n1655 ;
  assign n28312 = n720 & n15242 ;
  assign n28313 = ( n12615 & n26580 ) | ( n12615 & n28312 ) | ( n26580 & n28312 ) ;
  assign n28314 = ( n3854 & n14420 ) | ( n3854 & ~n24866 ) | ( n14420 & ~n24866 ) ;
  assign n28315 = n28314 ^ n4786 ^ 1'b0 ;
  assign n28316 = n17052 ^ n6065 ^ n496 ;
  assign n28318 = ( n319 & n5336 ) | ( n319 & n11159 ) | ( n5336 & n11159 ) ;
  assign n28317 = n11196 & n20298 ;
  assign n28319 = n28318 ^ n28317 ^ 1'b0 ;
  assign n28320 = ( n19881 & n28316 ) | ( n19881 & n28319 ) | ( n28316 & n28319 ) ;
  assign n28321 = n24717 & ~n24822 ;
  assign n28322 = n28321 ^ n25285 ^ 1'b0 ;
  assign n28323 = n26936 ^ n12523 ^ n5043 ;
  assign n28324 = n6009 ^ n5843 ^ n363 ;
  assign n28325 = n19458 & ~n28324 ;
  assign n28326 = ~n3215 & n28325 ;
  assign n28327 = ~n28323 & n28326 ;
  assign n28328 = n18036 ^ n10008 ^ n4880 ;
  assign n28329 = n27779 ^ n25106 ^ n2782 ;
  assign n28330 = n11462 ^ n4865 ^ 1'b0 ;
  assign n28331 = n19677 | n28330 ;
  assign n28332 = n28331 ^ n10435 ^ n3164 ;
  assign n28333 = n28332 ^ n16400 ^ n1115 ;
  assign n28334 = n18613 ^ n13663 ^ n10463 ;
  assign n28338 = ( n5024 & ~n15096 ) | ( n5024 & n26733 ) | ( ~n15096 & n26733 ) ;
  assign n28335 = n7677 | n24085 ;
  assign n28336 = n28335 ^ n2431 ^ 1'b0 ;
  assign n28337 = ~n1871 & n28336 ;
  assign n28339 = n28338 ^ n28337 ^ 1'b0 ;
  assign n28340 = n2556 & ~n23075 ;
  assign n28341 = ( ~n1098 & n3640 ) | ( ~n1098 & n6534 ) | ( n3640 & n6534 ) ;
  assign n28342 = ( n19731 & n28340 ) | ( n19731 & n28341 ) | ( n28340 & n28341 ) ;
  assign n28343 = n19843 ^ n6198 ^ 1'b0 ;
  assign n28344 = ~n28342 & n28343 ;
  assign n28345 = n21482 ^ n20489 ^ 1'b0 ;
  assign n28346 = n10292 ^ n9560 ^ 1'b0 ;
  assign n28347 = n7506 | n28346 ;
  assign n28348 = n6082 & ~n12380 ;
  assign n28349 = n28348 ^ n23454 ^ n17262 ;
  assign n28350 = ( n17682 & n28347 ) | ( n17682 & ~n28349 ) | ( n28347 & ~n28349 ) ;
  assign n28351 = ( ~n12068 & n15063 ) | ( ~n12068 & n28350 ) | ( n15063 & n28350 ) ;
  assign n28352 = n28260 ^ n19087 ^ n17041 ;
  assign n28353 = ( n4123 & n16254 ) | ( n4123 & n19254 ) | ( n16254 & n19254 ) ;
  assign n28354 = ( n1280 & n10701 ) | ( n1280 & n17240 ) | ( n10701 & n17240 ) ;
  assign n28355 = n28353 | n28354 ;
  assign n28356 = n16350 ^ n15149 ^ n10410 ;
  assign n28357 = ( ~n10898 & n11359 ) | ( ~n10898 & n16182 ) | ( n11359 & n16182 ) ;
  assign n28358 = ( ~n2233 & n5749 ) | ( ~n2233 & n28357 ) | ( n5749 & n28357 ) ;
  assign n28359 = n28358 ^ n10268 ^ n8123 ;
  assign n28360 = n5416 & n24959 ;
  assign n28361 = ~n9787 & n28360 ;
  assign n28362 = n28361 ^ n12547 ^ n7950 ;
  assign n28363 = n11181 ^ n5477 ^ n3032 ;
  assign n28364 = n15876 ^ n3966 ^ 1'b0 ;
  assign n28365 = ~n19141 & n28364 ;
  assign n28366 = n28365 ^ n7212 ^ 1'b0 ;
  assign n28367 = n2616 & ~n28366 ;
  assign n28368 = n28367 ^ n19648 ^ n14458 ;
  assign n28369 = ( n19104 & n28363 ) | ( n19104 & ~n28368 ) | ( n28363 & ~n28368 ) ;
  assign n28370 = n11741 ^ n5213 ^ 1'b0 ;
  assign n28371 = n4888 ^ n872 ^ 1'b0 ;
  assign n28372 = n19780 ^ n18623 ^ n2555 ;
  assign n28373 = n9657 & ~n16459 ;
  assign n28374 = n19164 ^ n6987 ^ n2998 ;
  assign n28375 = ~n3880 & n14152 ;
  assign n28376 = ( ~n24519 & n26754 ) | ( ~n24519 & n28375 ) | ( n26754 & n28375 ) ;
  assign n28377 = n18345 ^ n16416 ^ n12527 ;
  assign n28378 = n4637 & n28377 ;
  assign n28379 = n3335 & ~n11327 ;
  assign n28380 = ( n2825 & n7135 ) | ( n2825 & ~n28379 ) | ( n7135 & ~n28379 ) ;
  assign n28381 = n22347 ^ n10371 ^ 1'b0 ;
  assign n28382 = n1983 & n2931 ;
  assign n28383 = ( n5714 & n15502 ) | ( n5714 & n28382 ) | ( n15502 & n28382 ) ;
  assign n28384 = n28383 ^ n6420 ^ 1'b0 ;
  assign n28385 = n10715 | n28384 ;
  assign n28386 = n3407 | n16186 ;
  assign n28387 = n2023 & n28386 ;
  assign n28388 = n12322 & n28387 ;
  assign n28389 = n5946 | n11649 ;
  assign n28390 = n28389 ^ n18597 ^ 1'b0 ;
  assign n28391 = ( n3337 & n26740 ) | ( n3337 & n27466 ) | ( n26740 & n27466 ) ;
  assign n28392 = ( ~n3398 & n11415 ) | ( ~n3398 & n25943 ) | ( n11415 & n25943 ) ;
  assign n28393 = ( ~n7062 & n11426 ) | ( ~n7062 & n27275 ) | ( n11426 & n27275 ) ;
  assign n28394 = ( n6435 & n14267 ) | ( n6435 & ~n28393 ) | ( n14267 & ~n28393 ) ;
  assign n28395 = ( n12910 & ~n28392 ) | ( n12910 & n28394 ) | ( ~n28392 & n28394 ) ;
  assign n28396 = n16369 ^ n15657 ^ n5023 ;
  assign n28397 = n22269 ^ n14183 ^ 1'b0 ;
  assign n28398 = n28397 ^ n7780 ^ n4315 ;
  assign n28399 = ( ~n2583 & n28396 ) | ( ~n2583 & n28398 ) | ( n28396 & n28398 ) ;
  assign n28400 = ( n8389 & n14267 ) | ( n8389 & n14809 ) | ( n14267 & n14809 ) ;
  assign n28401 = n24228 ^ n20115 ^ 1'b0 ;
  assign n28403 = n17986 ^ n3667 ^ x122 ;
  assign n28404 = n28403 ^ n3413 ^ 1'b0 ;
  assign n28405 = ( n3231 & n11363 ) | ( n3231 & ~n28404 ) | ( n11363 & ~n28404 ) ;
  assign n28402 = n26156 ^ n1484 ^ 1'b0 ;
  assign n28406 = n28405 ^ n28402 ^ n264 ;
  assign n28408 = n20166 ^ n6905 ^ n1435 ;
  assign n28407 = n10472 ^ n7267 ^ 1'b0 ;
  assign n28409 = n28408 ^ n28407 ^ n7406 ;
  assign n28410 = n12149 ^ n3208 ^ 1'b0 ;
  assign n28411 = n28410 ^ n8578 ^ n8156 ;
  assign n28412 = ( ~n1278 & n13032 ) | ( ~n1278 & n24123 ) | ( n13032 & n24123 ) ;
  assign n28413 = ( n309 & n1528 ) | ( n309 & n5053 ) | ( n1528 & n5053 ) ;
  assign n28414 = n21471 & n28413 ;
  assign n28415 = ~n10057 & n28414 ;
  assign n28416 = n13828 | n28415 ;
  assign n28417 = n28412 | n28416 ;
  assign n28418 = n7333 & ~n27341 ;
  assign n28419 = n1586 & n1713 ;
  assign n28420 = n775 & n28419 ;
  assign n28422 = n12929 ^ n11623 ^ n4525 ;
  assign n28421 = n2808 | n11988 ;
  assign n28423 = n28422 ^ n28421 ^ 1'b0 ;
  assign n28424 = ( n20711 & ~n27152 ) | ( n20711 & n28423 ) | ( ~n27152 & n28423 ) ;
  assign n28429 = ( x39 & ~n13636 ) | ( x39 & n27951 ) | ( ~n13636 & n27951 ) ;
  assign n28425 = ( n10195 & n15822 ) | ( n10195 & ~n22532 ) | ( n15822 & ~n22532 ) ;
  assign n28426 = n28425 ^ n15168 ^ n10490 ;
  assign n28427 = n15523 ^ n4561 ^ 1'b0 ;
  assign n28428 = ~n28426 & n28427 ;
  assign n28430 = n28429 ^ n28428 ^ n24171 ;
  assign n28431 = n8135 & ~n13044 ;
  assign n28432 = n12842 & n28431 ;
  assign n28433 = n28432 ^ n12653 ^ n479 ;
  assign n28434 = n10746 ^ n4557 ^ 1'b0 ;
  assign n28435 = n28434 ^ n20644 ^ n5346 ;
  assign n28436 = n28435 ^ n23971 ^ 1'b0 ;
  assign n28437 = n19295 ^ n7190 ^ n1929 ;
  assign n28438 = ( n2906 & ~n23503 ) | ( n2906 & n23981 ) | ( ~n23503 & n23981 ) ;
  assign n28439 = ( n5181 & n16485 ) | ( n5181 & n28438 ) | ( n16485 & n28438 ) ;
  assign n28440 = n28439 ^ n20287 ^ n16422 ;
  assign n28441 = n20226 ^ n4216 ^ 1'b0 ;
  assign n28442 = n14286 & n28441 ;
  assign n28443 = n28442 ^ n1427 ^ n984 ;
  assign n28444 = n8273 | n10466 ;
  assign n28445 = n28444 ^ n5813 ^ 1'b0 ;
  assign n28446 = ( n6611 & n24868 ) | ( n6611 & ~n28445 ) | ( n24868 & ~n28445 ) ;
  assign n28447 = n28446 ^ n5933 ^ n5189 ;
  assign n28448 = ~n4809 & n12593 ;
  assign n28449 = ~n22971 & n28448 ;
  assign n28450 = n8839 ^ n709 ^ 1'b0 ;
  assign n28452 = n22708 ^ n3182 ^ 1'b0 ;
  assign n28453 = n12333 & n28452 ;
  assign n28454 = ~n13435 & n28453 ;
  assign n28455 = n28454 ^ n9382 ^ 1'b0 ;
  assign n28451 = n7309 | n28449 ;
  assign n28456 = n28455 ^ n28451 ^ 1'b0 ;
  assign n28457 = ( n9257 & n11990 ) | ( n9257 & n21790 ) | ( n11990 & n21790 ) ;
  assign n28458 = ( n2997 & n22698 ) | ( n2997 & n28457 ) | ( n22698 & n28457 ) ;
  assign n28459 = n21035 ^ n18609 ^ n1303 ;
  assign n28460 = ~n9215 & n25160 ;
  assign n28461 = n9143 & n28460 ;
  assign n28462 = n28461 ^ n24482 ^ 1'b0 ;
  assign n28463 = ( n4717 & n13836 ) | ( n4717 & n24527 ) | ( n13836 & n24527 ) ;
  assign n28464 = ( x90 & n10191 ) | ( x90 & ~n19252 ) | ( n10191 & ~n19252 ) ;
  assign n28465 = n28464 ^ n27383 ^ n15242 ;
  assign n28466 = n2073 | n2727 ;
  assign n28467 = n13729 & ~n18013 ;
  assign n28468 = n28467 ^ n22305 ^ n673 ;
  assign n28469 = ( n18532 & ~n28466 ) | ( n18532 & n28468 ) | ( ~n28466 & n28468 ) ;
  assign n28471 = ( ~n2626 & n15681 ) | ( ~n2626 & n16760 ) | ( n15681 & n16760 ) ;
  assign n28470 = n368 & n3386 ;
  assign n28472 = n28471 ^ n28470 ^ 1'b0 ;
  assign n28473 = n16565 ^ n7387 ^ 1'b0 ;
  assign n28474 = ~n11214 & n28473 ;
  assign n28475 = n26207 ^ n23279 ^ n5377 ;
  assign n28476 = n16238 ^ n15847 ^ n6579 ;
  assign n28477 = ~n9267 & n19200 ;
  assign n28478 = n28477 ^ n3513 ^ 1'b0 ;
  assign n28479 = n19106 ^ n9731 ^ n8495 ;
  assign n28480 = n2274 | n2699 ;
  assign n28481 = n24614 ^ n10537 ^ 1'b0 ;
  assign n28482 = ( n338 & n2076 ) | ( n338 & ~n28481 ) | ( n2076 & ~n28481 ) ;
  assign n28483 = ( n1958 & n7627 ) | ( n1958 & ~n7945 ) | ( n7627 & ~n7945 ) ;
  assign n28484 = ( n7548 & n11148 ) | ( n7548 & ~n11971 ) | ( n11148 & ~n11971 ) ;
  assign n28485 = n237 & ~n10409 ;
  assign n28486 = n28485 ^ n20045 ^ n15587 ;
  assign n28487 = n18535 ^ n17432 ^ n689 ;
  assign n28488 = n15002 ^ n9058 ^ 1'b0 ;
  assign n28489 = n11377 ^ n671 ^ 1'b0 ;
  assign n28490 = n27317 & ~n28489 ;
  assign n28491 = ( n10914 & n19545 ) | ( n10914 & n28490 ) | ( n19545 & n28490 ) ;
  assign n28497 = ( n7175 & n7426 ) | ( n7175 & ~n10177 ) | ( n7426 & ~n10177 ) ;
  assign n28496 = n13278 ^ n7367 ^ 1'b0 ;
  assign n28492 = n9316 ^ n8913 ^ n3900 ;
  assign n28493 = n12480 & ~n28492 ;
  assign n28494 = n28493 ^ n14348 ^ n6722 ;
  assign n28495 = ( n12301 & ~n15100 ) | ( n12301 & n28494 ) | ( ~n15100 & n28494 ) ;
  assign n28498 = n28497 ^ n28496 ^ n28495 ;
  assign n28499 = ( n1319 & ~n1705 ) | ( n1319 & n4414 ) | ( ~n1705 & n4414 ) ;
  assign n28500 = n24388 & ~n28499 ;
  assign n28501 = ( n12338 & n27790 ) | ( n12338 & n28500 ) | ( n27790 & n28500 ) ;
  assign n28502 = ( n5441 & ~n11653 ) | ( n5441 & n28501 ) | ( ~n11653 & n28501 ) ;
  assign n28503 = n11896 ^ n6042 ^ n1634 ;
  assign n28504 = ~n11000 & n28503 ;
  assign n28505 = n28504 ^ n8076 ^ 1'b0 ;
  assign n28506 = n28502 | n28505 ;
  assign n28507 = ( n17405 & n18306 ) | ( n17405 & ~n23348 ) | ( n18306 & ~n23348 ) ;
  assign n28508 = n28507 ^ n19762 ^ n17197 ;
  assign n28509 = n3279 | n10537 ;
  assign n28510 = n28508 & ~n28509 ;
  assign n28511 = n3695 ^ n1460 ^ x34 ;
  assign n28512 = n28511 ^ n19782 ^ n8295 ;
  assign n28513 = n9582 & n26189 ;
  assign n28514 = ( ~n3837 & n9974 ) | ( ~n3837 & n28513 ) | ( n9974 & n28513 ) ;
  assign n28516 = n16827 ^ n3767 ^ n2760 ;
  assign n28515 = n12663 ^ n12614 ^ n7788 ;
  assign n28517 = n28516 ^ n28515 ^ n8132 ;
  assign n28518 = ( n12083 & ~n15825 ) | ( n12083 & n28517 ) | ( ~n15825 & n28517 ) ;
  assign n28519 = ( x78 & ~n10198 ) | ( x78 & n28518 ) | ( ~n10198 & n28518 ) ;
  assign n28520 = ( n13536 & ~n14847 ) | ( n13536 & n24475 ) | ( ~n14847 & n24475 ) ;
  assign n28521 = ( n8954 & n28519 ) | ( n8954 & n28520 ) | ( n28519 & n28520 ) ;
  assign n28522 = ( n635 & ~n4997 ) | ( n635 & n9816 ) | ( ~n4997 & n9816 ) ;
  assign n28523 = n27311 ^ n20559 ^ 1'b0 ;
  assign n28524 = n15489 ^ n14187 ^ n4468 ;
  assign n28525 = ( ~n15866 & n28523 ) | ( ~n15866 & n28524 ) | ( n28523 & n28524 ) ;
  assign n28526 = n23368 ^ n13002 ^ 1'b0 ;
  assign n28527 = n878 & n28526 ;
  assign n28529 = n22275 ^ n15726 ^ n1874 ;
  assign n28528 = ( n12470 & n19286 ) | ( n12470 & n21235 ) | ( n19286 & n21235 ) ;
  assign n28530 = n28529 ^ n28528 ^ n1373 ;
  assign n28531 = n12869 ^ n3262 ^ n198 ;
  assign n28532 = n28531 ^ n10861 ^ n7600 ;
  assign n28533 = ( ~n1625 & n9229 ) | ( ~n1625 & n10010 ) | ( n9229 & n10010 ) ;
  assign n28534 = ( ~n3063 & n14335 ) | ( ~n3063 & n16422 ) | ( n14335 & n16422 ) ;
  assign n28535 = ( ~n8793 & n15417 ) | ( ~n8793 & n28534 ) | ( n15417 & n28534 ) ;
  assign n28536 = n25813 ^ n14234 ^ n8610 ;
  assign n28537 = ( n28533 & n28535 ) | ( n28533 & ~n28536 ) | ( n28535 & ~n28536 ) ;
  assign n28538 = n19461 ^ n17920 ^ n10380 ;
  assign n28539 = n17309 ^ n13012 ^ 1'b0 ;
  assign n28541 = ( n1411 & ~n14169 ) | ( n1411 & n15774 ) | ( ~n14169 & n15774 ) ;
  assign n28540 = n21208 ^ n16284 ^ n9987 ;
  assign n28542 = n28541 ^ n28540 ^ n27043 ;
  assign n28543 = n24702 ^ n4466 ^ n483 ;
  assign n28544 = ( n21396 & ~n27732 ) | ( n21396 & n28543 ) | ( ~n27732 & n28543 ) ;
  assign n28545 = n20725 ^ n691 ^ 1'b0 ;
  assign n28546 = ~n7148 & n28545 ;
  assign n28547 = n1866 & ~n2875 ;
  assign n28548 = n12402 & n28547 ;
  assign n28549 = n28548 ^ n26668 ^ 1'b0 ;
  assign n28550 = n4155 & n12414 ;
  assign n28551 = n18263 ^ n13388 ^ n3214 ;
  assign n28552 = ( ~n5427 & n25810 ) | ( ~n5427 & n28551 ) | ( n25810 & n28551 ) ;
  assign n28553 = n28550 | n28552 ;
  assign n28554 = n28549 | n28553 ;
  assign n28555 = ( n4976 & n10264 ) | ( n4976 & ~n17163 ) | ( n10264 & ~n17163 ) ;
  assign n28556 = n8764 ^ n4097 ^ n1365 ;
  assign n28557 = n10171 ^ n7747 ^ n7387 ;
  assign n28558 = ( ~n11114 & n28556 ) | ( ~n11114 & n28557 ) | ( n28556 & n28557 ) ;
  assign n28559 = ( n834 & n16632 ) | ( n834 & ~n18888 ) | ( n16632 & ~n18888 ) ;
  assign n28560 = n28559 ^ n19621 ^ n4878 ;
  assign n28561 = n10280 ^ n2042 ^ 1'b0 ;
  assign n28562 = ( n1255 & n2481 ) | ( n1255 & ~n5782 ) | ( n2481 & ~n5782 ) ;
  assign n28563 = n28562 ^ n22357 ^ n14348 ;
  assign n28564 = n9585 ^ n6309 ^ 1'b0 ;
  assign n28565 = n7051 & n28564 ;
  assign n28566 = ( n17149 & ~n19524 ) | ( n17149 & n25604 ) | ( ~n19524 & n25604 ) ;
  assign n28567 = ( n1805 & n4412 ) | ( n1805 & ~n28566 ) | ( n4412 & ~n28566 ) ;
  assign n28568 = ( n954 & n28565 ) | ( n954 & n28567 ) | ( n28565 & n28567 ) ;
  assign n28569 = ( n14072 & n15708 ) | ( n14072 & ~n28568 ) | ( n15708 & ~n28568 ) ;
  assign n28570 = n17846 ^ n16944 ^ n6641 ;
  assign n28571 = n22001 ^ n5018 ^ n3986 ;
  assign n28572 = ( n2880 & n24224 ) | ( n2880 & ~n28571 ) | ( n24224 & ~n28571 ) ;
  assign n28573 = ( n11674 & n18740 ) | ( n11674 & ~n28572 ) | ( n18740 & ~n28572 ) ;
  assign n28574 = n6838 | n28573 ;
  assign n28575 = n12068 | n28574 ;
  assign n28579 = n18669 ^ n305 ^ 1'b0 ;
  assign n28580 = n28579 ^ n20560 ^ n12562 ;
  assign n28578 = n9931 ^ n2374 ^ 1'b0 ;
  assign n28576 = ~n5552 & n23224 ;
  assign n28577 = n28576 ^ n26148 ^ 1'b0 ;
  assign n28581 = n28580 ^ n28578 ^ n28577 ;
  assign n28582 = ( n11592 & n16280 ) | ( n11592 & ~n16386 ) | ( n16280 & ~n16386 ) ;
  assign n28583 = n20490 ^ n4461 ^ 1'b0 ;
  assign n28584 = n15546 & ~n16587 ;
  assign n28585 = n28584 ^ n22669 ^ n19925 ;
  assign n28586 = n16067 ^ n13471 ^ n6910 ;
  assign n28588 = n10347 ^ n6802 ^ n1735 ;
  assign n28587 = n12256 ^ n9656 ^ 1'b0 ;
  assign n28589 = n28588 ^ n28587 ^ n19765 ;
  assign n28594 = ( ~n451 & n1919 ) | ( ~n451 & n5193 ) | ( n1919 & n5193 ) ;
  assign n28592 = ( n810 & n5437 ) | ( n810 & ~n11663 ) | ( n5437 & ~n11663 ) ;
  assign n28593 = n28592 ^ n5065 ^ n1063 ;
  assign n28590 = n21263 ^ n10622 ^ n6707 ;
  assign n28591 = n28590 ^ n8063 ^ 1'b0 ;
  assign n28595 = n28594 ^ n28593 ^ n28591 ;
  assign n28596 = ( n12103 & n16462 ) | ( n12103 & ~n28595 ) | ( n16462 & ~n28595 ) ;
  assign n28597 = ( n699 & ~n10761 ) | ( n699 & n28596 ) | ( ~n10761 & n28596 ) ;
  assign n28598 = ( n826 & n15121 ) | ( n826 & n16107 ) | ( n15121 & n16107 ) ;
  assign n28599 = ( n3950 & ~n5859 ) | ( n3950 & n12945 ) | ( ~n5859 & n12945 ) ;
  assign n28600 = n21524 ^ n19365 ^ n7976 ;
  assign n28601 = n16598 ^ n10004 ^ n3746 ;
  assign n28602 = n19768 ^ n7996 ^ x117 ;
  assign n28603 = n8782 ^ n6988 ^ n140 ;
  assign n28604 = n28603 ^ n9376 ^ n8516 ;
  assign n28605 = n28604 ^ n24175 ^ n11990 ;
  assign n28606 = ( n869 & n16419 ) | ( n869 & n24899 ) | ( n16419 & n24899 ) ;
  assign n28607 = ( n1994 & n14679 ) | ( n1994 & n28606 ) | ( n14679 & n28606 ) ;
  assign n28608 = ( n5074 & n14017 ) | ( n5074 & ~n25010 ) | ( n14017 & ~n25010 ) ;
  assign n28609 = ( n3053 & n21320 ) | ( n3053 & n28608 ) | ( n21320 & n28608 ) ;
  assign n28610 = n16951 ^ n7646 ^ n2418 ;
  assign n28611 = n28610 ^ n10740 ^ n9939 ;
  assign n28615 = n1336 & ~n9204 ;
  assign n28616 = n28615 ^ n9354 ^ 1'b0 ;
  assign n28612 = ( n1320 & ~n1686 ) | ( n1320 & n1823 ) | ( ~n1686 & n1823 ) ;
  assign n28613 = n28612 ^ n9887 ^ n5528 ;
  assign n28614 = ( n1589 & ~n9967 ) | ( n1589 & n28613 ) | ( ~n9967 & n28613 ) ;
  assign n28617 = n28616 ^ n28614 ^ n18433 ;
  assign n28618 = ~n24015 & n28617 ;
  assign n28619 = n28611 & n28618 ;
  assign n28620 = n23861 ^ n12663 ^ 1'b0 ;
  assign n28623 = ( n204 & n9124 ) | ( n204 & ~n19104 ) | ( n9124 & ~n19104 ) ;
  assign n28621 = n13215 | n18882 ;
  assign n28622 = n28621 ^ n14182 ^ 1'b0 ;
  assign n28624 = n28623 ^ n28622 ^ n6379 ;
  assign n28625 = n8023 & n11902 ;
  assign n28626 = ( n12914 & ~n22571 ) | ( n12914 & n28625 ) | ( ~n22571 & n28625 ) ;
  assign n28627 = n24276 ^ n23616 ^ n10699 ;
  assign n28628 = n28627 ^ n19661 ^ n15240 ;
  assign n28629 = n3462 & ~n24083 ;
  assign n28630 = n28629 ^ n21872 ^ 1'b0 ;
  assign n28631 = ( n8554 & n10273 ) | ( n8554 & n28630 ) | ( n10273 & n28630 ) ;
  assign n28632 = n16654 ^ n16624 ^ 1'b0 ;
  assign n28633 = n12712 ^ n2313 ^ 1'b0 ;
  assign n28634 = n1263 | n1830 ;
  assign n28635 = n1134 & ~n28634 ;
  assign n28636 = n14352 | n28635 ;
  assign n28637 = ( n19186 & n22724 ) | ( n19186 & ~n28636 ) | ( n22724 & ~n28636 ) ;
  assign n28638 = n7232 & n9840 ;
  assign n28639 = n2845 & n28638 ;
  assign n28640 = ( n5010 & n12711 ) | ( n5010 & ~n28639 ) | ( n12711 & ~n28639 ) ;
  assign n28641 = n16516 & ~n28640 ;
  assign n28642 = n19236 ^ n6688 ^ 1'b0 ;
  assign n28643 = ( n7047 & n8237 ) | ( n7047 & n11438 ) | ( n8237 & n11438 ) ;
  assign n28644 = ( n7068 & n12040 ) | ( n7068 & n17827 ) | ( n12040 & n17827 ) ;
  assign n28645 = n28644 ^ n8921 ^ 1'b0 ;
  assign n28648 = ( n4608 & n13351 ) | ( n4608 & ~n19707 ) | ( n13351 & ~n19707 ) ;
  assign n28646 = ~n6285 & n9236 ;
  assign n28647 = ~n2508 & n28646 ;
  assign n28649 = n28648 ^ n28647 ^ n184 ;
  assign n28650 = ( n28643 & n28645 ) | ( n28643 & n28649 ) | ( n28645 & n28649 ) ;
  assign n28651 = n19243 ^ n12621 ^ 1'b0 ;
  assign n28652 = n28651 ^ n22767 ^ n852 ;
  assign n28653 = ( n2211 & n26589 ) | ( n2211 & ~n28652 ) | ( n26589 & ~n28652 ) ;
  assign n28654 = n17090 & n22896 ;
  assign n28655 = n28654 ^ n23535 ^ n23246 ;
  assign n28656 = n6267 & n7795 ;
  assign n28657 = ( n3779 & n5007 ) | ( n3779 & n20934 ) | ( n5007 & n20934 ) ;
  assign n28658 = n6144 & ~n28657 ;
  assign n28659 = n28658 ^ n22166 ^ 1'b0 ;
  assign n28660 = ( n10676 & ~n19655 ) | ( n10676 & n25678 ) | ( ~n19655 & n25678 ) ;
  assign n28661 = n21611 ^ n16501 ^ n7860 ;
  assign n28662 = n8242 ^ n7143 ^ n222 ;
  assign n28663 = n9938 & ~n28662 ;
  assign n28666 = n12884 ^ n5968 ^ n1357 ;
  assign n28664 = ( n9621 & ~n9782 ) | ( n9621 & n11641 ) | ( ~n9782 & n11641 ) ;
  assign n28665 = n28664 ^ n17728 ^ n6059 ;
  assign n28667 = n28666 ^ n28665 ^ n10309 ;
  assign n28668 = n16163 | n25464 ;
  assign n28669 = n15721 ^ n12800 ^ n1675 ;
  assign n28670 = n28669 ^ n19985 ^ n6962 ;
  assign n28671 = n28670 ^ n19827 ^ n1917 ;
  assign n28672 = n12129 | n28671 ;
  assign n28673 = n24895 ^ n21617 ^ n8287 ;
  assign n28674 = ( ~n597 & n6183 ) | ( ~n597 & n28673 ) | ( n6183 & n28673 ) ;
  assign n28675 = ( n5707 & n9091 ) | ( n5707 & n15080 ) | ( n9091 & n15080 ) ;
  assign n28676 = n28675 ^ n22894 ^ n4795 ;
  assign n28677 = n9223 | n21111 ;
  assign n28678 = n1693 & ~n21664 ;
  assign n28679 = ~n7528 & n23948 ;
  assign n28680 = ( n13434 & n24432 ) | ( n13434 & ~n28679 ) | ( n24432 & ~n28679 ) ;
  assign n28681 = n27554 ^ n17492 ^ n9701 ;
  assign n28682 = n3903 & ~n13651 ;
  assign n28683 = ( n9594 & n10948 ) | ( n9594 & ~n16635 ) | ( n10948 & ~n16635 ) ;
  assign n28684 = ( n19639 & n28682 ) | ( n19639 & n28683 ) | ( n28682 & n28683 ) ;
  assign n28685 = n9501 ^ n1950 ^ 1'b0 ;
  assign n28686 = n28685 ^ n27833 ^ 1'b0 ;
  assign n28687 = n12780 | n28686 ;
  assign n28688 = ( n28681 & n28684 ) | ( n28681 & n28687 ) | ( n28684 & n28687 ) ;
  assign n28689 = ( n14002 & n16104 ) | ( n14002 & n17105 ) | ( n16104 & n17105 ) ;
  assign n28690 = n28689 ^ n3178 ^ 1'b0 ;
  assign n28691 = n14755 ^ n10266 ^ n9416 ;
  assign n28692 = n28691 ^ n20420 ^ 1'b0 ;
  assign n28693 = ( ~n6973 & n15125 ) | ( ~n6973 & n23521 ) | ( n15125 & n23521 ) ;
  assign n28694 = n28692 & ~n28693 ;
  assign n28695 = ~n13526 & n23128 ;
  assign n28696 = ~n2721 & n9599 ;
  assign n28697 = n27495 & ~n28696 ;
  assign n28698 = n28697 ^ n8249 ^ 1'b0 ;
  assign n28703 = ( n12287 & n12986 ) | ( n12287 & n21542 ) | ( n12986 & n21542 ) ;
  assign n28701 = n2071 ^ n196 ^ 1'b0 ;
  assign n28702 = n11363 | n28701 ;
  assign n28699 = n9041 | n26143 ;
  assign n28700 = n28699 ^ n1452 ^ 1'b0 ;
  assign n28704 = n28703 ^ n28702 ^ n28700 ;
  assign n28707 = n12184 ^ n8158 ^ n1610 ;
  assign n28705 = n25675 ^ n18789 ^ n11292 ;
  assign n28706 = n28705 ^ n22238 ^ n18274 ;
  assign n28708 = n28707 ^ n28706 ^ n2945 ;
  assign n28709 = n18743 ^ n16565 ^ 1'b0 ;
  assign n28710 = n24441 ^ n10508 ^ n8247 ;
  assign n28711 = n28710 ^ n26533 ^ n4597 ;
  assign n28721 = n5448 ^ n3155 ^ n1643 ;
  assign n28722 = ~n14319 & n28721 ;
  assign n28723 = n28722 ^ n14178 ^ 1'b0 ;
  assign n28712 = n1436 & n4951 ;
  assign n28713 = ( n2569 & ~n2654 ) | ( n2569 & n28712 ) | ( ~n2654 & n28712 ) ;
  assign n28714 = n11599 | n28713 ;
  assign n28715 = n28714 ^ n15298 ^ n1635 ;
  assign n28716 = ( n8541 & n12593 ) | ( n8541 & n18318 ) | ( n12593 & n18318 ) ;
  assign n28717 = ( n163 & ~n11707 ) | ( n163 & n28716 ) | ( ~n11707 & n28716 ) ;
  assign n28718 = n28717 ^ n26498 ^ n12542 ;
  assign n28719 = ( x27 & n28715 ) | ( x27 & n28718 ) | ( n28715 & n28718 ) ;
  assign n28720 = n1385 & n28719 ;
  assign n28724 = n28723 ^ n28720 ^ 1'b0 ;
  assign n28725 = n162 | n19432 ;
  assign n28726 = n24036 & ~n28725 ;
  assign n28727 = ( ~n4195 & n9428 ) | ( ~n4195 & n14173 ) | ( n9428 & n14173 ) ;
  assign n28728 = ( ~n13074 & n19392 ) | ( ~n13074 & n28727 ) | ( n19392 & n28727 ) ;
  assign n28729 = ( ~n1810 & n2876 ) | ( ~n1810 & n13102 ) | ( n2876 & n13102 ) ;
  assign n28730 = ( ~n7267 & n8594 ) | ( ~n7267 & n28729 ) | ( n8594 & n28729 ) ;
  assign n28731 = n28730 ^ n21605 ^ n19618 ;
  assign n28732 = n18070 ^ n13154 ^ n1438 ;
  assign n28733 = n13391 & n14561 ;
  assign n28734 = ( n23519 & n28144 ) | ( n23519 & ~n28733 ) | ( n28144 & ~n28733 ) ;
  assign n28735 = n12586 ^ n6199 ^ n5773 ;
  assign n28736 = n202 | n3538 ;
  assign n28737 = ( n2658 & n24193 ) | ( n2658 & n24659 ) | ( n24193 & n24659 ) ;
  assign n28738 = n9079 ^ n3233 ^ n2529 ;
  assign n28739 = ( ~n17945 & n27983 ) | ( ~n17945 & n28738 ) | ( n27983 & n28738 ) ;
  assign n28740 = n12931 | n28739 ;
  assign n28741 = n28737 & ~n28740 ;
  assign n28742 = ( n3636 & n10463 ) | ( n3636 & n19449 ) | ( n10463 & n19449 ) ;
  assign n28743 = n14629 & ~n28742 ;
  assign n28744 = n28743 ^ n7176 ^ 1'b0 ;
  assign n28745 = n25488 ^ n21634 ^ 1'b0 ;
  assign n28746 = n7157 & ~n28745 ;
  assign n28747 = ( ~n11234 & n13667 ) | ( ~n11234 & n24224 ) | ( n13667 & n24224 ) ;
  assign n28748 = ( n13876 & ~n27045 ) | ( n13876 & n28747 ) | ( ~n27045 & n28747 ) ;
  assign n28749 = ( n2596 & ~n5835 ) | ( n2596 & n16746 ) | ( ~n5835 & n16746 ) ;
  assign n28750 = n9235 & n9271 ;
  assign n28751 = n25138 ^ n13050 ^ n9023 ;
  assign n28752 = ( n9198 & n10661 ) | ( n9198 & n28751 ) | ( n10661 & n28751 ) ;
  assign n28753 = n28752 ^ n8893 ^ n3311 ;
  assign n28754 = ( n2220 & n18628 ) | ( n2220 & n20268 ) | ( n18628 & n20268 ) ;
  assign n28755 = n19919 ^ n6151 ^ 1'b0 ;
  assign n28756 = ~n24944 & n28755 ;
  assign n28757 = ( n1113 & n14501 ) | ( n1113 & ~n28756 ) | ( n14501 & ~n28756 ) ;
  assign n28758 = ~n2356 & n18291 ;
  assign n28759 = n28758 ^ n19355 ^ 1'b0 ;
  assign n28763 = n9964 ^ n2011 ^ n582 ;
  assign n28761 = n26102 ^ n16913 ^ 1'b0 ;
  assign n28762 = n25659 & n28761 ;
  assign n28764 = n28763 ^ n28762 ^ 1'b0 ;
  assign n28760 = n3079 | n10504 ;
  assign n28765 = n28764 ^ n28760 ^ 1'b0 ;
  assign n28766 = n20820 ^ n5399 ^ x117 ;
  assign n28767 = ( n10778 & n17898 ) | ( n10778 & ~n28766 ) | ( n17898 & ~n28766 ) ;
  assign n28768 = n20744 ^ n4222 ^ n2539 ;
  assign n28769 = n1575 | n13857 ;
  assign n28771 = ( n5417 & n10412 ) | ( n5417 & n15483 ) | ( n10412 & n15483 ) ;
  assign n28770 = ~n6581 & n18723 ;
  assign n28772 = n28771 ^ n28770 ^ n3308 ;
  assign n28773 = n2952 | n15012 ;
  assign n28774 = n28773 ^ n17850 ^ 1'b0 ;
  assign n28775 = n16043 ^ n8701 ^ n8109 ;
  assign n28776 = ( ~n25570 & n28774 ) | ( ~n25570 & n28775 ) | ( n28774 & n28775 ) ;
  assign n28777 = ( n706 & n28168 ) | ( n706 & ~n28776 ) | ( n28168 & ~n28776 ) ;
  assign n28778 = n19738 ^ n13587 ^ n7238 ;
  assign n28779 = ( n2186 & n8577 ) | ( n2186 & ~n15233 ) | ( n8577 & ~n15233 ) ;
  assign n28780 = ( n3692 & n4081 ) | ( n3692 & n7509 ) | ( n4081 & n7509 ) ;
  assign n28781 = n28780 ^ n23705 ^ n4935 ;
  assign n28782 = n11718 ^ n11267 ^ 1'b0 ;
  assign n28783 = n2450 & n28782 ;
  assign n28784 = ( n638 & n6721 ) | ( n638 & ~n28783 ) | ( n6721 & ~n28783 ) ;
  assign n28785 = ( n9804 & n27185 ) | ( n9804 & n28784 ) | ( n27185 & n28784 ) ;
  assign n28786 = n28785 ^ n3668 ^ 1'b0 ;
  assign n28787 = n17105 & ~n28786 ;
  assign n28788 = ( n523 & ~n3722 ) | ( n523 & n8149 ) | ( ~n3722 & n8149 ) ;
  assign n28789 = n28788 ^ n4413 ^ 1'b0 ;
  assign n28790 = n395 | n12795 ;
  assign n28791 = n11911 & ~n28790 ;
  assign n28792 = n28791 ^ n10198 ^ n6572 ;
  assign n28793 = ( ~n14567 & n28789 ) | ( ~n14567 & n28792 ) | ( n28789 & n28792 ) ;
  assign n28794 = n22507 ^ n20731 ^ n12284 ;
  assign n28795 = ( ~n5526 & n5782 ) | ( ~n5526 & n15261 ) | ( n5782 & n15261 ) ;
  assign n28796 = ( n2602 & ~n3535 ) | ( n2602 & n7566 ) | ( ~n3535 & n7566 ) ;
  assign n28797 = n28796 ^ n20983 ^ n13931 ;
  assign n28798 = n28797 ^ n5446 ^ n3434 ;
  assign n28799 = ( ~n18138 & n28795 ) | ( ~n18138 & n28798 ) | ( n28795 & n28798 ) ;
  assign n28800 = n13700 ^ n242 ^ 1'b0 ;
  assign n28801 = n28800 ^ n6383 ^ 1'b0 ;
  assign n28802 = ( n4167 & n7180 ) | ( n4167 & n21245 ) | ( n7180 & n21245 ) ;
  assign n28803 = n20250 ^ n12654 ^ n7270 ;
  assign n28804 = n8818 | n16051 ;
  assign n28805 = ( n1144 & n12663 ) | ( n1144 & n27061 ) | ( n12663 & n27061 ) ;
  assign n28806 = n9264 & ~n28805 ;
  assign n28807 = ~n9677 & n28806 ;
  assign n28808 = n22837 ^ n1724 ^ 1'b0 ;
  assign n28809 = n27092 ^ n22815 ^ 1'b0 ;
  assign n28810 = n28808 | n28809 ;
  assign n28811 = n11196 & n12848 ;
  assign n28812 = n3613 & n28811 ;
  assign n28813 = ( n166 & ~n8098 ) | ( n166 & n16917 ) | ( ~n8098 & n16917 ) ;
  assign n28814 = n22898 ^ n5001 ^ n1049 ;
  assign n28815 = ( n2477 & n28675 ) | ( n2477 & ~n28814 ) | ( n28675 & ~n28814 ) ;
  assign n28816 = n852 & ~n28815 ;
  assign n28817 = n4014 & n6084 ;
  assign n28818 = ( n1117 & n8152 ) | ( n1117 & ~n27869 ) | ( n8152 & ~n27869 ) ;
  assign n28819 = ( n8757 & n19896 ) | ( n8757 & ~n24313 ) | ( n19896 & ~n24313 ) ;
  assign n28820 = n2398 | n5417 ;
  assign n28821 = n28820 ^ n23711 ^ n23176 ;
  assign n28822 = n12748 ^ n6331 ^ n1431 ;
  assign n28823 = n28822 ^ n7397 ^ 1'b0 ;
  assign n28824 = ~n2093 & n2826 ;
  assign n28825 = n5058 & n28824 ;
  assign n28826 = ( n3319 & ~n4183 ) | ( n3319 & n12653 ) | ( ~n4183 & n12653 ) ;
  assign n28827 = ~n3118 & n28256 ;
  assign n28828 = n28826 & n28827 ;
  assign n28829 = ( ~n1804 & n4399 ) | ( ~n1804 & n18462 ) | ( n4399 & n18462 ) ;
  assign n28830 = ( n1910 & n3838 ) | ( n1910 & ~n18817 ) | ( n3838 & ~n18817 ) ;
  assign n28832 = n28168 ^ n22913 ^ n11335 ;
  assign n28831 = n11576 ^ n8550 ^ n7108 ;
  assign n28833 = n28832 ^ n28831 ^ 1'b0 ;
  assign n28834 = n26685 ^ n7872 ^ 1'b0 ;
  assign n28835 = n13131 | n28834 ;
  assign n28836 = ( n10614 & ~n13471 ) | ( n10614 & n28835 ) | ( ~n13471 & n28835 ) ;
  assign n28837 = ~n12625 & n15125 ;
  assign n28838 = ( n3900 & ~n15243 ) | ( n3900 & n24802 ) | ( ~n15243 & n24802 ) ;
  assign n28839 = n28838 ^ n18135 ^ n2705 ;
  assign n28840 = ( n6301 & n25586 ) | ( n6301 & n28839 ) | ( n25586 & n28839 ) ;
  assign n28841 = n17108 ^ n13995 ^ 1'b0 ;
  assign n28842 = n12026 | n28841 ;
  assign n28843 = n22230 | n28842 ;
  assign n28844 = n28843 ^ n24867 ^ n260 ;
  assign n28845 = ( n5028 & n15028 ) | ( n5028 & ~n28844 ) | ( n15028 & ~n28844 ) ;
  assign n28846 = ( n12018 & n13774 ) | ( n12018 & n21921 ) | ( n13774 & n21921 ) ;
  assign n28847 = n18037 & n28846 ;
  assign n28848 = n28847 ^ n17922 ^ 1'b0 ;
  assign n28849 = n28848 ^ n4456 ^ 1'b0 ;
  assign n28850 = ( ~n1138 & n1156 ) | ( ~n1138 & n15310 ) | ( n1156 & n15310 ) ;
  assign n28851 = ( ~n772 & n9673 ) | ( ~n772 & n23430 ) | ( n9673 & n23430 ) ;
  assign n28852 = ( n5162 & ~n12101 ) | ( n5162 & n28851 ) | ( ~n12101 & n28851 ) ;
  assign n28856 = ( n1282 & n8540 ) | ( n1282 & ~n19238 ) | ( n8540 & ~n19238 ) ;
  assign n28853 = n1329 | n17142 ;
  assign n28854 = n17757 & ~n28853 ;
  assign n28855 = n28854 ^ n17277 ^ n13491 ;
  assign n28857 = n28856 ^ n28855 ^ 1'b0 ;
  assign n28858 = ( n5631 & ~n19705 ) | ( n5631 & n23889 ) | ( ~n19705 & n23889 ) ;
  assign n28859 = ( n3908 & n28857 ) | ( n3908 & ~n28858 ) | ( n28857 & ~n28858 ) ;
  assign n28860 = ( n3091 & n11096 ) | ( n3091 & n14679 ) | ( n11096 & n14679 ) ;
  assign n28861 = ( ~n13286 & n17237 ) | ( ~n13286 & n28860 ) | ( n17237 & n28860 ) ;
  assign n28862 = ( ~n461 & n11212 ) | ( ~n461 & n26427 ) | ( n11212 & n26427 ) ;
  assign n28863 = n28862 ^ n12113 ^ 1'b0 ;
  assign n28864 = ( n12228 & n12943 ) | ( n12228 & n14364 ) | ( n12943 & n14364 ) ;
  assign n28865 = n28864 ^ n4255 ^ 1'b0 ;
  assign n28866 = ~n19618 & n28865 ;
  assign n28867 = n599 & n23364 ;
  assign n28868 = n28867 ^ n6358 ^ 1'b0 ;
  assign n28869 = n24720 ^ n13638 ^ 1'b0 ;
  assign n28870 = n15869 | n28869 ;
  assign n28871 = ( n236 & n5214 ) | ( n236 & n5484 ) | ( n5214 & n5484 ) ;
  assign n28872 = n28871 ^ n11745 ^ n6210 ;
  assign n28873 = n12022 & n28872 ;
  assign n28874 = n28873 ^ n26679 ^ 1'b0 ;
  assign n28875 = ( n440 & n24831 ) | ( n440 & n28874 ) | ( n24831 & n28874 ) ;
  assign n28876 = ( n15238 & n27982 ) | ( n15238 & n28875 ) | ( n27982 & n28875 ) ;
  assign n28879 = ( n2224 & ~n4969 ) | ( n2224 & n6029 ) | ( ~n4969 & n6029 ) ;
  assign n28877 = n753 & n5050 ;
  assign n28878 = n28877 ^ n23904 ^ 1'b0 ;
  assign n28880 = n28879 ^ n28878 ^ n22552 ;
  assign n28881 = n17169 ^ n9495 ^ n9367 ;
  assign n28882 = ( n21116 & n26624 ) | ( n21116 & ~n28881 ) | ( n26624 & ~n28881 ) ;
  assign n28883 = n16086 ^ n13066 ^ n3785 ;
  assign n28884 = ( n440 & ~n27348 ) | ( n440 & n28883 ) | ( ~n27348 & n28883 ) ;
  assign n28885 = n17729 ^ n10589 ^ 1'b0 ;
  assign n28886 = n28885 ^ n3262 ^ n1166 ;
  assign n28887 = ( n3512 & n27132 ) | ( n3512 & ~n27190 ) | ( n27132 & ~n27190 ) ;
  assign n28888 = n13992 & n26575 ;
  assign n28889 = ~n10645 & n17176 ;
  assign n28890 = n28889 ^ n171 ^ 1'b0 ;
  assign n28891 = n28890 ^ n4092 ^ n851 ;
  assign n28892 = n14848 ^ n9834 ^ n6451 ;
  assign n28893 = n15389 & ~n28892 ;
  assign n28894 = ~n6018 & n28893 ;
  assign n28895 = n17685 ^ n831 ^ 1'b0 ;
  assign n28896 = ~n3396 & n28895 ;
  assign n28897 = ( n13651 & n20511 ) | ( n13651 & n26922 ) | ( n20511 & n26922 ) ;
  assign n28898 = ( n13582 & n28838 ) | ( n13582 & ~n28897 ) | ( n28838 & ~n28897 ) ;
  assign n28899 = n25087 ^ n12390 ^ 1'b0 ;
  assign n28900 = ( n3692 & n16941 ) | ( n3692 & n28899 ) | ( n16941 & n28899 ) ;
  assign n28901 = n28900 ^ n15574 ^ 1'b0 ;
  assign n28902 = ( n14875 & n20006 ) | ( n14875 & n28901 ) | ( n20006 & n28901 ) ;
  assign n28903 = n13557 ^ n1329 ^ n245 ;
  assign n28904 = ( n3204 & n5619 ) | ( n3204 & n28903 ) | ( n5619 & n28903 ) ;
  assign n28905 = ( n4078 & n10771 ) | ( n4078 & n19977 ) | ( n10771 & n19977 ) ;
  assign n28906 = ( n9632 & n10522 ) | ( n9632 & ~n28905 ) | ( n10522 & ~n28905 ) ;
  assign n28907 = ~n3153 & n9255 ;
  assign n28908 = ~n10554 & n28907 ;
  assign n28909 = n22522 ^ n16428 ^ n740 ;
  assign n28910 = ~n28908 & n28909 ;
  assign n28911 = ~n2566 & n19228 ;
  assign n28912 = n26933 ^ n13521 ^ n3776 ;
  assign n28913 = n6159 ^ n3252 ^ n2295 ;
  assign n28914 = ( n14308 & n14567 ) | ( n14308 & n20744 ) | ( n14567 & n20744 ) ;
  assign n28915 = n28914 ^ n26345 ^ n7903 ;
  assign n28916 = ( n13067 & ~n28913 ) | ( n13067 & n28915 ) | ( ~n28913 & n28915 ) ;
  assign n28917 = n8842 ^ n8334 ^ 1'b0 ;
  assign n28918 = ~n6298 & n15478 ;
  assign n28919 = ~n168 & n28918 ;
  assign n28920 = ~n6432 & n22277 ;
  assign n28921 = n28920 ^ n20972 ^ 1'b0 ;
  assign n28922 = n27616 ^ n6181 ^ 1'b0 ;
  assign n28923 = n27106 & ~n28922 ;
  assign n28924 = n28923 ^ n24318 ^ n2305 ;
  assign n28925 = n5458 & n28924 ;
  assign n28926 = ~n18443 & n28925 ;
  assign n28928 = ( n733 & n9516 ) | ( n733 & n10761 ) | ( n9516 & n10761 ) ;
  assign n28927 = n18902 ^ n4924 ^ n1930 ;
  assign n28929 = n28928 ^ n28927 ^ n16217 ;
  assign n28930 = ( n14348 & n21421 ) | ( n14348 & n28929 ) | ( n21421 & n28929 ) ;
  assign n28931 = ( n3883 & n15071 ) | ( n3883 & ~n19387 ) | ( n15071 & ~n19387 ) ;
  assign n28932 = n2787 | n22940 ;
  assign n28933 = n28932 ^ n12095 ^ 1'b0 ;
  assign n28934 = n24408 ^ n10708 ^ n9840 ;
  assign n28935 = n4878 ^ n2107 ^ 1'b0 ;
  assign n28936 = ( n28933 & ~n28934 ) | ( n28933 & n28935 ) | ( ~n28934 & n28935 ) ;
  assign n28937 = n14357 & n19008 ;
  assign n28938 = n13035 ^ n3297 ^ n2128 ;
  assign n28939 = ( n1706 & n28937 ) | ( n1706 & ~n28938 ) | ( n28937 & ~n28938 ) ;
  assign n28940 = ( ~n4452 & n12811 ) | ( ~n4452 & n28939 ) | ( n12811 & n28939 ) ;
  assign n28941 = ( n10962 & ~n14567 ) | ( n10962 & n16354 ) | ( ~n14567 & n16354 ) ;
  assign n28942 = ~n3554 & n18487 ;
  assign n28943 = ~n13104 & n28942 ;
  assign n28944 = ( n6492 & ~n12063 ) | ( n6492 & n20066 ) | ( ~n12063 & n20066 ) ;
  assign n28946 = n8854 ^ n8234 ^ n995 ;
  assign n28945 = ( n15958 & ~n16132 ) | ( n15958 & n23973 ) | ( ~n16132 & n23973 ) ;
  assign n28947 = n28946 ^ n28945 ^ n25748 ;
  assign n28948 = n28947 ^ n23690 ^ 1'b0 ;
  assign n28949 = n13566 ^ n3719 ^ 1'b0 ;
  assign n28950 = n20174 ^ n16915 ^ n5808 ;
  assign n28951 = n28950 ^ n2715 ^ 1'b0 ;
  assign n28952 = ( n7600 & n13708 ) | ( n7600 & n25736 ) | ( n13708 & n25736 ) ;
  assign n28953 = n23156 ^ n22986 ^ n815 ;
  assign n28954 = ( n10519 & n19920 ) | ( n10519 & n28953 ) | ( n19920 & n28953 ) ;
  assign n28957 = n11826 ^ n1061 ^ 1'b0 ;
  assign n28955 = n7439 | n15377 ;
  assign n28956 = n28955 ^ n20736 ^ 1'b0 ;
  assign n28958 = n28957 ^ n28956 ^ n9164 ;
  assign n28959 = n17381 | n23742 ;
  assign n28960 = n28959 ^ n10684 ^ 1'b0 ;
  assign n28961 = n28960 ^ n13464 ^ 1'b0 ;
  assign n28962 = n23250 | n28961 ;
  assign n28963 = n22796 ^ n3833 ^ 1'b0 ;
  assign n28964 = ~n12690 & n28963 ;
  assign n28966 = n5640 & ~n20089 ;
  assign n28967 = n28966 ^ n25598 ^ n25435 ;
  assign n28965 = n5464 | n22990 ;
  assign n28968 = n28967 ^ n28965 ^ 1'b0 ;
  assign n28969 = n19476 ^ n6548 ^ 1'b0 ;
  assign n28971 = ( ~n5526 & n9034 ) | ( ~n5526 & n13083 ) | ( n9034 & n13083 ) ;
  assign n28970 = n6287 & n6784 ;
  assign n28972 = n28971 ^ n28970 ^ n362 ;
  assign n28973 = ( n2272 & n3865 ) | ( n2272 & ~n13740 ) | ( n3865 & ~n13740 ) ;
  assign n28974 = ~n18782 & n28973 ;
  assign n28976 = ( n3847 & n9961 ) | ( n3847 & ~n23599 ) | ( n9961 & ~n23599 ) ;
  assign n28975 = ( n1239 & n18413 ) | ( n1239 & n26863 ) | ( n18413 & n26863 ) ;
  assign n28977 = n28976 ^ n28975 ^ n10049 ;
  assign n28978 = ( n15578 & n28974 ) | ( n15578 & n28977 ) | ( n28974 & n28977 ) ;
  assign n28979 = n13308 ^ n12616 ^ n7898 ;
  assign n28980 = n28979 ^ n17532 ^ 1'b0 ;
  assign n28981 = ~n9930 & n28980 ;
  assign n28982 = n28981 ^ n27658 ^ 1'b0 ;
  assign n28984 = ( n176 & n16196 ) | ( n176 & n27681 ) | ( n16196 & n27681 ) ;
  assign n28985 = ( n6657 & n25739 ) | ( n6657 & ~n28984 ) | ( n25739 & ~n28984 ) ;
  assign n28983 = n21887 ^ n7998 ^ 1'b0 ;
  assign n28986 = n28985 ^ n28983 ^ n19695 ;
  assign n28989 = n25090 ^ n18270 ^ n11822 ;
  assign n28987 = ( n7660 & n15263 ) | ( n7660 & ~n27223 ) | ( n15263 & ~n27223 ) ;
  assign n28988 = ( n4183 & n18475 ) | ( n4183 & n28987 ) | ( n18475 & n28987 ) ;
  assign n28990 = n28989 ^ n28988 ^ n13830 ;
  assign n28991 = ( n3464 & n14101 ) | ( n3464 & n19721 ) | ( n14101 & n19721 ) ;
  assign n28992 = n6840 & ~n28991 ;
  assign n28993 = n28992 ^ n2065 ^ 1'b0 ;
  assign n28995 = ( x68 & ~n3943 ) | ( x68 & n12249 ) | ( ~n3943 & n12249 ) ;
  assign n28994 = n5164 ^ n4892 ^ n2937 ;
  assign n28996 = n28995 ^ n28994 ^ n343 ;
  assign n28997 = ~n14117 & n21708 ;
  assign n28998 = ( n1991 & ~n4266 ) | ( n1991 & n28997 ) | ( ~n4266 & n28997 ) ;
  assign n28999 = n9117 & n10875 ;
  assign n29000 = n2846 & n28999 ;
  assign n29001 = n29000 ^ n15995 ^ n5809 ;
  assign n29002 = n5478 ^ n1940 ^ 1'b0 ;
  assign n29003 = n9424 | n29002 ;
  assign n29004 = n29003 ^ n12076 ^ 1'b0 ;
  assign n29005 = ( n2024 & ~n2644 ) | ( n2024 & n20490 ) | ( ~n2644 & n20490 ) ;
  assign n29006 = n29005 ^ n24214 ^ n12643 ;
  assign n29007 = n3705 | n3885 ;
  assign n29008 = n29007 ^ n8003 ^ 1'b0 ;
  assign n29009 = ( n590 & ~n12600 ) | ( n590 & n29008 ) | ( ~n12600 & n29008 ) ;
  assign n29010 = ( n14337 & n22923 ) | ( n14337 & n29009 ) | ( n22923 & n29009 ) ;
  assign n29011 = n9462 & ~n11715 ;
  assign n29012 = ( ~n27963 & n29010 ) | ( ~n27963 & n29011 ) | ( n29010 & n29011 ) ;
  assign n29013 = ( n3803 & n11148 ) | ( n3803 & ~n17147 ) | ( n11148 & ~n17147 ) ;
  assign n29014 = n26909 ^ n26797 ^ n1331 ;
  assign n29015 = n29014 ^ n4424 ^ 1'b0 ;
  assign n29016 = n29015 ^ n28412 ^ n19192 ;
  assign n29017 = n29016 ^ n1693 ^ 1'b0 ;
  assign n29018 = ~n2881 & n29017 ;
  assign n29019 = ( n2731 & ~n2866 ) | ( n2731 & n12355 ) | ( ~n2866 & n12355 ) ;
  assign n29020 = n29019 ^ n6982 ^ 1'b0 ;
  assign n29021 = n5307 & ~n29020 ;
  assign n29022 = n29021 ^ n6904 ^ 1'b0 ;
  assign n29023 = ( n15266 & n21083 ) | ( n15266 & ~n21405 ) | ( n21083 & ~n21405 ) ;
  assign n29024 = n29023 ^ n25695 ^ n183 ;
  assign n29026 = n14654 ^ n915 ^ 1'b0 ;
  assign n29027 = ~n26937 & n29026 ;
  assign n29025 = n2335 & ~n2376 ;
  assign n29028 = n29027 ^ n29025 ^ n26206 ;
  assign n29029 = ~n8482 & n9153 ;
  assign n29030 = ( n16157 & n26143 ) | ( n16157 & n29029 ) | ( n26143 & n29029 ) ;
  assign n29031 = n7433 ^ n6738 ^ n5896 ;
  assign n29032 = n2360 & n29031 ;
  assign n29033 = n22861 & n29032 ;
  assign n29034 = ( n10657 & ~n18799 ) | ( n10657 & n29033 ) | ( ~n18799 & n29033 ) ;
  assign n29035 = ( n23939 & n26090 ) | ( n23939 & ~n29034 ) | ( n26090 & ~n29034 ) ;
  assign n29036 = n29035 ^ n14824 ^ 1'b0 ;
  assign n29037 = ( n348 & n5972 ) | ( n348 & ~n19672 ) | ( n5972 & ~n19672 ) ;
  assign n29040 = n2690 & ~n6901 ;
  assign n29041 = n29040 ^ n17744 ^ 1'b0 ;
  assign n29038 = n21491 ^ n10073 ^ n8683 ;
  assign n29039 = n29038 ^ n14677 ^ 1'b0 ;
  assign n29042 = n29041 ^ n29039 ^ n16383 ;
  assign n29043 = ( ~n10875 & n13190 ) | ( ~n10875 & n17586 ) | ( n13190 & n17586 ) ;
  assign n29044 = n12876 | n19510 ;
  assign n29045 = ( n5942 & ~n8508 ) | ( n5942 & n29044 ) | ( ~n8508 & n29044 ) ;
  assign n29046 = n10906 & ~n29045 ;
  assign n29047 = n22955 | n29046 ;
  assign n29048 = ( n3075 & n10508 ) | ( n3075 & n12874 ) | ( n10508 & n12874 ) ;
  assign n29049 = ( n3382 & n16928 ) | ( n3382 & ~n29048 ) | ( n16928 & ~n29048 ) ;
  assign n29050 = n22621 ^ n6590 ^ n3463 ;
  assign n29051 = n7738 ^ n6372 ^ 1'b0 ;
  assign n29052 = n29051 ^ n25137 ^ n293 ;
  assign n29053 = n4089 & n10516 ;
  assign n29056 = n8727 & n27951 ;
  assign n29057 = n29056 ^ n11107 ^ 1'b0 ;
  assign n29055 = n3120 & n3791 ;
  assign n29058 = n29057 ^ n29055 ^ 1'b0 ;
  assign n29054 = n28639 ^ n19245 ^ n5583 ;
  assign n29059 = n29058 ^ n29054 ^ n2642 ;
  assign n29060 = n16519 ^ n6273 ^ 1'b0 ;
  assign n29061 = n10119 | n29060 ;
  assign n29062 = ( n3711 & n5062 ) | ( n3711 & ~n23786 ) | ( n5062 & ~n23786 ) ;
  assign n29063 = ( ~n3944 & n8350 ) | ( ~n3944 & n29062 ) | ( n8350 & n29062 ) ;
  assign n29064 = n29063 ^ n10416 ^ n6582 ;
  assign n29065 = ( n26509 & ~n29061 ) | ( n26509 & n29064 ) | ( ~n29061 & n29064 ) ;
  assign n29066 = n10179 ^ n3135 ^ n2637 ;
  assign n29067 = n16814 ^ n8167 ^ n5394 ;
  assign n29068 = ( n1326 & ~n8449 ) | ( n1326 & n29067 ) | ( ~n8449 & n29067 ) ;
  assign n29069 = n29068 ^ n7393 ^ n4629 ;
  assign n29070 = ( n7054 & n29066 ) | ( n7054 & ~n29069 ) | ( n29066 & ~n29069 ) ;
  assign n29071 = n3731 ^ n3104 ^ n2560 ;
  assign n29072 = n29071 ^ n15435 ^ n7425 ;
  assign n29077 = n12976 ^ n235 ^ 1'b0 ;
  assign n29078 = n29077 ^ n22508 ^ n13077 ;
  assign n29073 = n8176 ^ n5752 ^ n2670 ;
  assign n29074 = n29073 ^ n6113 ^ n2411 ;
  assign n29075 = ( n9328 & n9986 ) | ( n9328 & ~n12344 ) | ( n9986 & ~n12344 ) ;
  assign n29076 = ( ~n2138 & n29074 ) | ( ~n2138 & n29075 ) | ( n29074 & n29075 ) ;
  assign n29079 = n29078 ^ n29076 ^ n8621 ;
  assign n29080 = n7732 & n29079 ;
  assign n29081 = n11967 & n29080 ;
  assign n29083 = ( ~n9027 & n9271 ) | ( ~n9027 & n13279 ) | ( n9271 & n13279 ) ;
  assign n29084 = ( n781 & ~n18744 ) | ( n781 & n21497 ) | ( ~n18744 & n21497 ) ;
  assign n29085 = n29084 ^ n19257 ^ 1'b0 ;
  assign n29086 = n29083 & n29085 ;
  assign n29082 = n801 & n19013 ;
  assign n29087 = n29086 ^ n29082 ^ 1'b0 ;
  assign n29088 = ( n10381 & ~n14596 ) | ( n10381 & n18384 ) | ( ~n14596 & n18384 ) ;
  assign n29089 = ( n1091 & n13651 ) | ( n1091 & n19508 ) | ( n13651 & n19508 ) ;
  assign n29090 = n11075 & ~n16150 ;
  assign n29091 = n29090 ^ n25609 ^ n23729 ;
  assign n29092 = ~n1567 & n29091 ;
  assign n29093 = n19317 ^ n16334 ^ n9860 ;
  assign n29094 = ( n4248 & ~n8147 ) | ( n4248 & n29093 ) | ( ~n8147 & n29093 ) ;
  assign n29095 = ( n12208 & n16470 ) | ( n12208 & n29094 ) | ( n16470 & n29094 ) ;
  assign n29096 = n24925 ^ n22286 ^ n4299 ;
  assign n29097 = ( ~n3124 & n5309 ) | ( ~n3124 & n22900 ) | ( n5309 & n22900 ) ;
  assign n29100 = n7698 ^ n5518 ^ n2685 ;
  assign n29098 = n9585 & ~n25100 ;
  assign n29099 = ( n5451 & n28254 ) | ( n5451 & n29098 ) | ( n28254 & n29098 ) ;
  assign n29101 = n29100 ^ n29099 ^ n3233 ;
  assign n29102 = n14166 | n15010 ;
  assign n29103 = n29102 ^ n20814 ^ 1'b0 ;
  assign n29104 = n5573 & ~n28036 ;
  assign n29105 = ~n4778 & n29104 ;
  assign n29106 = n11112 ^ n1822 ^ 1'b0 ;
  assign n29107 = n29106 ^ n24903 ^ n12410 ;
  assign n29108 = n29107 ^ n9628 ^ 1'b0 ;
  assign n29109 = n29105 | n29108 ;
  assign n29110 = n24915 ^ n22436 ^ n21104 ;
  assign n29111 = ( n582 & n2173 ) | ( n582 & n11301 ) | ( n2173 & n11301 ) ;
  assign n29112 = ( n771 & ~n24190 ) | ( n771 & n29111 ) | ( ~n24190 & n29111 ) ;
  assign n29113 = n1153 & n11650 ;
  assign n29114 = ( n6519 & n17695 ) | ( n6519 & ~n29113 ) | ( n17695 & ~n29113 ) ;
  assign n29115 = n8270 | n17986 ;
  assign n29116 = ( n6793 & ~n12900 ) | ( n6793 & n29115 ) | ( ~n12900 & n29115 ) ;
  assign n29117 = n17756 & ~n22195 ;
  assign n29118 = n29117 ^ n7029 ^ 1'b0 ;
  assign n29119 = n29118 ^ n10039 ^ n7305 ;
  assign n29120 = ~n10834 & n24107 ;
  assign n29121 = n29120 ^ n5150 ^ 1'b0 ;
  assign n29122 = n665 | n17051 ;
  assign n29123 = n29122 ^ n12123 ^ 1'b0 ;
  assign n29124 = n9858 | n12091 ;
  assign n29125 = n29123 | n29124 ;
  assign n29126 = ( n29119 & n29121 ) | ( n29119 & n29125 ) | ( n29121 & n29125 ) ;
  assign n29127 = ( n26106 & n26977 ) | ( n26106 & n29126 ) | ( n26977 & n29126 ) ;
  assign n29128 = n3031 ^ n1326 ^ 1'b0 ;
  assign n29129 = ( ~n8676 & n12238 ) | ( ~n8676 & n12767 ) | ( n12238 & n12767 ) ;
  assign n29130 = ( n7309 & ~n27426 ) | ( n7309 & n29129 ) | ( ~n27426 & n29129 ) ;
  assign n29131 = ( n2702 & ~n11114 ) | ( n2702 & n11567 ) | ( ~n11114 & n11567 ) ;
  assign n29132 = n27882 ^ n4840 ^ 1'b0 ;
  assign n29133 = n13123 | n29132 ;
  assign n29134 = n26747 ^ n4445 ^ n3122 ;
  assign n29135 = n29134 ^ n18252 ^ n9258 ;
  assign n29136 = n29135 ^ n28785 ^ n12200 ;
  assign n29137 = n29136 ^ n23512 ^ n23176 ;
  assign n29138 = n11532 | n13371 ;
  assign n29139 = ( n10030 & n13469 ) | ( n10030 & ~n29138 ) | ( n13469 & ~n29138 ) ;
  assign n29140 = ( n7225 & ~n11707 ) | ( n7225 & n29139 ) | ( ~n11707 & n29139 ) ;
  assign n29145 = ( n2008 & n10512 ) | ( n2008 & ~n13481 ) | ( n10512 & ~n13481 ) ;
  assign n29144 = n4611 | n9705 ;
  assign n29146 = n29145 ^ n29144 ^ 1'b0 ;
  assign n29141 = n14736 ^ n5342 ^ 1'b0 ;
  assign n29142 = n29141 ^ n11984 ^ n6349 ;
  assign n29143 = ( n6058 & ~n7001 ) | ( n6058 & n29142 ) | ( ~n7001 & n29142 ) ;
  assign n29147 = n29146 ^ n29143 ^ n27333 ;
  assign n29148 = n11237 | n15549 ;
  assign n29149 = n1710 & n29148 ;
  assign n29150 = n16066 ^ n6741 ^ 1'b0 ;
  assign n29151 = n29150 ^ n17613 ^ n3540 ;
  assign n29152 = n13460 ^ n3285 ^ 1'b0 ;
  assign n29153 = n29152 ^ n9399 ^ n2869 ;
  assign n29154 = n29153 ^ n7987 ^ n7842 ;
  assign n29155 = ( n6659 & n12354 ) | ( n6659 & n22709 ) | ( n12354 & n22709 ) ;
  assign n29156 = ( n3967 & n10803 ) | ( n3967 & ~n10809 ) | ( n10803 & ~n10809 ) ;
  assign n29157 = n17586 ^ n1970 ^ 1'b0 ;
  assign n29158 = ~n20496 & n29157 ;
  assign n29159 = n29158 ^ n4935 ^ 1'b0 ;
  assign n29160 = n29156 & n29159 ;
  assign n29161 = n26625 | n28313 ;
  assign n29162 = n21864 ^ n11088 ^ 1'b0 ;
  assign n29163 = ( n6812 & ~n7483 ) | ( n6812 & n10334 ) | ( ~n7483 & n10334 ) ;
  assign n29164 = n11473 ^ n6253 ^ n3593 ;
  assign n29165 = n26404 ^ n19508 ^ n9608 ;
  assign n29166 = n17302 ^ n9032 ^ n5559 ;
  assign n29167 = ~n23802 & n29166 ;
  assign n29168 = n17376 ^ n11720 ^ n873 ;
  assign n29169 = ( n2025 & n11450 ) | ( n2025 & ~n19232 ) | ( n11450 & ~n19232 ) ;
  assign n29170 = n29169 ^ n29057 ^ n9750 ;
  assign n29171 = ( n1674 & n18290 ) | ( n1674 & ~n29170 ) | ( n18290 & ~n29170 ) ;
  assign n29172 = n24883 ^ n2079 ^ 1'b0 ;
  assign n29173 = n14391 ^ n150 ^ 1'b0 ;
  assign n29174 = n18013 | n29173 ;
  assign n29175 = n10168 & ~n24409 ;
  assign n29176 = n18048 ^ n1286 ^ n563 ;
  assign n29177 = n10783 ^ n4400 ^ n2160 ;
  assign n29178 = ( n10420 & n22213 ) | ( n10420 & n23610 ) | ( n22213 & n23610 ) ;
  assign n29179 = ( ~n2333 & n3201 ) | ( ~n2333 & n7933 ) | ( n3201 & n7933 ) ;
  assign n29180 = n7429 & n12872 ;
  assign n29181 = n21542 & n29180 ;
  assign n29183 = n16928 ^ n4264 ^ n1433 ;
  assign n29182 = n17955 ^ n15369 ^ n1929 ;
  assign n29184 = n29183 ^ n29182 ^ n5906 ;
  assign n29185 = ( n808 & n11404 ) | ( n808 & ~n16988 ) | ( n11404 & ~n16988 ) ;
  assign n29186 = n29185 ^ n2735 ^ 1'b0 ;
  assign n29187 = n21937 | n29186 ;
  assign n29188 = ( n5734 & n29184 ) | ( n5734 & ~n29187 ) | ( n29184 & ~n29187 ) ;
  assign n29189 = n14851 ^ n5186 ^ 1'b0 ;
  assign n29190 = n11494 ^ n4491 ^ 1'b0 ;
  assign n29191 = ~n21762 & n29190 ;
  assign n29192 = ~n5950 & n14829 ;
  assign n29193 = n12762 & n29192 ;
  assign n29194 = ( n2880 & n3328 ) | ( n2880 & n12550 ) | ( n3328 & n12550 ) ;
  assign n29195 = ( ~n12193 & n16820 ) | ( ~n12193 & n29194 ) | ( n16820 & n29194 ) ;
  assign n29196 = ( n4163 & n14570 ) | ( n4163 & ~n20266 ) | ( n14570 & ~n20266 ) ;
  assign n29197 = ( n8253 & n18626 ) | ( n8253 & ~n29196 ) | ( n18626 & ~n29196 ) ;
  assign n29199 = ( n2206 & n7292 ) | ( n2206 & ~n14222 ) | ( n7292 & ~n14222 ) ;
  assign n29198 = n13624 & n15970 ;
  assign n29200 = n29199 ^ n29198 ^ 1'b0 ;
  assign n29201 = ( n14412 & ~n29197 ) | ( n14412 & n29200 ) | ( ~n29197 & n29200 ) ;
  assign n29202 = ( n4432 & n10185 ) | ( n4432 & n20028 ) | ( n10185 & n20028 ) ;
  assign n29203 = n13480 ^ n1791 ^ x31 ;
  assign n29204 = n7863 ^ n6921 ^ n2614 ;
  assign n29205 = ( n8634 & n29203 ) | ( n8634 & n29204 ) | ( n29203 & n29204 ) ;
  assign n29206 = ( n15020 & n22255 ) | ( n15020 & n29205 ) | ( n22255 & n29205 ) ;
  assign n29207 = n26092 ^ n16251 ^ n7868 ;
  assign n29208 = n5121 ^ n3590 ^ n974 ;
  assign n29209 = ( ~n13932 & n17965 ) | ( ~n13932 & n29208 ) | ( n17965 & n29208 ) ;
  assign n29210 = n29209 ^ n12785 ^ n5825 ;
  assign n29211 = n8137 & n9941 ;
  assign n29212 = ( ~n7735 & n12029 ) | ( ~n7735 & n29199 ) | ( n12029 & n29199 ) ;
  assign n29213 = n9451 | n15148 ;
  assign n29214 = n29213 ^ n5049 ^ 1'b0 ;
  assign n29215 = n326 | n14005 ;
  assign n29216 = n29215 ^ n3653 ^ 1'b0 ;
  assign n29217 = n29214 & ~n29216 ;
  assign n29218 = ( n732 & n6516 ) | ( n732 & ~n7261 ) | ( n6516 & ~n7261 ) ;
  assign n29219 = ~n2028 & n29218 ;
  assign n29220 = ~n26873 & n29219 ;
  assign n29221 = ( n2297 & ~n16704 ) | ( n2297 & n29220 ) | ( ~n16704 & n29220 ) ;
  assign n29222 = ( n575 & ~n4029 ) | ( n575 & n29221 ) | ( ~n4029 & n29221 ) ;
  assign n29223 = n29222 ^ n5398 ^ 1'b0 ;
  assign n29224 = n18540 & ~n29223 ;
  assign n29227 = n16508 ^ n8936 ^ 1'b0 ;
  assign n29228 = n16979 & n29227 ;
  assign n29229 = n29228 ^ n22351 ^ 1'b0 ;
  assign n29225 = n16799 ^ n1402 ^ n1391 ;
  assign n29226 = ( n3221 & n26822 ) | ( n3221 & ~n29225 ) | ( n26822 & ~n29225 ) ;
  assign n29230 = n29229 ^ n29226 ^ n16121 ;
  assign n29233 = ( n8185 & n11462 ) | ( n8185 & n21801 ) | ( n11462 & n21801 ) ;
  assign n29231 = n1791 & ~n7008 ;
  assign n29232 = n15952 & n29231 ;
  assign n29234 = n29233 ^ n29232 ^ 1'b0 ;
  assign n29235 = n29234 ^ n7891 ^ n4866 ;
  assign n29236 = n20683 ^ n19997 ^ n4354 ;
  assign n29237 = ( n20233 & n21930 ) | ( n20233 & ~n29236 ) | ( n21930 & ~n29236 ) ;
  assign n29239 = n23939 ^ n16467 ^ n11373 ;
  assign n29238 = ( n7824 & n10502 ) | ( n7824 & n21739 ) | ( n10502 & n21739 ) ;
  assign n29240 = n29239 ^ n29238 ^ n26855 ;
  assign n29241 = n24437 ^ n10881 ^ 1'b0 ;
  assign n29242 = n6576 & n29241 ;
  assign n29243 = n29242 ^ n13782 ^ n8885 ;
  assign n29244 = n13938 & n15080 ;
  assign n29245 = ( n3935 & ~n21856 ) | ( n3935 & n29244 ) | ( ~n21856 & n29244 ) ;
  assign n29246 = n15355 | n25085 ;
  assign n29247 = n29246 ^ n18325 ^ 1'b0 ;
  assign n29248 = n18846 ^ n16679 ^ n309 ;
  assign n29249 = ~n10093 & n29248 ;
  assign n29250 = ~n3785 & n29249 ;
  assign n29251 = n3648 ^ n2459 ^ 1'b0 ;
  assign n29252 = n25133 & n29251 ;
  assign n29253 = ( n12218 & n17690 ) | ( n12218 & ~n29252 ) | ( n17690 & ~n29252 ) ;
  assign n29254 = ( n7528 & n8838 ) | ( n7528 & n23363 ) | ( n8838 & n23363 ) ;
  assign n29255 = n29254 ^ n21693 ^ n18510 ;
  assign n29256 = n14880 ^ n7839 ^ n2576 ;
  assign n29257 = n24374 ^ n19628 ^ 1'b0 ;
  assign n29258 = n17912 & n29257 ;
  assign n29259 = ( ~x118 & n18203 ) | ( ~x118 & n29258 ) | ( n18203 & n29258 ) ;
  assign n29260 = n9038 ^ n7068 ^ n5953 ;
  assign n29261 = n26293 ^ n21449 ^ 1'b0 ;
  assign n29262 = n7965 ^ n5587 ^ n2525 ;
  assign n29263 = n29262 ^ n4281 ^ 1'b0 ;
  assign n29264 = n15208 & ~n29263 ;
  assign n29265 = n24960 ^ n11701 ^ n1224 ;
  assign n29266 = ~n6813 & n16570 ;
  assign n29267 = n29265 & n29266 ;
  assign n29268 = n22864 & n29267 ;
  assign n29269 = ( n10502 & n13909 ) | ( n10502 & ~n20535 ) | ( n13909 & ~n20535 ) ;
  assign n29272 = ( n7516 & n19990 ) | ( n7516 & n28347 ) | ( n19990 & n28347 ) ;
  assign n29270 = n9207 ^ n1870 ^ 1'b0 ;
  assign n29271 = n13948 | n29270 ;
  assign n29273 = n29272 ^ n29271 ^ n23017 ;
  assign n29274 = ( x63 & n683 ) | ( x63 & ~n10828 ) | ( n683 & ~n10828 ) ;
  assign n29275 = n21693 ^ n8797 ^ n1554 ;
  assign n29276 = ( n29242 & n29274 ) | ( n29242 & ~n29275 ) | ( n29274 & ~n29275 ) ;
  assign n29277 = n20871 & n29276 ;
  assign n29279 = n4626 & ~n14682 ;
  assign n29278 = n16573 ^ n11657 ^ 1'b0 ;
  assign n29280 = n29279 ^ n29278 ^ n27958 ;
  assign n29281 = ( n6979 & n12609 ) | ( n6979 & n13825 ) | ( n12609 & n13825 ) ;
  assign n29282 = n4096 ^ n3982 ^ n714 ;
  assign n29283 = n29282 ^ n9254 ^ n6983 ;
  assign n29284 = n22690 ^ n11232 ^ n8212 ;
  assign n29285 = n29274 ^ n23687 ^ n23361 ;
  assign n29286 = ( n15445 & n20090 ) | ( n15445 & n20874 ) | ( n20090 & n20874 ) ;
  assign n29287 = ~n9121 & n29286 ;
  assign n29288 = n29287 ^ n1037 ^ 1'b0 ;
  assign n29289 = n29288 ^ n22265 ^ 1'b0 ;
  assign n29290 = ~n29285 & n29289 ;
  assign n29291 = n25441 ^ n23497 ^ n6802 ;
  assign n29293 = n9192 & n10125 ;
  assign n29292 = n24603 ^ n17837 ^ n4331 ;
  assign n29294 = n29293 ^ n29292 ^ n25818 ;
  assign n29295 = n10559 & n11256 ;
  assign n29296 = n29295 ^ n8211 ^ 1'b0 ;
  assign n29297 = ( ~n5866 & n26890 ) | ( ~n5866 & n29296 ) | ( n26890 & n29296 ) ;
  assign n29298 = n7303 ^ n4844 ^ 1'b0 ;
  assign n29299 = ~n17153 & n29298 ;
  assign n29300 = ( n6071 & n21174 ) | ( n6071 & n29299 ) | ( n21174 & n29299 ) ;
  assign n29301 = ( n1918 & ~n17480 ) | ( n1918 & n22226 ) | ( ~n17480 & n22226 ) ;
  assign n29302 = n3328 & n19452 ;
  assign n29303 = n29302 ^ n5579 ^ 1'b0 ;
  assign n29304 = n29303 ^ n23404 ^ n4741 ;
  assign n29305 = ( n15420 & n29301 ) | ( n15420 & ~n29304 ) | ( n29301 & ~n29304 ) ;
  assign n29306 = ( n13500 & n14931 ) | ( n13500 & ~n21375 ) | ( n14931 & ~n21375 ) ;
  assign n29307 = n20258 ^ n17259 ^ 1'b0 ;
  assign n29308 = ( n1928 & n20491 ) | ( n1928 & ~n25186 ) | ( n20491 & ~n25186 ) ;
  assign n29309 = ( n1417 & n3713 ) | ( n1417 & ~n29308 ) | ( n3713 & ~n29308 ) ;
  assign n29310 = n29309 ^ n8745 ^ n209 ;
  assign n29311 = n29310 ^ n15985 ^ n7518 ;
  assign n29312 = n11152 ^ n2797 ^ x67 ;
  assign n29313 = n19517 ^ n501 ^ 1'b0 ;
  assign n29314 = n29312 & ~n29313 ;
  assign n29315 = n25445 ^ n3713 ^ n799 ;
  assign n29316 = n16129 ^ n7219 ^ 1'b0 ;
  assign n29317 = n29316 ^ n6345 ^ n1117 ;
  assign n29318 = n5274 ^ n5232 ^ n5113 ;
  assign n29319 = n23565 ^ n18267 ^ n7108 ;
  assign n29320 = n3306 ^ n886 ^ 1'b0 ;
  assign n29321 = ~n12251 & n29320 ;
  assign n29322 = ( n17441 & n23616 ) | ( n17441 & n29321 ) | ( n23616 & n29321 ) ;
  assign n29323 = n29322 ^ n18641 ^ n9787 ;
  assign n29324 = ~n5701 & n16303 ;
  assign n29325 = n20084 ^ n4540 ^ 1'b0 ;
  assign n29326 = n3151 | n29325 ;
  assign n29327 = ( n2015 & ~n5473 ) | ( n2015 & n16163 ) | ( ~n5473 & n16163 ) ;
  assign n29328 = n29327 ^ n27608 ^ 1'b0 ;
  assign n29329 = n2696 ^ n1890 ^ 1'b0 ;
  assign n29330 = n29328 & ~n29329 ;
  assign n29331 = n2124 | n26803 ;
  assign n29332 = n14503 | n29331 ;
  assign n29333 = n28955 ^ n26345 ^ 1'b0 ;
  assign n29334 = ( n17880 & n27050 ) | ( n17880 & n29333 ) | ( n27050 & n29333 ) ;
  assign n29335 = ( ~n13808 & n26537 ) | ( ~n13808 & n29334 ) | ( n26537 & n29334 ) ;
  assign n29336 = n15455 ^ n15190 ^ n11649 ;
  assign n29337 = n29336 ^ n27064 ^ n25373 ;
  assign n29338 = ( n16471 & ~n27318 ) | ( n16471 & n28622 ) | ( ~n27318 & n28622 ) ;
  assign n29339 = ( n9253 & n12475 ) | ( n9253 & ~n16636 ) | ( n12475 & ~n16636 ) ;
  assign n29340 = n22421 ^ n14213 ^ n393 ;
  assign n29341 = ( n20643 & ~n23716 ) | ( n20643 & n29340 ) | ( ~n23716 & n29340 ) ;
  assign n29342 = n11801 ^ n8513 ^ n575 ;
  assign n29343 = n1715 & n2584 ;
  assign n29344 = n29343 ^ n19714 ^ 1'b0 ;
  assign n29345 = n23808 ^ n1035 ^ 1'b0 ;
  assign n29346 = n13754 | n29345 ;
  assign n29347 = n468 | n5551 ;
  assign n29348 = n29347 ^ n7309 ^ 1'b0 ;
  assign n29349 = n19121 ^ n6616 ^ n4705 ;
  assign n29350 = n24820 ^ n18718 ^ n13948 ;
  assign n29351 = n6777 ^ n4801 ^ 1'b0 ;
  assign n29352 = n21226 & n29351 ;
  assign n29353 = n11891 ^ n10103 ^ 1'b0 ;
  assign n29354 = n8688 | n29353 ;
  assign n29355 = n29354 ^ n16356 ^ 1'b0 ;
  assign n29356 = n19801 & ~n29355 ;
  assign n29357 = ( n18857 & ~n24205 ) | ( n18857 & n29356 ) | ( ~n24205 & n29356 ) ;
  assign n29358 = ( ~n29350 & n29352 ) | ( ~n29350 & n29357 ) | ( n29352 & n29357 ) ;
  assign n29359 = n8860 | n25091 ;
  assign n29360 = n1940 | n29359 ;
  assign n29361 = ~n13081 & n13606 ;
  assign n29362 = n1554 & ~n29361 ;
  assign n29363 = n29362 ^ n18097 ^ 1'b0 ;
  assign n29364 = n29363 ^ n19279 ^ n16618 ;
  assign n29370 = n9584 & ~n14358 ;
  assign n29371 = n21606 & n29370 ;
  assign n29367 = ~n564 & n1701 ;
  assign n29368 = ~n6976 & n29367 ;
  assign n29366 = n7202 | n26251 ;
  assign n29369 = n29368 ^ n29366 ^ 1'b0 ;
  assign n29365 = n2991 & ~n13588 ;
  assign n29372 = n29371 ^ n29369 ^ n29365 ;
  assign n29373 = n27480 ^ n18018 ^ n12315 ;
  assign n29374 = n23114 ^ n10013 ^ 1'b0 ;
  assign n29375 = ( ~n4743 & n10554 ) | ( ~n4743 & n11707 ) | ( n10554 & n11707 ) ;
  assign n29376 = n29375 ^ n17363 ^ n12192 ;
  assign n29377 = n9585 ^ n4029 ^ n1247 ;
  assign n29380 = ( n4102 & n10813 ) | ( n4102 & ~n24372 ) | ( n10813 & ~n24372 ) ;
  assign n29378 = ( n9104 & ~n16988 ) | ( n9104 & n27452 ) | ( ~n16988 & n27452 ) ;
  assign n29379 = n29378 ^ n9466 ^ x16 ;
  assign n29381 = n29380 ^ n29379 ^ n18564 ;
  assign n29382 = n5316 & ~n24129 ;
  assign n29383 = n29382 ^ n10813 ^ n2276 ;
  assign n29384 = n11320 ^ n11263 ^ n721 ;
  assign n29385 = n29384 ^ n27440 ^ n11021 ;
  assign n29386 = n25911 ^ n25025 ^ n6384 ;
  assign n29387 = n13180 ^ n3215 ^ n3050 ;
  assign n29388 = ( n9258 & ~n23580 ) | ( n9258 & n29387 ) | ( ~n23580 & n29387 ) ;
  assign n29389 = ( ~n372 & n4888 ) | ( ~n372 & n14069 ) | ( n4888 & n14069 ) ;
  assign n29390 = n29389 ^ n11748 ^ n6234 ;
  assign n29391 = ( ~n5531 & n7028 ) | ( ~n5531 & n16335 ) | ( n7028 & n16335 ) ;
  assign n29392 = n29391 ^ n13785 ^ 1'b0 ;
  assign n29393 = ~n26493 & n29392 ;
  assign n29394 = n2446 & n3477 ;
  assign n29395 = ~n25381 & n29394 ;
  assign n29396 = n12498 ^ n8787 ^ 1'b0 ;
  assign n29397 = n6119 | n29396 ;
  assign n29398 = n8098 | n14728 ;
  assign n29399 = n29398 ^ n24280 ^ n23776 ;
  assign n29400 = ( n3156 & ~n14412 ) | ( n3156 & n20907 ) | ( ~n14412 & n20907 ) ;
  assign n29401 = ( ~n1063 & n2150 ) | ( ~n1063 & n3392 ) | ( n2150 & n3392 ) ;
  assign n29402 = ( n1541 & ~n2742 ) | ( n1541 & n29401 ) | ( ~n2742 & n29401 ) ;
  assign n29403 = ( n2074 & n11260 ) | ( n2074 & ~n19128 ) | ( n11260 & ~n19128 ) ;
  assign n29404 = n29403 ^ n13532 ^ n2754 ;
  assign n29405 = ( n558 & ~n7690 ) | ( n558 & n27927 ) | ( ~n7690 & n27927 ) ;
  assign n29406 = n25245 ^ n7645 ^ n5384 ;
  assign n29407 = n454 & n16438 ;
  assign n29408 = ~n12923 & n29407 ;
  assign n29409 = n29408 ^ n14154 ^ n6091 ;
  assign n29410 = n6463 & ~n16652 ;
  assign n29411 = n29410 ^ n13614 ^ 1'b0 ;
  assign n29412 = n17061 ^ n5423 ^ n2719 ;
  assign n29413 = ( n3520 & n9292 ) | ( n3520 & n24598 ) | ( n9292 & n24598 ) ;
  assign n29414 = n8921 & ~n21652 ;
  assign n29415 = n25996 & n29414 ;
  assign n29416 = n15495 ^ n12918 ^ n4269 ;
  assign n29417 = ( n29413 & n29415 ) | ( n29413 & n29416 ) | ( n29415 & n29416 ) ;
  assign n29418 = ( n5987 & n16209 ) | ( n5987 & n16916 ) | ( n16209 & n16916 ) ;
  assign n29419 = ( n6325 & n8313 ) | ( n6325 & n14310 ) | ( n8313 & n14310 ) ;
  assign n29420 = ( n4598 & n18609 ) | ( n4598 & ~n29419 ) | ( n18609 & ~n29419 ) ;
  assign n29421 = n29420 ^ n20451 ^ n10328 ;
  assign n29422 = n12666 & ~n29421 ;
  assign n29423 = ~n8445 & n28976 ;
  assign n29424 = n20002 & n29423 ;
  assign n29425 = n7059 & ~n15882 ;
  assign n29426 = ~n12594 & n29425 ;
  assign n29427 = n1944 & n15274 ;
  assign n29428 = n29427 ^ n27795 ^ 1'b0 ;
  assign n29429 = n28076 ^ n18526 ^ n18452 ;
  assign n29430 = ( n157 & n3904 ) | ( n157 & ~n8755 ) | ( n3904 & ~n8755 ) ;
  assign n29431 = n29430 ^ n24828 ^ n4129 ;
  assign n29432 = n1008 & ~n7991 ;
  assign n29433 = n29432 ^ n14205 ^ 1'b0 ;
  assign n29434 = ( ~n27379 & n29431 ) | ( ~n27379 & n29433 ) | ( n29431 & n29433 ) ;
  assign n29438 = n8631 ^ n5381 ^ 1'b0 ;
  assign n29435 = n12499 ^ n7030 ^ n1630 ;
  assign n29436 = ( n1137 & n2874 ) | ( n1137 & n29435 ) | ( n2874 & n29435 ) ;
  assign n29437 = n21628 & ~n29436 ;
  assign n29439 = n29438 ^ n29437 ^ n24389 ;
  assign n29440 = n24183 ^ n16507 ^ n9889 ;
  assign n29441 = ( ~n7698 & n16481 ) | ( ~n7698 & n29440 ) | ( n16481 & n29440 ) ;
  assign n29442 = n28587 ^ n16649 ^ n1569 ;
  assign n29443 = ( n6515 & n8073 ) | ( n6515 & ~n10099 ) | ( n8073 & ~n10099 ) ;
  assign n29444 = n29443 ^ n12773 ^ n6841 ;
  assign n29445 = ( ~n2050 & n22676 ) | ( ~n2050 & n28994 ) | ( n22676 & n28994 ) ;
  assign n29446 = ( n674 & n2722 ) | ( n674 & n28288 ) | ( n2722 & n28288 ) ;
  assign n29447 = n17480 ^ n2433 ^ 1'b0 ;
  assign n29448 = ~n8863 & n29447 ;
  assign n29450 = ~n4767 & n27280 ;
  assign n29449 = n3136 | n9600 ;
  assign n29451 = n29450 ^ n29449 ^ n16146 ;
  assign n29453 = n9725 ^ n1469 ^ 1'b0 ;
  assign n29454 = ( n837 & n4009 ) | ( n837 & ~n29453 ) | ( n4009 & ~n29453 ) ;
  assign n29455 = n10299 & ~n29454 ;
  assign n29456 = ~n9969 & n29455 ;
  assign n29452 = n14963 ^ n1309 ^ 1'b0 ;
  assign n29457 = n29456 ^ n29452 ^ n21660 ;
  assign n29458 = ( n9611 & ~n25712 ) | ( n9611 & n25875 ) | ( ~n25712 & n25875 ) ;
  assign n29459 = n19994 ^ n15835 ^ n4389 ;
  assign n29460 = ( ~n11516 & n29458 ) | ( ~n11516 & n29459 ) | ( n29458 & n29459 ) ;
  assign n29461 = ~n2220 & n26825 ;
  assign n29462 = ( ~n8538 & n20350 ) | ( ~n8538 & n24085 ) | ( n20350 & n24085 ) ;
  assign n29463 = n2144 & n12313 ;
  assign n29464 = n29463 ^ n23440 ^ n10609 ;
  assign n29465 = ( ~n8109 & n11073 ) | ( ~n8109 & n29464 ) | ( n11073 & n29464 ) ;
  assign n29467 = n3066 ^ n2496 ^ 1'b0 ;
  assign n29466 = n25182 ^ n20607 ^ n5047 ;
  assign n29468 = n29467 ^ n29466 ^ n6556 ;
  assign n29470 = n8171 ^ n4480 ^ 1'b0 ;
  assign n29471 = ~n2172 & n29470 ;
  assign n29472 = n29471 ^ n12060 ^ n11402 ;
  assign n29469 = n11762 | n22329 ;
  assign n29473 = n29472 ^ n29469 ^ 1'b0 ;
  assign n29474 = ( n5186 & ~n15257 ) | ( n5186 & n29473 ) | ( ~n15257 & n29473 ) ;
  assign n29475 = n6889 | n14574 ;
  assign n29476 = n6153 & n11444 ;
  assign n29477 = n29476 ^ n11757 ^ 1'b0 ;
  assign n29478 = n29475 & n29477 ;
  assign n29479 = n29478 ^ n18437 ^ 1'b0 ;
  assign n29480 = n10708 & ~n13681 ;
  assign n29481 = n29480 ^ n17321 ^ 1'b0 ;
  assign n29482 = n4300 ^ n3355 ^ x28 ;
  assign n29483 = ( ~n2279 & n5176 ) | ( ~n2279 & n29482 ) | ( n5176 & n29482 ) ;
  assign n29484 = n14670 ^ n6117 ^ n4024 ;
  assign n29485 = n14451 ^ n5942 ^ n4011 ;
  assign n29486 = n29485 ^ n24733 ^ n5850 ;
  assign n29487 = ( n8130 & ~n12048 ) | ( n8130 & n21455 ) | ( ~n12048 & n21455 ) ;
  assign n29488 = n13088 & ~n15090 ;
  assign n29489 = n29488 ^ n10658 ^ 1'b0 ;
  assign n29490 = n29489 ^ n22126 ^ n4444 ;
  assign n29491 = n29490 ^ n5784 ^ n5502 ;
  assign n29492 = ( n598 & n2089 ) | ( n598 & n13116 ) | ( n2089 & n13116 ) ;
  assign n29493 = ( n4913 & n18213 ) | ( n4913 & ~n29492 ) | ( n18213 & ~n29492 ) ;
  assign n29494 = ( n10001 & n14126 ) | ( n10001 & ~n21686 ) | ( n14126 & ~n21686 ) ;
  assign n29495 = n2695 | n29494 ;
  assign n29496 = n29495 ^ n1418 ^ n172 ;
  assign n29497 = n3511 | n25970 ;
  assign n29498 = n7619 | n29497 ;
  assign n29501 = ( n6851 & n7616 ) | ( n6851 & ~n8514 ) | ( n7616 & ~n8514 ) ;
  assign n29499 = ~n2334 & n4381 ;
  assign n29500 = n21469 & n29499 ;
  assign n29502 = n29501 ^ n29500 ^ n16096 ;
  assign n29503 = n29502 ^ n25586 ^ n2032 ;
  assign n29504 = n29503 ^ n8274 ^ 1'b0 ;
  assign n29505 = n3798 & ~n29504 ;
  assign n29506 = n15265 ^ n13890 ^ n4869 ;
  assign n29507 = n29506 ^ n25479 ^ 1'b0 ;
  assign n29508 = ~n22465 & n29507 ;
  assign n29512 = x25 & n2931 ;
  assign n29513 = n29512 ^ n12635 ^ 1'b0 ;
  assign n29510 = n22204 ^ n14072 ^ n5164 ;
  assign n29511 = n29510 ^ n27999 ^ n27658 ;
  assign n29509 = n17034 ^ n1089 ^ 1'b0 ;
  assign n29514 = n29513 ^ n29511 ^ n29509 ;
  assign n29515 = n9884 | n14614 ;
  assign n29516 = n20931 & n29515 ;
  assign n29517 = n10731 ^ n4735 ^ n1276 ;
  assign n29518 = n26243 ^ n21989 ^ n3216 ;
  assign n29519 = ( ~n10351 & n29517 ) | ( ~n10351 & n29518 ) | ( n29517 & n29518 ) ;
  assign n29520 = ( n17742 & n29516 ) | ( n17742 & ~n29519 ) | ( n29516 & ~n29519 ) ;
  assign n29521 = n7226 ^ n501 ^ 1'b0 ;
  assign n29522 = n2649 & n29521 ;
  assign n29523 = n29522 ^ n24857 ^ n7396 ;
  assign n29524 = ( n16158 & n16701 ) | ( n16158 & ~n22088 ) | ( n16701 & ~n22088 ) ;
  assign n29525 = ( n9116 & ~n22837 ) | ( n9116 & n29524 ) | ( ~n22837 & n29524 ) ;
  assign n29530 = ( n1045 & n2499 ) | ( n1045 & ~n3948 ) | ( n2499 & ~n3948 ) ;
  assign n29526 = n8646 & n16713 ;
  assign n29527 = n29526 ^ n6396 ^ n1889 ;
  assign n29528 = ( ~n1894 & n27784 ) | ( ~n1894 & n29527 ) | ( n27784 & n29527 ) ;
  assign n29529 = ( n17157 & ~n23010 ) | ( n17157 & n29528 ) | ( ~n23010 & n29528 ) ;
  assign n29531 = n29530 ^ n29529 ^ n9100 ;
  assign n29532 = ( n6883 & n9864 ) | ( n6883 & n10136 ) | ( n9864 & n10136 ) ;
  assign n29533 = ( n2626 & ~n3423 ) | ( n2626 & n29532 ) | ( ~n3423 & n29532 ) ;
  assign n29534 = n29533 ^ n29034 ^ n19142 ;
  assign n29535 = ( x73 & ~n13245 ) | ( x73 & n18892 ) | ( ~n13245 & n18892 ) ;
  assign n29537 = ( n6960 & n7472 ) | ( n6960 & n7884 ) | ( n7472 & n7884 ) ;
  assign n29538 = n29537 ^ n8864 ^ n3528 ;
  assign n29536 = ( n4038 & ~n4058 ) | ( n4038 & n28009 ) | ( ~n4058 & n28009 ) ;
  assign n29539 = n29538 ^ n29536 ^ n10622 ;
  assign n29540 = n29539 ^ n24417 ^ 1'b0 ;
  assign n29541 = n14828 ^ n1934 ^ 1'b0 ;
  assign n29542 = n17336 & ~n22023 ;
  assign n29543 = n29542 ^ n333 ^ 1'b0 ;
  assign n29545 = n16563 ^ n8451 ^ 1'b0 ;
  assign n29546 = n14515 & ~n29545 ;
  assign n29544 = ( n9526 & n12340 ) | ( n9526 & ~n15292 ) | ( n12340 & ~n15292 ) ;
  assign n29547 = n29546 ^ n29544 ^ n11872 ;
  assign n29548 = n25112 ^ n21489 ^ n6654 ;
  assign n29549 = n29548 ^ n11612 ^ n2432 ;
  assign n29550 = n29549 ^ n22001 ^ n4208 ;
  assign n29551 = n14974 ^ n13674 ^ n7608 ;
  assign n29552 = n29551 ^ n14832 ^ n3709 ;
  assign n29555 = n16473 ^ n1109 ^ 1'b0 ;
  assign n29553 = n8160 | n12160 ;
  assign n29554 = n4883 & ~n29553 ;
  assign n29556 = n29555 ^ n29554 ^ n12366 ;
  assign n29557 = n1772 & n13581 ;
  assign n29558 = ( n6956 & n25389 ) | ( n6956 & n29557 ) | ( n25389 & n29557 ) ;
  assign n29559 = n857 & ~n10901 ;
  assign n29560 = n29559 ^ n8168 ^ 1'b0 ;
  assign n29561 = n9489 ^ n6777 ^ 1'b0 ;
  assign n29562 = n22155 & n29561 ;
  assign n29563 = n11356 ^ n5613 ^ n4639 ;
  assign n29564 = n9745 | n24146 ;
  assign n29565 = n20420 & ~n29564 ;
  assign n29566 = n29565 ^ n16384 ^ 1'b0 ;
  assign n29567 = n22238 ^ n22143 ^ n6797 ;
  assign n29568 = n29567 ^ n8165 ^ n3543 ;
  assign n29569 = ( ~n1874 & n17333 ) | ( ~n1874 & n29568 ) | ( n17333 & n29568 ) ;
  assign n29570 = n12517 ^ n9541 ^ n4326 ;
  assign n29571 = n29570 ^ n24930 ^ n13810 ;
  assign n29572 = ( ~n8522 & n14991 ) | ( ~n8522 & n24310 ) | ( n14991 & n24310 ) ;
  assign n29573 = ( n25160 & n28348 ) | ( n25160 & n29572 ) | ( n28348 & n29572 ) ;
  assign n29574 = n28379 ^ n2862 ^ n2131 ;
  assign n29575 = ( n13516 & n16527 ) | ( n13516 & n21619 ) | ( n16527 & n21619 ) ;
  assign n29576 = n8120 & ~n29575 ;
  assign n29577 = n13577 & n29576 ;
  assign n29578 = n29577 ^ n29205 ^ n14230 ;
  assign n29579 = n17061 ^ n10441 ^ n10001 ;
  assign n29580 = ~n10475 & n14230 ;
  assign n29581 = ~n24291 & n29580 ;
  assign n29582 = ( n13713 & n24838 ) | ( n13713 & n29016 ) | ( n24838 & n29016 ) ;
  assign n29583 = n4332 ^ n2151 ^ n1456 ;
  assign n29584 = n29583 ^ n21039 ^ n8321 ;
  assign n29585 = ( n717 & n8010 ) | ( n717 & n22652 ) | ( n8010 & n22652 ) ;
  assign n29586 = ( n12030 & ~n17804 ) | ( n12030 & n29585 ) | ( ~n17804 & n29585 ) ;
  assign n29587 = ( n6069 & ~n12865 ) | ( n6069 & n17869 ) | ( ~n12865 & n17869 ) ;
  assign n29588 = n29587 ^ n9869 ^ n9864 ;
  assign n29589 = ( n7559 & n7910 ) | ( n7559 & ~n18564 ) | ( n7910 & ~n18564 ) ;
  assign n29590 = ~n3207 & n15507 ;
  assign n29591 = n7798 & n28097 ;
  assign n29592 = n29555 ^ n25920 ^ n22884 ;
  assign n29593 = ( n12125 & n29591 ) | ( n12125 & ~n29592 ) | ( n29591 & ~n29592 ) ;
  assign n29594 = n3013 & ~n7152 ;
  assign n29595 = n29594 ^ n5526 ^ 1'b0 ;
  assign n29596 = n10626 ^ n6500 ^ 1'b0 ;
  assign n29597 = ~n17242 & n29596 ;
  assign n29598 = n29597 ^ n12801 ^ 1'b0 ;
  assign n29599 = n6035 | n28001 ;
  assign n29600 = n29598 | n29599 ;
  assign n29601 = n5961 ^ n2015 ^ 1'b0 ;
  assign n29602 = n29601 ^ n5632 ^ n2930 ;
  assign n29603 = ( n5113 & ~n6393 ) | ( n5113 & n28625 ) | ( ~n6393 & n28625 ) ;
  assign n29604 = n18159 ^ n14090 ^ 1'b0 ;
  assign n29605 = n2810 & n29604 ;
  assign n29606 = n29605 ^ n18368 ^ n1478 ;
  assign n29607 = ( n5710 & n6995 ) | ( n5710 & n28504 ) | ( n6995 & n28504 ) ;
  assign n29608 = n29607 ^ n23859 ^ n9231 ;
  assign n29609 = n28752 ^ n22195 ^ 1'b0 ;
  assign n29610 = n14183 ^ n11430 ^ n8576 ;
  assign n29611 = ( n4043 & n6184 ) | ( n4043 & ~n12696 ) | ( n6184 & ~n12696 ) ;
  assign n29612 = ( n11290 & n15104 ) | ( n11290 & n20745 ) | ( n15104 & n20745 ) ;
  assign n29613 = n27337 ^ n16379 ^ 1'b0 ;
  assign n29614 = ( n5112 & n8367 ) | ( n5112 & n29613 ) | ( n8367 & n29613 ) ;
  assign n29615 = n7327 & n16431 ;
  assign n29616 = n29615 ^ n3701 ^ 1'b0 ;
  assign n29617 = n29616 ^ n9271 ^ n3306 ;
  assign n29618 = n6277 & n26390 ;
  assign n29619 = n28848 ^ n10008 ^ 1'b0 ;
  assign n29620 = n25210 ^ n15514 ^ 1'b0 ;
  assign n29621 = n4491 | n29620 ;
  assign n29622 = n29621 ^ n23772 ^ n9917 ;
  assign n29623 = ( n1638 & ~n11015 ) | ( n1638 & n29622 ) | ( ~n11015 & n29622 ) ;
  assign n29624 = n26620 ^ n26353 ^ n17213 ;
  assign n29625 = n26487 & ~n29624 ;
  assign n29626 = ~n19276 & n29625 ;
  assign n29627 = n15913 ^ n7013 ^ 1'b0 ;
  assign n29628 = n9757 ^ n2387 ^ n2286 ;
  assign n29629 = n29628 ^ n14020 ^ n760 ;
  assign n29630 = ( n3200 & n5314 ) | ( n3200 & ~n22410 ) | ( n5314 & ~n22410 ) ;
  assign n29631 = n29629 | n29630 ;
  assign n29632 = n5692 | n29334 ;
  assign n29633 = n26864 ^ n7269 ^ n3240 ;
  assign n29634 = n29633 ^ n9801 ^ n7093 ;
  assign n29635 = n18682 ^ n15000 ^ n11249 ;
  assign n29636 = ( n3563 & n9526 ) | ( n3563 & ~n12023 ) | ( n9526 & ~n12023 ) ;
  assign n29637 = n18213 & ~n29636 ;
  assign n29638 = n1701 | n29637 ;
  assign n29639 = ( ~n2610 & n4504 ) | ( ~n2610 & n13125 ) | ( n4504 & n13125 ) ;
  assign n29640 = ( ~n1507 & n15517 ) | ( ~n1507 & n29639 ) | ( n15517 & n29639 ) ;
  assign n29641 = n24314 ^ n19944 ^ 1'b0 ;
  assign n29642 = n29640 & ~n29641 ;
  assign n29643 = ( n7284 & n8861 ) | ( n7284 & ~n15441 ) | ( n8861 & ~n15441 ) ;
  assign n29644 = n13666 ^ n2037 ^ n1802 ;
  assign n29645 = ( n6800 & n20335 ) | ( n6800 & n29644 ) | ( n20335 & n29644 ) ;
  assign n29648 = n1280 & n12263 ;
  assign n29646 = n7274 | n14803 ;
  assign n29647 = n5876 | n29646 ;
  assign n29649 = n29648 ^ n29647 ^ n15429 ;
  assign n29650 = n29649 ^ n8220 ^ n6827 ;
  assign n29651 = ( n23361 & n25946 ) | ( n23361 & ~n29650 ) | ( n25946 & ~n29650 ) ;
  assign n29652 = n3977 & ~n8205 ;
  assign n29653 = n29652 ^ n8578 ^ 1'b0 ;
  assign n29654 = n6433 | n26254 ;
  assign n29655 = ( n1495 & n24708 ) | ( n1495 & n29654 ) | ( n24708 & n29654 ) ;
  assign n29656 = ( n25961 & ~n29653 ) | ( n25961 & n29655 ) | ( ~n29653 & n29655 ) ;
  assign n29657 = n29029 ^ n25264 ^ n7741 ;
  assign n29658 = ( n5625 & n6005 ) | ( n5625 & ~n29657 ) | ( n6005 & ~n29657 ) ;
  assign n29659 = n29658 ^ n18945 ^ n751 ;
  assign n29660 = n22364 ^ n16325 ^ n4934 ;
  assign n29666 = n3118 ^ n2414 ^ 1'b0 ;
  assign n29667 = ~n29513 & n29666 ;
  assign n29668 = n11257 ^ n8763 ^ 1'b0 ;
  assign n29669 = n29667 & n29668 ;
  assign n29663 = ( ~x126 & n1705 ) | ( ~x126 & n12231 ) | ( n1705 & n12231 ) ;
  assign n29661 = n432 & n18379 ;
  assign n29662 = n5766 | n29661 ;
  assign n29664 = n29663 ^ n29662 ^ 1'b0 ;
  assign n29665 = n29664 ^ n10511 ^ 1'b0 ;
  assign n29670 = n29669 ^ n29665 ^ n1868 ;
  assign n29671 = ( n7730 & n11640 ) | ( n7730 & ~n26392 ) | ( n11640 & ~n26392 ) ;
  assign n29672 = n7119 & n29671 ;
  assign n29673 = ( ~n776 & n6868 ) | ( ~n776 & n9143 ) | ( n6868 & n9143 ) ;
  assign n29674 = n29673 ^ n29619 ^ 1'b0 ;
  assign n29675 = n29672 | n29674 ;
  assign n29676 = n27849 ^ n6652 ^ n2808 ;
  assign n29681 = ( n2794 & n4725 ) | ( n2794 & ~n15090 ) | ( n4725 & ~n15090 ) ;
  assign n29677 = n28844 ^ n21240 ^ 1'b0 ;
  assign n29678 = n8991 | n29677 ;
  assign n29679 = n2456 ^ n178 ^ 1'b0 ;
  assign n29680 = ~n29678 & n29679 ;
  assign n29682 = n29681 ^ n29680 ^ 1'b0 ;
  assign n29683 = ~n29676 & n29682 ;
  assign n29684 = n18211 & ~n21719 ;
  assign n29685 = n29684 ^ n21179 ^ 1'b0 ;
  assign n29686 = ( ~n6331 & n13117 ) | ( ~n6331 & n21789 ) | ( n13117 & n21789 ) ;
  assign n29687 = n29686 ^ n15097 ^ n11087 ;
  assign n29688 = n29687 ^ n26987 ^ n1481 ;
  assign n29689 = n7698 ^ n4156 ^ n3372 ;
  assign n29690 = n18739 ^ n13199 ^ n4479 ;
  assign n29691 = ( n1799 & n29689 ) | ( n1799 & n29690 ) | ( n29689 & n29690 ) ;
  assign n29692 = n16384 ^ n12101 ^ n6092 ;
  assign n29693 = n12948 ^ n9564 ^ n3784 ;
  assign n29694 = n16876 ^ n8113 ^ n6242 ;
  assign n29695 = n29694 ^ n2021 ^ 1'b0 ;
  assign n29696 = ( n20330 & ~n21417 ) | ( n20330 & n24146 ) | ( ~n21417 & n24146 ) ;
  assign n29697 = n1378 & ~n3884 ;
  assign n29698 = n29697 ^ n582 ^ 1'b0 ;
  assign n29699 = ( n3995 & n6812 ) | ( n3995 & ~n29698 ) | ( n6812 & ~n29698 ) ;
  assign n29700 = n29699 ^ n25784 ^ 1'b0 ;
  assign n29701 = n13761 ^ n8407 ^ n2328 ;
  assign n29702 = n29701 ^ n17648 ^ n908 ;
  assign n29703 = n18425 ^ n16380 ^ n1241 ;
  assign n29704 = ( n1894 & n29702 ) | ( n1894 & ~n29703 ) | ( n29702 & ~n29703 ) ;
  assign n29705 = ( n7323 & n16617 ) | ( n7323 & n28340 ) | ( n16617 & n28340 ) ;
  assign n29706 = n14973 & n29705 ;
  assign n29707 = n12063 & n29706 ;
  assign n29710 = n10774 ^ n10427 ^ 1'b0 ;
  assign n29711 = n29710 ^ n21001 ^ n19438 ;
  assign n29708 = ( n2405 & ~n13825 ) | ( n2405 & n13971 ) | ( ~n13825 & n13971 ) ;
  assign n29709 = n27716 | n29708 ;
  assign n29712 = n29711 ^ n29709 ^ 1'b0 ;
  assign n29713 = n22886 ^ n14169 ^ 1'b0 ;
  assign n29714 = n323 & n19146 ;
  assign n29715 = n29714 ^ n26698 ^ n11523 ;
  assign n29716 = n21641 ^ n20662 ^ 1'b0 ;
  assign n29717 = n21843 ^ n13596 ^ n10274 ;
  assign n29718 = n167 & n23231 ;
  assign n29719 = n29718 ^ n21765 ^ 1'b0 ;
  assign n29720 = n29719 ^ n18256 ^ n13814 ;
  assign n29721 = n26929 ^ n10681 ^ n6157 ;
  assign n29722 = n29075 ^ n6460 ^ n6180 ;
  assign n29723 = n29722 ^ n13026 ^ n7128 ;
  assign n29724 = ( n1842 & n2689 ) | ( n1842 & n8316 ) | ( n2689 & n8316 ) ;
  assign n29725 = n29724 ^ n24152 ^ n11619 ;
  assign n29726 = n9547 ^ n4137 ^ 1'b0 ;
  assign n29727 = n6931 & ~n29726 ;
  assign n29728 = n26756 & n29727 ;
  assign n29729 = n29725 & n29728 ;
  assign n29730 = n13841 ^ n11984 ^ 1'b0 ;
  assign n29731 = n10185 ^ x21 ^ 1'b0 ;
  assign n29732 = n29730 & n29731 ;
  assign n29733 = n14329 & ~n25342 ;
  assign n29734 = n2094 & ~n19299 ;
  assign n29735 = ~n29733 & n29734 ;
  assign n29736 = ( ~n3094 & n20368 ) | ( ~n3094 & n23981 ) | ( n20368 & n23981 ) ;
  assign n29737 = n27422 ^ n5597 ^ n5010 ;
  assign n29738 = n29736 | n29737 ;
  assign n29739 = n29738 ^ n13278 ^ n6149 ;
  assign n29740 = n29739 ^ n14109 ^ n10522 ;
  assign n29741 = n18398 ^ n12775 ^ n2947 ;
  assign n29742 = n11274 | n16857 ;
  assign n29743 = n29742 ^ n428 ^ 1'b0 ;
  assign n29744 = ( ~n9898 & n24634 ) | ( ~n9898 & n29743 ) | ( n24634 & n29743 ) ;
  assign n29745 = n26978 ^ n15823 ^ n5904 ;
  assign n29746 = n25897 ^ n16460 ^ n4732 ;
  assign n29747 = n29746 ^ n4203 ^ n1628 ;
  assign n29748 = n28976 ^ n17427 ^ n1999 ;
  assign n29749 = n29748 ^ n15464 ^ n3467 ;
  assign n29750 = n5296 & ~n29057 ;
  assign n29751 = n27009 ^ n24530 ^ 1'b0 ;
  assign n29752 = n29750 & n29751 ;
  assign n29753 = n20609 ^ n16613 ^ n8823 ;
  assign n29754 = n29753 ^ n19273 ^ 1'b0 ;
  assign n29755 = n7473 & ~n10735 ;
  assign n29756 = ~n16888 & n29755 ;
  assign n29757 = n29743 ^ n22145 ^ n2945 ;
  assign n29758 = n29757 ^ n13946 ^ n11067 ;
  assign n29759 = ( ~n1145 & n1831 ) | ( ~n1145 & n12017 ) | ( n1831 & n12017 ) ;
  assign n29760 = n29759 ^ n21179 ^ n21150 ;
  assign n29761 = ( ~n8662 & n15363 ) | ( ~n8662 & n29760 ) | ( n15363 & n29760 ) ;
  assign n29763 = n5664 & n6922 ;
  assign n29764 = ~n2831 & n29763 ;
  assign n29762 = n11939 ^ n10195 ^ x79 ;
  assign n29765 = n29764 ^ n29762 ^ n22424 ;
  assign n29766 = n29686 ^ n19609 ^ n7260 ;
  assign n29767 = n17352 ^ n17318 ^ n3929 ;
  assign n29768 = ( n1982 & n2558 ) | ( n1982 & n15099 ) | ( n2558 & n15099 ) ;
  assign n29772 = n21760 ^ n7817 ^ 1'b0 ;
  assign n29773 = n29772 ^ n21682 ^ n5886 ;
  assign n29769 = n14652 ^ n6165 ^ n5676 ;
  assign n29770 = n26047 ^ n3940 ^ n397 ;
  assign n29771 = ( ~n8597 & n29769 ) | ( ~n8597 & n29770 ) | ( n29769 & n29770 ) ;
  assign n29774 = n29773 ^ n29771 ^ n21664 ;
  assign n29775 = ( n3246 & n6905 ) | ( n3246 & ~n23994 ) | ( n6905 & ~n23994 ) ;
  assign n29776 = n18080 ^ n14770 ^ x70 ;
  assign n29777 = n11044 & ~n29776 ;
  assign n29778 = n29777 ^ n22564 ^ 1'b0 ;
  assign n29779 = n19377 ^ n10785 ^ n167 ;
  assign n29780 = n5531 ^ n2837 ^ 1'b0 ;
  assign n29781 = n8753 ^ n7526 ^ n3731 ;
  assign n29782 = n29781 ^ n21966 ^ n19542 ;
  assign n29783 = n12143 ^ n263 ^ 1'b0 ;
  assign n29784 = n10238 | n29783 ;
  assign n29785 = ~n9792 & n18542 ;
  assign n29786 = n29785 ^ n25757 ^ 1'b0 ;
  assign n29787 = n29784 | n29786 ;
  assign n29788 = n23104 ^ n15503 ^ n5585 ;
  assign n29789 = n27452 ^ n24517 ^ n11844 ;
  assign n29790 = n9569 ^ n7954 ^ n4465 ;
  assign n29791 = n29790 ^ n24342 ^ n22849 ;
  assign n29792 = n29791 ^ n13736 ^ n12898 ;
  assign n29793 = n29792 ^ n6133 ^ n2577 ;
  assign n29794 = n8893 | n26186 ;
  assign n29795 = n29794 ^ n1715 ^ 1'b0 ;
  assign n29796 = n29795 ^ n18551 ^ n196 ;
  assign n29797 = n29796 ^ n5763 ^ n1263 ;
  assign n29798 = n6857 & n26494 ;
  assign n29799 = n5204 & n29798 ;
  assign n29800 = ~n4368 & n15855 ;
  assign n29801 = n29800 ^ n16380 ^ 1'b0 ;
  assign n29802 = n4228 & ~n29801 ;
  assign n29803 = n29799 & n29802 ;
  assign n29804 = n12728 ^ n3136 ^ n2722 ;
  assign n29805 = n29804 ^ n22695 ^ n1052 ;
  assign n29806 = ( n995 & n4378 ) | ( n995 & ~n7898 ) | ( n4378 & ~n7898 ) ;
  assign n29807 = n29806 ^ n6133 ^ n3585 ;
  assign n29808 = ( n5049 & n29805 ) | ( n5049 & ~n29807 ) | ( n29805 & ~n29807 ) ;
  assign n29809 = n29808 ^ n17278 ^ 1'b0 ;
  assign n29811 = n14453 ^ n5506 ^ n4878 ;
  assign n29812 = n29811 ^ n17012 ^ n2515 ;
  assign n29810 = n24074 ^ n4539 ^ n2233 ;
  assign n29813 = n29812 ^ n29810 ^ n4793 ;
  assign n29822 = n2966 & ~n6903 ;
  assign n29823 = ~n3012 & n29822 ;
  assign n29820 = n9412 ^ n9227 ^ n1594 ;
  assign n29821 = n29820 ^ n13913 ^ n4295 ;
  assign n29816 = n3108 | n4633 ;
  assign n29817 = n29816 ^ n2771 ^ 1'b0 ;
  assign n29814 = n4004 | n16791 ;
  assign n29815 = n29814 ^ n5407 ^ 1'b0 ;
  assign n29818 = n29817 ^ n29815 ^ n4021 ;
  assign n29819 = ( ~n3488 & n13223 ) | ( ~n3488 & n29818 ) | ( n13223 & n29818 ) ;
  assign n29824 = n29823 ^ n29821 ^ n29819 ;
  assign n29825 = n5652 | n20984 ;
  assign n29826 = n25541 ^ n11514 ^ n8647 ;
  assign n29827 = n26033 ^ n3114 ^ n2277 ;
  assign n29828 = n25487 ^ n4205 ^ 1'b0 ;
  assign n29829 = ~n3642 & n29828 ;
  assign n29830 = n1541 & ~n27747 ;
  assign n29831 = n29830 ^ n19448 ^ 1'b0 ;
  assign n29832 = ~n4406 & n23763 ;
  assign n29833 = n29832 ^ n4129 ^ 1'b0 ;
  assign n29834 = n27258 ^ n26830 ^ n6095 ;
  assign n29835 = n14533 & ~n29834 ;
  assign n29836 = n1007 | n29835 ;
  assign n29837 = n29833 | n29836 ;
  assign n29839 = ( n4917 & n10560 ) | ( n4917 & ~n21023 ) | ( n10560 & ~n21023 ) ;
  assign n29838 = ( ~n8003 & n9207 ) | ( ~n8003 & n13653 ) | ( n9207 & n13653 ) ;
  assign n29840 = n29839 ^ n29838 ^ 1'b0 ;
  assign n29841 = n22138 ^ n2415 ^ 1'b0 ;
  assign n29842 = n3395 & n29841 ;
  assign n29843 = n29842 ^ n22156 ^ n5841 ;
  assign n29844 = n18349 ^ n17046 ^ n12036 ;
  assign n29845 = n22215 ^ n7236 ^ 1'b0 ;
  assign n29846 = n6036 | n9575 ;
  assign n29847 = n29846 ^ n2661 ^ 1'b0 ;
  assign n29848 = n26000 ^ n8433 ^ 1'b0 ;
  assign n29849 = ~n29847 & n29848 ;
  assign n29850 = ( ~n19674 & n23724 ) | ( ~n19674 & n29849 ) | ( n23724 & n29849 ) ;
  assign n29851 = ( n2810 & n6613 ) | ( n2810 & n9454 ) | ( n6613 & n9454 ) ;
  assign n29852 = ( n4296 & ~n6229 ) | ( n4296 & n8709 ) | ( ~n6229 & n8709 ) ;
  assign n29853 = n18976 ^ n10404 ^ n8743 ;
  assign n29854 = n14973 & ~n29853 ;
  assign n29855 = n29854 ^ n20408 ^ 1'b0 ;
  assign n29856 = ~n4273 & n20736 ;
  assign n29857 = n4824 & n29856 ;
  assign n29858 = ~n13033 & n14451 ;
  assign n29859 = n29858 ^ n1266 ^ 1'b0 ;
  assign n29860 = n9890 & ~n27348 ;
  assign n29861 = n1530 & n29860 ;
  assign n29862 = n29861 ^ n4786 ^ 1'b0 ;
  assign n29863 = ~n20646 & n29862 ;
  assign n29864 = ( n5971 & n24315 ) | ( n5971 & n29863 ) | ( n24315 & n29863 ) ;
  assign n29865 = n7846 ^ n5785 ^ n2984 ;
  assign n29866 = ( n11052 & n17330 ) | ( n11052 & n21096 ) | ( n17330 & n21096 ) ;
  assign n29867 = ( n5661 & ~n7224 ) | ( n5661 & n29866 ) | ( ~n7224 & n29866 ) ;
  assign n29868 = ( n6225 & n29865 ) | ( n6225 & n29867 ) | ( n29865 & n29867 ) ;
  assign n29869 = n4200 ^ n1423 ^ 1'b0 ;
  assign n29870 = n9354 & ~n29869 ;
  assign n29871 = ~n6200 & n14845 ;
  assign n29872 = n29871 ^ n10550 ^ 1'b0 ;
  assign n29873 = ( n12848 & ~n28044 ) | ( n12848 & n29872 ) | ( ~n28044 & n29872 ) ;
  assign n29874 = ( n2344 & ~n29870 ) | ( n2344 & n29873 ) | ( ~n29870 & n29873 ) ;
  assign n29875 = n7021 ^ n6283 ^ n1996 ;
  assign n29876 = n7783 & ~n29526 ;
  assign n29877 = ~n1760 & n29876 ;
  assign n29878 = ( n23152 & ~n29875 ) | ( n23152 & n29877 ) | ( ~n29875 & n29877 ) ;
  assign n29879 = n11181 ^ n5207 ^ n2103 ;
  assign n29880 = n29879 ^ n24500 ^ n9985 ;
  assign n29881 = ( n5217 & n5642 ) | ( n5217 & ~n29880 ) | ( n5642 & ~n29880 ) ;
  assign n29882 = n21224 ^ n1936 ^ n538 ;
  assign n29883 = n26533 ^ n20179 ^ n1350 ;
  assign n29885 = ( n5413 & ~n16195 ) | ( n5413 & n18730 ) | ( ~n16195 & n18730 ) ;
  assign n29886 = n1869 | n10738 ;
  assign n29887 = n29885 | n29886 ;
  assign n29884 = ( n1182 & ~n3294 ) | ( n1182 & n11071 ) | ( ~n3294 & n11071 ) ;
  assign n29888 = n29887 ^ n29884 ^ n8338 ;
  assign n29889 = n26843 ^ n23307 ^ n14777 ;
  assign n29890 = n16677 ^ n13988 ^ 1'b0 ;
  assign n29891 = ~n29889 & n29890 ;
  assign n29892 = n21368 ^ n7451 ^ 1'b0 ;
  assign n29893 = n21244 ^ n7546 ^ 1'b0 ;
  assign n29894 = n29892 & ~n29893 ;
  assign n29895 = n27179 ^ n18155 ^ n16917 ;
  assign n29896 = n5407 ^ n1733 ^ 1'b0 ;
  assign n29897 = ( n9254 & n19410 ) | ( n9254 & n29896 ) | ( n19410 & n29896 ) ;
  assign n29898 = ( n3026 & ~n20647 ) | ( n3026 & n20987 ) | ( ~n20647 & n20987 ) ;
  assign n29899 = ( n961 & n13600 ) | ( n961 & n29898 ) | ( n13600 & n29898 ) ;
  assign n29900 = n24824 ^ n20067 ^ n10329 ;
  assign n29901 = ( ~n7894 & n29805 ) | ( ~n7894 & n29900 ) | ( n29805 & n29900 ) ;
  assign n29902 = n15675 ^ n12290 ^ 1'b0 ;
  assign n29903 = ( ~n178 & n12263 ) | ( ~n178 & n29902 ) | ( n12263 & n29902 ) ;
  assign n29904 = ( ~n4108 & n15409 ) | ( ~n4108 & n29903 ) | ( n15409 & n29903 ) ;
  assign n29905 = n18866 ^ n14848 ^ n7007 ;
  assign n29906 = ( ~n4381 & n8264 ) | ( ~n4381 & n9935 ) | ( n8264 & n9935 ) ;
  assign n29907 = n9850 ^ n1473 ^ 1'b0 ;
  assign n29908 = n27099 ^ n21778 ^ n10446 ;
  assign n29909 = ( n7620 & n8632 ) | ( n7620 & ~n22607 ) | ( n8632 & ~n22607 ) ;
  assign n29910 = ( n717 & ~n10023 ) | ( n717 & n11113 ) | ( ~n10023 & n11113 ) ;
  assign n29911 = n23324 ^ n9351 ^ n3619 ;
  assign n29914 = n13800 ^ n3062 ^ n1588 ;
  assign n29912 = n5031 | n6647 ;
  assign n29913 = n13058 | n29912 ;
  assign n29915 = n29914 ^ n29913 ^ n15078 ;
  assign n29916 = n1797 | n4642 ;
  assign n29917 = ( ~n9466 & n20712 ) | ( ~n9466 & n29916 ) | ( n20712 & n29916 ) ;
  assign n29918 = n29917 ^ n18400 ^ 1'b0 ;
  assign n29919 = n29918 ^ n13143 ^ n4930 ;
  assign n29920 = n3262 & n17094 ;
  assign n29921 = n29920 ^ n5024 ^ 1'b0 ;
  assign n29922 = n6813 & ~n29921 ;
  assign n29923 = n9949 & n26718 ;
  assign n29924 = ~n305 & n29923 ;
  assign n29925 = n27129 ^ n21611 ^ 1'b0 ;
  assign n29926 = ~n12217 & n29925 ;
  assign n29927 = n17005 ^ n6697 ^ 1'b0 ;
  assign n29928 = ( n11140 & ~n25311 ) | ( n11140 & n29927 ) | ( ~n25311 & n29927 ) ;
  assign n29929 = ( n3140 & n20625 ) | ( n3140 & n29928 ) | ( n20625 & n29928 ) ;
  assign n29930 = n7908 & n16651 ;
  assign n29931 = ( n22250 & n27515 ) | ( n22250 & ~n29930 ) | ( n27515 & ~n29930 ) ;
  assign n29932 = ( n1139 & ~n11853 ) | ( n1139 & n29931 ) | ( ~n11853 & n29931 ) ;
  assign n29933 = ( x52 & n3299 ) | ( x52 & ~n7950 ) | ( n3299 & ~n7950 ) ;
  assign n29934 = ( n648 & n14568 ) | ( n648 & ~n26844 ) | ( n14568 & ~n26844 ) ;
  assign n29935 = ( n6759 & n13102 ) | ( n6759 & ~n20087 ) | ( n13102 & ~n20087 ) ;
  assign n29936 = n29935 ^ n13924 ^ n9191 ;
  assign n29937 = n24841 ^ n13731 ^ n6963 ;
  assign n29938 = ( ~n15348 & n29936 ) | ( ~n15348 & n29937 ) | ( n29936 & n29937 ) ;
  assign n29939 = n9359 ^ n4323 ^ 1'b0 ;
  assign n29940 = n29939 ^ n20326 ^ n9637 ;
  assign n29941 = ( n16215 & ~n29681 ) | ( n16215 & n29940 ) | ( ~n29681 & n29940 ) ;
  assign n29942 = n10878 ^ n1045 ^ x26 ;
  assign n29943 = ~n21062 & n29942 ;
  assign n29944 = n29943 ^ n26000 ^ 1'b0 ;
  assign n29945 = n27492 ^ n3190 ^ 1'b0 ;
  assign n29946 = n7930 | n21114 ;
  assign n29947 = n29946 ^ n23960 ^ 1'b0 ;
  assign n29948 = ( n9552 & ~n14381 ) | ( n9552 & n24423 ) | ( ~n14381 & n24423 ) ;
  assign n29949 = ( x29 & ~n1884 ) | ( x29 & n29948 ) | ( ~n1884 & n29948 ) ;
  assign n29950 = ( n8265 & ~n20173 ) | ( n8265 & n24942 ) | ( ~n20173 & n24942 ) ;
  assign n29951 = n7816 ^ n6337 ^ n3769 ;
  assign n29952 = n29950 | n29951 ;
  assign n29953 = n7773 | n29952 ;
  assign n29956 = n26863 ^ n8447 ^ n3480 ;
  assign n29954 = n12208 & ~n15381 ;
  assign n29955 = n15671 & n29954 ;
  assign n29957 = n29956 ^ n29955 ^ n22585 ;
  assign n29964 = n11649 ^ n3737 ^ 1'b0 ;
  assign n29958 = n25189 ^ n22452 ^ n616 ;
  assign n29959 = n29958 ^ n9288 ^ n1930 ;
  assign n29960 = ( x71 & n9496 ) | ( x71 & ~n26153 ) | ( n9496 & ~n26153 ) ;
  assign n29961 = n1395 & ~n28338 ;
  assign n29962 = ~n2232 & n29961 ;
  assign n29963 = ( n29959 & n29960 ) | ( n29959 & n29962 ) | ( n29960 & n29962 ) ;
  assign n29965 = n29964 ^ n29963 ^ n16067 ;
  assign n29966 = n12455 ^ n4882 ^ 1'b0 ;
  assign n29967 = ~n12428 & n29966 ;
  assign n29968 = n29967 ^ n9588 ^ 1'b0 ;
  assign n29969 = n29968 ^ n25433 ^ n2530 ;
  assign n29970 = n29969 ^ n4021 ^ 1'b0 ;
  assign n29971 = n21748 & ~n29970 ;
  assign n29972 = ( n7290 & n29965 ) | ( n7290 & ~n29971 ) | ( n29965 & ~n29971 ) ;
  assign n29973 = n24442 & n28797 ;
  assign n29974 = ( n4207 & n9384 ) | ( n4207 & n10802 ) | ( n9384 & n10802 ) ;
  assign n29975 = ( n2417 & n17007 ) | ( n2417 & ~n29974 ) | ( n17007 & ~n29974 ) ;
  assign n29976 = n14989 ^ n8287 ^ n2492 ;
  assign n29977 = ( n2624 & n15121 ) | ( n2624 & ~n29976 ) | ( n15121 & ~n29976 ) ;
  assign n29979 = n2100 | n10052 ;
  assign n29980 = n29979 ^ n11877 ^ 1'b0 ;
  assign n29978 = ( ~n10185 & n24930 ) | ( ~n10185 & n25909 ) | ( n24930 & n25909 ) ;
  assign n29981 = n29980 ^ n29978 ^ n6967 ;
  assign n29982 = n12289 & ~n20176 ;
  assign n29983 = n29982 ^ n18022 ^ 1'b0 ;
  assign n29984 = n23703 ^ n7976 ^ 1'b0 ;
  assign n29985 = n25532 & ~n29984 ;
  assign n29986 = ~n10396 & n19248 ;
  assign n29987 = n28533 ^ n12393 ^ n8435 ;
  assign n29988 = n29987 ^ n20409 ^ n277 ;
  assign n29989 = n11596 & ~n19857 ;
  assign n29990 = n29989 ^ n26409 ^ n1978 ;
  assign n29991 = ( n1572 & n14300 ) | ( n1572 & n27156 ) | ( n14300 & n27156 ) ;
  assign n29992 = ( n6454 & ~n13199 ) | ( n6454 & n17121 ) | ( ~n13199 & n17121 ) ;
  assign n29993 = ( x126 & ~n4924 ) | ( x126 & n9752 ) | ( ~n4924 & n9752 ) ;
  assign n29994 = ( ~n1206 & n29992 ) | ( ~n1206 & n29993 ) | ( n29992 & n29993 ) ;
  assign n29995 = ( n1493 & ~n9202 ) | ( n1493 & n29994 ) | ( ~n9202 & n29994 ) ;
  assign n29996 = ( n2286 & ~n29991 ) | ( n2286 & n29995 ) | ( ~n29991 & n29995 ) ;
  assign n29997 = ( ~n11645 & n20118 ) | ( ~n11645 & n21036 ) | ( n20118 & n21036 ) ;
  assign n29998 = n7240 ^ n3820 ^ 1'b0 ;
  assign n29999 = n7819 & n29998 ;
  assign n30000 = n29999 ^ n17218 ^ n14138 ;
  assign n30001 = n1462 & n12438 ;
  assign n30002 = ~n17452 & n30001 ;
  assign n30003 = n30002 ^ n28934 ^ n16531 ;
  assign n30004 = ( ~n484 & n11491 ) | ( ~n484 & n29653 ) | ( n11491 & n29653 ) ;
  assign n30005 = n30004 ^ n6395 ^ 1'b0 ;
  assign n30006 = n4690 | n30005 ;
  assign n30007 = n2064 ^ n1549 ^ n1326 ;
  assign n30008 = n30007 ^ n29183 ^ n11900 ;
  assign n30009 = n14829 ^ n7371 ^ n3107 ;
  assign n30010 = n30009 ^ n24066 ^ n13480 ;
  assign n30011 = ( n6417 & n30008 ) | ( n6417 & ~n30010 ) | ( n30008 & ~n30010 ) ;
  assign n30012 = n13617 & ~n24634 ;
  assign n30013 = n29424 ^ n25458 ^ n13347 ;
  assign n30014 = ( n6462 & n13388 ) | ( n6462 & ~n19683 ) | ( n13388 & ~n19683 ) ;
  assign n30015 = ( n20887 & n27412 ) | ( n20887 & ~n30014 ) | ( n27412 & ~n30014 ) ;
  assign n30016 = ( n10597 & n11328 ) | ( n10597 & ~n30015 ) | ( n11328 & ~n30015 ) ;
  assign n30017 = ( n4432 & ~n24349 ) | ( n4432 & n30016 ) | ( ~n24349 & n30016 ) ;
  assign n30022 = n11728 & ~n12085 ;
  assign n30023 = ( n11194 & n14906 ) | ( n11194 & n30022 ) | ( n14906 & n30022 ) ;
  assign n30019 = n21077 ^ n1456 ^ 1'b0 ;
  assign n30018 = ~n3759 & n13832 ;
  assign n30020 = n30019 ^ n30018 ^ 1'b0 ;
  assign n30021 = n30020 ^ n15013 ^ n4302 ;
  assign n30024 = n30023 ^ n30021 ^ n21000 ;
  assign n30025 = ( n902 & ~n9626 ) | ( n902 & n18058 ) | ( ~n9626 & n18058 ) ;
  assign n30026 = ( n1621 & n12110 ) | ( n1621 & n23846 ) | ( n12110 & n23846 ) ;
  assign n30027 = ( n29853 & n30025 ) | ( n29853 & n30026 ) | ( n30025 & n30026 ) ;
  assign n30028 = ( n9297 & n19825 ) | ( n9297 & n30027 ) | ( n19825 & n30027 ) ;
  assign n30029 = n10158 & n20136 ;
  assign n30030 = n30029 ^ n9222 ^ n8410 ;
  assign n30031 = n16853 & n29733 ;
  assign n30032 = ~n21641 & n30031 ;
  assign n30033 = ( n2850 & n5656 ) | ( n2850 & ~n9685 ) | ( n5656 & ~n9685 ) ;
  assign n30034 = ( n6255 & n23919 ) | ( n6255 & ~n30033 ) | ( n23919 & ~n30033 ) ;
  assign n30035 = ( n11975 & ~n30032 ) | ( n11975 & n30034 ) | ( ~n30032 & n30034 ) ;
  assign n30036 = ~n974 & n30035 ;
  assign n30037 = n30036 ^ n16364 ^ 1'b0 ;
  assign n30038 = n22469 & n29032 ;
  assign n30039 = n8255 & n30038 ;
  assign n30040 = n16120 | n16467 ;
  assign n30041 = n30040 ^ n19408 ^ 1'b0 ;
  assign n30042 = ( n8220 & n10125 ) | ( n8220 & n19517 ) | ( n10125 & n19517 ) ;
  assign n30043 = n17409 ^ n13581 ^ n1230 ;
  assign n30044 = n30043 ^ n24476 ^ n7873 ;
  assign n30045 = ( n2640 & n15592 ) | ( n2640 & n29279 ) | ( n15592 & n29279 ) ;
  assign n30046 = ( n1049 & n3424 ) | ( n1049 & n11935 ) | ( n3424 & n11935 ) ;
  assign n30047 = ( n2036 & n3397 ) | ( n2036 & n4350 ) | ( n3397 & n4350 ) ;
  assign n30048 = ( n1652 & n18023 ) | ( n1652 & n30047 ) | ( n18023 & n30047 ) ;
  assign n30049 = ( n3268 & n11616 ) | ( n3268 & ~n28410 ) | ( n11616 & ~n28410 ) ;
  assign n30050 = ( n4651 & n21129 ) | ( n4651 & ~n30049 ) | ( n21129 & ~n30049 ) ;
  assign n30051 = n27716 ^ n15708 ^ n11694 ;
  assign n30052 = n3840 & ~n8313 ;
  assign n30053 = ( ~n5921 & n16527 ) | ( ~n5921 & n27228 ) | ( n16527 & n27228 ) ;
  assign n30054 = ( n12866 & n18126 ) | ( n12866 & ~n30053 ) | ( n18126 & ~n30053 ) ;
  assign n30055 = n6543 | n30054 ;
  assign n30056 = n30055 ^ n13428 ^ 1'b0 ;
  assign n30057 = ~n1215 & n16364 ;
  assign n30058 = n30057 ^ n27784 ^ 1'b0 ;
  assign n30059 = n25077 ^ n24432 ^ n21539 ;
  assign n30060 = n4667 ^ n3538 ^ n1405 ;
  assign n30061 = n19121 ^ n4696 ^ 1'b0 ;
  assign n30062 = ( ~n7054 & n30060 ) | ( ~n7054 & n30061 ) | ( n30060 & n30061 ) ;
  assign n30063 = n8870 ^ n367 ^ x39 ;
  assign n30064 = n29285 & n30063 ;
  assign n30065 = ( n12040 & ~n30008 ) | ( n12040 & n30064 ) | ( ~n30008 & n30064 ) ;
  assign n30066 = ( n2766 & n10525 ) | ( n2766 & n26748 ) | ( n10525 & n26748 ) ;
  assign n30067 = n30066 ^ n7931 ^ n4023 ;
  assign n30068 = n2455 & ~n5718 ;
  assign n30069 = n30068 ^ n3175 ^ 1'b0 ;
  assign n30070 = n18438 ^ n12223 ^ n561 ;
  assign n30071 = ( n28718 & ~n30069 ) | ( n28718 & n30070 ) | ( ~n30069 & n30070 ) ;
  assign n30072 = ( ~n7917 & n11510 ) | ( ~n7917 & n27784 ) | ( n11510 & n27784 ) ;
  assign n30073 = n16261 & n18106 ;
  assign n30074 = ( n9415 & n14098 ) | ( n9415 & n30073 ) | ( n14098 & n30073 ) ;
  assign n30075 = ~n30072 & n30074 ;
  assign n30076 = n11264 & n15266 ;
  assign n30077 = n30076 ^ n7261 ^ 1'b0 ;
  assign n30078 = n30077 ^ n23335 ^ n4890 ;
  assign n30079 = n30078 ^ n14250 ^ 1'b0 ;
  assign n30080 = ~n27179 & n30079 ;
  assign n30081 = ( n16283 & n18390 ) | ( n16283 & n26328 ) | ( n18390 & n26328 ) ;
  assign n30082 = n30081 ^ n10463 ^ n3157 ;
  assign n30083 = ( n450 & n9733 ) | ( n450 & n30082 ) | ( n9733 & n30082 ) ;
  assign n30084 = ( n8063 & n10333 ) | ( n8063 & n30083 ) | ( n10333 & n30083 ) ;
  assign n30085 = n18452 ^ n6427 ^ 1'b0 ;
  assign n30086 = ( n4211 & n10239 ) | ( n4211 & ~n22712 ) | ( n10239 & ~n22712 ) ;
  assign n30087 = ( ~n12196 & n17740 ) | ( ~n12196 & n18440 ) | ( n17740 & n18440 ) ;
  assign n30088 = n30087 ^ n24984 ^ n2754 ;
  assign n30090 = n1460 & ~n13659 ;
  assign n30091 = ~n2085 & n30090 ;
  assign n30089 = ( n1045 & ~n9511 ) | ( n1045 & n19162 ) | ( ~n9511 & n19162 ) ;
  assign n30092 = n30091 ^ n30089 ^ 1'b0 ;
  assign n30093 = ( n4553 & n13275 ) | ( n4553 & ~n25905 ) | ( n13275 & ~n25905 ) ;
  assign n30094 = ( n22508 & n28536 ) | ( n22508 & n30093 ) | ( n28536 & n30093 ) ;
  assign n30095 = ( ~n2276 & n2395 ) | ( ~n2276 & n25077 ) | ( n2395 & n25077 ) ;
  assign n30096 = n9783 & ~n20829 ;
  assign n30097 = n30096 ^ n10610 ^ n7353 ;
  assign n30098 = ( ~n2331 & n30095 ) | ( ~n2331 & n30097 ) | ( n30095 & n30097 ) ;
  assign n30099 = ( n7792 & n24244 ) | ( n7792 & ~n30098 ) | ( n24244 & ~n30098 ) ;
  assign n30100 = n26067 ^ n4299 ^ n3990 ;
  assign n30101 = ( n5822 & n21854 ) | ( n5822 & ~n24146 ) | ( n21854 & ~n24146 ) ;
  assign n30102 = n4432 & ~n30101 ;
  assign n30103 = n30102 ^ n5429 ^ 1'b0 ;
  assign n30104 = n12184 & ~n19459 ;
  assign n30105 = n25393 ^ n12727 ^ 1'b0 ;
  assign n30106 = ~n9195 & n30105 ;
  assign n30108 = ( n1570 & n2147 ) | ( n1570 & ~n26920 ) | ( n2147 & ~n26920 ) ;
  assign n30109 = n17716 ^ n9339 ^ 1'b0 ;
  assign n30110 = n30108 | n30109 ;
  assign n30111 = n30110 ^ n29408 ^ n5972 ;
  assign n30107 = n27367 ^ n3835 ^ n1601 ;
  assign n30112 = n30111 ^ n30107 ^ 1'b0 ;
  assign n30113 = n13808 | n15146 ;
  assign n30114 = ( n4739 & ~n16369 ) | ( n4739 & n30113 ) | ( ~n16369 & n30113 ) ;
  assign n30115 = n24452 ^ n11578 ^ n10221 ;
  assign n30116 = ( n16719 & n22053 ) | ( n16719 & ~n30115 ) | ( n22053 & ~n30115 ) ;
  assign n30117 = ( n4843 & n13927 ) | ( n4843 & n29031 ) | ( n13927 & n29031 ) ;
  assign n30118 = n3773 & ~n4522 ;
  assign n30119 = ~n3142 & n30118 ;
  assign n30120 = n30119 ^ n8618 ^ n1467 ;
  assign n30121 = n17085 ^ n3927 ^ n886 ;
  assign n30122 = n14617 ^ n12970 ^ n2816 ;
  assign n30123 = n4252 ^ n2916 ^ n2089 ;
  assign n30124 = n11611 ^ n6685 ^ 1'b0 ;
  assign n30125 = ~n30123 & n30124 ;
  assign n30126 = n15126 ^ n2183 ^ 1'b0 ;
  assign n30127 = n30125 & ~n30126 ;
  assign n30128 = n1737 | n7024 ;
  assign n30129 = n11925 | n20080 ;
  assign n30130 = n22331 ^ n20202 ^ 1'b0 ;
  assign n30131 = n18185 ^ n18103 ^ 1'b0 ;
  assign n30132 = ( n3403 & ~n27237 ) | ( n3403 & n30131 ) | ( ~n27237 & n30131 ) ;
  assign n30133 = ( n1344 & n27010 ) | ( n1344 & n30132 ) | ( n27010 & n30132 ) ;
  assign n30140 = n402 & n2907 ;
  assign n30141 = n30140 ^ n7151 ^ 1'b0 ;
  assign n30142 = n30141 ^ n29093 ^ n1610 ;
  assign n30143 = ( n6216 & n16258 ) | ( n6216 & n30142 ) | ( n16258 & n30142 ) ;
  assign n30144 = ( n18018 & n24441 ) | ( n18018 & ~n30143 ) | ( n24441 & ~n30143 ) ;
  assign n30138 = n10378 ^ n3503 ^ 1'b0 ;
  assign n30134 = n7276 ^ n6715 ^ n3294 ;
  assign n30135 = n30134 ^ n14044 ^ n753 ;
  assign n30136 = n30135 ^ n23554 ^ n6293 ;
  assign n30137 = n22269 & n30136 ;
  assign n30139 = n30138 ^ n30137 ^ 1'b0 ;
  assign n30145 = n30144 ^ n30139 ^ n19571 ;
  assign n30152 = ( ~n10803 & n24342 ) | ( ~n10803 & n26159 ) | ( n24342 & n26159 ) ;
  assign n30146 = n24276 ^ n5693 ^ n258 ;
  assign n30147 = n3004 ^ n940 ^ n439 ;
  assign n30148 = n30147 ^ n11589 ^ n3915 ;
  assign n30149 = n30148 ^ n12355 ^ n1539 ;
  assign n30150 = n30149 ^ n9587 ^ n1864 ;
  assign n30151 = ( n13350 & n30146 ) | ( n13350 & ~n30150 ) | ( n30146 & ~n30150 ) ;
  assign n30153 = n30152 ^ n30151 ^ n24554 ;
  assign n30154 = n7636 | n18036 ;
  assign n30155 = n30154 ^ n3564 ^ n801 ;
  assign n30156 = ( n14984 & n28627 ) | ( n14984 & ~n30155 ) | ( n28627 & ~n30155 ) ;
  assign n30157 = ( n19177 & ~n19215 ) | ( n19177 & n30156 ) | ( ~n19215 & n30156 ) ;
  assign n30158 = ( n4643 & ~n18097 ) | ( n4643 & n25663 ) | ( ~n18097 & n25663 ) ;
  assign n30159 = ( n13617 & n17318 ) | ( n13617 & ~n29903 ) | ( n17318 & ~n29903 ) ;
  assign n30160 = ( ~n16115 & n21397 ) | ( ~n16115 & n30159 ) | ( n21397 & n30159 ) ;
  assign n30161 = n24149 ^ n23819 ^ n15049 ;
  assign n30162 = ( ~n30158 & n30160 ) | ( ~n30158 & n30161 ) | ( n30160 & n30161 ) ;
  assign n30163 = n17781 ^ n1694 ^ 1'b0 ;
  assign n30164 = n25749 & n30163 ;
  assign n30165 = n3480 & n22059 ;
  assign n30166 = n10563 ^ n7967 ^ n526 ;
  assign n30167 = ( n16711 & ~n19374 ) | ( n16711 & n30166 ) | ( ~n19374 & n30166 ) ;
  assign n30168 = n16672 ^ n5978 ^ n4695 ;
  assign n30169 = n24525 ^ n23896 ^ n11855 ;
  assign n30170 = n13022 ^ n12340 ^ n8429 ;
  assign n30171 = ( n3845 & n18046 ) | ( n3845 & n30170 ) | ( n18046 & n30170 ) ;
  assign n30172 = n12696 ^ n8989 ^ n4248 ;
  assign n30177 = ( ~n2903 & n4376 ) | ( ~n2903 & n17657 ) | ( n4376 & n17657 ) ;
  assign n30178 = n30177 ^ n20614 ^ n3855 ;
  assign n30173 = n19930 ^ n7329 ^ n5306 ;
  assign n30174 = n7112 & n23364 ;
  assign n30175 = n30174 ^ n14966 ^ n4098 ;
  assign n30176 = ( n14454 & n30173 ) | ( n14454 & n30175 ) | ( n30173 & n30175 ) ;
  assign n30179 = n30178 ^ n30176 ^ 1'b0 ;
  assign n30180 = ( n5774 & n14687 ) | ( n5774 & n23097 ) | ( n14687 & n23097 ) ;
  assign n30181 = ~n299 & n3362 ;
  assign n30182 = n30181 ^ n22837 ^ n15058 ;
  assign n30183 = n19937 ^ n10367 ^ 1'b0 ;
  assign n30184 = n10145 & ~n30183 ;
  assign n30185 = n30184 ^ n4291 ^ 1'b0 ;
  assign n30186 = n30182 | n30185 ;
  assign n30187 = n30186 ^ n5827 ^ 1'b0 ;
  assign n30188 = n3365 & n30187 ;
  assign n30189 = n30180 & n30188 ;
  assign n30190 = n25598 ^ n7654 ^ n3877 ;
  assign n30191 = n23700 & ~n30190 ;
  assign n30192 = ~n27662 & n30191 ;
  assign n30193 = n2313 ^ n849 ^ n337 ;
  assign n30194 = ~n10569 & n30193 ;
  assign n30195 = ( n6966 & ~n13553 ) | ( n6966 & n18610 ) | ( ~n13553 & n18610 ) ;
  assign n30196 = n22133 & n30195 ;
  assign n30197 = ~n30194 & n30196 ;
  assign n30198 = n12775 ^ n8998 ^ 1'b0 ;
  assign n30199 = n19146 & n30198 ;
  assign n30200 = n30199 ^ n14125 ^ x6 ;
  assign n30201 = n3349 & ~n10122 ;
  assign n30202 = ~n30200 & n30201 ;
  assign n30203 = ( n11905 & n13950 ) | ( n11905 & n14218 ) | ( n13950 & n14218 ) ;
  assign n30204 = n30203 ^ n26170 ^ n6855 ;
  assign n30205 = n28548 ^ n8775 ^ n7154 ;
  assign n30206 = ( ~n1810 & n4813 ) | ( ~n1810 & n17675 ) | ( n4813 & n17675 ) ;
  assign n30207 = n14018 & ~n20797 ;
  assign n30208 = n30207 ^ n2309 ^ 1'b0 ;
  assign n30209 = ( n1384 & n27849 ) | ( n1384 & ~n30208 ) | ( n27849 & ~n30208 ) ;
  assign n30215 = n23491 ^ n22185 ^ n8573 ;
  assign n30216 = ( ~n1452 & n19936 ) | ( ~n1452 & n30215 ) | ( n19936 & n30215 ) ;
  assign n30210 = ( n3726 & n7322 ) | ( n3726 & ~n9170 ) | ( n7322 & ~n9170 ) ;
  assign n30211 = ( n5837 & ~n7513 ) | ( n5837 & n8041 ) | ( ~n7513 & n8041 ) ;
  assign n30212 = ~n14245 & n30211 ;
  assign n30213 = n5451 & n30212 ;
  assign n30214 = n30210 & ~n30213 ;
  assign n30217 = n30216 ^ n30214 ^ n27980 ;
  assign n30218 = n8392 ^ n6583 ^ n3085 ;
  assign n30219 = n30218 ^ n21959 ^ n214 ;
  assign n30220 = ( n3614 & n7174 ) | ( n3614 & ~n8087 ) | ( n7174 & ~n8087 ) ;
  assign n30221 = ( ~n4780 & n21733 ) | ( ~n4780 & n30220 ) | ( n21733 & n30220 ) ;
  assign n30222 = n30221 ^ n3750 ^ 1'b0 ;
  assign n30223 = n27750 | n29454 ;
  assign n30224 = n9395 | n30223 ;
  assign n30225 = n29138 ^ n16558 ^ n8803 ;
  assign n30226 = n15466 & n30225 ;
  assign n30227 = n11335 & n30226 ;
  assign n30228 = ( n5783 & n11624 ) | ( n5783 & ~n27239 ) | ( n11624 & ~n27239 ) ;
  assign n30229 = n30228 ^ n6737 ^ 1'b0 ;
  assign n30230 = n10322 ^ n8969 ^ n3316 ;
  assign n30231 = n6747 ^ n4693 ^ n918 ;
  assign n30232 = ( ~n12301 & n16187 ) | ( ~n12301 & n26651 ) | ( n16187 & n26651 ) ;
  assign n30233 = ( ~n1167 & n2699 ) | ( ~n1167 & n10454 ) | ( n2699 & n10454 ) ;
  assign n30234 = ( n5344 & ~n7428 ) | ( n5344 & n30233 ) | ( ~n7428 & n30233 ) ;
  assign n30235 = ( n8130 & ~n23519 ) | ( n8130 & n28900 ) | ( ~n23519 & n28900 ) ;
  assign n30236 = ( n5036 & n16813 ) | ( n5036 & n28248 ) | ( n16813 & n28248 ) ;
  assign n30237 = ( ~n3126 & n14848 ) | ( ~n3126 & n26685 ) | ( n14848 & n26685 ) ;
  assign n30238 = n906 & ~n28094 ;
  assign n30239 = ~n26821 & n30238 ;
  assign n30240 = n8630 ^ n6687 ^ n6529 ;
  assign n30241 = n10250 ^ n5112 ^ n1220 ;
  assign n30242 = n30241 ^ n17080 ^ n3829 ;
  assign n30243 = ( n11761 & n17242 ) | ( n11761 & n30242 ) | ( n17242 & n30242 ) ;
  assign n30244 = n4289 ^ n1740 ^ 1'b0 ;
  assign n30245 = n8388 | n30244 ;
  assign n30246 = n6416 | n19635 ;
  assign n30247 = ( n21750 & n23195 ) | ( n21750 & n30246 ) | ( n23195 & n30246 ) ;
  assign n30248 = n30245 | n30247 ;
  assign n30249 = n30248 ^ n6085 ^ 1'b0 ;
  assign n30250 = n29266 ^ n28318 ^ n18411 ;
  assign n30251 = ( n3015 & n13672 ) | ( n3015 & ~n24042 ) | ( n13672 & ~n24042 ) ;
  assign n30252 = ( n1990 & ~n5452 ) | ( n1990 & n19407 ) | ( ~n5452 & n19407 ) ;
  assign n30253 = ( n1412 & n6409 ) | ( n1412 & n13054 ) | ( n6409 & n13054 ) ;
  assign n30254 = n28007 ^ n21471 ^ n2769 ;
  assign n30255 = ( n18823 & n24699 ) | ( n18823 & n30254 ) | ( n24699 & n30254 ) ;
  assign n30256 = n10023 | n26527 ;
  assign n30257 = n30256 ^ n25439 ^ 1'b0 ;
  assign n30258 = n16886 ^ n10516 ^ n7417 ;
  assign n30259 = ( n1803 & n8907 ) | ( n1803 & n18831 ) | ( n8907 & n18831 ) ;
  assign n30260 = ( ~n21170 & n28970 ) | ( ~n21170 & n30259 ) | ( n28970 & n30259 ) ;
  assign n30261 = n28648 ^ n15182 ^ n633 ;
  assign n30262 = n30261 ^ n28727 ^ n4544 ;
  assign n30263 = n30262 ^ n2570 ^ n959 ;
  assign n30264 = ( n5876 & n27578 ) | ( n5876 & n29861 ) | ( n27578 & n29861 ) ;
  assign n30265 = ( n5950 & n12821 ) | ( n5950 & ~n21370 ) | ( n12821 & ~n21370 ) ;
  assign n30266 = ~n21330 & n26969 ;
  assign n30267 = n6987 ^ n1750 ^ n1664 ;
  assign n30268 = ~n8123 & n15886 ;
  assign n30269 = n30268 ^ n15776 ^ n11382 ;
  assign n30270 = ( n24072 & n30267 ) | ( n24072 & ~n30269 ) | ( n30267 & ~n30269 ) ;
  assign n30271 = ( n2818 & ~n10920 ) | ( n2818 & n30270 ) | ( ~n10920 & n30270 ) ;
  assign n30272 = ( n2131 & n2412 ) | ( n2131 & n4185 ) | ( n2412 & n4185 ) ;
  assign n30273 = n8159 ^ x110 ^ 1'b0 ;
  assign n30274 = n30272 & ~n30273 ;
  assign n30275 = ~n17441 & n22916 ;
  assign n30276 = n30275 ^ n5693 ^ 1'b0 ;
  assign n30277 = n22137 ^ n11342 ^ n3184 ;
  assign n30278 = n30277 ^ n3493 ^ 1'b0 ;
  assign n30285 = ( n2613 & n5015 ) | ( n2613 & n10904 ) | ( n5015 & n10904 ) ;
  assign n30286 = n30285 ^ n582 ^ 1'b0 ;
  assign n30287 = ( n8256 & n18416 ) | ( n8256 & n30286 ) | ( n18416 & n30286 ) ;
  assign n30283 = ( n14807 & n15997 ) | ( n14807 & n17505 ) | ( n15997 & n17505 ) ;
  assign n30284 = ( n9121 & ~n17775 ) | ( n9121 & n30283 ) | ( ~n17775 & n30283 ) ;
  assign n30279 = n20510 ^ n8848 ^ n790 ;
  assign n30280 = ( n7897 & n16340 ) | ( n7897 & ~n30279 ) | ( n16340 & ~n30279 ) ;
  assign n30281 = n30280 ^ n6713 ^ 1'b0 ;
  assign n30282 = n4144 & ~n30281 ;
  assign n30288 = n30287 ^ n30284 ^ n30282 ;
  assign n30289 = n14820 ^ n8205 ^ n5915 ;
  assign n30290 = n13128 ^ n1477 ^ 1'b0 ;
  assign n30291 = n8570 | n30290 ;
  assign n30292 = ( n14820 & n30289 ) | ( n14820 & ~n30291 ) | ( n30289 & ~n30291 ) ;
  assign n30293 = n30292 ^ n4332 ^ n2620 ;
  assign n30294 = n28785 | n30293 ;
  assign n30296 = n12205 ^ n2727 ^ 1'b0 ;
  assign n30295 = ( n6087 & n15572 ) | ( n6087 & n20698 ) | ( n15572 & n20698 ) ;
  assign n30297 = n30296 ^ n30295 ^ x45 ;
  assign n30298 = n23276 ^ n14615 ^ n457 ;
  assign n30299 = ( n2544 & ~n16726 ) | ( n2544 & n25077 ) | ( ~n16726 & n25077 ) ;
  assign n30300 = ~n18628 & n29401 ;
  assign n30301 = ( n8658 & ~n23414 ) | ( n8658 & n30300 ) | ( ~n23414 & n30300 ) ;
  assign n30302 = n3191 & n18491 ;
  assign n30303 = ( n577 & ~n20057 ) | ( n577 & n30302 ) | ( ~n20057 & n30302 ) ;
  assign n30304 = n22331 ^ n11687 ^ 1'b0 ;
  assign n30305 = n440 & n30304 ;
  assign n30306 = n15009 ^ n7831 ^ 1'b0 ;
  assign n30307 = n21470 & n30306 ;
  assign n30308 = n21118 ^ n5761 ^ n4751 ;
  assign n30309 = n30308 ^ n20931 ^ n4668 ;
  assign n30310 = n20808 & ~n30309 ;
  assign n30311 = n585 & n30310 ;
  assign n30312 = ( n977 & n27087 ) | ( n977 & ~n28707 ) | ( n27087 & ~n28707 ) ;
  assign n30315 = n27154 ^ n14679 ^ n13058 ;
  assign n30316 = ( ~n2898 & n9686 ) | ( ~n2898 & n30315 ) | ( n9686 & n30315 ) ;
  assign n30314 = n7057 ^ n2890 ^ 1'b0 ;
  assign n30313 = n10623 ^ n551 ^ 1'b0 ;
  assign n30317 = n30316 ^ n30314 ^ n30313 ;
  assign n30318 = n23559 ^ n23335 ^ n8577 ;
  assign n30319 = n25342 ^ n16827 ^ n3570 ;
  assign n30320 = n30319 ^ n27063 ^ 1'b0 ;
  assign n30321 = ( n14232 & n16909 ) | ( n14232 & n30320 ) | ( n16909 & n30320 ) ;
  assign n30322 = n20359 & ~n27154 ;
  assign n30323 = n15332 ^ n5047 ^ n149 ;
  assign n30326 = n510 & ~n3537 ;
  assign n30327 = n30326 ^ n22667 ^ 1'b0 ;
  assign n30324 = n18689 ^ n8000 ^ n3613 ;
  assign n30325 = n24145 & ~n30324 ;
  assign n30328 = n30327 ^ n30325 ^ n10748 ;
  assign n30329 = n30125 ^ n6812 ^ n2825 ;
  assign n30330 = n26639 ^ n24636 ^ n5452 ;
  assign n30331 = n7468 & ~n30330 ;
  assign n30332 = n11077 ^ n9198 ^ 1'b0 ;
  assign n30333 = ~n7329 & n30332 ;
  assign n30334 = ~n414 & n30333 ;
  assign n30335 = n30334 ^ n18776 ^ 1'b0 ;
  assign n30336 = ~n5901 & n20899 ;
  assign n30337 = ~n24399 & n30336 ;
  assign n30338 = ( n15543 & ~n27332 ) | ( n15543 & n30337 ) | ( ~n27332 & n30337 ) ;
  assign n30339 = n17406 ^ n15450 ^ n11417 ;
  assign n30342 = n5989 ^ n3593 ^ n2165 ;
  assign n30340 = n20769 ^ n3271 ^ n2335 ;
  assign n30341 = n30340 ^ n11985 ^ n9943 ;
  assign n30343 = n30342 ^ n30341 ^ n23221 ;
  assign n30344 = n12310 ^ n12296 ^ n6529 ;
  assign n30345 = ~n8831 & n20555 ;
  assign n30346 = n30345 ^ n2331 ^ 1'b0 ;
  assign n30347 = ( ~n12029 & n30344 ) | ( ~n12029 & n30346 ) | ( n30344 & n30346 ) ;
  assign n30348 = n30347 ^ n2794 ^ n438 ;
  assign n30349 = n12267 ^ n7514 ^ n7028 ;
  assign n30350 = ( n4936 & n8109 ) | ( n4936 & ~n15635 ) | ( n8109 & ~n15635 ) ;
  assign n30351 = n30350 ^ n14897 ^ n7668 ;
  assign n30352 = n6920 ^ n6823 ^ n3190 ;
  assign n30353 = ( n2115 & ~n11404 ) | ( n2115 & n13451 ) | ( ~n11404 & n13451 ) ;
  assign n30354 = ( n6649 & n9243 ) | ( n6649 & n30353 ) | ( n9243 & n30353 ) ;
  assign n30355 = n30354 ^ n2818 ^ 1'b0 ;
  assign n30356 = ~n3893 & n30355 ;
  assign n30357 = n15234 & ~n29005 ;
  assign n30358 = n10901 & n30357 ;
  assign n30359 = n30358 ^ n6929 ^ 1'b0 ;
  assign n30360 = n27364 & n30359 ;
  assign n30361 = n16816 ^ n10751 ^ 1'b0 ;
  assign n30362 = n18388 | n30361 ;
  assign n30365 = ( ~n861 & n18396 ) | ( ~n861 & n21364 ) | ( n18396 & n21364 ) ;
  assign n30363 = n25707 ^ n18844 ^ 1'b0 ;
  assign n30364 = ~n12398 & n30363 ;
  assign n30366 = n30365 ^ n30364 ^ n16463 ;
  assign n30367 = n26525 ^ n24101 ^ n4712 ;
  assign n30368 = n30367 ^ n19641 ^ n3160 ;
  assign n30369 = n23728 ^ n13805 ^ n10776 ;
  assign n30372 = ( n10416 & ~n11910 ) | ( n10416 & n23167 ) | ( ~n11910 & n23167 ) ;
  assign n30373 = ( n21738 & n22184 ) | ( n21738 & n30372 ) | ( n22184 & n30372 ) ;
  assign n30370 = n196 & ~n11271 ;
  assign n30371 = n30370 ^ n24712 ^ n2199 ;
  assign n30374 = n30373 ^ n30371 ^ n12150 ;
  assign n30375 = n19926 ^ n18375 ^ n13931 ;
  assign n30376 = n16580 ^ n8640 ^ n5474 ;
  assign n30378 = n15225 ^ n10855 ^ 1'b0 ;
  assign n30377 = ~n17341 & n19880 ;
  assign n30379 = n30378 ^ n30377 ^ 1'b0 ;
  assign n30380 = n27669 ^ n12749 ^ n6386 ;
  assign n30381 = n30380 ^ n27707 ^ 1'b0 ;
  assign n30382 = n23153 | n30381 ;
  assign n30383 = ~n4156 & n9531 ;
  assign n30384 = n30383 ^ n18814 ^ n4700 ;
  assign n30385 = n21069 ^ n10103 ^ 1'b0 ;
  assign n30386 = ~n30384 & n30385 ;
  assign n30387 = n6380 | n8866 ;
  assign n30388 = n30387 ^ n11707 ^ n3110 ;
  assign n30391 = n23424 ^ n19705 ^ n7290 ;
  assign n30389 = n3386 & n8661 ;
  assign n30390 = ( n14012 & n19831 ) | ( n14012 & n30389 ) | ( n19831 & n30389 ) ;
  assign n30392 = n30391 ^ n30390 ^ n30047 ;
  assign n30393 = n30392 ^ n25924 ^ n13144 ;
  assign n30394 = n11861 ^ n6928 ^ n3336 ;
  assign n30395 = x42 & n3299 ;
  assign n30396 = n3458 | n4418 ;
  assign n30397 = n30396 ^ n12616 ^ n1827 ;
  assign n30398 = ( ~n2908 & n9113 ) | ( ~n2908 & n30397 ) | ( n9113 & n30397 ) ;
  assign n30399 = n30398 ^ n26477 ^ n26003 ;
  assign n30400 = ( n30394 & n30395 ) | ( n30394 & n30399 ) | ( n30395 & n30399 ) ;
  assign n30401 = n27255 ^ n15911 ^ n5964 ;
  assign n30402 = n5513 ^ n3451 ^ n2954 ;
  assign n30403 = ( n3152 & ~n11311 ) | ( n3152 & n30402 ) | ( ~n11311 & n30402 ) ;
  assign n30404 = ~n26584 & n30403 ;
  assign n30405 = n15096 ^ n9753 ^ 1'b0 ;
  assign n30406 = ( n10579 & ~n23673 ) | ( n10579 & n30405 ) | ( ~n23673 & n30405 ) ;
  assign n30407 = ~n7625 & n16377 ;
  assign n30408 = n30407 ^ n14561 ^ 1'b0 ;
  assign n30409 = ( n317 & ~n6903 ) | ( n317 & n30408 ) | ( ~n6903 & n30408 ) ;
  assign n30410 = n17102 ^ n10064 ^ 1'b0 ;
  assign n30411 = n26527 | n30410 ;
  assign n30412 = ( n13848 & ~n18838 ) | ( n13848 & n19884 ) | ( ~n18838 & n19884 ) ;
  assign n30413 = n30412 ^ n12239 ^ 1'b0 ;
  assign n30414 = n28643 ^ n10587 ^ n2230 ;
  assign n30415 = n28279 ^ n9620 ^ 1'b0 ;
  assign n30416 = n28260 ^ n18464 ^ 1'b0 ;
  assign n30417 = ( n3100 & n10089 ) | ( n3100 & ~n30416 ) | ( n10089 & ~n30416 ) ;
  assign n30418 = ( n3423 & n14011 ) | ( n3423 & n20126 ) | ( n14011 & n20126 ) ;
  assign n30419 = n21307 ^ n9622 ^ n6426 ;
  assign n30420 = ( n2417 & n11573 ) | ( n2417 & n13650 ) | ( n11573 & n13650 ) ;
  assign n30421 = n165 | n3882 ;
  assign n30422 = n5837 & ~n30421 ;
  assign n30423 = n30422 ^ n14315 ^ n5019 ;
  assign n30424 = n1385 & n5006 ;
  assign n30425 = ~n30423 & n30424 ;
  assign n30426 = n18814 ^ n2949 ^ 1'b0 ;
  assign n30427 = n222 | n30426 ;
  assign n30428 = n17176 ^ n12245 ^ 1'b0 ;
  assign n30429 = n892 & ~n30428 ;
  assign n30430 = ( ~n15152 & n19875 ) | ( ~n15152 & n20890 ) | ( n19875 & n20890 ) ;
  assign n30431 = ( n1109 & ~n7622 ) | ( n1109 & n30430 ) | ( ~n7622 & n30430 ) ;
  assign n30432 = n4221 | n9325 ;
  assign n30433 = n30431 | n30432 ;
  assign n30434 = ~n21364 & n30433 ;
  assign n30435 = ~n30429 & n30434 ;
  assign n30436 = n1187 & ~n9263 ;
  assign n30437 = n6419 & n30436 ;
  assign n30438 = ( ~n10093 & n14554 ) | ( ~n10093 & n30437 ) | ( n14554 & n30437 ) ;
  assign n30439 = n2010 ^ n302 ^ 1'b0 ;
  assign n30440 = n30439 ^ n7779 ^ n2156 ;
  assign n30441 = n5044 ^ n3716 ^ 1'b0 ;
  assign n30442 = n21656 & ~n30441 ;
  assign n30443 = ( n13601 & n30440 ) | ( n13601 & n30442 ) | ( n30440 & n30442 ) ;
  assign n30444 = ( ~n3385 & n9450 ) | ( ~n3385 & n10813 ) | ( n9450 & n10813 ) ;
  assign n30445 = n30444 ^ n9041 ^ 1'b0 ;
  assign n30446 = ( n2025 & ~n11583 ) | ( n2025 & n30445 ) | ( ~n11583 & n30445 ) ;
  assign n30447 = n15726 ^ n12380 ^ n172 ;
  assign n30451 = ( n1012 & n5840 ) | ( n1012 & n9595 ) | ( n5840 & n9595 ) ;
  assign n30448 = n2011 | n3706 ;
  assign n30449 = n30448 ^ n9736 ^ 1'b0 ;
  assign n30450 = n30449 ^ n6995 ^ n3244 ;
  assign n30452 = n30451 ^ n30450 ^ n6057 ;
  assign n30453 = ( ~n5697 & n6591 ) | ( ~n5697 & n23338 ) | ( n6591 & n23338 ) ;
  assign n30454 = ( ~n1789 & n5293 ) | ( ~n1789 & n17816 ) | ( n5293 & n17816 ) ;
  assign n30455 = ~n11736 & n30454 ;
  assign n30456 = n30455 ^ n6285 ^ 1'b0 ;
  assign n30457 = n30456 ^ n15251 ^ n7295 ;
  assign n30458 = ( n3436 & ~n8251 ) | ( n3436 & n30457 ) | ( ~n8251 & n30457 ) ;
  assign n30459 = ~n488 & n30458 ;
  assign n30460 = ~n29771 & n30459 ;
  assign n30461 = n12461 | n28639 ;
  assign n30462 = n13079 & ~n30461 ;
  assign n30463 = ( n2156 & n18044 ) | ( n2156 & n21350 ) | ( n18044 & n21350 ) ;
  assign n30464 = n7119 ^ n2049 ^ 1'b0 ;
  assign n30465 = ~n11510 & n30464 ;
  assign n30466 = n30465 ^ n12798 ^ n4798 ;
  assign n30467 = n20788 ^ n3292 ^ n3257 ;
  assign n30468 = n30467 ^ n23802 ^ n3584 ;
  assign n30469 = n2471 & n2501 ;
  assign n30470 = n30469 ^ n21787 ^ 1'b0 ;
  assign n30471 = n30470 ^ n4935 ^ n3100 ;
  assign n30472 = n17992 ^ n12367 ^ n5749 ;
  assign n30473 = ( ~n16082 & n29077 ) | ( ~n16082 & n30472 ) | ( n29077 & n30472 ) ;
  assign n30474 = ( n7124 & n30471 ) | ( n7124 & n30473 ) | ( n30471 & n30473 ) ;
  assign n30475 = n18603 ^ n3614 ^ 1'b0 ;
  assign n30476 = ( ~n4816 & n15532 ) | ( ~n4816 & n30475 ) | ( n15532 & n30475 ) ;
  assign n30477 = n30476 ^ n29948 ^ n11819 ;
  assign n30478 = n18329 ^ n15681 ^ n13213 ;
  assign n30479 = ( ~n29639 & n30151 ) | ( ~n29639 & n30478 ) | ( n30151 & n30478 ) ;
  assign n30480 = ~n16555 & n16634 ;
  assign n30482 = ( n13755 & n14158 ) | ( n13755 & ~n15128 ) | ( n14158 & ~n15128 ) ;
  assign n30481 = ( n1992 & n2249 ) | ( n1992 & n22967 ) | ( n2249 & n22967 ) ;
  assign n30483 = n30482 ^ n30481 ^ n3972 ;
  assign n30484 = ( x124 & n654 ) | ( x124 & ~n12141 ) | ( n654 & ~n12141 ) ;
  assign n30485 = ( x44 & ~n25530 ) | ( x44 & n30484 ) | ( ~n25530 & n30484 ) ;
  assign n30486 = ~n6908 & n7183 ;
  assign n30487 = ( n9957 & n10753 ) | ( n9957 & n22931 ) | ( n10753 & n22931 ) ;
  assign n30488 = n30487 ^ n30358 ^ 1'b0 ;
  assign n30489 = n1538 & n10145 ;
  assign n30490 = n30489 ^ n18671 ^ n3297 ;
  assign n30491 = n15489 ^ n9498 ^ n8199 ;
  assign n30492 = ( n4177 & n5993 ) | ( n4177 & ~n30491 ) | ( n5993 & ~n30491 ) ;
  assign n30498 = ( ~n4870 & n7325 ) | ( ~n4870 & n23860 ) | ( n7325 & n23860 ) ;
  assign n30493 = n427 & n4190 ;
  assign n30494 = n3252 & n30493 ;
  assign n30495 = n30494 ^ n9847 ^ n4313 ;
  assign n30496 = n17277 & ~n30495 ;
  assign n30497 = n30496 ^ n21849 ^ n9346 ;
  assign n30499 = n30498 ^ n30497 ^ n383 ;
  assign n30500 = n23973 ^ n391 ^ 1'b0 ;
  assign n30501 = n18671 ^ n6086 ^ 1'b0 ;
  assign n30502 = n30500 & n30501 ;
  assign n30503 = n30502 ^ n18468 ^ n2767 ;
  assign n30505 = n2532 | n4735 ;
  assign n30504 = ( n4421 & n5319 ) | ( n4421 & n16082 ) | ( n5319 & n16082 ) ;
  assign n30506 = n30505 ^ n30504 ^ n7856 ;
  assign n30507 = n30506 ^ n14829 ^ n14285 ;
  assign n30508 = n8361 ^ n1378 ^ 1'b0 ;
  assign n30509 = ~n22186 & n30508 ;
  assign n30510 = n28565 ^ n20179 ^ n2813 ;
  assign n30511 = n3008 & n19466 ;
  assign n30512 = n30511 ^ n7354 ^ 1'b0 ;
  assign n30513 = n8989 & n30512 ;
  assign n30514 = n30510 & n30513 ;
  assign n30521 = ( ~n2504 & n7367 ) | ( ~n2504 & n22151 ) | ( n7367 & n22151 ) ;
  assign n30517 = n9449 & ~n29181 ;
  assign n30518 = ~n24885 & n30517 ;
  assign n30515 = ( n1518 & ~n5357 ) | ( n1518 & n7354 ) | ( ~n5357 & n7354 ) ;
  assign n30516 = n20865 | n30515 ;
  assign n30519 = n30518 ^ n30516 ^ n1453 ;
  assign n30520 = n11924 & ~n30519 ;
  assign n30522 = n30521 ^ n30520 ^ 1'b0 ;
  assign n30523 = ( n9359 & ~n20973 ) | ( n9359 & n22469 ) | ( ~n20973 & n22469 ) ;
  assign n30524 = ( n5974 & n18438 ) | ( n5974 & n30523 ) | ( n18438 & n30523 ) ;
  assign n30525 = n17213 ^ n1129 ^ 1'b0 ;
  assign n30526 = n12101 & ~n30525 ;
  assign n30527 = n30526 ^ n28789 ^ 1'b0 ;
  assign n30528 = n23986 ^ n17928 ^ n4926 ;
  assign n30529 = n28383 ^ n20713 ^ n5160 ;
  assign n30530 = ( n6570 & n11513 ) | ( n6570 & ~n14460 ) | ( n11513 & ~n14460 ) ;
  assign n30531 = ~n25046 & n30530 ;
  assign n30532 = ~n6713 & n27667 ;
  assign n30533 = ( n20067 & n28885 ) | ( n20067 & ~n30532 ) | ( n28885 & ~n30532 ) ;
  assign n30534 = ( ~n12499 & n15619 ) | ( ~n12499 & n15988 ) | ( n15619 & n15988 ) ;
  assign n30535 = n17516 | n24205 ;
  assign n30536 = n30535 ^ n18675 ^ 1'b0 ;
  assign n30537 = ( n23766 & n26406 ) | ( n23766 & n30536 ) | ( n26406 & n30536 ) ;
  assign n30538 = ~n917 & n4127 ;
  assign n30539 = n30538 ^ n3356 ^ 1'b0 ;
  assign n30540 = n7615 | n7715 ;
  assign n30541 = n30539 & ~n30540 ;
  assign n30542 = n30541 ^ n2515 ^ 1'b0 ;
  assign n30543 = n24684 ^ n9366 ^ 1'b0 ;
  assign n30544 = n30542 & n30543 ;
  assign n30546 = n10193 | n23771 ;
  assign n30547 = n30546 ^ n5137 ^ 1'b0 ;
  assign n30548 = ( n5221 & n9400 ) | ( n5221 & n30547 ) | ( n9400 & n30547 ) ;
  assign n30545 = n7905 | n18706 ;
  assign n30549 = n30548 ^ n30545 ^ 1'b0 ;
  assign n30550 = ~n16739 & n22324 ;
  assign n30551 = ~n3385 & n30550 ;
  assign n30552 = n30551 ^ n15772 ^ n14887 ;
  assign n30553 = n3884 | n7453 ;
  assign n30554 = n517 & ~n30553 ;
  assign n30555 = ( n6147 & n22690 ) | ( n6147 & n30554 ) | ( n22690 & n30554 ) ;
  assign n30556 = n5760 ^ n3576 ^ n1667 ;
  assign n30557 = n3118 ^ n1707 ^ 1'b0 ;
  assign n30558 = ~n30556 & n30557 ;
  assign n30559 = ( n14284 & n18078 ) | ( n14284 & ~n30558 ) | ( n18078 & ~n30558 ) ;
  assign n30561 = n7741 & n13697 ;
  assign n30562 = n23646 & n30561 ;
  assign n30560 = n19813 & n26947 ;
  assign n30563 = n30562 ^ n30560 ^ 1'b0 ;
  assign n30564 = n30563 ^ n15652 ^ n6165 ;
  assign n30565 = ( n8467 & ~n13538 ) | ( n8467 & n24024 ) | ( ~n13538 & n24024 ) ;
  assign n30566 = n15578 ^ n4852 ^ 1'b0 ;
  assign n30569 = n8870 & ~n9170 ;
  assign n30570 = ( n8602 & ~n21647 ) | ( n8602 & n30569 ) | ( ~n21647 & n30569 ) ;
  assign n30567 = n4326 & ~n9653 ;
  assign n30568 = n30567 ^ n1939 ^ 1'b0 ;
  assign n30571 = n30570 ^ n30568 ^ n3561 ;
  assign n30572 = n12185 & ~n30571 ;
  assign n30573 = n13455 | n15216 ;
  assign n30574 = n27764 & ~n30573 ;
  assign n30575 = n14459 | n17170 ;
  assign n30576 = n30575 ^ n10146 ^ 1'b0 ;
  assign n30577 = n22229 ^ n10776 ^ n10296 ;
  assign n30578 = ( n16466 & n25496 ) | ( n16466 & ~n30577 ) | ( n25496 & ~n30577 ) ;
  assign n30579 = ( ~n4403 & n8431 ) | ( ~n4403 & n24129 ) | ( n8431 & n24129 ) ;
  assign n30580 = ( n4998 & n6499 ) | ( n4998 & ~n18414 ) | ( n6499 & ~n18414 ) ;
  assign n30581 = n30580 ^ n5774 ^ 1'b0 ;
  assign n30582 = n30581 ^ n9665 ^ n4205 ;
  assign n30583 = ( n21364 & n30579 ) | ( n21364 & ~n30582 ) | ( n30579 & ~n30582 ) ;
  assign n30584 = n11496 ^ n2516 ^ n567 ;
  assign n30585 = ( n6322 & ~n6802 ) | ( n6322 & n26633 ) | ( ~n6802 & n26633 ) ;
  assign n30586 = ( n23819 & ~n30584 ) | ( n23819 & n30585 ) | ( ~n30584 & n30585 ) ;
  assign n30587 = ( n1544 & n20197 ) | ( n1544 & n27416 ) | ( n20197 & n27416 ) ;
  assign n30588 = n30587 ^ n18319 ^ n4796 ;
  assign n30589 = ( n1308 & n5858 ) | ( n1308 & ~n27432 ) | ( n5858 & ~n27432 ) ;
  assign n30590 = n25124 ^ n9018 ^ n4735 ;
  assign n30591 = n30590 ^ n29820 ^ n19148 ;
  assign n30592 = n24310 ^ n18452 ^ n9982 ;
  assign n30593 = n5786 & n18150 ;
  assign n30594 = n30593 ^ n25245 ^ 1'b0 ;
  assign n30595 = n30203 ^ n24576 ^ n3744 ;
  assign n30596 = ( n4882 & n12602 ) | ( n4882 & ~n20267 ) | ( n12602 & ~n20267 ) ;
  assign n30597 = n20745 | n30596 ;
  assign n30598 = ( n17047 & n19993 ) | ( n17047 & n30597 ) | ( n19993 & n30597 ) ;
  assign n30599 = n5701 & n14109 ;
  assign n30600 = n30599 ^ n28347 ^ n22662 ;
  assign n30601 = ( n4356 & ~n20783 ) | ( n4356 & n27008 ) | ( ~n20783 & n27008 ) ;
  assign n30602 = n21770 ^ n17941 ^ n15149 ;
  assign n30603 = n16230 ^ n16134 ^ n7195 ;
  assign n30604 = n9972 ^ n8081 ^ n3121 ;
  assign n30605 = ( n3013 & ~n3820 ) | ( n3013 & n30604 ) | ( ~n3820 & n30604 ) ;
  assign n30606 = n30605 ^ n25579 ^ n21416 ;
  assign n30608 = n4683 & ~n13921 ;
  assign n30609 = n30608 ^ n29413 ^ 1'b0 ;
  assign n30607 = n1493 & ~n7008 ;
  assign n30610 = n30609 ^ n30607 ^ n15525 ;
  assign n30611 = ( ~n5190 & n8219 ) | ( ~n5190 & n18667 ) | ( n8219 & n18667 ) ;
  assign n30612 = n30611 ^ n27932 ^ 1'b0 ;
  assign n30613 = n4370 | n30612 ;
  assign n30614 = ( ~n4731 & n24435 ) | ( ~n4731 & n28275 ) | ( n24435 & n28275 ) ;
  assign n30615 = ~n29424 & n30614 ;
  assign n30616 = n14357 & n30615 ;
  assign n30617 = ~n10368 & n10813 ;
  assign n30618 = ~n19277 & n30617 ;
  assign n30619 = ( n4015 & ~n11001 ) | ( n4015 & n14686 ) | ( ~n11001 & n14686 ) ;
  assign n30620 = n30619 ^ n19437 ^ n18023 ;
  assign n30621 = ( n2656 & n13887 ) | ( n2656 & ~n14050 ) | ( n13887 & ~n14050 ) ;
  assign n30622 = ( n9627 & n13435 ) | ( n9627 & ~n30621 ) | ( n13435 & ~n30621 ) ;
  assign n30623 = ( n5140 & ~n13266 ) | ( n5140 & n18563 ) | ( ~n13266 & n18563 ) ;
  assign n30624 = n24861 ^ n12616 ^ n6071 ;
  assign n30625 = n12694 & ~n28626 ;
  assign n30626 = n7228 ^ n6302 ^ n6067 ;
  assign n30627 = n18160 ^ n5494 ^ n1765 ;
  assign n30628 = n30627 ^ n22007 ^ 1'b0 ;
  assign n30629 = ( ~n2079 & n10127 ) | ( ~n2079 & n29046 ) | ( n10127 & n29046 ) ;
  assign n30630 = n20994 ^ n15543 ^ 1'b0 ;
  assign n30632 = n15381 ^ n3173 ^ n1909 ;
  assign n30631 = ( n13629 & ~n22758 ) | ( n13629 & n23369 ) | ( ~n22758 & n23369 ) ;
  assign n30633 = n30632 ^ n30631 ^ n28302 ;
  assign n30634 = n21965 ^ n3376 ^ x53 ;
  assign n30635 = n16691 ^ n14755 ^ n5631 ;
  assign n30636 = n21245 ^ n2892 ^ n2394 ;
  assign n30640 = ( n5379 & ~n8989 ) | ( n5379 & n16909 ) | ( ~n8989 & n16909 ) ;
  assign n30637 = n20998 ^ n10110 ^ 1'b0 ;
  assign n30638 = ~n15822 & n30637 ;
  assign n30639 = ( ~n6343 & n8351 ) | ( ~n6343 & n30638 ) | ( n8351 & n30638 ) ;
  assign n30641 = n30640 ^ n30639 ^ n4823 ;
  assign n30642 = n22328 ^ n3208 ^ n899 ;
  assign n30643 = ~n10738 & n19644 ;
  assign n30644 = ~n1967 & n30643 ;
  assign n30645 = ~n1926 & n9974 ;
  assign n30646 = n30645 ^ n7101 ^ 1'b0 ;
  assign n30647 = n26579 ^ n3907 ^ n3256 ;
  assign n30648 = n30647 ^ n2747 ^ 1'b0 ;
  assign n30649 = ~n26997 & n30648 ;
  assign n30650 = n4828 ^ n3396 ^ n936 ;
  assign n30651 = ( n2068 & n6208 ) | ( n2068 & n6443 ) | ( n6208 & n6443 ) ;
  assign n30652 = ( ~n10025 & n29950 ) | ( ~n10025 & n30651 ) | ( n29950 & n30651 ) ;
  assign n30653 = n16359 ^ n10938 ^ n5702 ;
  assign n30654 = n23367 ^ n19999 ^ n18847 ;
  assign n30655 = n9943 ^ n3061 ^ 1'b0 ;
  assign n30656 = n30655 ^ n14641 ^ n1848 ;
  assign n30657 = n25902 ^ n16238 ^ 1'b0 ;
  assign n30658 = n30657 ^ n14222 ^ n2783 ;
  assign n30659 = n18224 ^ n14313 ^ n9891 ;
  assign n30660 = ( n1991 & n7687 ) | ( n1991 & n22304 ) | ( n7687 & n22304 ) ;
  assign n30662 = ( ~n4773 & n9091 ) | ( ~n4773 & n17209 ) | ( n9091 & n17209 ) ;
  assign n30661 = ~n1810 & n3328 ;
  assign n30663 = n30662 ^ n30661 ^ 1'b0 ;
  assign n30664 = ~n3130 & n22768 ;
  assign n30665 = n30664 ^ n17774 ^ 1'b0 ;
  assign n30666 = n6643 | n18589 ;
  assign n30667 = n30666 ^ n15635 ^ 1'b0 ;
  assign n30668 = n23207 ^ n11109 ^ n4627 ;
  assign n30669 = n30668 ^ n5408 ^ n5227 ;
  assign n30670 = n26718 ^ n19800 ^ 1'b0 ;
  assign n30671 = n11388 & ~n30670 ;
  assign n30672 = n30671 ^ n9495 ^ n1638 ;
  assign n30674 = ( n696 & n4740 ) | ( n696 & ~n10839 ) | ( n4740 & ~n10839 ) ;
  assign n30673 = ( ~n3714 & n10594 ) | ( ~n3714 & n13340 ) | ( n10594 & n13340 ) ;
  assign n30675 = n30674 ^ n30673 ^ n5683 ;
  assign n30676 = n12893 ^ n8537 ^ n7902 ;
  assign n30677 = n28134 ^ n20466 ^ n10472 ;
  assign n30678 = ( n8451 & n15581 ) | ( n8451 & ~n20609 ) | ( n15581 & ~n20609 ) ;
  assign n30679 = ( n23518 & n27466 ) | ( n23518 & ~n30678 ) | ( n27466 & ~n30678 ) ;
  assign n30680 = n7406 | n15687 ;
  assign n30681 = ( ~n7246 & n30465 ) | ( ~n7246 & n30680 ) | ( n30465 & n30680 ) ;
  assign n30682 = n16660 ^ n10048 ^ 1'b0 ;
  assign n30683 = n1695 & n30682 ;
  assign n30684 = n30683 ^ n3581 ^ 1'b0 ;
  assign n30685 = n4186 & ~n5968 ;
  assign n30686 = n10517 | n23620 ;
  assign n30687 = n30686 ^ n7922 ^ 1'b0 ;
  assign n30688 = n30687 ^ n18995 ^ n1183 ;
  assign n30693 = ( n2100 & n5926 ) | ( n2100 & ~n24961 ) | ( n5926 & ~n24961 ) ;
  assign n30689 = n7320 & ~n19258 ;
  assign n30690 = n30689 ^ n19923 ^ 1'b0 ;
  assign n30691 = n30690 ^ n1591 ^ 1'b0 ;
  assign n30692 = ~n17080 & n30691 ;
  assign n30694 = n30693 ^ n30692 ^ n7156 ;
  assign n30695 = ( n2422 & n2529 ) | ( n2422 & n4619 ) | ( n2529 & n4619 ) ;
  assign n30696 = n30695 ^ n25527 ^ n3515 ;
  assign n30697 = ( ~n16747 & n16790 ) | ( ~n16747 & n28528 ) | ( n16790 & n28528 ) ;
  assign n30698 = n20959 ^ n7814 ^ n2609 ;
  assign n30700 = n15887 ^ n9599 ^ n5522 ;
  assign n30699 = n4504 & ~n16445 ;
  assign n30701 = n30700 ^ n30699 ^ 1'b0 ;
  assign n30702 = ( ~n11130 & n28577 ) | ( ~n11130 & n30701 ) | ( n28577 & n30701 ) ;
  assign n30703 = n6626 ^ n5799 ^ n2297 ;
  assign n30704 = ( n5576 & ~n7274 ) | ( n5576 & n30703 ) | ( ~n7274 & n30703 ) ;
  assign n30705 = n28960 ^ n27747 ^ n19394 ;
  assign n30706 = n30705 ^ n15907 ^ n9552 ;
  assign n30707 = n18164 ^ n17982 ^ n10462 ;
  assign n30708 = ~n14139 & n30707 ;
  assign n30709 = ~n13833 & n30708 ;
  assign n30710 = n1901 & ~n29368 ;
  assign n30711 = n1380 & n2913 ;
  assign n30712 = n30711 ^ n15225 ^ 1'b0 ;
  assign n30713 = ( ~n14507 & n17308 ) | ( ~n14507 & n30259 ) | ( n17308 & n30259 ) ;
  assign n30714 = ( n211 & ~n3357 ) | ( n211 & n3524 ) | ( ~n3357 & n3524 ) ;
  assign n30715 = ( n9738 & ~n28412 ) | ( n9738 & n30714 ) | ( ~n28412 & n30714 ) ;
  assign n30716 = ( n24009 & n30487 ) | ( n24009 & ~n30715 ) | ( n30487 & ~n30715 ) ;
  assign n30717 = ( n19258 & ~n30713 ) | ( n19258 & n30716 ) | ( ~n30713 & n30716 ) ;
  assign n30718 = ( n1290 & ~n13496 ) | ( n1290 & n21851 ) | ( ~n13496 & n21851 ) ;
  assign n30719 = n30718 ^ n19108 ^ n168 ;
  assign n30720 = n21471 ^ n20078 ^ n18447 ;
  assign n30721 = n30720 ^ n11057 ^ n4529 ;
  assign n30722 = ( n16587 & ~n23690 ) | ( n16587 & n30505 ) | ( ~n23690 & n30505 ) ;
  assign n30723 = n30722 ^ n25530 ^ n21719 ;
  assign n30724 = ( n20372 & ~n23618 ) | ( n20372 & n27498 ) | ( ~n23618 & n27498 ) ;
  assign n30725 = ( n6885 & ~n16249 ) | ( n6885 & n28190 ) | ( ~n16249 & n28190 ) ;
  assign n30726 = n5024 ^ n2958 ^ 1'b0 ;
  assign n30727 = n30726 ^ n20089 ^ n5597 ;
  assign n30728 = ( n7878 & ~n14571 ) | ( n7878 & n25906 ) | ( ~n14571 & n25906 ) ;
  assign n30729 = n30728 ^ n8339 ^ 1'b0 ;
  assign n30730 = n13848 & ~n30729 ;
  assign n30731 = ~n8639 & n30730 ;
  assign n30732 = ( n30725 & ~n30727 ) | ( n30725 & n30731 ) | ( ~n30727 & n30731 ) ;
  assign n30733 = n1972 & ~n26309 ;
  assign n30734 = n6980 ^ n4204 ^ n782 ;
  assign n30735 = n30734 ^ n10934 ^ n1679 ;
  assign n30736 = n30735 ^ n7006 ^ n2840 ;
  assign n30737 = ( n18701 & n21095 ) | ( n18701 & n26633 ) | ( n21095 & n26633 ) ;
  assign n30738 = n16848 ^ n15706 ^ 1'b0 ;
  assign n30739 = ~n30737 & n30738 ;
  assign n30740 = n2058 ^ n724 ^ 1'b0 ;
  assign n30741 = n27582 | n30740 ;
  assign n30742 = ~n4301 & n25496 ;
  assign n30743 = n30742 ^ n4527 ^ 1'b0 ;
  assign n30744 = ( ~n2388 & n25018 ) | ( ~n2388 & n29023 ) | ( n25018 & n29023 ) ;
  assign n30745 = n24711 ^ n10544 ^ n7976 ;
  assign n30746 = n28640 ^ n13650 ^ n1332 ;
  assign n30747 = n30746 ^ n19016 ^ 1'b0 ;
  assign n30748 = n9300 & n12850 ;
  assign n30749 = ( n7592 & n12227 ) | ( n7592 & n27071 ) | ( n12227 & n27071 ) ;
  assign n30750 = ( ~n7428 & n10187 ) | ( ~n7428 & n22469 ) | ( n10187 & n22469 ) ;
  assign n30751 = ( n6961 & n20947 ) | ( n6961 & ~n22611 ) | ( n20947 & ~n22611 ) ;
  assign n30752 = n3959 & ~n18422 ;
  assign n30753 = n7633 & n30752 ;
  assign n30754 = ( n500 & ~n15319 ) | ( n500 & n30753 ) | ( ~n15319 & n30753 ) ;
  assign n30755 = ( n2637 & n28892 ) | ( n2637 & n30754 ) | ( n28892 & n30754 ) ;
  assign n30756 = n17560 ^ n5088 ^ n1929 ;
  assign n30757 = n30756 ^ n21833 ^ 1'b0 ;
  assign n30758 = ~n28775 & n30757 ;
  assign n30759 = n9864 | n17781 ;
  assign n30760 = n5286 & ~n30759 ;
  assign n30761 = ( n9618 & n23258 ) | ( n9618 & n30760 ) | ( n23258 & n30760 ) ;
  assign n30762 = n30761 ^ n9429 ^ 1'b0 ;
  assign n30763 = n12172 & n30762 ;
  assign n30764 = ( n809 & n8684 ) | ( n809 & n8820 ) | ( n8684 & n8820 ) ;
  assign n30765 = n20224 & ~n26263 ;
  assign n30766 = ~n2849 & n30765 ;
  assign n30767 = ( n8944 & n30764 ) | ( n8944 & ~n30766 ) | ( n30764 & ~n30766 ) ;
  assign n30769 = n21243 ^ n12159 ^ n6239 ;
  assign n30768 = n22351 ^ n14504 ^ n13448 ;
  assign n30770 = n30769 ^ n30768 ^ n22738 ;
  assign n30771 = ( n7260 & n9408 ) | ( n7260 & ~n11361 ) | ( n9408 & ~n11361 ) ;
  assign n30772 = n6532 | n25794 ;
  assign n30773 = ( n306 & ~n25500 ) | ( n306 & n30772 ) | ( ~n25500 & n30772 ) ;
  assign n30774 = n24548 ^ n17312 ^ n442 ;
  assign n30775 = n528 & n15266 ;
  assign n30776 = n1492 | n24588 ;
  assign n30777 = n30776 ^ n23281 ^ 1'b0 ;
  assign n30778 = ( n29750 & n30775 ) | ( n29750 & n30777 ) | ( n30775 & n30777 ) ;
  assign n30779 = n9668 ^ n5148 ^ 1'b0 ;
  assign n30780 = ( ~n13994 & n21790 ) | ( ~n13994 & n30779 ) | ( n21790 & n30779 ) ;
  assign n30781 = n27081 ^ n23869 ^ n5972 ;
  assign n30782 = n11507 & n18184 ;
  assign n30783 = n7903 & n30782 ;
  assign n30784 = ~n8642 & n27577 ;
  assign n30785 = ~n24558 & n30784 ;
  assign n30786 = n945 & n5724 ;
  assign n30787 = n5251 & n30786 ;
  assign n30788 = n23921 ^ n22830 ^ n7303 ;
  assign n30789 = n30788 ^ n28696 ^ n11872 ;
  assign n30790 = ( n3144 & ~n6729 ) | ( n3144 & n7561 ) | ( ~n6729 & n7561 ) ;
  assign n30791 = n30790 ^ n16820 ^ n1015 ;
  assign n30792 = ( n6199 & n11755 ) | ( n6199 & n18087 ) | ( n11755 & n18087 ) ;
  assign n30793 = n21766 ^ n5471 ^ n1872 ;
  assign n30794 = n16501 ^ n5592 ^ n1485 ;
  assign n30795 = n16948 ^ n6233 ^ x3 ;
  assign n30796 = n22668 ^ n15076 ^ n9430 ;
  assign n30797 = ( n3301 & n5763 ) | ( n3301 & n17943 ) | ( n5763 & n17943 ) ;
  assign n30798 = n21067 ^ n2222 ^ n413 ;
  assign n30799 = n29810 ^ n19536 ^ 1'b0 ;
  assign n30800 = ~n30798 & n30799 ;
  assign n30801 = n29062 ^ n20863 ^ n5146 ;
  assign n30802 = n12794 ^ n10764 ^ n7486 ;
  assign n30803 = ( n5425 & n26944 ) | ( n5425 & n30802 ) | ( n26944 & n30802 ) ;
  assign n30804 = ( n9940 & ~n18792 ) | ( n9940 & n28588 ) | ( ~n18792 & n28588 ) ;
  assign n30805 = n20874 ^ n5468 ^ n2216 ;
  assign n30806 = n23595 ^ n11066 ^ n9382 ;
  assign n30807 = ( n9068 & n21730 ) | ( n9068 & n23257 ) | ( n21730 & n23257 ) ;
  assign n30808 = ( n4321 & n11573 ) | ( n4321 & ~n18209 ) | ( n11573 & ~n18209 ) ;
  assign n30809 = n30808 ^ n7205 ^ n2163 ;
  assign n30810 = n30807 & n30809 ;
  assign n30811 = ( n6303 & n9495 ) | ( n6303 & n21118 ) | ( n9495 & n21118 ) ;
  assign n30812 = n30811 ^ n12075 ^ n3792 ;
  assign n30813 = n26812 ^ n25041 ^ 1'b0 ;
  assign n30814 = n27632 ^ n4001 ^ 1'b0 ;
  assign n30815 = n16580 | n30814 ;
  assign n30816 = ~n9570 & n27948 ;
  assign n30817 = n30816 ^ n3450 ^ 1'b0 ;
  assign n30818 = n26469 ^ n15274 ^ x38 ;
  assign n30819 = ( ~n4622 & n28280 ) | ( ~n4622 & n30818 ) | ( n28280 & n30818 ) ;
  assign n30820 = n21611 ^ n17119 ^ 1'b0 ;
  assign n30821 = ~n30819 & n30820 ;
  assign n30822 = n16359 | n22701 ;
  assign n30823 = n18756 ^ n17738 ^ 1'b0 ;
  assign n30824 = n16575 ^ n11170 ^ n6845 ;
  assign n30825 = n30824 ^ n8412 ^ n889 ;
  assign n30826 = n4763 | n7528 ;
  assign n30827 = n30826 ^ n19010 ^ n11074 ;
  assign n30828 = n5882 | n7559 ;
  assign n30829 = n3485 | n30828 ;
  assign n30830 = ( n3244 & n6658 ) | ( n3244 & ~n22490 ) | ( n6658 & ~n22490 ) ;
  assign n30831 = n1620 & n13946 ;
  assign n30832 = n30831 ^ n12786 ^ n5281 ;
  assign n30833 = n30832 ^ n18403 ^ 1'b0 ;
  assign n30834 = ~n9600 & n17229 ;
  assign n30835 = n5710 ^ n5674 ^ n3050 ;
  assign n30836 = n12765 & n17259 ;
  assign n30837 = ~n6083 & n30836 ;
  assign n30838 = ( n16597 & n30835 ) | ( n16597 & ~n30837 ) | ( n30835 & ~n30837 ) ;
  assign n30839 = ( n8519 & ~n11496 ) | ( n8519 & n17310 ) | ( ~n11496 & n17310 ) ;
  assign n30840 = n30839 ^ n11156 ^ n1380 ;
  assign n30841 = n27565 ^ n23187 ^ n18998 ;
  assign n30842 = n21096 ^ n18976 ^ 1'b0 ;
  assign n30846 = n20900 ^ n3054 ^ 1'b0 ;
  assign n30847 = n24058 | n30846 ;
  assign n30843 = ( ~n11161 & n24399 ) | ( ~n11161 & n27662 ) | ( n24399 & n27662 ) ;
  assign n30844 = n30843 ^ n7953 ^ n3866 ;
  assign n30845 = n25173 | n30844 ;
  assign n30848 = n30847 ^ n30845 ^ n18077 ;
  assign n30849 = n30848 ^ n23432 ^ n1876 ;
  assign n30850 = ( n19256 & n30842 ) | ( n19256 & ~n30849 ) | ( n30842 & ~n30849 ) ;
  assign n30851 = n11306 ^ n10577 ^ n6940 ;
  assign n30852 = n15040 ^ n13183 ^ 1'b0 ;
  assign n30853 = ( ~n20127 & n30851 ) | ( ~n20127 & n30852 ) | ( n30851 & n30852 ) ;
  assign n30854 = n10316 ^ n5812 ^ n3671 ;
  assign n30855 = ~n29357 & n30854 ;
  assign n30856 = ( n5376 & ~n9444 ) | ( n5376 & n14786 ) | ( ~n9444 & n14786 ) ;
  assign n30857 = n30856 ^ n7703 ^ 1'b0 ;
  assign n30858 = n9804 & n30857 ;
  assign n30859 = n7244 | n23440 ;
  assign n30860 = n9329 | n30859 ;
  assign n30861 = ( n3782 & n17460 ) | ( n3782 & n26310 ) | ( n17460 & n26310 ) ;
  assign n30862 = n21535 ^ n21166 ^ n12992 ;
  assign n30863 = n23617 ^ n19437 ^ n7689 ;
  assign n30864 = ( n2041 & ~n2794 ) | ( n2041 & n12211 ) | ( ~n2794 & n12211 ) ;
  assign n30865 = n3156 & n12495 ;
  assign n30866 = n27971 & n30865 ;
  assign n30867 = ( n6931 & ~n21966 ) | ( n6931 & n30866 ) | ( ~n21966 & n30866 ) ;
  assign n30868 = n12573 | n30867 ;
  assign n30869 = n30674 ^ n11839 ^ 1'b0 ;
  assign n30870 = n16711 & ~n30869 ;
  assign n30871 = ( n17452 & ~n18274 ) | ( n17452 & n30870 ) | ( ~n18274 & n30870 ) ;
  assign n30872 = n30871 ^ n3899 ^ 1'b0 ;
  assign n30873 = ~n6415 & n29705 ;
  assign n30874 = n30873 ^ n1163 ^ 1'b0 ;
  assign n30875 = n17019 | n30874 ;
  assign n30876 = n24500 & ~n30875 ;
  assign n30877 = n2570 & n19662 ;
  assign n30878 = n30877 ^ n19530 ^ 1'b0 ;
  assign n30879 = n4982 & ~n15363 ;
  assign n30880 = ~n27317 & n30879 ;
  assign n30881 = ( ~n5595 & n13128 ) | ( ~n5595 & n13992 ) | ( n13128 & n13992 ) ;
  assign n30882 = n30881 ^ n14247 ^ n7534 ;
  assign n30883 = ( n3096 & n6959 ) | ( n3096 & n15269 ) | ( n6959 & n15269 ) ;
  assign n30884 = ( n2965 & ~n20093 ) | ( n2965 & n30883 ) | ( ~n20093 & n30883 ) ;
  assign n30885 = n30884 ^ n22012 ^ n18829 ;
  assign n30886 = ( x106 & n13169 ) | ( x106 & n30885 ) | ( n13169 & n30885 ) ;
  assign n30887 = n26062 ^ n24399 ^ n15826 ;
  assign n30891 = ( ~n1674 & n5972 ) | ( ~n1674 & n7665 ) | ( n5972 & n7665 ) ;
  assign n30890 = ( n9059 & n15638 ) | ( n9059 & ~n23684 ) | ( n15638 & ~n23684 ) ;
  assign n30888 = n6749 ^ n4210 ^ n1203 ;
  assign n30889 = ( n2361 & n9207 ) | ( n2361 & ~n30888 ) | ( n9207 & ~n30888 ) ;
  assign n30892 = n30891 ^ n30890 ^ n30889 ;
  assign n30893 = ( ~n3982 & n17857 ) | ( ~n3982 & n18911 ) | ( n17857 & n18911 ) ;
  assign n30894 = n17758 | n30893 ;
  assign n30895 = n17778 ^ n8255 ^ n4421 ;
  assign n30896 = ( n10867 & n11257 ) | ( n10867 & n13221 ) | ( n11257 & n13221 ) ;
  assign n30897 = n22272 ^ n18973 ^ n1774 ;
  assign n30898 = ( n10771 & ~n30896 ) | ( n10771 & n30897 ) | ( ~n30896 & n30897 ) ;
  assign n30900 = n1449 & n11653 ;
  assign n30901 = n30900 ^ n805 ^ 1'b0 ;
  assign n30899 = n2208 | n7531 ;
  assign n30902 = n30901 ^ n30899 ^ 1'b0 ;
  assign n30903 = n18694 | n28626 ;
  assign n30904 = n30902 | n30903 ;
  assign n30905 = n9116 | n11354 ;
  assign n30906 = n30905 ^ n12646 ^ 1'b0 ;
  assign n30907 = ~n1253 & n6634 ;
  assign n30908 = n9970 & ~n11088 ;
  assign n30909 = n30908 ^ n14615 ^ 1'b0 ;
  assign n30910 = ( n21778 & ~n30907 ) | ( n21778 & n30909 ) | ( ~n30907 & n30909 ) ;
  assign n30911 = n13491 ^ n3140 ^ n567 ;
  assign n30912 = n30911 ^ n10603 ^ n3220 ;
  assign n30913 = n20795 ^ n20615 ^ n9638 ;
  assign n30914 = ( ~n4289 & n12237 ) | ( ~n4289 & n30913 ) | ( n12237 & n30913 ) ;
  assign n30915 = ( ~n3518 & n5388 ) | ( ~n3518 & n29435 ) | ( n5388 & n29435 ) ;
  assign n30916 = n5793 ^ n5635 ^ 1'b0 ;
  assign n30917 = n9478 | n30916 ;
  assign n30918 = n30917 ^ n7437 ^ n4185 ;
  assign n30919 = ( n1790 & n18843 ) | ( n1790 & ~n30769 ) | ( n18843 & ~n30769 ) ;
  assign n30920 = ( n30915 & n30918 ) | ( n30915 & ~n30919 ) | ( n30918 & ~n30919 ) ;
  assign n30921 = n25839 ^ n11278 ^ n1001 ;
  assign n30922 = ( n11583 & n12200 ) | ( n11583 & ~n27196 ) | ( n12200 & ~n27196 ) ;
  assign n30923 = n30922 ^ n26358 ^ n5928 ;
  assign n30924 = n30923 ^ n18337 ^ n14593 ;
  assign n30925 = ( n903 & ~n11451 ) | ( n903 & n13453 ) | ( ~n11451 & n13453 ) ;
  assign n30926 = n30387 ^ n11451 ^ n5003 ;
  assign n30927 = n21979 ^ n14107 ^ n5977 ;
  assign n30928 = n30927 ^ n7835 ^ 1'b0 ;
  assign n30929 = n5735 ^ n5348 ^ 1'b0 ;
  assign n30930 = ~n3085 & n30929 ;
  assign n30931 = ( ~n5948 & n7588 ) | ( ~n5948 & n11199 ) | ( n7588 & n11199 ) ;
  assign n30932 = ( n1869 & n23781 ) | ( n1869 & ~n25186 ) | ( n23781 & ~n25186 ) ;
  assign n30933 = ( n3757 & n18235 ) | ( n3757 & ~n30932 ) | ( n18235 & ~n30932 ) ;
  assign n30934 = ( n10753 & n30931 ) | ( n10753 & n30933 ) | ( n30931 & n30933 ) ;
  assign n30935 = ( n790 & n7255 ) | ( n790 & ~n30934 ) | ( n7255 & ~n30934 ) ;
  assign n30936 = ( ~n3688 & n6007 ) | ( ~n3688 & n16606 ) | ( n6007 & n16606 ) ;
  assign n30938 = ( ~n497 & n4755 ) | ( ~n497 & n14833 ) | ( n4755 & n14833 ) ;
  assign n30937 = n161 & n7975 ;
  assign n30939 = n30938 ^ n30937 ^ 1'b0 ;
  assign n30940 = ~n548 & n30939 ;
  assign n30941 = ( n11920 & ~n14993 ) | ( n11920 & n24964 ) | ( ~n14993 & n24964 ) ;
  assign n30942 = ( n511 & ~n17116 ) | ( n511 & n30941 ) | ( ~n17116 & n30941 ) ;
  assign n30943 = ~n2430 & n13810 ;
  assign n30944 = n8605 ^ n5358 ^ n509 ;
  assign n30945 = n23763 & n25529 ;
  assign n30946 = ( n3901 & n4473 ) | ( n3901 & ~n27577 ) | ( n4473 & ~n27577 ) ;
  assign n30951 = n20318 & ~n26236 ;
  assign n30947 = n26010 ^ n25802 ^ n15302 ;
  assign n30948 = n30373 ^ n28279 ^ n6776 ;
  assign n30949 = ( n5852 & n27852 ) | ( n5852 & n30948 ) | ( n27852 & n30948 ) ;
  assign n30950 = ~n30947 & n30949 ;
  assign n30952 = n30951 ^ n30950 ^ 1'b0 ;
  assign n30953 = n29199 ^ n5735 ^ 1'b0 ;
  assign n30955 = n18001 ^ n5766 ^ n1719 ;
  assign n30956 = n30955 ^ n10351 ^ n6651 ;
  assign n30957 = n30956 ^ n11105 ^ 1'b0 ;
  assign n30958 = n30957 ^ n18865 ^ n16671 ;
  assign n30954 = n26561 ^ n14458 ^ n534 ;
  assign n30959 = n30958 ^ n30954 ^ 1'b0 ;
  assign n30960 = n30953 | n30959 ;
  assign n30961 = n19390 ^ n5424 ^ n2028 ;
  assign n30962 = n9392 ^ n7565 ^ n1638 ;
  assign n30963 = n30962 ^ n16378 ^ n15860 ;
  assign n30964 = n22408 ^ n9931 ^ n2842 ;
  assign n30965 = ( n1377 & n29791 ) | ( n1377 & n30964 ) | ( n29791 & n30964 ) ;
  assign n30966 = n24828 ^ n3045 ^ n1410 ;
  assign n30967 = n30966 ^ n17199 ^ n516 ;
  assign n30968 = n20874 ^ n20760 ^ n7481 ;
  assign n30969 = n19901 ^ n14559 ^ n11222 ;
  assign n30970 = ( n1516 & ~n8906 ) | ( n1516 & n23019 ) | ( ~n8906 & n23019 ) ;
  assign n30971 = n30970 ^ n13152 ^ x1 ;
  assign n30972 = n4011 ^ n3685 ^ 1'b0 ;
  assign n30973 = n2897 | n30972 ;
  assign n30974 = n1759 & n9822 ;
  assign n30975 = n30973 & n30974 ;
  assign n30976 = n15591 | n30975 ;
  assign n30977 = n30976 ^ n8019 ^ 1'b0 ;
  assign n30978 = n7008 & ~n15484 ;
  assign n30979 = ( n16814 & ~n30888 ) | ( n16814 & n30978 ) | ( ~n30888 & n30978 ) ;
  assign n30980 = ( ~n1575 & n2890 ) | ( ~n1575 & n14183 ) | ( n2890 & n14183 ) ;
  assign n30981 = n13747 & n30980 ;
  assign n30982 = n30979 & n30981 ;
  assign n30983 = n28254 ^ n6231 ^ n6092 ;
  assign n30986 = n7222 | n11205 ;
  assign n30987 = n30986 ^ n5648 ^ 1'b0 ;
  assign n30988 = n30987 ^ n4174 ^ n439 ;
  assign n30984 = n6739 ^ n3967 ^ 1'b0 ;
  assign n30985 = n14353 | n30984 ;
  assign n30989 = n30988 ^ n30985 ^ n15925 ;
  assign n30990 = ~n4125 & n10759 ;
  assign n30991 = n9347 & n30990 ;
  assign n30992 = ( n14271 & n25435 ) | ( n14271 & ~n30991 ) | ( n25435 & ~n30991 ) ;
  assign n30993 = ( n1655 & n4156 ) | ( n1655 & n11118 ) | ( n4156 & n11118 ) ;
  assign n30994 = n27078 ^ n10544 ^ n3222 ;
  assign n30995 = ~n30993 & n30994 ;
  assign n30996 = ~n997 & n11436 ;
  assign n30997 = ( n4148 & n9935 ) | ( n4148 & n30996 ) | ( n9935 & n30996 ) ;
  assign n30998 = ( n7124 & n21268 ) | ( n7124 & n24028 ) | ( n21268 & n24028 ) ;
  assign n30999 = n20589 ^ n19809 ^ 1'b0 ;
  assign n31000 = n30277 | n30999 ;
  assign n31001 = n3856 ^ n1813 ^ n1063 ;
  assign n31002 = n31001 ^ n28403 ^ n1724 ;
  assign n31003 = n5164 & n31002 ;
  assign n31004 = n31003 ^ n19714 ^ 1'b0 ;
  assign n31005 = n17640 ^ n5874 ^ n2726 ;
  assign n31006 = n13506 | n31005 ;
  assign n31007 = n1743 & ~n31006 ;
  assign n31008 = n17569 ^ n614 ^ x117 ;
  assign n31009 = n22741 ^ n21052 ^ n17802 ;
  assign n31010 = n31009 ^ n22913 ^ n8301 ;
  assign n31011 = ( n3875 & n10652 ) | ( n3875 & ~n20781 ) | ( n10652 & ~n20781 ) ;
  assign n31012 = n31011 ^ n11948 ^ n3971 ;
  assign n31013 = ( n479 & n1526 ) | ( n479 & n11064 ) | ( n1526 & n11064 ) ;
  assign n31014 = ( n14571 & ~n18398 ) | ( n14571 & n31013 ) | ( ~n18398 & n31013 ) ;
  assign n31015 = ( n13067 & n27282 ) | ( n13067 & ~n31014 ) | ( n27282 & ~n31014 ) ;
  assign n31016 = n31015 ^ n9151 ^ n1122 ;
  assign n31017 = n31016 ^ n2761 ^ n158 ;
  assign n31019 = ( n5226 & n8863 ) | ( n5226 & n19158 ) | ( n8863 & n19158 ) ;
  assign n31018 = n27523 ^ n26530 ^ n7125 ;
  assign n31020 = n31019 ^ n31018 ^ n434 ;
  assign n31021 = n31020 ^ n26827 ^ n10856 ;
  assign n31022 = ( n3273 & n6233 ) | ( n3273 & ~n13289 ) | ( n6233 & ~n13289 ) ;
  assign n31023 = n31022 ^ n6730 ^ n399 ;
  assign n31024 = n28002 ^ n15484 ^ n214 ;
  assign n31025 = n2801 & n24441 ;
  assign n31026 = n24586 & n31025 ;
  assign n31027 = n736 & n4651 ;
  assign n31028 = ( n5512 & n12084 ) | ( n5512 & n29522 ) | ( n12084 & n29522 ) ;
  assign n31029 = n31028 ^ n2896 ^ 1'b0 ;
  assign n31030 = n31027 | n31029 ;
  assign n31031 = n1080 & ~n7798 ;
  assign n31032 = ( n4573 & ~n28788 ) | ( n4573 & n31031 ) | ( ~n28788 & n31031 ) ;
  assign n31033 = n7780 ^ n4398 ^ 1'b0 ;
  assign n31034 = n5532 | n31033 ;
  assign n31035 = n31032 & ~n31034 ;
  assign n31036 = n17015 ^ n5013 ^ n1180 ;
  assign n31037 = ~n19800 & n31036 ;
  assign n31038 = n15110 & ~n31037 ;
  assign n31039 = n16708 & ~n29951 ;
  assign n31040 = n9951 & n24869 ;
  assign n31041 = n2107 & n31040 ;
  assign n31042 = n31041 ^ n22347 ^ 1'b0 ;
  assign n31044 = n15476 ^ n6147 ^ 1'b0 ;
  assign n31043 = n15151 ^ n12237 ^ n6241 ;
  assign n31045 = n31044 ^ n31043 ^ n23969 ;
  assign n31046 = n17220 ^ n9321 ^ n7538 ;
  assign n31047 = ( n10606 & n21268 ) | ( n10606 & ~n31046 ) | ( n21268 & ~n31046 ) ;
  assign n31048 = n11330 & ~n21264 ;
  assign n31049 = n31048 ^ n27379 ^ n6439 ;
  assign n31050 = ( n4396 & ~n28216 ) | ( n4396 & n31049 ) | ( ~n28216 & n31049 ) ;
  assign n31051 = n8099 ^ n4193 ^ 1'b0 ;
  assign n31052 = n5513 & n31051 ;
  assign n31053 = n8241 & n16927 ;
  assign n31054 = n31053 ^ n16563 ^ 1'b0 ;
  assign n31055 = ~n2249 & n14344 ;
  assign n31056 = ~n24861 & n31055 ;
  assign n31057 = n11281 | n19164 ;
  assign n31058 = ( ~n13824 & n20643 ) | ( ~n13824 & n23810 ) | ( n20643 & n23810 ) ;
  assign n31059 = ( n295 & n31057 ) | ( n295 & n31058 ) | ( n31057 & n31058 ) ;
  assign n31060 = ( n1025 & ~n2170 ) | ( n1025 & n20049 ) | ( ~n2170 & n20049 ) ;
  assign n31061 = ( n2350 & n10424 ) | ( n2350 & ~n13351 ) | ( n10424 & ~n13351 ) ;
  assign n31062 = ( n6731 & ~n20769 ) | ( n6731 & n31061 ) | ( ~n20769 & n31061 ) ;
  assign n31063 = ( ~n6817 & n15708 ) | ( ~n6817 & n31062 ) | ( n15708 & n31062 ) ;
  assign n31064 = ( n19290 & ~n21627 ) | ( n19290 & n31063 ) | ( ~n21627 & n31063 ) ;
  assign n31065 = ( x37 & n14976 ) | ( x37 & n30705 ) | ( n14976 & n30705 ) ;
  assign n31066 = ( n11022 & n11534 ) | ( n11022 & ~n16839 ) | ( n11534 & ~n16839 ) ;
  assign n31069 = n23731 ^ n15799 ^ n7818 ;
  assign n31067 = n21095 ^ n13123 ^ n9236 ;
  assign n31068 = n31067 ^ n18483 ^ n1021 ;
  assign n31070 = n31069 ^ n31068 ^ 1'b0 ;
  assign n31071 = ( ~n2618 & n6083 ) | ( ~n2618 & n23823 ) | ( n6083 & n23823 ) ;
  assign n31072 = ( ~n3221 & n4838 ) | ( ~n3221 & n31071 ) | ( n4838 & n31071 ) ;
  assign n31073 = ( n1464 & n5756 ) | ( n1464 & ~n15833 ) | ( n5756 & ~n15833 ) ;
  assign n31074 = n31073 ^ n5209 ^ n3150 ;
  assign n31075 = ~n3839 & n31074 ;
  assign n31076 = ~n31072 & n31075 ;
  assign n31077 = n13712 ^ n11098 ^ 1'b0 ;
  assign n31078 = n27500 & n31077 ;
  assign n31079 = n12587 ^ n8679 ^ 1'b0 ;
  assign n31080 = n24850 | n31079 ;
  assign n31081 = n28300 ^ n11109 ^ 1'b0 ;
  assign n31082 = ( n2495 & n3566 ) | ( n2495 & n4016 ) | ( n3566 & n4016 ) ;
  assign n31083 = ( ~n2066 & n12372 ) | ( ~n2066 & n31082 ) | ( n12372 & n31082 ) ;
  assign n31084 = n31083 ^ n26718 ^ n2940 ;
  assign n31085 = n31084 ^ n5288 ^ n2231 ;
  assign n31086 = ( n7681 & n8342 ) | ( n7681 & ~n20411 ) | ( n8342 & ~n20411 ) ;
  assign n31087 = n26353 ^ n18507 ^ n7217 ;
  assign n31088 = ( ~n4064 & n15892 ) | ( ~n4064 & n31087 ) | ( n15892 & n31087 ) ;
  assign n31089 = ( n20040 & ~n31086 ) | ( n20040 & n31088 ) | ( ~n31086 & n31088 ) ;
  assign n31090 = n21770 ^ n21344 ^ n1709 ;
  assign n31091 = n31090 ^ n23328 ^ n19842 ;
  assign n31092 = n31091 ^ n11278 ^ n4171 ;
  assign n31093 = n30957 ^ n9258 ^ 1'b0 ;
  assign n31094 = ( ~n5132 & n16147 ) | ( ~n5132 & n17991 ) | ( n16147 & n17991 ) ;
  assign n31095 = n31094 ^ n23209 ^ n1374 ;
  assign n31096 = ( n380 & n5703 ) | ( n380 & ~n14207 ) | ( n5703 & ~n14207 ) ;
  assign n31097 = n11280 ^ n6915 ^ n6075 ;
  assign n31098 = ( ~n24586 & n31096 ) | ( ~n24586 & n31097 ) | ( n31096 & n31097 ) ;
  assign n31099 = n10307 & ~n26493 ;
  assign n31100 = n6570 & n31099 ;
  assign n31101 = ~n9268 & n18837 ;
  assign n31102 = ~n4895 & n31101 ;
  assign n31103 = ( n3149 & n14793 ) | ( n3149 & n31102 ) | ( n14793 & n31102 ) ;
  assign n31106 = ( ~n2997 & n6059 ) | ( ~n2997 & n9913 ) | ( n6059 & n9913 ) ;
  assign n31104 = ( n6371 & n21872 ) | ( n6371 & n25574 ) | ( n21872 & n25574 ) ;
  assign n31105 = ( n17224 & n21437 ) | ( n17224 & n31104 ) | ( n21437 & n31104 ) ;
  assign n31107 = n31106 ^ n31105 ^ n13084 ;
  assign n31108 = ~n2915 & n13156 ;
  assign n31109 = ~n29583 & n31108 ;
  assign n31110 = n6255 ^ n3812 ^ n201 ;
  assign n31111 = ( n720 & n2790 ) | ( n720 & ~n31110 ) | ( n2790 & ~n31110 ) ;
  assign n31112 = ( n7551 & n31109 ) | ( n7551 & n31111 ) | ( n31109 & n31111 ) ;
  assign n31114 = ( n3026 & n15496 ) | ( n3026 & ~n26299 ) | ( n15496 & ~n26299 ) ;
  assign n31113 = n4041 | n12625 ;
  assign n31115 = n31114 ^ n31113 ^ 1'b0 ;
  assign n31116 = ( n21177 & n23456 ) | ( n21177 & ~n31115 ) | ( n23456 & ~n31115 ) ;
  assign n31117 = ( n21306 & ~n25721 ) | ( n21306 & n28640 ) | ( ~n25721 & n28640 ) ;
  assign n31118 = ( ~n7849 & n9959 ) | ( ~n7849 & n31117 ) | ( n9959 & n31117 ) ;
  assign n31119 = n31118 ^ n30922 ^ n25109 ;
  assign n31120 = n22008 ^ n7175 ^ n3586 ;
  assign n31121 = n3726 | n19691 ;
  assign n31122 = n31121 ^ n27861 ^ 1'b0 ;
  assign n31123 = n31122 ^ n24238 ^ n3953 ;
  assign n31124 = n13131 & ~n14922 ;
  assign n31125 = n8575 & n28386 ;
  assign n31126 = n31125 ^ n18363 ^ 1'b0 ;
  assign n31127 = ( n4710 & n7493 ) | ( n4710 & n18117 ) | ( n7493 & n18117 ) ;
  assign n31128 = n31127 ^ n3595 ^ n1380 ;
  assign n31129 = n31128 ^ n29054 ^ 1'b0 ;
  assign n31130 = n4146 & ~n8883 ;
  assign n31131 = ~n3416 & n31130 ;
  assign n31132 = n31131 ^ n18621 ^ n2858 ;
  assign n31133 = ( ~n25041 & n27580 ) | ( ~n25041 & n30364 ) | ( n27580 & n30364 ) ;
  assign n31134 = n3213 & n13114 ;
  assign n31135 = n31134 ^ n15839 ^ n6670 ;
  assign n31136 = ( ~n8250 & n27757 ) | ( ~n8250 & n31135 ) | ( n27757 & n31135 ) ;
  assign n31137 = ( n10541 & n11099 ) | ( n10541 & ~n31136 ) | ( n11099 & ~n31136 ) ;
  assign n31140 = ( n2369 & n3435 ) | ( n2369 & ~n3497 ) | ( n3435 & ~n3497 ) ;
  assign n31141 = ~n4113 & n31140 ;
  assign n31142 = n13412 & n31141 ;
  assign n31143 = n31142 ^ n4486 ^ n2142 ;
  assign n31138 = n16597 | n17144 ;
  assign n31139 = n14130 | n31138 ;
  assign n31144 = n31143 ^ n31139 ^ 1'b0 ;
  assign n31145 = ( n11802 & n13715 ) | ( n11802 & n20419 ) | ( n13715 & n20419 ) ;
  assign n31146 = n11635 ^ n8695 ^ n5454 ;
  assign n31147 = ( n1320 & n1937 ) | ( n1320 & ~n31146 ) | ( n1937 & ~n31146 ) ;
  assign n31148 = ( n1742 & n19698 ) | ( n1742 & n31147 ) | ( n19698 & n31147 ) ;
  assign n31150 = ( n2485 & n4148 ) | ( n2485 & ~n22421 ) | ( n4148 & ~n22421 ) ;
  assign n31149 = ( n1706 & n16195 ) | ( n1706 & ~n19931 ) | ( n16195 & ~n19931 ) ;
  assign n31151 = n31150 ^ n31149 ^ n13944 ;
  assign n31152 = n3968 | n13955 ;
  assign n31153 = n31152 ^ n24185 ^ 1'b0 ;
  assign n31154 = ~n19882 & n27100 ;
  assign n31155 = n12994 & n31154 ;
  assign n31156 = ( n3419 & ~n25593 ) | ( n3419 & n31155 ) | ( ~n25593 & n31155 ) ;
  assign n31157 = n14272 ^ n8826 ^ 1'b0 ;
  assign n31158 = n31156 & n31157 ;
  assign n31159 = n4525 & ~n7249 ;
  assign n31160 = n4620 ^ n3943 ^ 1'b0 ;
  assign n31161 = ( n1538 & n7600 ) | ( n1538 & ~n25890 ) | ( n7600 & ~n25890 ) ;
  assign n31162 = n7503 | n22953 ;
  assign n31163 = n31162 ^ n7199 ^ n6481 ;
  assign n31164 = ( n5889 & n23395 ) | ( n5889 & n26920 ) | ( n23395 & n26920 ) ;
  assign n31165 = n31164 ^ n30885 ^ n30651 ;
  assign n31167 = ( n1901 & n13247 ) | ( n1901 & n20105 ) | ( n13247 & n20105 ) ;
  assign n31168 = n31167 ^ n23071 ^ n12369 ;
  assign n31166 = n16614 ^ n6390 ^ n5306 ;
  assign n31169 = n31168 ^ n31166 ^ n16273 ;
  assign n31170 = n26908 & n31169 ;
  assign n31171 = ( n1253 & n1653 ) | ( n1253 & n30422 ) | ( n1653 & n30422 ) ;
  assign n31172 = n19146 ^ n1025 ^ 1'b0 ;
  assign n31173 = n7145 | n20013 ;
  assign n31174 = n9043 & ~n31173 ;
  assign n31175 = ( n11927 & n31172 ) | ( n11927 & n31174 ) | ( n31172 & n31174 ) ;
  assign n31176 = ( n6255 & n17744 ) | ( n6255 & ~n31175 ) | ( n17744 & ~n31175 ) ;
  assign n31177 = n25189 ^ n21716 ^ n11639 ;
  assign n31178 = n31177 ^ n13173 ^ n10280 ;
  assign n31179 = ( n347 & n3433 ) | ( n347 & n31178 ) | ( n3433 & n31178 ) ;
  assign n31180 = n31179 ^ n13160 ^ n4395 ;
  assign n31181 = n31180 ^ n27554 ^ n9590 ;
  assign n31182 = n31181 ^ n20828 ^ n6801 ;
  assign n31183 = n2346 & n18239 ;
  assign n31184 = ~n1827 & n31183 ;
  assign n31185 = n23583 ^ n7724 ^ n491 ;
  assign n31186 = n31185 ^ n27630 ^ 1'b0 ;
  assign n31187 = n6721 ^ n4885 ^ 1'b0 ;
  assign n31188 = n11436 ^ n6917 ^ 1'b0 ;
  assign n31189 = n6807 | n7905 ;
  assign n31190 = n31189 ^ n5218 ^ 1'b0 ;
  assign n31191 = n31190 ^ n27494 ^ n23525 ;
  assign n31192 = n17405 ^ n17022 ^ n7340 ;
  assign n31193 = ( ~n9450 & n15768 ) | ( ~n9450 & n21649 ) | ( n15768 & n21649 ) ;
  assign n31194 = n7070 | n24605 ;
  assign n31195 = n5926 | n31194 ;
  assign n31196 = n3777 & ~n24043 ;
  assign n31197 = n31196 ^ n24886 ^ 1'b0 ;
  assign n31198 = ( n7153 & n31195 ) | ( n7153 & ~n31197 ) | ( n31195 & ~n31197 ) ;
  assign n31199 = ( n8029 & n17154 ) | ( n8029 & ~n19787 ) | ( n17154 & ~n19787 ) ;
  assign n31200 = n31199 ^ n11477 ^ x64 ;
  assign n31201 = n8014 ^ n7198 ^ n2376 ;
  assign n31202 = n11161 & n17191 ;
  assign n31203 = n21545 ^ n4440 ^ 1'b0 ;
  assign n31204 = n31202 | n31203 ;
  assign n31205 = n20250 ^ n9599 ^ n6647 ;
  assign n31206 = n31205 ^ n3000 ^ 1'b0 ;
  assign n31207 = n5076 & n9828 ;
  assign n31208 = ( ~n7040 & n15201 ) | ( ~n7040 & n31207 ) | ( n15201 & n31207 ) ;
  assign n31209 = ~n3924 & n4964 ;
  assign n31210 = n31209 ^ n451 ^ 1'b0 ;
  assign n31211 = n31210 ^ n8677 ^ n3430 ;
  assign n31212 = ( n796 & n10809 ) | ( n796 & n21737 ) | ( n10809 & n21737 ) ;
  assign n31213 = ( ~n9146 & n15043 ) | ( ~n9146 & n17496 ) | ( n15043 & n17496 ) ;
  assign n31214 = ( n11379 & n31212 ) | ( n11379 & n31213 ) | ( n31212 & n31213 ) ;
  assign n31215 = ( n8847 & n15279 ) | ( n8847 & ~n20760 ) | ( n15279 & ~n20760 ) ;
  assign n31216 = ( n7201 & n27041 ) | ( n7201 & ~n31215 ) | ( n27041 & ~n31215 ) ;
  assign n31217 = n3903 ^ n3407 ^ n2120 ;
  assign n31219 = n6475 & ~n9772 ;
  assign n31220 = n31219 ^ n289 ^ 1'b0 ;
  assign n31221 = n31220 ^ n8900 ^ 1'b0 ;
  assign n31218 = n16455 ^ n11810 ^ n5928 ;
  assign n31222 = n31221 ^ n31218 ^ n24270 ;
  assign n31223 = x112 & ~n4528 ;
  assign n31224 = n31223 ^ n20729 ^ 1'b0 ;
  assign n31225 = n31224 ^ n28502 ^ n9266 ;
  assign n31226 = ( n197 & ~n6887 ) | ( n197 & n25483 ) | ( ~n6887 & n25483 ) ;
  assign n31227 = n31226 ^ n20888 ^ n1350 ;
  assign n31228 = n9082 | n15759 ;
  assign n31229 = n31228 ^ n10378 ^ n1497 ;
  assign n31230 = ~n9616 & n31229 ;
  assign n31231 = n31230 ^ n18718 ^ 1'b0 ;
  assign n31232 = n4659 | n14801 ;
  assign n31233 = n31232 ^ n5026 ^ 1'b0 ;
  assign n31234 = ( n17337 & n21657 ) | ( n17337 & ~n27645 ) | ( n21657 & ~n27645 ) ;
  assign n31235 = ( n3620 & n8822 ) | ( n3620 & n21035 ) | ( n8822 & n21035 ) ;
  assign n31236 = n423 & ~n31235 ;
  assign n31237 = ( ~n17334 & n29963 ) | ( ~n17334 & n31236 ) | ( n29963 & n31236 ) ;
  assign n31238 = ( ~n5734 & n19148 ) | ( ~n5734 & n26336 ) | ( n19148 & n26336 ) ;
  assign n31239 = n8519 ^ n5624 ^ n4102 ;
  assign n31240 = ( n2291 & ~n17256 ) | ( n2291 & n31239 ) | ( ~n17256 & n31239 ) ;
  assign n31241 = n12833 ^ n12380 ^ 1'b0 ;
  assign n31242 = ~n28766 & n31241 ;
  assign n31243 = ( n13832 & n23606 ) | ( n13832 & ~n31242 ) | ( n23606 & ~n31242 ) ;
  assign n31246 = n9286 & n26595 ;
  assign n31247 = n23559 & n31246 ;
  assign n31244 = n17403 ^ n8336 ^ n7011 ;
  assign n31245 = n31244 ^ n10239 ^ n8296 ;
  assign n31248 = n31247 ^ n31245 ^ n3485 ;
  assign n31249 = ( n922 & n1780 ) | ( n922 & ~n8568 ) | ( n1780 & ~n8568 ) ;
  assign n31250 = ~n3560 & n7958 ;
  assign n31251 = n4717 & n31250 ;
  assign n31252 = ( n9864 & n31249 ) | ( n9864 & ~n31251 ) | ( n31249 & ~n31251 ) ;
  assign n31254 = n6904 ^ n5682 ^ n2619 ;
  assign n31253 = n18732 ^ n12019 ^ n5209 ;
  assign n31255 = n31254 ^ n31253 ^ n18166 ;
  assign n31256 = ~n7948 & n26467 ;
  assign n31257 = n31256 ^ n26217 ^ 1'b0 ;
  assign n31258 = n27460 ^ n6702 ^ n445 ;
  assign n31259 = ( n865 & n31257 ) | ( n865 & n31258 ) | ( n31257 & n31258 ) ;
  assign n31260 = n31259 ^ n3997 ^ 1'b0 ;
  assign n31261 = ( n13138 & n16067 ) | ( n13138 & ~n29622 ) | ( n16067 & ~n29622 ) ;
  assign n31262 = n31261 ^ n13626 ^ n2396 ;
  assign n31263 = ( n13117 & n30827 ) | ( n13117 & ~n31262 ) | ( n30827 & ~n31262 ) ;
  assign n31264 = n11578 ^ n7997 ^ 1'b0 ;
  assign n31265 = ( n6460 & n30470 ) | ( n6460 & ~n31264 ) | ( n30470 & ~n31264 ) ;
  assign n31266 = n30831 ^ n9304 ^ n5906 ;
  assign n31267 = n17853 ^ n9930 ^ n8319 ;
  assign n31268 = n8176 & n23021 ;
  assign n31269 = n28529 ^ n24715 ^ n2596 ;
  assign n31270 = ( n10426 & ~n31268 ) | ( n10426 & n31269 ) | ( ~n31268 & n31269 ) ;
  assign n31271 = n25468 ^ n22871 ^ n6150 ;
  assign n31272 = ( n2677 & n6759 ) | ( n2677 & ~n14034 ) | ( n6759 & ~n14034 ) ;
  assign n31273 = n31272 ^ n28548 ^ n15566 ;
  assign n31274 = ~n154 & n2748 ;
  assign n31275 = ~n10979 & n31274 ;
  assign n31276 = n21743 ^ n18006 ^ n9470 ;
  assign n31277 = n31276 ^ n4465 ^ n3105 ;
  assign n31279 = n9935 | n10645 ;
  assign n31278 = n19906 ^ n15825 ^ n1485 ;
  assign n31280 = n31279 ^ n31278 ^ n26092 ;
  assign n31281 = n22873 ^ n19603 ^ n18870 ;
  assign n31282 = ( n191 & ~n12500 ) | ( n191 & n28664 ) | ( ~n12500 & n28664 ) ;
  assign n31283 = ( n6084 & n31281 ) | ( n6084 & ~n31282 ) | ( n31281 & ~n31282 ) ;
  assign n31284 = ( n2093 & ~n2998 ) | ( n2093 & n10998 ) | ( ~n2998 & n10998 ) ;
  assign n31285 = ( n11424 & n17086 ) | ( n11424 & ~n26480 ) | ( n17086 & ~n26480 ) ;
  assign n31293 = n4637 | n9367 ;
  assign n31294 = n6797 | n31293 ;
  assign n31291 = n12670 ^ n5933 ^ 1'b0 ;
  assign n31286 = n25580 ^ n19252 ^ n15888 ;
  assign n31287 = ( n6945 & n13932 ) | ( n6945 & n31286 ) | ( n13932 & n31286 ) ;
  assign n31288 = ~n11867 & n31287 ;
  assign n31289 = ~n5514 & n31288 ;
  assign n31290 = n31289 ^ n23904 ^ n11217 ;
  assign n31292 = n31291 ^ n31290 ^ 1'b0 ;
  assign n31295 = n31294 ^ n31292 ^ n9044 ;
  assign n31296 = ( n5080 & n5489 ) | ( n5080 & n7644 ) | ( n5489 & n7644 ) ;
  assign n31297 = ( n145 & n8165 ) | ( n145 & ~n31296 ) | ( n8165 & ~n31296 ) ;
  assign n31298 = n19104 ^ n9686 ^ n6554 ;
  assign n31299 = ( n2821 & n8970 ) | ( n2821 & ~n31298 ) | ( n8970 & ~n31298 ) ;
  assign n31300 = n2760 ^ n2042 ^ 1'b0 ;
  assign n31301 = n6725 & n13385 ;
  assign n31303 = n15930 ^ n11055 ^ n3170 ;
  assign n31304 = ( n9321 & n9484 ) | ( n9321 & ~n31303 ) | ( n9484 & ~n31303 ) ;
  assign n31305 = ( n3213 & n18044 ) | ( n3213 & ~n31304 ) | ( n18044 & ~n31304 ) ;
  assign n31302 = ~n12512 & n30827 ;
  assign n31306 = n31305 ^ n31302 ^ 1'b0 ;
  assign n31307 = ( n2511 & n8854 ) | ( n2511 & ~n17799 ) | ( n8854 & ~n17799 ) ;
  assign n31308 = n31307 ^ n18440 ^ n896 ;
  assign n31309 = n31308 ^ n30512 ^ n2504 ;
  assign n31310 = ( n17153 & n20255 ) | ( n17153 & n28226 ) | ( n20255 & n28226 ) ;
  assign n31311 = ~n6984 & n14936 ;
  assign n31312 = n31311 ^ n13920 ^ n4101 ;
  assign n31313 = n27296 ^ n17603 ^ 1'b0 ;
  assign n31314 = n1675 ^ n1515 ^ 1'b0 ;
  assign n31315 = ~n1841 & n31314 ;
  assign n31316 = ( n2841 & ~n25267 ) | ( n2841 & n31315 ) | ( ~n25267 & n31315 ) ;
  assign n31317 = n287 & ~n19382 ;
  assign n31318 = ( ~n2637 & n5165 ) | ( ~n2637 & n14125 ) | ( n5165 & n14125 ) ;
  assign n31319 = n15459 ^ n11267 ^ n7804 ;
  assign n31321 = n30655 ^ n21209 ^ n18656 ;
  assign n31320 = n2612 & n26594 ;
  assign n31322 = n31321 ^ n31320 ^ 1'b0 ;
  assign n31323 = n28948 ^ n24032 ^ 1'b0 ;
  assign n31324 = n21594 & ~n31323 ;
  assign n31325 = ( n6863 & n21054 ) | ( n6863 & n24129 ) | ( n21054 & n24129 ) ;
  assign n31326 = ( n3937 & ~n8132 ) | ( n3937 & n16164 ) | ( ~n8132 & n16164 ) ;
  assign n31327 = ( n2355 & n9967 ) | ( n2355 & ~n11973 ) | ( n9967 & ~n11973 ) ;
  assign n31328 = ( n20530 & n23684 ) | ( n20530 & n31327 ) | ( n23684 & n31327 ) ;
  assign n31329 = n14897 ^ n5582 ^ 1'b0 ;
  assign n31330 = ( n2338 & n5696 ) | ( n2338 & n6194 ) | ( n5696 & n6194 ) ;
  assign n31331 = n31330 ^ n26124 ^ n3776 ;
  assign n31332 = ( n11322 & ~n13692 ) | ( n11322 & n20681 ) | ( ~n13692 & n20681 ) ;
  assign n31333 = ( n3182 & n10883 ) | ( n3182 & n26978 ) | ( n10883 & n26978 ) ;
  assign n31334 = n3464 | n7775 ;
  assign n31335 = n31334 ^ n4101 ^ 1'b0 ;
  assign n31336 = n28072 ^ n27616 ^ n18507 ;
  assign n31337 = ( n8129 & n9637 ) | ( n8129 & ~n12474 ) | ( n9637 & ~n12474 ) ;
  assign n31338 = n31337 ^ n25031 ^ n456 ;
  assign n31339 = n31338 ^ n30451 ^ 1'b0 ;
  assign n31340 = ~n9614 & n31339 ;
  assign n31341 = n27689 ^ n17963 ^ 1'b0 ;
  assign n31342 = n11956 & ~n31341 ;
  assign n31343 = n16854 & n31342 ;
  assign n31344 = n31343 ^ n11612 ^ 1'b0 ;
  assign n31345 = ( ~n31336 & n31340 ) | ( ~n31336 & n31344 ) | ( n31340 & n31344 ) ;
  assign n31346 = ( n4491 & ~n9866 ) | ( n4491 & n15995 ) | ( ~n9866 & n15995 ) ;
  assign n31347 = n28122 ^ n19316 ^ n1755 ;
  assign n31348 = ( n2077 & ~n2563 ) | ( n2077 & n9618 ) | ( ~n2563 & n9618 ) ;
  assign n31349 = n31348 ^ n24798 ^ n1152 ;
  assign n31350 = ( n12377 & n19531 ) | ( n12377 & ~n31349 ) | ( n19531 & ~n31349 ) ;
  assign n31351 = n24965 | n30033 ;
  assign n31352 = n28934 ^ n16255 ^ 1'b0 ;
  assign n31353 = n31352 ^ n7860 ^ n5289 ;
  assign n31354 = ( n2478 & n2725 ) | ( n2478 & ~n27927 ) | ( n2725 & ~n27927 ) ;
  assign n31355 = n11745 ^ x124 ^ 1'b0 ;
  assign n31356 = n8588 ^ n8313 ^ n3164 ;
  assign n31357 = n31356 ^ n30365 ^ n5061 ;
  assign n31358 = ( n14445 & n15390 ) | ( n14445 & ~n22634 ) | ( n15390 & ~n22634 ) ;
  assign n31359 = n31357 & n31358 ;
  assign n31360 = n3174 ^ x55 ^ 1'b0 ;
  assign n31361 = n6660 | n31360 ;
  assign n31362 = ( n3917 & n20056 ) | ( n3917 & ~n24414 ) | ( n20056 & ~n24414 ) ;
  assign n31363 = n31362 ^ n7198 ^ 1'b0 ;
  assign n31364 = n1063 | n30190 ;
  assign n31365 = n31005 ^ n23801 ^ n822 ;
  assign n31366 = n856 ^ n752 ^ 1'b0 ;
  assign n31367 = x42 & n31366 ;
  assign n31368 = n31367 ^ n29913 ^ n9787 ;
  assign n31369 = n31368 ^ n5161 ^ 1'b0 ;
  assign n31370 = ( n4472 & n22152 ) | ( n4472 & ~n31369 ) | ( n22152 & ~n31369 ) ;
  assign n31371 = ( n5822 & n26598 ) | ( n5822 & ~n28323 ) | ( n26598 & ~n28323 ) ;
  assign n31372 = ( n3385 & n5885 ) | ( n3385 & ~n21222 ) | ( n5885 & ~n21222 ) ;
  assign n31373 = n25182 ^ n16121 ^ 1'b0 ;
  assign n31374 = ( n3225 & ~n25678 ) | ( n3225 & n31373 ) | ( ~n25678 & n31373 ) ;
  assign n31376 = ( n2921 & n4892 ) | ( n2921 & n7005 ) | ( n4892 & n7005 ) ;
  assign n31375 = ~n7078 & n19835 ;
  assign n31377 = n31376 ^ n31375 ^ 1'b0 ;
  assign n31378 = n15868 ^ n14998 ^ n8234 ;
  assign n31379 = n27414 ^ n1998 ^ 1'b0 ;
  assign n31380 = n31378 & n31379 ;
  assign n31382 = ( n24131 & ~n27591 ) | ( n24131 & n30584 ) | ( ~n27591 & n30584 ) ;
  assign n31381 = n26924 ^ n22594 ^ n6226 ;
  assign n31383 = n31382 ^ n31381 ^ n24103 ;
  assign n31386 = n6060 ^ n799 ^ 1'b0 ;
  assign n31387 = ~n624 & n31386 ;
  assign n31388 = ( n2818 & n4435 ) | ( n2818 & n27611 ) | ( n4435 & n27611 ) ;
  assign n31389 = ( n20638 & ~n31387 ) | ( n20638 & n31388 ) | ( ~n31387 & n31388 ) ;
  assign n31384 = n1911 & ~n3353 ;
  assign n31385 = ~n7397 & n31384 ;
  assign n31390 = n31389 ^ n31385 ^ n7810 ;
  assign n31391 = n23205 ^ n19822 ^ 1'b0 ;
  assign n31392 = n9443 & ~n14059 ;
  assign n31393 = n5860 & n22676 ;
  assign n31394 = ( n869 & n27703 ) | ( n869 & ~n31393 ) | ( n27703 & ~n31393 ) ;
  assign n31395 = n31394 ^ n15741 ^ n1907 ;
  assign n31396 = ( n4208 & n15403 ) | ( n4208 & n15521 ) | ( n15403 & n15521 ) ;
  assign n31397 = n31396 ^ n9303 ^ n4774 ;
  assign n31398 = ( ~n4714 & n8507 ) | ( ~n4714 & n31397 ) | ( n8507 & n31397 ) ;
  assign n31399 = n21532 ^ n13135 ^ n2515 ;
  assign n31400 = ( n4816 & ~n9010 ) | ( n4816 & n22208 ) | ( ~n9010 & n22208 ) ;
  assign n31401 = ~n9864 & n17881 ;
  assign n31402 = n31401 ^ n29286 ^ 1'b0 ;
  assign n31403 = n2861 & ~n23705 ;
  assign n31404 = n31403 ^ n9372 ^ 1'b0 ;
  assign n31405 = ( ~n11638 & n19154 ) | ( ~n11638 & n19375 ) | ( n19154 & n19375 ) ;
  assign n31406 = n20885 & n22583 ;
  assign n31407 = ~n868 & n24610 ;
  assign n31408 = n31406 & n31407 ;
  assign n31409 = ~n31405 & n31408 ;
  assign n31410 = n24379 ^ n12390 ^ n11198 ;
  assign n31411 = ( n5122 & ~n7976 ) | ( n5122 & n10626 ) | ( ~n7976 & n10626 ) ;
  assign n31412 = n31411 ^ n14364 ^ n3878 ;
  assign n31413 = ( n13834 & ~n15042 ) | ( n13834 & n26420 ) | ( ~n15042 & n26420 ) ;
  assign n31414 = ~n7494 & n26243 ;
  assign n31415 = n31414 ^ n16897 ^ n12770 ;
  assign n31416 = n29672 ^ n28176 ^ n3405 ;
  assign n31417 = n31416 ^ n30551 ^ n18053 ;
  assign n31418 = n13838 ^ n11819 ^ n11083 ;
  assign n31419 = n7693 | n31418 ;
  assign n31420 = n30380 ^ n6941 ^ 1'b0 ;
  assign n31421 = n31420 ^ n14108 ^ n7741 ;
  assign n31422 = n30753 ^ n28044 ^ n25905 ;
  assign n31423 = n18961 ^ n2218 ^ 1'b0 ;
  assign n31424 = n31422 | n31423 ;
  assign n31425 = ~n16558 & n21289 ;
  assign n31426 = n18833 & n31425 ;
  assign n31427 = n25293 ^ n17016 ^ n11096 ;
  assign n31428 = n9371 & ~n31427 ;
  assign n31429 = ( n1420 & n9140 ) | ( n1420 & n13824 ) | ( n9140 & n13824 ) ;
  assign n31430 = n8957 ^ n6148 ^ n4323 ;
  assign n31431 = ( n13273 & ~n31429 ) | ( n13273 & n31430 ) | ( ~n31429 & n31430 ) ;
  assign n31432 = ( n11834 & n21606 ) | ( n11834 & n31431 ) | ( n21606 & n31431 ) ;
  assign n31433 = ( n11992 & n14603 ) | ( n11992 & ~n19862 ) | ( n14603 & ~n19862 ) ;
  assign n31434 = ~n612 & n7108 ;
  assign n31435 = n31434 ^ n23460 ^ n20656 ;
  assign n31436 = n22410 ^ n7525 ^ n360 ;
  assign n31437 = n24106 ^ n8753 ^ 1'b0 ;
  assign n31438 = n31436 & ~n31437 ;
  assign n31439 = ( n9416 & n18804 ) | ( n9416 & ~n31438 ) | ( n18804 & ~n31438 ) ;
  assign n31440 = ( n3060 & n5908 ) | ( n3060 & n11653 ) | ( n5908 & n11653 ) ;
  assign n31441 = n25180 ^ n17941 ^ n11787 ;
  assign n31442 = n26685 ^ n8904 ^ n6124 ;
  assign n31443 = n12481 ^ n1144 ^ 1'b0 ;
  assign n31444 = ~n11485 & n31443 ;
  assign n31445 = n1401 & ~n9889 ;
  assign n31446 = n6852 & n31445 ;
  assign n31447 = n25547 | n31446 ;
  assign n31448 = n11918 & ~n31447 ;
  assign n31449 = n22016 ^ n9507 ^ 1'b0 ;
  assign n31450 = ~n23119 & n31449 ;
  assign n31451 = n28516 ^ n10942 ^ n6835 ;
  assign n31452 = n31451 ^ n12889 ^ n321 ;
  assign n31453 = n22937 ^ n20615 ^ n7560 ;
  assign n31454 = n19569 ^ n3093 ^ 1'b0 ;
  assign n31455 = n29875 ^ n3146 ^ 1'b0 ;
  assign n31456 = n31454 & n31455 ;
  assign n31457 = ( n23154 & n31453 ) | ( n23154 & ~n31456 ) | ( n31453 & ~n31456 ) ;
  assign n31458 = ( n4350 & n8220 ) | ( n4350 & n31457 ) | ( n8220 & n31457 ) ;
  assign n31459 = n7730 ^ n4494 ^ n954 ;
  assign n31460 = n31459 ^ n23473 ^ n22455 ;
  assign n31461 = n24837 ^ n9772 ^ 1'b0 ;
  assign n31462 = n12631 & ~n31461 ;
  assign n31463 = n31462 ^ n15770 ^ n7397 ;
  assign n31464 = ( ~n5141 & n11750 ) | ( ~n5141 & n31463 ) | ( n11750 & n31463 ) ;
  assign n31465 = n11559 & ~n30047 ;
  assign n31466 = n25681 | n31465 ;
  assign n31467 = n27136 ^ n14532 ^ n7849 ;
  assign n31468 = ( n3559 & n14922 ) | ( n3559 & n28453 ) | ( n14922 & n28453 ) ;
  assign n31469 = ( n3084 & ~n31467 ) | ( n3084 & n31468 ) | ( ~n31467 & n31468 ) ;
  assign n31470 = n31469 ^ n15467 ^ 1'b0 ;
  assign n31471 = n5182 & ~n5799 ;
  assign n31472 = n31471 ^ n10265 ^ 1'b0 ;
  assign n31473 = ( n16318 & n19739 ) | ( n16318 & ~n31472 ) | ( n19739 & ~n31472 ) ;
  assign n31474 = ( ~n3926 & n29453 ) | ( ~n3926 & n31473 ) | ( n29453 & n31473 ) ;
  assign n31475 = n14516 ^ n6654 ^ n1380 ;
  assign n31476 = n26571 ^ n18532 ^ 1'b0 ;
  assign n31477 = n9998 & n31476 ;
  assign n31478 = n9891 ^ n6635 ^ n759 ;
  assign n31479 = n31478 ^ n9461 ^ 1'b0 ;
  assign n31480 = ~n22598 & n31479 ;
  assign n31481 = n17208 ^ n6226 ^ n2310 ;
  assign n31482 = ( n13498 & n26003 ) | ( n13498 & n31481 ) | ( n26003 & n31481 ) ;
  assign n31483 = n31482 ^ n13359 ^ n554 ;
  assign n31484 = ( n3115 & n12852 ) | ( n3115 & ~n21971 ) | ( n12852 & ~n21971 ) ;
  assign n31485 = n16822 ^ n10946 ^ n7241 ;
  assign n31486 = n31485 ^ n25499 ^ n580 ;
  assign n31487 = n11949 ^ n8988 ^ n1527 ;
  assign n31488 = n31487 ^ n12730 ^ n296 ;
  assign n31489 = n12032 & ~n15040 ;
  assign n31490 = n31488 & n31489 ;
  assign n31491 = n22047 ^ n11994 ^ 1'b0 ;
  assign n31492 = ~n31490 & n31491 ;
  assign n31493 = ( n12705 & n14579 ) | ( n12705 & n31492 ) | ( n14579 & n31492 ) ;
  assign n31495 = n16505 ^ n2170 ^ x72 ;
  assign n31494 = n20785 ^ n18256 ^ n10772 ;
  assign n31496 = n31495 ^ n31494 ^ n25366 ;
  assign n31499 = n20273 ^ n8410 ^ n652 ;
  assign n31500 = n1967 & n11786 ;
  assign n31501 = ~n31499 & n31500 ;
  assign n31502 = n2049 | n31501 ;
  assign n31497 = n9113 | n21132 ;
  assign n31498 = n12456 | n31497 ;
  assign n31503 = n31502 ^ n31498 ^ n28515 ;
  assign n31509 = n18665 ^ n4688 ^ n2023 ;
  assign n31506 = ( ~n4218 & n5175 ) | ( ~n4218 & n10987 ) | ( n5175 & n10987 ) ;
  assign n31507 = ( n3967 & n23891 ) | ( n3967 & ~n31506 ) | ( n23891 & ~n31506 ) ;
  assign n31508 = n31507 ^ n23781 ^ n3279 ;
  assign n31504 = n1409 | n23879 ;
  assign n31505 = n31504 ^ n20015 ^ 1'b0 ;
  assign n31510 = n31509 ^ n31508 ^ n31505 ;
  assign n31511 = n21144 ^ n17024 ^ n10761 ;
  assign n31512 = n1633 | n19148 ;
  assign n31513 = n1551 | n31512 ;
  assign n31514 = ( ~n2706 & n11895 ) | ( ~n2706 & n28036 ) | ( n11895 & n28036 ) ;
  assign n31515 = ( n8275 & ~n12656 ) | ( n8275 & n22208 ) | ( ~n12656 & n22208 ) ;
  assign n31516 = ( n2293 & n13715 ) | ( n2293 & ~n25047 ) | ( n13715 & ~n25047 ) ;
  assign n31517 = n31516 ^ n12682 ^ n1822 ;
  assign n31518 = ( n2299 & n15334 ) | ( n2299 & ~n18934 ) | ( n15334 & ~n18934 ) ;
  assign n31519 = ( n2733 & n5733 ) | ( n2733 & n31518 ) | ( n5733 & n31518 ) ;
  assign n31520 = n19273 ^ n17321 ^ 1'b0 ;
  assign n31521 = ( n12643 & ~n21988 ) | ( n12643 & n30948 ) | ( ~n21988 & n30948 ) ;
  assign n31522 = n685 & n12185 ;
  assign n31523 = ( ~n13420 & n29823 ) | ( ~n13420 & n31522 ) | ( n29823 & n31522 ) ;
  assign n31524 = n21427 ^ n14568 ^ 1'b0 ;
  assign n31525 = n4471 & n31524 ;
  assign n31526 = n2425 & ~n7449 ;
  assign n31527 = n31526 ^ n3640 ^ 1'b0 ;
  assign n31528 = ~n10056 & n31527 ;
  assign n31529 = ( n8658 & n9328 ) | ( n8658 & n11664 ) | ( n9328 & n11664 ) ;
  assign n31530 = n12113 ^ n6281 ^ n5006 ;
  assign n31531 = ( n13813 & n28640 ) | ( n13813 & n31530 ) | ( n28640 & n31530 ) ;
  assign n31532 = n31531 ^ n29170 ^ n9652 ;
  assign n31533 = ( ~n2132 & n6548 ) | ( ~n2132 & n12659 ) | ( n6548 & n12659 ) ;
  assign n31534 = ( n9253 & ~n9614 ) | ( n9253 & n14310 ) | ( ~n9614 & n14310 ) ;
  assign n31535 = n31534 ^ n17300 ^ n12308 ;
  assign n31536 = n31535 ^ n22555 ^ 1'b0 ;
  assign n31537 = n31533 & n31536 ;
  assign n31538 = ( n17308 & ~n31532 ) | ( n17308 & n31537 ) | ( ~n31532 & n31537 ) ;
  assign n31539 = ( ~n3230 & n7051 ) | ( ~n3230 & n7654 ) | ( n7051 & n7654 ) ;
  assign n31540 = n12905 ^ n10695 ^ 1'b0 ;
  assign n31541 = n11170 & ~n31540 ;
  assign n31542 = ( n19778 & n20833 ) | ( n19778 & n29750 ) | ( n20833 & n29750 ) ;
  assign n31543 = ( ~n8515 & n9214 ) | ( ~n8515 & n29522 ) | ( n9214 & n29522 ) ;
  assign n31544 = n1959 & n17219 ;
  assign n31545 = n15968 & n31544 ;
  assign n31546 = ( n8451 & n31543 ) | ( n8451 & n31545 ) | ( n31543 & n31545 ) ;
  assign n31547 = ( ~n4271 & n7309 ) | ( ~n4271 & n16501 ) | ( n7309 & n16501 ) ;
  assign n31548 = ( n17410 & n17937 ) | ( n17410 & n31547 ) | ( n17937 & n31547 ) ;
  assign n31549 = n28800 ^ n25364 ^ n19915 ;
  assign n31550 = ( n29387 & n31548 ) | ( n29387 & n31549 ) | ( n31548 & n31549 ) ;
  assign n31551 = n28937 ^ n7792 ^ 1'b0 ;
  assign n31552 = x114 & ~n18920 ;
  assign n31553 = n31552 ^ n10766 ^ 1'b0 ;
  assign n31554 = n20311 ^ n19494 ^ n986 ;
  assign n31555 = n31554 ^ n21018 ^ n17133 ;
  assign n31556 = n31555 ^ n27681 ^ n14026 ;
  assign n31557 = n23772 ^ n6380 ^ 1'b0 ;
  assign n31558 = ~n6358 & n31557 ;
  assign n31559 = n6702 ^ n881 ^ 1'b0 ;
  assign n31560 = ~n17924 & n29769 ;
  assign n31561 = n31559 & n31560 ;
  assign n31562 = ( n21698 & n31558 ) | ( n21698 & ~n31561 ) | ( n31558 & ~n31561 ) ;
  assign n31563 = ( n23518 & n28119 ) | ( n23518 & n31562 ) | ( n28119 & n31562 ) ;
  assign n31564 = n4764 ^ n4162 ^ 1'b0 ;
  assign n31565 = n31564 ^ n6071 ^ n4771 ;
  assign n31566 = ~n11990 & n13471 ;
  assign n31567 = n8994 & n31566 ;
  assign n31568 = n31567 ^ n25405 ^ n19408 ;
  assign n31569 = ( n6965 & ~n31565 ) | ( n6965 & n31568 ) | ( ~n31565 & n31568 ) ;
  assign n31570 = n29655 ^ n2893 ^ 1'b0 ;
  assign n31571 = ~n7788 & n10860 ;
  assign n31572 = n14040 ^ n12342 ^ n5733 ;
  assign n31573 = n9650 ^ n4300 ^ 1'b0 ;
  assign n31574 = n10751 | n31573 ;
  assign n31575 = n25439 ^ n22718 ^ n5799 ;
  assign n31576 = ( n22473 & ~n31574 ) | ( n22473 & n31575 ) | ( ~n31574 & n31575 ) ;
  assign n31577 = ( n19685 & n23824 ) | ( n19685 & ~n31576 ) | ( n23824 & ~n31576 ) ;
  assign n31578 = ( n20622 & ~n25929 ) | ( n20622 & n30848 ) | ( ~n25929 & n30848 ) ;
  assign n31579 = ( ~n3244 & n16745 ) | ( ~n3244 & n31578 ) | ( n16745 & n31578 ) ;
  assign n31580 = ( n7956 & ~n18968 ) | ( n7956 & n26244 ) | ( ~n18968 & n26244 ) ;
  assign n31581 = n3972 & n9518 ;
  assign n31582 = ( n3449 & n13415 ) | ( n3449 & ~n31581 ) | ( n13415 & ~n31581 ) ;
  assign n31583 = n31582 ^ n12645 ^ 1'b0 ;
  assign n31584 = n31580 & n31583 ;
  assign n31585 = ( ~n5146 & n20820 ) | ( ~n5146 & n21227 ) | ( n20820 & n21227 ) ;
  assign n31586 = n5253 & ~n31585 ;
  assign n31587 = ( n2405 & n24685 ) | ( n2405 & ~n31586 ) | ( n24685 & ~n31586 ) ;
  assign n31588 = n7444 ^ n5107 ^ n4648 ;
  assign n31589 = n4521 | n31588 ;
  assign n31590 = n31587 | n31589 ;
  assign n31591 = n24897 ^ n8810 ^ n1952 ;
  assign n31592 = n4355 ^ n4190 ^ n854 ;
  assign n31593 = n31592 ^ n16644 ^ n3782 ;
  assign n31594 = ~n10617 & n15483 ;
  assign n31595 = ~n31593 & n31594 ;
  assign n31596 = ( n1959 & n4837 ) | ( n1959 & n31595 ) | ( n4837 & n31595 ) ;
  assign n31597 = ( n10101 & ~n13774 ) | ( n10101 & n15234 ) | ( ~n13774 & n15234 ) ;
  assign n31598 = n10691 & n27190 ;
  assign n31603 = n22207 ^ n9067 ^ n3442 ;
  assign n31602 = ( ~n436 & n16189 ) | ( ~n436 & n20094 ) | ( n16189 & n20094 ) ;
  assign n31599 = ( ~n7607 & n9577 ) | ( ~n7607 & n19724 ) | ( n9577 & n19724 ) ;
  assign n31600 = n595 | n9977 ;
  assign n31601 = ( n6422 & n31599 ) | ( n6422 & ~n31600 ) | ( n31599 & ~n31600 ) ;
  assign n31604 = n31603 ^ n31602 ^ n31601 ;
  assign n31605 = n26997 ^ n12180 ^ n11699 ;
  assign n31606 = n31605 ^ n8156 ^ 1'b0 ;
  assign n31607 = ( n4158 & ~n9257 ) | ( n4158 & n19083 ) | ( ~n9257 & n19083 ) ;
  assign n31608 = ( n404 & n18148 ) | ( n404 & n22410 ) | ( n18148 & n22410 ) ;
  assign n31609 = n26589 ^ n11020 ^ 1'b0 ;
  assign n31610 = n25878 & n31609 ;
  assign n31611 = n6018 | n27141 ;
  assign n31612 = n23851 | n31611 ;
  assign n31613 = n19434 ^ n7719 ^ 1'b0 ;
  assign n31614 = ~n25419 & n31613 ;
  assign n31615 = ( ~n5660 & n10892 ) | ( ~n5660 & n16799 ) | ( n10892 & n16799 ) ;
  assign n31616 = n12268 ^ n10734 ^ n9686 ;
  assign n31617 = n16898 | n20839 ;
  assign n31618 = n10784 & n16174 ;
  assign n31619 = n18138 & n31618 ;
  assign n31620 = ( n13357 & n23207 ) | ( n13357 & n31619 ) | ( n23207 & n31619 ) ;
  assign n31621 = n20245 & n29475 ;
  assign n31622 = ~n8844 & n16033 ;
  assign n31623 = n22364 ^ n7902 ^ 1'b0 ;
  assign n31624 = ( n31576 & ~n31622 ) | ( n31576 & n31623 ) | ( ~n31622 & n31623 ) ;
  assign n31625 = n26910 ^ n19102 ^ n16380 ;
  assign n31626 = n18196 ^ n4387 ^ 1'b0 ;
  assign n31627 = ( n26202 & n28739 ) | ( n26202 & n31626 ) | ( n28739 & n31626 ) ;
  assign n31628 = n2845 | n11384 ;
  assign n31629 = n31628 ^ n8670 ^ 1'b0 ;
  assign n31630 = ~n1160 & n31629 ;
  assign n31631 = n28835 & n31630 ;
  assign n31632 = ( n4368 & n9646 ) | ( n4368 & n28966 ) | ( n9646 & n28966 ) ;
  assign n31633 = n27220 ^ n14725 ^ n5924 ;
  assign n31634 = n31420 ^ n10048 ^ 1'b0 ;
  assign n31635 = ( ~n1071 & n16977 ) | ( ~n1071 & n29035 ) | ( n16977 & n29035 ) ;
  assign n31636 = n20721 ^ n10464 ^ n5360 ;
  assign n31637 = n6736 & n9552 ;
  assign n31638 = ( n4861 & n18799 ) | ( n4861 & n31637 ) | ( n18799 & n31637 ) ;
  assign n31639 = ~n1697 & n15281 ;
  assign n31640 = n833 & n15866 ;
  assign n31641 = n20936 & n31640 ;
  assign n31642 = n6205 & ~n31641 ;
  assign n31643 = n18619 & n31642 ;
  assign n31644 = ( n6315 & n12270 ) | ( n6315 & n12637 ) | ( n12270 & n12637 ) ;
  assign n31645 = n11757 ^ n5813 ^ 1'b0 ;
  assign n31646 = ~n31644 & n31645 ;
  assign n31647 = ( ~n10927 & n31643 ) | ( ~n10927 & n31646 ) | ( n31643 & n31646 ) ;
  assign n31648 = ~n11253 & n31352 ;
  assign n31649 = n6244 & n31648 ;
  assign n31650 = ( n332 & ~n1388 ) | ( n332 & n20157 ) | ( ~n1388 & n20157 ) ;
  assign n31651 = n3475 | n31650 ;
  assign n31652 = n3340 | n31651 ;
  assign n31653 = n28325 ^ n10727 ^ 1'b0 ;
  assign n31654 = ( n14205 & n14367 ) | ( n14205 & ~n20662 ) | ( n14367 & ~n20662 ) ;
  assign n31655 = n17374 ^ n3944 ^ 1'b0 ;
  assign n31656 = n31655 ^ n20862 ^ n10089 ;
  assign n31657 = ( n6967 & n12074 ) | ( n6967 & n12611 ) | ( n12074 & n12611 ) ;
  assign n31658 = n9051 | n12237 ;
  assign n31659 = n6493 & ~n31658 ;
  assign n31660 = ( ~n13750 & n31657 ) | ( ~n13750 & n31659 ) | ( n31657 & n31659 ) ;
  assign n31661 = n27614 ^ n13088 ^ n6571 ;
  assign n31662 = ( n14568 & ~n17169 ) | ( n14568 & n30933 ) | ( ~n17169 & n30933 ) ;
  assign n31663 = n29228 ^ n12427 ^ n8121 ;
  assign n31664 = n31663 ^ n7967 ^ n6067 ;
  assign n31665 = n24144 & n31094 ;
  assign n31666 = n29766 & n30769 ;
  assign n31667 = ~n10580 & n31666 ;
  assign n31668 = n12804 & ~n17730 ;
  assign n31669 = ~n3508 & n31668 ;
  assign n31670 = n10155 ^ n6439 ^ n5773 ;
  assign n31671 = ( n2297 & ~n4091 ) | ( n2297 & n13552 ) | ( ~n4091 & n13552 ) ;
  assign n31672 = n20676 ^ n13113 ^ n10062 ;
  assign n31673 = ( n31670 & ~n31671 ) | ( n31670 & n31672 ) | ( ~n31671 & n31672 ) ;
  assign n31674 = ~n6356 & n10589 ;
  assign n31675 = n31674 ^ n16442 ^ n5709 ;
  assign n31676 = n31675 ^ n8811 ^ 1'b0 ;
  assign n31677 = n9545 ^ n3967 ^ n947 ;
  assign n31678 = ~n1361 & n6345 ;
  assign n31679 = ( n12918 & n28550 ) | ( n12918 & ~n31678 ) | ( n28550 & ~n31678 ) ;
  assign n31680 = n3218 & ~n5614 ;
  assign n31681 = n31680 ^ n25538 ^ 1'b0 ;
  assign n31682 = ( n15229 & n26322 ) | ( n15229 & ~n31681 ) | ( n26322 & ~n31681 ) ;
  assign n31683 = n9240 ^ n1165 ^ 1'b0 ;
  assign n31684 = n9212 & n31683 ;
  assign n31685 = ( n2402 & n15689 ) | ( n2402 & ~n31684 ) | ( n15689 & ~n31684 ) ;
  assign n31686 = ( n8825 & ~n19000 ) | ( n8825 & n20764 ) | ( ~n19000 & n20764 ) ;
  assign n31687 = ( n5962 & n28261 ) | ( n5962 & ~n31686 ) | ( n28261 & ~n31686 ) ;
  assign n31688 = n24883 ^ n18130 ^ 1'b0 ;
  assign n31689 = ( n22790 & n25774 ) | ( n22790 & n31688 ) | ( n25774 & n31688 ) ;
  assign n31690 = n7902 & ~n12956 ;
  assign n31691 = ~n2709 & n31690 ;
  assign n31692 = n2047 & ~n9447 ;
  assign n31693 = n8925 & n31692 ;
  assign n31694 = n25445 | n31693 ;
  assign n31695 = n31694 ^ n12770 ^ 1'b0 ;
  assign n31696 = n3060 | n8012 ;
  assign n31697 = n31696 ^ n7215 ^ 1'b0 ;
  assign n31698 = n18893 ^ n15636 ^ n683 ;
  assign n31699 = n31698 ^ n11912 ^ 1'b0 ;
  assign n31700 = ( n5981 & n15833 ) | ( n5981 & n31699 ) | ( n15833 & n31699 ) ;
  assign n31701 = n31700 ^ n30471 ^ n3635 ;
  assign n31702 = n31701 ^ n20024 ^ n7236 ;
  assign n31703 = n28687 ^ n2789 ^ 1'b0 ;
  assign n31704 = n30632 ^ n5073 ^ n2810 ;
  assign n31705 = n31704 ^ n11306 ^ n7622 ;
  assign n31706 = ( ~n6989 & n20442 ) | ( ~n6989 & n31705 ) | ( n20442 & n31705 ) ;
  assign n31707 = n28468 ^ n25543 ^ 1'b0 ;
  assign n31708 = n5578 ^ n4014 ^ 1'b0 ;
  assign n31709 = n31708 ^ n29215 ^ n253 ;
  assign n31710 = n8472 & ~n8785 ;
  assign n31711 = ~n9817 & n31710 ;
  assign n31712 = ( n2010 & ~n2532 ) | ( n2010 & n31711 ) | ( ~n2532 & n31711 ) ;
  assign n31713 = n3042 & ~n12883 ;
  assign n31714 = ( ~n2234 & n16422 ) | ( ~n2234 & n31713 ) | ( n16422 & n31713 ) ;
  assign n31715 = n22845 ^ n18075 ^ n14364 ;
  assign n31716 = n31715 ^ n7945 ^ 1'b0 ;
  assign n31719 = n19668 ^ n11255 ^ n5088 ;
  assign n31717 = n25985 ^ n21513 ^ n12746 ;
  assign n31718 = ~n7036 & n31717 ;
  assign n31720 = n31719 ^ n31718 ^ 1'b0 ;
  assign n31721 = n1709 | n4089 ;
  assign n31722 = n3542 & ~n31721 ;
  assign n31723 = ( n19829 & ~n28675 ) | ( n19829 & n31722 ) | ( ~n28675 & n31722 ) ;
  assign n31724 = n31723 ^ n22347 ^ n3407 ;
  assign n31725 = n26784 ^ n26047 ^ n11845 ;
  assign n31726 = ( n3563 & n10327 ) | ( n3563 & ~n15341 ) | ( n10327 & ~n15341 ) ;
  assign n31727 = n31726 ^ n2653 ^ 1'b0 ;
  assign n31728 = n11607 ^ n3057 ^ n1919 ;
  assign n31729 = n31728 ^ n4344 ^ n3576 ;
  assign n31730 = ( ~n7903 & n20529 ) | ( ~n7903 & n23463 ) | ( n20529 & n23463 ) ;
  assign n31731 = n29792 ^ n15392 ^ n14747 ;
  assign n31732 = ( ~n3356 & n23190 ) | ( ~n3356 & n24480 ) | ( n23190 & n24480 ) ;
  assign n31733 = n5730 | n9545 ;
  assign n31734 = n1004 & ~n31733 ;
  assign n31735 = n31734 ^ n5304 ^ 1'b0 ;
  assign n31736 = n25544 | n31735 ;
  assign n31737 = n26183 ^ n6119 ^ 1'b0 ;
  assign n31738 = n31736 | n31737 ;
  assign n31739 = ( n12961 & n17374 ) | ( n12961 & ~n18106 ) | ( n17374 & ~n18106 ) ;
  assign n31740 = n31739 ^ n4911 ^ 1'b0 ;
  assign n31741 = n3964 ^ n2137 ^ 1'b0 ;
  assign n31742 = n31741 ^ n4153 ^ 1'b0 ;
  assign n31743 = n20643 | n31742 ;
  assign n31744 = ( n6024 & ~n8678 ) | ( n6024 & n29536 ) | ( ~n8678 & n29536 ) ;
  assign n31745 = n388 | n2372 ;
  assign n31746 = n31745 ^ n24724 ^ n17140 ;
  assign n31747 = ~n7326 & n19458 ;
  assign n31748 = n13345 & ~n19073 ;
  assign n31749 = ~n31747 & n31748 ;
  assign n31750 = n25297 & ~n31749 ;
  assign n31751 = n9265 | n17391 ;
  assign n31752 = ( n6506 & n27438 ) | ( n6506 & n31751 ) | ( n27438 & n31751 ) ;
  assign n31753 = n22965 ^ n9059 ^ n5573 ;
  assign n31754 = ( n13378 & n31752 ) | ( n13378 & ~n31753 ) | ( n31752 & ~n31753 ) ;
  assign n31755 = n282 & ~n17878 ;
  assign n31756 = n31755 ^ n27440 ^ 1'b0 ;
  assign n31757 = ( n16462 & n17474 ) | ( n16462 & ~n31756 ) | ( n17474 & ~n31756 ) ;
  assign n31758 = ( ~n1745 & n21784 ) | ( ~n1745 & n31340 ) | ( n21784 & n31340 ) ;
  assign n31759 = ( n308 & n2934 ) | ( n308 & n11696 ) | ( n2934 & n11696 ) ;
  assign n31760 = ( ~n8375 & n17363 ) | ( ~n8375 & n31759 ) | ( n17363 & n31759 ) ;
  assign n31761 = n22073 ^ n7985 ^ n1265 ;
  assign n31762 = n31761 ^ n25926 ^ n22978 ;
  assign n31763 = n23766 ^ n16667 ^ 1'b0 ;
  assign n31764 = n13811 & n31763 ;
  assign n31765 = ( n645 & n6123 ) | ( n645 & n29799 ) | ( n6123 & n29799 ) ;
  assign n31766 = n31765 ^ n9728 ^ 1'b0 ;
  assign n31767 = n10813 ^ n5640 ^ n2660 ;
  assign n31768 = n31767 ^ n21125 ^ n10347 ;
  assign n31769 = n31768 ^ n15338 ^ 1'b0 ;
  assign n31770 = n22525 ^ n10838 ^ n5476 ;
  assign n31771 = n10170 & n21355 ;
  assign n31772 = ( ~n5630 & n24853 ) | ( ~n5630 & n29987 ) | ( n24853 & n29987 ) ;
  assign n31773 = n8084 ^ n6091 ^ n5484 ;
  assign n31776 = ( ~n3915 & n5559 ) | ( ~n3915 & n8282 ) | ( n5559 & n8282 ) ;
  assign n31777 = ( n5310 & n13507 ) | ( n5310 & ~n31776 ) | ( n13507 & ~n31776 ) ;
  assign n31778 = ( n530 & n4914 ) | ( n530 & ~n31777 ) | ( n4914 & ~n31777 ) ;
  assign n31774 = ( n9960 & n13283 ) | ( n9960 & ~n19690 ) | ( n13283 & ~n19690 ) ;
  assign n31775 = ( ~n17934 & n18584 ) | ( ~n17934 & n31774 ) | ( n18584 & n31774 ) ;
  assign n31779 = n31778 ^ n31775 ^ n24244 ;
  assign n31780 = n15867 ^ n2050 ^ n277 ;
  assign n31781 = ( n9434 & n11595 ) | ( n9434 & ~n19922 ) | ( n11595 & ~n19922 ) ;
  assign n31782 = ( n1822 & n15802 ) | ( n1822 & n31781 ) | ( n15802 & n31781 ) ;
  assign n31783 = n31782 ^ n27775 ^ n11016 ;
  assign n31784 = n7754 & n13688 ;
  assign n31785 = ~n9942 & n31784 ;
  assign n31786 = ( n7620 & n11645 ) | ( n7620 & ~n16885 ) | ( n11645 & ~n16885 ) ;
  assign n31787 = n21108 ^ n14795 ^ n9005 ;
  assign n31788 = ( n7796 & ~n31786 ) | ( n7796 & n31787 ) | ( ~n31786 & n31787 ) ;
  assign n31789 = n1228 & ~n18475 ;
  assign n31790 = n31788 & n31789 ;
  assign n31791 = n7389 ^ n5290 ^ 1'b0 ;
  assign n31792 = n7399 & n31791 ;
  assign n31793 = n29430 ^ n19544 ^ 1'b0 ;
  assign n31794 = ( ~n244 & n3259 ) | ( ~n244 & n20418 ) | ( n3259 & n20418 ) ;
  assign n31795 = n30954 ^ n10749 ^ 1'b0 ;
  assign n31796 = ( n5683 & n18342 ) | ( n5683 & n19780 ) | ( n18342 & n19780 ) ;
  assign n31797 = n14515 ^ n12745 ^ 1'b0 ;
  assign n31798 = ( ~n16765 & n17467 ) | ( ~n16765 & n18656 ) | ( n17467 & n18656 ) ;
  assign n31799 = ( n2901 & n3867 ) | ( n2901 & n14063 ) | ( n3867 & n14063 ) ;
  assign n31800 = ( ~n11038 & n31798 ) | ( ~n11038 & n31799 ) | ( n31798 & n31799 ) ;
  assign n31801 = n9058 ^ n8321 ^ 1'b0 ;
  assign n31802 = n8302 | n31801 ;
  assign n31803 = ( n31797 & n31800 ) | ( n31797 & ~n31802 ) | ( n31800 & ~n31802 ) ;
  assign n31804 = n24903 ^ n10669 ^ 1'b0 ;
  assign n31805 = ( n10795 & n18034 ) | ( n10795 & n31804 ) | ( n18034 & n31804 ) ;
  assign n31806 = ( n528 & ~n1826 ) | ( n528 & n2770 ) | ( ~n1826 & n2770 ) ;
  assign n31807 = n31487 ^ n27863 ^ n14842 ;
  assign n31808 = ( ~n2702 & n24277 ) | ( ~n2702 & n31807 ) | ( n24277 & n31807 ) ;
  assign n31809 = n31073 ^ n4799 ^ 1'b0 ;
  assign n31810 = n16238 | n31809 ;
  assign n31811 = n15689 ^ n325 ^ 1'b0 ;
  assign n31812 = ~n9417 & n31811 ;
  assign n31813 = ( n8798 & n9726 ) | ( n8798 & n27582 ) | ( n9726 & n27582 ) ;
  assign n31814 = ( n3823 & n13507 ) | ( n3823 & ~n31813 ) | ( n13507 & ~n31813 ) ;
  assign n31815 = n5367 & ~n24993 ;
  assign n31817 = n23795 ^ n17598 ^ n16186 ;
  assign n31816 = n10622 ^ n7963 ^ n7429 ;
  assign n31818 = n31817 ^ n31816 ^ n11664 ;
  assign n31819 = ( n20579 & n23009 ) | ( n20579 & n31150 ) | ( n23009 & n31150 ) ;
  assign n31820 = ( n4080 & n6649 ) | ( n4080 & n16906 ) | ( n6649 & n16906 ) ;
  assign n31821 = n752 & ~n5005 ;
  assign n31822 = ( n28500 & n31820 ) | ( n28500 & n31821 ) | ( n31820 & n31821 ) ;
  assign n31823 = ( n915 & n5388 ) | ( n915 & ~n17580 ) | ( n5388 & ~n17580 ) ;
  assign n31824 = n19093 ^ n11681 ^ 1'b0 ;
  assign n31825 = n22518 | n31824 ;
  assign n31826 = n18985 | n31825 ;
  assign n31827 = n31826 ^ n8265 ^ 1'b0 ;
  assign n31828 = ( n5023 & n16186 ) | ( n5023 & ~n31827 ) | ( n16186 & ~n31827 ) ;
  assign n31829 = n31828 ^ n28183 ^ n2717 ;
  assign n31830 = ( x26 & n1357 ) | ( x26 & n4962 ) | ( n1357 & n4962 ) ;
  assign n31831 = n31830 ^ n3344 ^ 1'b0 ;
  assign n31832 = n21245 | n31831 ;
  assign n31833 = ( n3670 & n5656 ) | ( n3670 & n8237 ) | ( n5656 & n8237 ) ;
  assign n31834 = ~n13601 & n31833 ;
  assign n31835 = ~n27383 & n31834 ;
  assign n31836 = n24053 ^ n14627 ^ n8888 ;
  assign n31839 = n19683 ^ n6868 ^ n3135 ;
  assign n31840 = n31839 ^ n14665 ^ n2536 ;
  assign n31837 = ( n2709 & n9772 ) | ( n2709 & ~n14382 ) | ( n9772 & ~n14382 ) ;
  assign n31838 = ( n1125 & n2380 ) | ( n1125 & n31837 ) | ( n2380 & n31837 ) ;
  assign n31841 = n31840 ^ n31838 ^ n1121 ;
  assign n31842 = n13857 ^ n432 ^ 1'b0 ;
  assign n31843 = ( n3047 & ~n16139 ) | ( n3047 & n31842 ) | ( ~n16139 & n31842 ) ;
  assign n31844 = ( n16686 & n22489 ) | ( n16686 & n31843 ) | ( n22489 & n31843 ) ;
  assign n31845 = ( ~n1790 & n22711 ) | ( ~n1790 & n31844 ) | ( n22711 & n31844 ) ;
  assign n31846 = n22715 ^ n18192 ^ n8563 ;
  assign n31847 = n22348 & n31846 ;
  assign n31848 = n31118 ^ n12949 ^ n9532 ;
  assign n31849 = ( n14821 & n21976 ) | ( n14821 & n25321 ) | ( n21976 & n25321 ) ;
  assign n31850 = ( n1481 & ~n30178 ) | ( n1481 & n31849 ) | ( ~n30178 & n31849 ) ;
  assign n31851 = n26832 ^ n20031 ^ n4839 ;
  assign n31852 = n1460 & n30296 ;
  assign n31853 = n31852 ^ n10394 ^ 1'b0 ;
  assign n31854 = n31853 ^ n16083 ^ n5181 ;
  assign n31855 = ~n6036 & n27980 ;
  assign n31856 = n31855 ^ n27728 ^ 1'b0 ;
  assign n31857 = n2171 ^ n1053 ^ 1'b0 ;
  assign n31858 = ~n8041 & n31857 ;
  assign n31859 = n5056 ^ n2365 ^ 1'b0 ;
  assign n31860 = n22328 ^ n19599 ^ n404 ;
  assign n31861 = n31860 ^ n24506 ^ n21021 ;
  assign n31862 = n25427 ^ n15381 ^ n12442 ;
  assign n31863 = ( n15020 & n15671 ) | ( n15020 & ~n31862 ) | ( n15671 & ~n31862 ) ;
  assign n31864 = ( ~n9392 & n9817 ) | ( ~n9392 & n12265 ) | ( n9817 & n12265 ) ;
  assign n31865 = ( n2557 & n4168 ) | ( n2557 & ~n16031 ) | ( n4168 & ~n16031 ) ;
  assign n31866 = n31865 ^ n29466 ^ n5838 ;
  assign n31867 = n15020 & n18099 ;
  assign n31868 = ~n31866 & n31867 ;
  assign n31869 = n31868 ^ n12801 ^ n2540 ;
  assign n31870 = n27916 ^ n16998 ^ n15065 ;
  assign n31871 = n11544 ^ n11535 ^ 1'b0 ;
  assign n31872 = n31871 ^ n16558 ^ n15272 ;
  assign n31873 = n26448 ^ n25064 ^ n16173 ;
  assign n31874 = n24762 ^ n4066 ^ 1'b0 ;
  assign n31875 = n11456 & n31874 ;
  assign n31876 = n3150 & n27150 ;
  assign n31877 = ~n31875 & n31876 ;
  assign n31878 = n28363 ^ n18555 ^ n13560 ;
  assign n31879 = n31878 ^ n21916 ^ 1'b0 ;
  assign n31880 = n6613 & ~n31879 ;
  assign n31881 = n26869 ^ n3079 ^ 1'b0 ;
  assign n31882 = n25201 ^ n9958 ^ 1'b0 ;
  assign n31883 = n31882 ^ n23840 ^ n4752 ;
  assign n31885 = n11272 & ~n17300 ;
  assign n31886 = n6650 & n31885 ;
  assign n31884 = n28900 ^ n27547 ^ 1'b0 ;
  assign n31887 = n31886 ^ n31884 ^ n7620 ;
  assign n31888 = n23321 ^ n15512 ^ n11563 ;
  assign n31889 = n31888 ^ n3614 ^ n3433 ;
  assign n31892 = ( n14421 & n28241 ) | ( n14421 & n28984 ) | ( n28241 & n28984 ) ;
  assign n31890 = n7565 | n16105 ;
  assign n31891 = n13036 & ~n31890 ;
  assign n31893 = n31892 ^ n31891 ^ 1'b0 ;
  assign n31894 = n23458 ^ n184 ^ 1'b0 ;
  assign n31895 = n13516 & n31894 ;
  assign n31896 = n23888 ^ n20697 ^ n11487 ;
  assign n31897 = ( n6677 & ~n31895 ) | ( n6677 & n31896 ) | ( ~n31895 & n31896 ) ;
  assign n31898 = ( n7811 & n7939 ) | ( n7811 & ~n17492 ) | ( n7939 & ~n17492 ) ;
  assign n31899 = n26894 ^ n20940 ^ n6374 ;
  assign n31900 = n2388 | n16855 ;
  assign n31901 = n21955 ^ n17471 ^ 1'b0 ;
  assign n31902 = ~n29034 & n31901 ;
  assign n31903 = ( n692 & n7354 ) | ( n692 & n10279 ) | ( n7354 & n10279 ) ;
  assign n31904 = n31903 ^ n29511 ^ n815 ;
  assign n31905 = n629 & ~n7080 ;
  assign n31906 = n31905 ^ n4301 ^ 1'b0 ;
  assign n31907 = n31906 ^ n25739 ^ n1201 ;
  assign n31908 = ( ~n12426 & n16147 ) | ( ~n12426 & n31907 ) | ( n16147 & n31907 ) ;
  assign n31909 = n31548 ^ n30166 ^ n18925 ;
  assign n31910 = n24715 ^ n21095 ^ n13049 ;
  assign n31911 = n31910 ^ n4417 ^ n1186 ;
  assign n31912 = n8350 ^ n4914 ^ n2878 ;
  assign n31913 = n15958 ^ n13031 ^ n7445 ;
  assign n31914 = ( n28548 & n31912 ) | ( n28548 & n31913 ) | ( n31912 & n31913 ) ;
  assign n31915 = n3648 & ~n22302 ;
  assign n31916 = n31915 ^ n5736 ^ 1'b0 ;
  assign n31917 = n31916 ^ n28132 ^ n2832 ;
  assign n31918 = n8352 & ~n31917 ;
  assign n31919 = ~n2572 & n10650 ;
  assign n31920 = n31919 ^ n4692 ^ 1'b0 ;
  assign n31921 = ( n2706 & ~n20244 ) | ( n2706 & n31920 ) | ( ~n20244 & n31920 ) ;
  assign n31922 = ~n831 & n2577 ;
  assign n31923 = ( ~n629 & n11297 ) | ( ~n629 & n31922 ) | ( n11297 & n31922 ) ;
  assign n31924 = ( n9227 & n17821 ) | ( n9227 & n31923 ) | ( n17821 & n31923 ) ;
  assign n31925 = ( n6794 & n12616 ) | ( n6794 & ~n23789 ) | ( n12616 & ~n23789 ) ;
  assign n31926 = n31925 ^ n28644 ^ n20971 ;
  assign n31927 = n31926 ^ n24402 ^ 1'b0 ;
  assign n31928 = n11751 & n31927 ;
  assign n31929 = ~n5268 & n13471 ;
  assign n31930 = n31478 ^ n29016 ^ n5381 ;
  assign n31931 = n10694 | n22848 ;
  assign n31932 = n28412 ^ n27631 ^ n7011 ;
  assign n31933 = n31932 ^ n6701 ^ 1'b0 ;
  assign n31934 = ~n28764 & n31933 ;
  assign n31935 = ( ~n1206 & n4354 ) | ( ~n1206 & n9065 ) | ( n4354 & n9065 ) ;
  assign n31936 = ( n7233 & ~n9570 ) | ( n7233 & n31935 ) | ( ~n9570 & n31935 ) ;
  assign n31937 = n31936 ^ n25810 ^ 1'b0 ;
  assign n31938 = n31937 ^ n22075 ^ n15018 ;
  assign n31939 = n22207 ^ n9441 ^ n2037 ;
  assign n31940 = n4581 | n19178 ;
  assign n31941 = n31939 & ~n31940 ;
  assign n31942 = n31941 ^ n15911 ^ n5034 ;
  assign n31943 = n13236 & ~n31942 ;
  assign n31945 = ( n2112 & n7232 ) | ( n2112 & n7914 ) | ( n7232 & n7914 ) ;
  assign n31946 = n31945 ^ n2998 ^ 1'b0 ;
  assign n31944 = n24502 & n26987 ;
  assign n31947 = n31946 ^ n31944 ^ n4323 ;
  assign n31948 = n22407 ^ n3375 ^ 1'b0 ;
  assign n31949 = ( n28403 & n30032 ) | ( n28403 & n31948 ) | ( n30032 & n31948 ) ;
  assign n31950 = ( ~n5583 & n28193 ) | ( ~n5583 & n31949 ) | ( n28193 & n31949 ) ;
  assign n31951 = n19906 ^ n17298 ^ n7903 ;
  assign n31952 = n31951 ^ n17759 ^ n14557 ;
  assign n31953 = n25095 ^ n14196 ^ n8907 ;
  assign n31954 = n12504 ^ n2944 ^ 1'b0 ;
  assign n31955 = n550 | n31954 ;
  assign n31956 = ( ~n3276 & n28497 ) | ( ~n3276 & n31955 ) | ( n28497 & n31955 ) ;
  assign n31957 = ~n5090 & n13054 ;
  assign n31958 = n31957 ^ n31838 ^ 1'b0 ;
  assign n31959 = n17644 ^ n16723 ^ n920 ;
  assign n31960 = ( n8077 & n9345 ) | ( n8077 & n31840 ) | ( n9345 & n31840 ) ;
  assign n31961 = ( ~n22965 & n31959 ) | ( ~n22965 & n31960 ) | ( n31959 & n31960 ) ;
  assign n31962 = n7682 & ~n11122 ;
  assign n31963 = ~n5708 & n31962 ;
  assign n31964 = n31963 ^ n7407 ^ n1294 ;
  assign n31965 = ( n3593 & n11494 ) | ( n3593 & n23967 ) | ( n11494 & n23967 ) ;
  assign n31966 = n23158 ^ n13232 ^ 1'b0 ;
  assign n31967 = n3068 & ~n8064 ;
  assign n31968 = n31967 ^ n3151 ^ 1'b0 ;
  assign n31969 = ~n14995 & n20530 ;
  assign n31970 = ( n1258 & n5045 ) | ( n1258 & ~n25416 ) | ( n5045 & ~n25416 ) ;
  assign n31971 = ( n6268 & ~n12515 ) | ( n6268 & n12637 ) | ( ~n12515 & n12637 ) ;
  assign n31972 = n31971 ^ n22246 ^ n16447 ;
  assign n31973 = ( n7820 & ~n17081 ) | ( n7820 & n29678 ) | ( ~n17081 & n29678 ) ;
  assign n31974 = n9274 & n15401 ;
  assign n31975 = ( n8850 & ~n15953 ) | ( n8850 & n22304 ) | ( ~n15953 & n22304 ) ;
  assign n31976 = ( n14362 & n14532 ) | ( n14362 & ~n15015 ) | ( n14532 & ~n15015 ) ;
  assign n31977 = n3755 & ~n13051 ;
  assign n31978 = ( n541 & n31587 ) | ( n541 & ~n31977 ) | ( n31587 & ~n31977 ) ;
  assign n31979 = n29094 ^ n17679 ^ 1'b0 ;
  assign n31980 = x46 & ~n31979 ;
  assign n31981 = n2849 & ~n14858 ;
  assign n31982 = n20304 & n31981 ;
  assign n31983 = n23317 ^ n16120 ^ n8455 ;
  assign n31984 = n22705 ^ n20338 ^ n15450 ;
  assign n31985 = n23317 ^ n1498 ^ n1030 ;
  assign n31986 = ( ~n3760 & n13407 ) | ( ~n3760 & n31985 ) | ( n13407 & n31985 ) ;
  assign n31987 = n27400 ^ n13015 ^ n12158 ;
  assign n31988 = ( n9005 & ~n22554 ) | ( n9005 & n31987 ) | ( ~n22554 & n31987 ) ;
  assign n31989 = n28007 ^ n18917 ^ n5242 ;
  assign n31990 = ( n5232 & n12730 ) | ( n5232 & ~n31989 ) | ( n12730 & ~n31989 ) ;
  assign n31993 = n12660 & ~n19434 ;
  assign n31994 = n31993 ^ n17012 ^ 1'b0 ;
  assign n31991 = ( ~n3904 & n8319 ) | ( ~n3904 & n9276 ) | ( n8319 & n9276 ) ;
  assign n31992 = n31991 ^ n19916 ^ 1'b0 ;
  assign n31995 = n31994 ^ n31992 ^ 1'b0 ;
  assign n31996 = n31995 ^ n21900 ^ n6679 ;
  assign n31997 = ( n1469 & n17071 ) | ( n1469 & ~n27330 ) | ( n17071 & ~n27330 ) ;
  assign n31998 = n16657 ^ n4535 ^ 1'b0 ;
  assign n31999 = ( ~n16384 & n24598 ) | ( ~n16384 & n31998 ) | ( n24598 & n31998 ) ;
  assign n32000 = n28860 ^ n25077 ^ n16863 ;
  assign n32001 = n11863 ^ x111 ^ 1'b0 ;
  assign n32002 = n32000 & ~n32001 ;
  assign n32003 = n1025 & ~n1143 ;
  assign n32004 = n32003 ^ n22260 ^ 1'b0 ;
  assign n32005 = ( n9309 & n15106 ) | ( n9309 & ~n16598 ) | ( n15106 & ~n16598 ) ;
  assign n32006 = ( n5206 & n13634 ) | ( n5206 & n19390 ) | ( n13634 & n19390 ) ;
  assign n32007 = ( n8354 & ~n32005 ) | ( n8354 & n32006 ) | ( ~n32005 & n32006 ) ;
  assign n32008 = n3702 | n32007 ;
  assign n32009 = n11806 & ~n32008 ;
  assign n32010 = n22853 ^ n16913 ^ n9975 ;
  assign n32011 = n27322 ^ n5662 ^ 1'b0 ;
  assign n32012 = n21397 ^ n20565 ^ n1912 ;
  assign n32013 = n32012 ^ n13870 ^ n10282 ;
  assign n32015 = n14550 ^ n11568 ^ n9022 ;
  assign n32014 = n239 & n21984 ;
  assign n32016 = n32015 ^ n32014 ^ n1134 ;
  assign n32017 = n32016 ^ n9975 ^ n2759 ;
  assign n32018 = n9366 | n9701 ;
  assign n32019 = n32018 ^ n9761 ^ n2212 ;
  assign n32020 = n32019 ^ n7024 ^ n702 ;
  assign n32022 = n15409 ^ n11933 ^ n10136 ;
  assign n32021 = ( n17560 & ~n18506 ) | ( n17560 & n19920 ) | ( ~n18506 & n19920 ) ;
  assign n32023 = n32022 ^ n32021 ^ n16082 ;
  assign n32024 = ( n5923 & ~n8422 ) | ( n5923 & n15390 ) | ( ~n8422 & n15390 ) ;
  assign n32025 = n32024 ^ n29955 ^ n14890 ;
  assign n32026 = n16958 ^ n8077 ^ n3572 ;
  assign n32027 = n31565 ^ n9596 ^ n4667 ;
  assign n32028 = ( n3849 & n15496 ) | ( n3849 & ~n32027 ) | ( n15496 & ~n32027 ) ;
  assign n32029 = n7670 & n32028 ;
  assign n32030 = n32029 ^ n12382 ^ 1'b0 ;
  assign n32031 = ( n7091 & n9030 ) | ( n7091 & n14449 ) | ( n9030 & n14449 ) ;
  assign n32032 = n32031 ^ n31708 ^ n18452 ;
  assign n32033 = n3129 & n23608 ;
  assign n32034 = n32033 ^ n12663 ^ 1'b0 ;
  assign n32035 = n32034 ^ n20475 ^ n12145 ;
  assign n32036 = n27169 ^ n16787 ^ n9851 ;
  assign n32037 = ( n3228 & n4626 ) | ( n3228 & n32036 ) | ( n4626 & n32036 ) ;
  assign n32038 = ( n1908 & n4891 ) | ( n1908 & ~n20875 ) | ( n4891 & ~n20875 ) ;
  assign n32039 = n17275 ^ n12367 ^ n2234 ;
  assign n32040 = n32039 ^ n10294 ^ n1786 ;
  assign n32041 = ( n13434 & ~n32038 ) | ( n13434 & n32040 ) | ( ~n32038 & n32040 ) ;
  assign n32042 = ( n968 & n2897 ) | ( n968 & n13396 ) | ( n2897 & n13396 ) ;
  assign n32043 = n1979 & n20352 ;
  assign n32044 = n5162 & n32043 ;
  assign n32045 = ( n7261 & ~n18890 ) | ( n7261 & n32044 ) | ( ~n18890 & n32044 ) ;
  assign n32046 = n20874 ^ n8017 ^ 1'b0 ;
  assign n32047 = n16967 ^ n14239 ^ n9722 ;
  assign n32048 = n662 & ~n20809 ;
  assign n32049 = n32048 ^ n30450 ^ n12400 ;
  assign n32051 = n13299 ^ n11033 ^ 1'b0 ;
  assign n32052 = n19582 & ~n32051 ;
  assign n32050 = ~n8645 & n22938 ;
  assign n32053 = n32052 ^ n32050 ^ 1'b0 ;
  assign n32055 = ( n14717 & n14789 ) | ( n14717 & n25025 ) | ( n14789 & n25025 ) ;
  assign n32056 = ( n17147 & n22158 ) | ( n17147 & ~n32055 ) | ( n22158 & ~n32055 ) ;
  assign n32054 = n6431 & n16199 ;
  assign n32057 = n32056 ^ n32054 ^ 1'b0 ;
  assign n32058 = n1138 | n19237 ;
  assign n32059 = n26914 ^ n25310 ^ n16508 ;
  assign n32060 = n14353 ^ n13954 ^ n10035 ;
  assign n32061 = ( n10499 & n12856 ) | ( n10499 & n32060 ) | ( n12856 & n32060 ) ;
  assign n32062 = n32061 ^ n31422 ^ n5160 ;
  assign n32063 = ( n1747 & n14920 ) | ( n1747 & ~n32062 ) | ( n14920 & ~n32062 ) ;
  assign n32064 = n13572 ^ n11726 ^ n3648 ;
  assign n32065 = ~n6293 & n24315 ;
  assign n32066 = ~n23801 & n32065 ;
  assign n32067 = n3847 & ~n24947 ;
  assign n32068 = n6640 | n24650 ;
  assign n32069 = n6285 & ~n32068 ;
  assign n32070 = n32069 ^ n9176 ^ 1'b0 ;
  assign n32071 = n6215 | n32070 ;
  assign n32072 = n32067 | n32071 ;
  assign n32073 = n32066 & ~n32072 ;
  assign n32074 = ( n2146 & ~n32064 ) | ( n2146 & n32073 ) | ( ~n32064 & n32073 ) ;
  assign n32076 = ( n3477 & n7733 ) | ( n3477 & ~n9295 ) | ( n7733 & ~n9295 ) ;
  assign n32077 = ( n2028 & n28375 ) | ( n2028 & n32076 ) | ( n28375 & n32076 ) ;
  assign n32075 = n31830 ^ n9410 ^ 1'b0 ;
  assign n32078 = n32077 ^ n32075 ^ n4717 ;
  assign n32079 = ( n4246 & ~n6172 ) | ( n4246 & n6972 ) | ( ~n6172 & n6972 ) ;
  assign n32080 = ( n16067 & ~n24890 ) | ( n16067 & n32079 ) | ( ~n24890 & n32079 ) ;
  assign n32081 = ( n16726 & n24739 ) | ( n16726 & ~n28202 ) | ( n24739 & ~n28202 ) ;
  assign n32082 = ( ~n8910 & n9980 ) | ( ~n8910 & n30521 ) | ( n9980 & n30521 ) ;
  assign n32083 = n4248 ^ n1521 ^ 1'b0 ;
  assign n32084 = n2965 & ~n7283 ;
  assign n32085 = n32084 ^ n30454 ^ 1'b0 ;
  assign n32086 = ( n19940 & ~n32083 ) | ( n19940 & n32085 ) | ( ~n32083 & n32085 ) ;
  assign n32087 = n31616 & ~n32086 ;
  assign n32088 = n32087 ^ n27703 ^ 1'b0 ;
  assign n32089 = n2082 | n9367 ;
  assign n32090 = n11638 | n32089 ;
  assign n32091 = ( ~n1818 & n4089 ) | ( ~n1818 & n23235 ) | ( n4089 & n23235 ) ;
  assign n32092 = n32091 ^ n3909 ^ 1'b0 ;
  assign n32093 = n5266 & ~n32092 ;
  assign n32094 = n30154 ^ n21090 ^ 1'b0 ;
  assign n32095 = n13814 & ~n32094 ;
  assign n32096 = n32095 ^ n28396 ^ n7183 ;
  assign n32097 = ( n3023 & n3999 ) | ( n3023 & n7746 ) | ( n3999 & n7746 ) ;
  assign n32098 = n25464 ^ n3570 ^ 1'b0 ;
  assign n32099 = ~n18217 & n32098 ;
  assign n32100 = ( ~n546 & n10915 ) | ( ~n546 & n32099 ) | ( n10915 & n32099 ) ;
  assign n32101 = n28121 ^ n21458 ^ 1'b0 ;
  assign n32102 = ~n17365 & n26995 ;
  assign n32103 = ( x37 & n14533 ) | ( x37 & n30147 ) | ( n14533 & n30147 ) ;
  assign n32104 = ( ~n13042 & n14656 ) | ( ~n13042 & n32103 ) | ( n14656 & n32103 ) ;
  assign n32105 = n32104 ^ n16325 ^ n12029 ;
  assign n32106 = ( n1170 & ~n9301 ) | ( n1170 & n18282 ) | ( ~n9301 & n18282 ) ;
  assign n32107 = n29119 ^ n23974 ^ n21304 ;
  assign n32108 = n21077 ^ n19645 ^ n2895 ;
  assign n32109 = n32108 ^ n30412 ^ n22978 ;
  assign n32110 = ( n31296 & n32107 ) | ( n31296 & ~n32109 ) | ( n32107 & ~n32109 ) ;
  assign n32111 = n5895 ^ n996 ^ 1'b0 ;
  assign n32112 = n20539 & ~n32111 ;
  assign n32113 = n29506 ^ n7189 ^ 1'b0 ;
  assign n32114 = n9237 & n32113 ;
  assign n32115 = n32091 ^ n11840 ^ x121 ;
  assign n32116 = n32115 ^ n14030 ^ n2868 ;
  assign n32120 = ( ~n4876 & n13723 ) | ( ~n4876 & n14431 ) | ( n13723 & n14431 ) ;
  assign n32117 = n22987 ^ n1531 ^ 1'b0 ;
  assign n32118 = n5306 & ~n32117 ;
  assign n32119 = ( n12013 & n25993 ) | ( n12013 & n32118 ) | ( n25993 & n32118 ) ;
  assign n32121 = n32120 ^ n32119 ^ n30923 ;
  assign n32123 = n4806 ^ n4193 ^ n385 ;
  assign n32122 = ~n6310 & n29100 ;
  assign n32124 = n32123 ^ n32122 ^ 1'b0 ;
  assign n32125 = n32124 ^ n25082 ^ n9354 ;
  assign n32126 = n32125 ^ n17465 ^ 1'b0 ;
  assign n32127 = n21823 ^ n12869 ^ n6819 ;
  assign n32129 = n30245 ^ n5787 ^ n634 ;
  assign n32130 = n32129 ^ n29214 ^ n17652 ;
  assign n32128 = ( n16886 & n19976 ) | ( n16886 & ~n22784 ) | ( n19976 & ~n22784 ) ;
  assign n32131 = n32130 ^ n32128 ^ n26003 ;
  assign n32132 = n12521 ^ n11790 ^ n937 ;
  assign n32133 = ( n399 & n22406 ) | ( n399 & n32132 ) | ( n22406 & n32132 ) ;
  assign n32134 = n16747 ^ n1618 ^ n677 ;
  assign n32135 = n19417 ^ n12395 ^ n3895 ;
  assign n32136 = ( n5355 & n32015 ) | ( n5355 & n32135 ) | ( n32015 & n32135 ) ;
  assign n32137 = n5405 & n12228 ;
  assign n32138 = n3344 & n32137 ;
  assign n32139 = n24630 ^ n9557 ^ 1'b0 ;
  assign n32140 = x117 & ~n32139 ;
  assign n32141 = n3876 & ~n6283 ;
  assign n32142 = ( n4238 & n20187 ) | ( n4238 & ~n26233 ) | ( n20187 & ~n26233 ) ;
  assign n32143 = ( n16420 & n18590 ) | ( n16420 & n32142 ) | ( n18590 & n32142 ) ;
  assign n32144 = ( ~n19161 & n32141 ) | ( ~n19161 & n32143 ) | ( n32141 & n32143 ) ;
  assign n32145 = n32144 ^ n28035 ^ n12193 ;
  assign n32146 = n12664 | n32145 ;
  assign n32147 = ( n7674 & n11255 ) | ( n7674 & ~n12691 ) | ( n11255 & ~n12691 ) ;
  assign n32148 = ( n7271 & ~n12510 ) | ( n7271 & n27013 ) | ( ~n12510 & n27013 ) ;
  assign n32149 = ( ~n17145 & n17582 ) | ( ~n17145 & n30994 ) | ( n17582 & n30994 ) ;
  assign n32150 = n11020 ^ n5940 ^ 1'b0 ;
  assign n32151 = ~n3229 & n32150 ;
  assign n32152 = ( n1462 & ~n5331 ) | ( n1462 & n32151 ) | ( ~n5331 & n32151 ) ;
  assign n32153 = n11165 ^ n1289 ^ 1'b0 ;
  assign n32154 = ( n5668 & ~n9822 ) | ( n5668 & n32153 ) | ( ~n9822 & n32153 ) ;
  assign n32155 = n25050 ^ n23575 ^ n7604 ;
  assign n32156 = n32155 ^ n9610 ^ 1'b0 ;
  assign n32157 = ( ~n6465 & n7981 ) | ( ~n6465 & n9708 ) | ( n7981 & n9708 ) ;
  assign n32158 = ( ~n13031 & n15799 ) | ( ~n13031 & n32157 ) | ( n15799 & n32157 ) ;
  assign n32159 = ( ~n1641 & n4661 ) | ( ~n1641 & n29450 ) | ( n4661 & n29450 ) ;
  assign n32160 = n32159 ^ n4193 ^ 1'b0 ;
  assign n32161 = n11526 ^ n6097 ^ 1'b0 ;
  assign n32162 = n32160 & n32161 ;
  assign n32163 = ( n11426 & n32158 ) | ( n11426 & n32162 ) | ( n32158 & n32162 ) ;
  assign n32164 = ~n11412 & n14081 ;
  assign n32165 = n6215 & n32164 ;
  assign n32166 = n29294 ^ n24018 ^ 1'b0 ;
  assign n32167 = ~n24306 & n32166 ;
  assign n32168 = ( ~n16011 & n18969 ) | ( ~n16011 & n28596 ) | ( n18969 & n28596 ) ;
  assign n32169 = ( ~n2209 & n13637 ) | ( ~n2209 & n17249 ) | ( n13637 & n17249 ) ;
  assign n32170 = n32169 ^ n25318 ^ n3005 ;
  assign n32171 = n20666 ^ n13720 ^ n8522 ;
  assign n32172 = ( n2154 & n3823 ) | ( n2154 & ~n24588 ) | ( n3823 & ~n24588 ) ;
  assign n32173 = n32172 ^ n23471 ^ n2615 ;
  assign n32174 = ( n6175 & ~n31922 ) | ( n6175 & n32173 ) | ( ~n31922 & n32173 ) ;
  assign n32175 = n18652 ^ n7968 ^ n4917 ;
  assign n32176 = n32175 ^ n30246 ^ n22275 ;
  assign n32177 = ( n1024 & ~n16101 ) | ( n1024 & n28938 ) | ( ~n16101 & n28938 ) ;
  assign n32180 = ( ~n2458 & n29158 ) | ( ~n2458 & n30927 ) | ( n29158 & n30927 ) ;
  assign n32181 = n32180 ^ n6928 ^ 1'b0 ;
  assign n32179 = n6776 & n21412 ;
  assign n32182 = n32181 ^ n32179 ^ 1'b0 ;
  assign n32178 = n21894 ^ n20887 ^ n18195 ;
  assign n32183 = n32182 ^ n32178 ^ n7943 ;
  assign n32184 = ( n8896 & n11100 ) | ( n8896 & n26698 ) | ( n11100 & n26698 ) ;
  assign n32185 = n14288 ^ n3004 ^ 1'b0 ;
  assign n32186 = n23215 | n32185 ;
  assign n32187 = n2930 ^ n761 ^ 1'b0 ;
  assign n32188 = ~n5973 & n32187 ;
  assign n32189 = ~n152 & n29286 ;
  assign n32190 = ~n26012 & n32189 ;
  assign n32195 = ( ~n3513 & n10322 ) | ( ~n3513 & n13317 ) | ( n10322 & n13317 ) ;
  assign n32192 = n8302 | n25347 ;
  assign n32193 = n32192 ^ n26513 ^ 1'b0 ;
  assign n32191 = n17125 | n24186 ;
  assign n32194 = n32193 ^ n32191 ^ 1'b0 ;
  assign n32196 = n32195 ^ n32194 ^ n15368 ;
  assign n32197 = n14078 | n30004 ;
  assign n32198 = n10421 | n32197 ;
  assign n32199 = ( ~x62 & n17941 ) | ( ~x62 & n32198 ) | ( n17941 & n32198 ) ;
  assign n32200 = n13038 ^ n2217 ^ 1'b0 ;
  assign n32201 = n24820 ^ n21117 ^ n16356 ;
  assign n32202 = ( n17920 & n32200 ) | ( n17920 & n32201 ) | ( n32200 & n32201 ) ;
  assign n32203 = n29719 ^ n224 ^ 1'b0 ;
  assign n32204 = n28413 ^ n11363 ^ n4437 ;
  assign n32205 = ( n326 & n7152 ) | ( n326 & n16213 ) | ( n7152 & n16213 ) ;
  assign n32206 = ( n6755 & n23669 ) | ( n6755 & ~n32205 ) | ( n23669 & ~n32205 ) ;
  assign n32207 = n19084 ^ n11929 ^ n5742 ;
  assign n32208 = n28899 ^ n711 ^ 1'b0 ;
  assign n32209 = n732 & n32208 ;
  assign n32210 = n17806 & n32209 ;
  assign n32211 = n32210 ^ n5653 ^ 1'b0 ;
  assign n32212 = n14060 | n32211 ;
  assign n32213 = n10315 & ~n32212 ;
  assign n32214 = ( ~n6508 & n21557 ) | ( ~n6508 & n32213 ) | ( n21557 & n32213 ) ;
  assign n32215 = n10028 & n15497 ;
  assign n32216 = ~n11101 & n32215 ;
  assign n32217 = n25210 ^ n16667 ^ 1'b0 ;
  assign n32218 = n15398 & ~n32217 ;
  assign n32219 = ( n1901 & n6944 ) | ( n1901 & ~n16888 ) | ( n6944 & ~n16888 ) ;
  assign n32220 = n20157 ^ n18551 ^ 1'b0 ;
  assign n32221 = n32219 | n32220 ;
  assign n32222 = n27452 ^ n5373 ^ n2825 ;
  assign n32223 = n8144 | n26756 ;
  assign n32224 = n10869 & ~n17539 ;
  assign n32225 = n32224 ^ n22585 ^ n2428 ;
  assign n32226 = ( n5542 & ~n5603 ) | ( n5542 & n6144 ) | ( ~n5603 & n6144 ) ;
  assign n32227 = n32226 ^ n28237 ^ n11786 ;
  assign n32228 = n4344 | n27755 ;
  assign n32229 = n14789 & ~n32228 ;
  assign n32230 = ( n9354 & ~n10348 ) | ( n9354 & n32229 ) | ( ~n10348 & n32229 ) ;
  assign n32231 = n3320 | n8282 ;
  assign n32232 = n5150 & ~n11269 ;
  assign n32233 = n27779 ^ n842 ^ 1'b0 ;
  assign n32234 = ( n2135 & ~n5142 ) | ( n2135 & n24318 ) | ( ~n5142 & n24318 ) ;
  assign n32235 = n5342 & ~n32234 ;
  assign n32236 = n32235 ^ n26155 ^ 1'b0 ;
  assign n32237 = ( ~n4731 & n6829 ) | ( ~n4731 & n14325 ) | ( n6829 & n14325 ) ;
  assign n32238 = n29526 ^ n14131 ^ 1'b0 ;
  assign n32239 = n32237 & ~n32238 ;
  assign n32240 = ~n9075 & n20875 ;
  assign n32241 = n25951 ^ n12930 ^ n5752 ;
  assign n32242 = n32241 ^ n18766 ^ n769 ;
  assign n32243 = n32242 ^ n26513 ^ n5554 ;
  assign n32244 = n21453 ^ n16015 ^ n11879 ;
  assign n32247 = ~n4114 & n11665 ;
  assign n32245 = n8203 | n10714 ;
  assign n32246 = n32245 ^ n3170 ^ 1'b0 ;
  assign n32248 = n32247 ^ n32246 ^ n24591 ;
  assign n32249 = n25870 ^ n11596 ^ n8559 ;
  assign n32250 = ( n11832 & n13171 ) | ( n11832 & n32249 ) | ( n13171 & n32249 ) ;
  assign n32251 = n4645 & n32250 ;
  assign n32252 = n11044 & n26731 ;
  assign n32253 = n27961 & ~n32252 ;
  assign n32254 = n27785 ^ n10102 ^ n2708 ;
  assign n32255 = n2527 & n19018 ;
  assign n32256 = n32255 ^ n7322 ^ 1'b0 ;
  assign n32257 = n32256 ^ n29356 ^ n21888 ;
  assign n32258 = ( n3070 & ~n4952 ) | ( n3070 & n5808 ) | ( ~n4952 & n5808 ) ;
  assign n32259 = n12202 & n32258 ;
  assign n32260 = n13150 & n32259 ;
  assign n32261 = n1641 & ~n12780 ;
  assign n32262 = n8051 & n32261 ;
  assign n32263 = n3067 & n31528 ;
  assign n32264 = n32263 ^ n30431 ^ 1'b0 ;
  assign n32265 = n6894 & ~n24298 ;
  assign n32266 = n32265 ^ n30870 ^ n28517 ;
  assign n32267 = ( n10973 & ~n23515 ) | ( n10973 & n30571 ) | ( ~n23515 & n30571 ) ;
  assign n32268 = ( n4728 & ~n5351 ) | ( n4728 & n25652 ) | ( ~n5351 & n25652 ) ;
  assign n32269 = n32268 ^ n7328 ^ n5631 ;
  assign n32270 = n15956 ^ n4409 ^ n2585 ;
  assign n32271 = ( n5548 & n16550 ) | ( n5548 & ~n32270 ) | ( n16550 & ~n32270 ) ;
  assign n32272 = n23047 ^ n3210 ^ x55 ;
  assign n32275 = n18976 & n22122 ;
  assign n32273 = ( n3603 & n17715 ) | ( n3603 & n29781 ) | ( n17715 & n29781 ) ;
  assign n32274 = ( ~n7528 & n10981 ) | ( ~n7528 & n32273 ) | ( n10981 & n32273 ) ;
  assign n32276 = n32275 ^ n32274 ^ n6007 ;
  assign n32277 = ( n8629 & n15467 ) | ( n8629 & n20720 ) | ( n15467 & n20720 ) ;
  assign n32278 = ~n550 & n12082 ;
  assign n32279 = ( ~n21389 & n28065 ) | ( ~n21389 & n32278 ) | ( n28065 & n32278 ) ;
  assign n32280 = n22213 ^ n9316 ^ n8485 ;
  assign n32281 = n6567 & n32280 ;
  assign n32282 = n12591 & ~n32281 ;
  assign n32283 = ~n24164 & n32282 ;
  assign n32284 = n863 & n30949 ;
  assign n32285 = ~n9372 & n32284 ;
  assign n32286 = n3525 ^ n2145 ^ 1'b0 ;
  assign n32287 = n32286 ^ n13699 ^ 1'b0 ;
  assign n32288 = ~n16387 & n32287 ;
  assign n32289 = n32288 ^ n17708 ^ n4511 ;
  assign n32290 = n15020 & ~n32289 ;
  assign n32291 = n32290 ^ n7986 ^ 1'b0 ;
  assign n32292 = n32198 ^ n29757 ^ x65 ;
  assign n32293 = n17883 ^ n10651 ^ 1'b0 ;
  assign n32294 = n6715 ^ n3320 ^ n1854 ;
  assign n32295 = ( n15151 & ~n15751 ) | ( n15151 & n32067 ) | ( ~n15751 & n32067 ) ;
  assign n32296 = n16171 ^ n2258 ^ 1'b0 ;
  assign n32297 = n32296 ^ n32178 ^ n706 ;
  assign n32298 = n8931 ^ n4668 ^ 1'b0 ;
  assign n32299 = n11035 | n32298 ;
  assign n32300 = n32299 ^ n24032 ^ n634 ;
  assign n32301 = n31868 ^ n25848 ^ x75 ;
  assign n32302 = n9561 ^ n8411 ^ n7152 ;
  assign n32303 = n32302 ^ n17982 ^ n12617 ;
  assign n32304 = n14487 ^ n8617 ^ 1'b0 ;
  assign n32305 = n16638 & n32304 ;
  assign n32306 = ( n16787 & ~n25575 ) | ( n16787 & n28738 ) | ( ~n25575 & n28738 ) ;
  assign n32307 = n21626 ^ n6085 ^ 1'b0 ;
  assign n32308 = n31939 | n32307 ;
  assign n32309 = ( n18252 & n22679 ) | ( n18252 & ~n32308 ) | ( n22679 & ~n32308 ) ;
  assign n32310 = n26540 ^ n11519 ^ n5308 ;
  assign n32311 = n12149 ^ n2656 ^ 1'b0 ;
  assign n32312 = n30848 ^ n21555 ^ n18433 ;
  assign n32313 = n8065 ^ n2432 ^ x51 ;
  assign n32314 = n32313 ^ n13509 ^ 1'b0 ;
  assign n32315 = n7034 ^ n3363 ^ 1'b0 ;
  assign n32316 = n3413 & ~n32315 ;
  assign n32317 = n32316 ^ n3318 ^ 1'b0 ;
  assign n32319 = n11212 ^ n7437 ^ n2036 ;
  assign n32320 = n32319 ^ n10053 ^ n2233 ;
  assign n32321 = ( n14169 & ~n18404 ) | ( n14169 & n32320 ) | ( ~n18404 & n32320 ) ;
  assign n32318 = n10897 | n27156 ;
  assign n32322 = n32321 ^ n32318 ^ 1'b0 ;
  assign n32323 = ( n3263 & n32317 ) | ( n3263 & ~n32322 ) | ( n32317 & ~n32322 ) ;
  assign n32324 = ( ~n12163 & n12181 ) | ( ~n12163 & n23965 ) | ( n12181 & n23965 ) ;
  assign n32325 = n25751 ^ n14260 ^ n5329 ;
  assign n32326 = n16649 & n32325 ;
  assign n32327 = n6751 | n10059 ;
  assign n32328 = n11366 & ~n32327 ;
  assign n32329 = n30571 ^ n25074 ^ n20626 ;
  assign n32330 = n9841 ^ n9750 ^ 1'b0 ;
  assign n32331 = n11134 ^ n6433 ^ 1'b0 ;
  assign n32334 = ( n2248 & ~n3633 ) | ( n2248 & n12800 ) | ( ~n3633 & n12800 ) ;
  assign n32332 = ~n4804 & n18913 ;
  assign n32333 = n32332 ^ n31224 ^ n15937 ;
  assign n32335 = n32334 ^ n32333 ^ n12085 ;
  assign n32336 = n20096 ^ n5926 ^ 1'b0 ;
  assign n32337 = n31228 ^ n27367 ^ n2843 ;
  assign n32338 = ( ~n22568 & n32336 ) | ( ~n22568 & n32337 ) | ( n32336 & n32337 ) ;
  assign n32339 = n12929 & ~n19846 ;
  assign n32340 = n32339 ^ n30590 ^ n3525 ;
  assign n32341 = n3745 ^ n1778 ^ 1'b0 ;
  assign n32342 = n19731 ^ n8681 ^ 1'b0 ;
  assign n32343 = n19780 | n32342 ;
  assign n32344 = ( n6106 & n32341 ) | ( n6106 & n32343 ) | ( n32341 & n32343 ) ;
  assign n32345 = n32344 ^ n10355 ^ n7689 ;
  assign n32346 = ( n8469 & n14991 ) | ( n8469 & ~n31595 ) | ( n14991 & ~n31595 ) ;
  assign n32347 = n11847 ^ n10819 ^ n921 ;
  assign n32348 = ( n8339 & n32343 ) | ( n8339 & ~n32347 ) | ( n32343 & ~n32347 ) ;
  assign n32349 = ~n20316 & n22951 ;
  assign n32350 = ~n32348 & n32349 ;
  assign n32351 = n3530 | n26399 ;
  assign n32352 = n32351 ^ n24389 ^ 1'b0 ;
  assign n32353 = ( n462 & n13218 ) | ( n462 & ~n25125 ) | ( n13218 & ~n25125 ) ;
  assign n32354 = ( n8419 & n8605 ) | ( n8419 & n12290 ) | ( n8605 & n12290 ) ;
  assign n32355 = n32354 ^ n1306 ^ 1'b0 ;
  assign n32359 = ( n380 & n6992 ) | ( n380 & n31530 ) | ( n6992 & n31530 ) ;
  assign n32360 = n32359 ^ n16899 ^ 1'b0 ;
  assign n32356 = ~n1864 & n4678 ;
  assign n32357 = n32356 ^ n162 ^ 1'b0 ;
  assign n32358 = ( n8710 & ~n11359 ) | ( n8710 & n32357 ) | ( ~n11359 & n32357 ) ;
  assign n32361 = n32360 ^ n32358 ^ n15456 ;
  assign n32362 = n7921 & ~n19739 ;
  assign n32363 = n32362 ^ n8348 ^ 1'b0 ;
  assign n32364 = ( n17039 & ~n22664 ) | ( n17039 & n32363 ) | ( ~n22664 & n32363 ) ;
  assign n32365 = ~n8465 & n24671 ;
  assign n32366 = n31229 ^ n13139 ^ n1395 ;
  assign n32367 = ( n3787 & ~n17107 ) | ( n3787 & n32366 ) | ( ~n17107 & n32366 ) ;
  assign n32369 = ( x102 & ~n11769 ) | ( x102 & n13654 ) | ( ~n11769 & n13654 ) ;
  assign n32368 = n23536 ^ n9489 ^ n6650 ;
  assign n32370 = n32369 ^ n32368 ^ n6409 ;
  assign n32371 = ( n3709 & n5835 ) | ( n3709 & n10059 ) | ( n5835 & n10059 ) ;
  assign n32372 = ~n8311 & n10108 ;
  assign n32373 = n32372 ^ n22257 ^ n7516 ;
  assign n32374 = ( n1448 & ~n8094 ) | ( n1448 & n21836 ) | ( ~n8094 & n21836 ) ;
  assign n32375 = ( n881 & n17256 ) | ( n881 & n32374 ) | ( n17256 & n32374 ) ;
  assign n32376 = n7026 & n32375 ;
  assign n32377 = n32373 & n32376 ;
  assign n32378 = n12291 ^ n444 ^ 1'b0 ;
  assign n32379 = n27608 & n32378 ;
  assign n32380 = n6403 & n21793 ;
  assign n32381 = n32380 ^ n2188 ^ 1'b0 ;
  assign n32382 = n12519 & ~n28081 ;
  assign n32383 = n32382 ^ n29044 ^ n12658 ;
  assign n32384 = n25635 ^ n11958 ^ 1'b0 ;
  assign n32385 = n32384 ^ n25512 ^ n1456 ;
  assign n32386 = ( ~n12180 & n18034 ) | ( ~n12180 & n32385 ) | ( n18034 & n32385 ) ;
  assign n32387 = n6299 ^ n2724 ^ n177 ;
  assign n32388 = n32387 ^ n30451 ^ n23515 ;
  assign n32389 = n21482 | n24828 ;
  assign n32390 = n32389 ^ n5155 ^ 1'b0 ;
  assign n32391 = n27318 ^ n4482 ^ n4468 ;
  assign n32392 = ( n4030 & n32390 ) | ( n4030 & n32391 ) | ( n32390 & n32391 ) ;
  assign n32393 = n20733 | n28590 ;
  assign n32394 = n32393 ^ n15464 ^ 1'b0 ;
  assign n32395 = ~n2704 & n6571 ;
  assign n32396 = ( n20261 & n32394 ) | ( n20261 & n32395 ) | ( n32394 & n32395 ) ;
  assign n32397 = n12117 ^ n2893 ^ 1'b0 ;
  assign n32398 = ~n3342 & n5875 ;
  assign n32399 = n15958 & n32398 ;
  assign n32400 = ( n862 & ~n4480 ) | ( n862 & n32399 ) | ( ~n4480 & n32399 ) ;
  assign n32401 = n4016 & n7058 ;
  assign n32402 = ~n16917 & n32401 ;
  assign n32403 = ( n11707 & n32400 ) | ( n11707 & ~n32402 ) | ( n32400 & ~n32402 ) ;
  assign n32404 = n32403 ^ n26446 ^ n20150 ;
  assign n32405 = n32067 ^ n20605 ^ n13764 ;
  assign n32406 = n32405 ^ n18177 ^ n8789 ;
  assign n32407 = ( n1869 & n2746 ) | ( n1869 & ~n8511 ) | ( n2746 & ~n8511 ) ;
  assign n32408 = n14304 & n32407 ;
  assign n32409 = n32408 ^ n5730 ^ 1'b0 ;
  assign n32410 = n17073 ^ n894 ^ 1'b0 ;
  assign n32411 = x58 & n32410 ;
  assign y0 = x10 ;
  assign y1 = x15 ;
  assign y2 = x21 ;
  assign y3 = x30 ;
  assign y4 = x42 ;
  assign y5 = x54 ;
  assign y6 = x66 ;
  assign y7 = x79 ;
  assign y8 = x93 ;
  assign y9 = x110 ;
  assign y10 = x111 ;
  assign y11 = x113 ;
  assign y12 = x114 ;
  assign y13 = x120 ;
  assign y14 = n131 ;
  assign y15 = ~1'b0 ;
  assign y16 = ~n136 ;
  assign y17 = ~n138 ;
  assign y18 = ~n139 ;
  assign y19 = ~n143 ;
  assign y20 = n144 ;
  assign y21 = ~n147 ;
  assign y22 = n150 ;
  assign y23 = ~n152 ;
  assign y24 = n153 ;
  assign y25 = ~n162 ;
  assign y26 = n174 ;
  assign y27 = ~n178 ;
  assign y28 = ~n179 ;
  assign y29 = ~n191 ;
  assign y30 = ~n199 ;
  assign y31 = n201 ;
  assign y32 = ~n205 ;
  assign y33 = ~n219 ;
  assign y34 = n228 ;
  assign y35 = ~n235 ;
  assign y36 = ~n238 ;
  assign y37 = n242 ;
  assign y38 = n248 ;
  assign y39 = ~n255 ;
  assign y40 = n261 ;
  assign y41 = ~n266 ;
  assign y42 = n278 ;
  assign y43 = n280 ;
  assign y44 = n282 ;
  assign y45 = n289 ;
  assign y46 = n292 ;
  assign y47 = n294 ;
  assign y48 = ~1'b0 ;
  assign y49 = n304 ;
  assign y50 = n314 ;
  assign y51 = ~n319 ;
  assign y52 = ~n320 ;
  assign y53 = ~n325 ;
  assign y54 = ~n334 ;
  assign y55 = ~n337 ;
  assign y56 = ~n339 ;
  assign y57 = n346 ;
  assign y58 = ~n354 ;
  assign y59 = n368 ;
  assign y60 = n375 ;
  assign y61 = n386 ;
  assign y62 = ~1'b0 ;
  assign y63 = ~n395 ;
  assign y64 = ~n397 ;
  assign y65 = n407 ;
  assign y66 = n409 ;
  assign y67 = ~1'b0 ;
  assign y68 = n410 ;
  assign y69 = ~n414 ;
  assign y70 = ~n418 ;
  assign y71 = ~n421 ;
  assign y72 = n426 ;
  assign y73 = n440 ;
  assign y74 = n448 ;
  assign y75 = n459 ;
  assign y76 = n464 ;
  assign y77 = n465 ;
  assign y78 = ~1'b0 ;
  assign y79 = ~n468 ;
  assign y80 = ~n488 ;
  assign y81 = ~n500 ;
  assign y82 = ~n501 ;
  assign y83 = ~n505 ;
  assign y84 = ~n508 ;
  assign y85 = ~n515 ;
  assign y86 = ~n549 ;
  assign y87 = ~n562 ;
  assign y88 = ~n572 ;
  assign y89 = ~n579 ;
  assign y90 = ~n598 ;
  assign y91 = n599 ;
  assign y92 = ~n605 ;
  assign y93 = ~n618 ;
  assign y94 = ~n636 ;
  assign y95 = n643 ;
  assign y96 = n646 ;
  assign y97 = ~n659 ;
  assign y98 = n662 ;
  assign y99 = ~n665 ;
  assign y100 = ~1'b0 ;
  assign y101 = n678 ;
  assign y102 = ~n681 ;
  assign y103 = n692 ;
  assign y104 = ~n694 ;
  assign y105 = n695 ;
  assign y106 = n708 ;
  assign y107 = ~n711 ;
  assign y108 = n712 ;
  assign y109 = n714 ;
  assign y110 = n719 ;
  assign y111 = ~n737 ;
  assign y112 = n753 ;
  assign y113 = ~1'b0 ;
  assign y114 = n756 ;
  assign y115 = n761 ;
  assign y116 = n765 ;
  assign y117 = n770 ;
  assign y118 = n773 ;
  assign y119 = ~n775 ;
  assign y120 = ~n778 ;
  assign y121 = ~n788 ;
  assign y122 = n797 ;
  assign y123 = n800 ;
  assign y124 = n801 ;
  assign y125 = ~n804 ;
  assign y126 = ~n805 ;
  assign y127 = n806 ;
  assign y128 = n810 ;
  assign y129 = n817 ;
  assign y130 = n833 ;
  assign y131 = ~n835 ;
  assign y132 = n840 ;
  assign y133 = ~n842 ;
  assign y134 = n854 ;
  assign y135 = n857 ;
  assign y136 = n862 ;
  assign y137 = n863 ;
  assign y138 = n864 ;
  assign y139 = ~n868 ;
  assign y140 = ~n872 ;
  assign y141 = n876 ;
  assign y142 = n879 ;
  assign y143 = ~n883 ;
  assign y144 = ~n887 ;
  assign y145 = ~n891 ;
  assign y146 = ~n893 ;
  assign y147 = ~n901 ;
  assign y148 = n906 ;
  assign y149 = ~n909 ;
  assign y150 = n913 ;
  assign y151 = ~n916 ;
  assign y152 = ~n917 ;
  assign y153 = n930 ;
  assign y154 = ~1'b0 ;
  assign y155 = ~n932 ;
  assign y156 = ~n940 ;
  assign y157 = ~n948 ;
  assign y158 = n949 ;
  assign y159 = n952 ;
  assign y160 = n953 ;
  assign y161 = n960 ;
  assign y162 = ~n974 ;
  assign y163 = n990 ;
  assign y164 = n997 ;
  assign y165 = n1003 ;
  assign y166 = ~n1007 ;
  assign y167 = ~n1011 ;
  assign y168 = n1018 ;
  assign y169 = n1025 ;
  assign y170 = ~n1031 ;
  assign y171 = ~n1035 ;
  assign y172 = ~n1039 ;
  assign y173 = ~1'b0 ;
  assign y174 = ~1'b0 ;
  assign y175 = n1042 ;
  assign y176 = ~n1053 ;
  assign y177 = ~n1056 ;
  assign y178 = n1058 ;
  assign y179 = ~n1059 ;
  assign y180 = ~n1064 ;
  assign y181 = ~n1068 ;
  assign y182 = ~1'b0 ;
  assign y183 = n1086 ;
  assign y184 = n1088 ;
  assign y185 = n1107 ;
  assign y186 = n1110 ;
  assign y187 = ~n1112 ;
  assign y188 = ~n1114 ;
  assign y189 = ~n1115 ;
  assign y190 = n1135 ;
  assign y191 = ~1'b0 ;
  assign y192 = n1144 ;
  assign y193 = ~n1145 ;
  assign y194 = ~1'b0 ;
  assign y195 = ~n1160 ;
  assign y196 = ~n1181 ;
  assign y197 = n1187 ;
  assign y198 = ~n1189 ;
  assign y199 = n1195 ;
  assign y200 = n1207 ;
  assign y201 = ~1'b0 ;
  assign y202 = ~n1215 ;
  assign y203 = ~n1218 ;
  assign y204 = n1219 ;
  assign y205 = n1222 ;
  assign y206 = n1228 ;
  assign y207 = n1229 ;
  assign y208 = ~1'b0 ;
  assign y209 = ~n1230 ;
  assign y210 = ~n1237 ;
  assign y211 = n1243 ;
  assign y212 = ~n1245 ;
  assign y213 = n1250 ;
  assign y214 = ~n1254 ;
  assign y215 = n1268 ;
  assign y216 = n1271 ;
  assign y217 = ~n1278 ;
  assign y218 = n1283 ;
  assign y219 = ~n1284 ;
  assign y220 = ~n1290 ;
  assign y221 = n1300 ;
  assign y222 = n1309 ;
  assign y223 = ~n1315 ;
  assign y224 = ~1'b0 ;
  assign y225 = ~n1322 ;
  assign y226 = ~n1325 ;
  assign y227 = ~n1328 ;
  assign y228 = n1338 ;
  assign y229 = n1342 ;
  assign y230 = ~n1343 ;
  assign y231 = ~n1349 ;
  assign y232 = ~n1361 ;
  assign y233 = n1378 ;
  assign y234 = n1382 ;
  assign y235 = n1385 ;
  assign y236 = ~n1386 ;
  assign y237 = n1387 ;
  assign y238 = n1394 ;
  assign y239 = ~1'b0 ;
  assign y240 = ~n1397 ;
  assign y241 = ~1'b0 ;
  assign y242 = ~n1409 ;
  assign y243 = ~n1414 ;
  assign y244 = ~n1084 ;
  assign y245 = n1415 ;
  assign y246 = ~n1435 ;
  assign y247 = ~n1448 ;
  assign y248 = ~n1457 ;
  assign y249 = ~n1458 ;
  assign y250 = ~n1466 ;
  assign y251 = n1471 ;
  assign y252 = n1475 ;
  assign y253 = n1477 ;
  assign y254 = n1482 ;
  assign y255 = ~n1492 ;
  assign y256 = n1508 ;
  assign y257 = ~n1511 ;
  assign y258 = ~n1527 ;
  assign y259 = n1531 ;
  assign y260 = n1537 ;
  assign y261 = n1541 ;
  assign y262 = ~n1552 ;
  assign y263 = n1576 ;
  assign y264 = n1579 ;
  assign y265 = n1582 ;
  assign y266 = n1591 ;
  assign y267 = ~n1604 ;
  assign y268 = ~n1606 ;
  assign y269 = ~n1625 ;
  assign y270 = n1641 ;
  assign y271 = ~n1644 ;
  assign y272 = n1648 ;
  assign y273 = n1665 ;
  assign y274 = ~n1670 ;
  assign y275 = ~n1672 ;
  assign y276 = ~n1675 ;
  assign y277 = ~n1680 ;
  assign y278 = ~n1682 ;
  assign y279 = ~n1687 ;
  assign y280 = n1690 ;
  assign y281 = n1693 ;
  assign y282 = ~n1694 ;
  assign y283 = n1695 ;
  assign y284 = n1701 ;
  assign y285 = ~n1707 ;
  assign y286 = n1708 ;
  assign y287 = n1711 ;
  assign y288 = n1719 ;
  assign y289 = ~n1729 ;
  assign y290 = ~n1731 ;
  assign y291 = ~n1732 ;
  assign y292 = ~n1733 ;
  assign y293 = n1735 ;
  assign y294 = ~n1736 ;
  assign y295 = ~n1737 ;
  assign y296 = n1751 ;
  assign y297 = ~n1757 ;
  assign y298 = n1759 ;
  assign y299 = n1767 ;
  assign y300 = ~n1779 ;
  assign y301 = n1783 ;
  assign y302 = ~1'b0 ;
  assign y303 = n1791 ;
  assign y304 = ~n1794 ;
  assign y305 = ~n1797 ;
  assign y306 = n1803 ;
  assign y307 = n1820 ;
  assign y308 = ~n1841 ;
  assign y309 = ~n1844 ;
  assign y310 = n1850 ;
  assign y311 = n1866 ;
  assign y312 = n1870 ;
  assign y313 = ~n1871 ;
  assign y314 = n1873 ;
  assign y315 = n1879 ;
  assign y316 = ~n1901 ;
  assign y317 = ~1'b0 ;
  assign y318 = n1913 ;
  assign y319 = ~n1916 ;
  assign y320 = n1922 ;
  assign y321 = ~1'b0 ;
  assign y322 = ~n1926 ;
  assign y323 = n1930 ;
  assign y324 = ~n1933 ;
  assign y325 = n1944 ;
  assign y326 = ~n1948 ;
  assign y327 = ~n1968 ;
  assign y328 = ~n1977 ;
  assign y329 = n1979 ;
  assign y330 = n1985 ;
  assign y331 = n1992 ;
  assign y332 = ~n1997 ;
  assign y333 = ~n1999 ;
  assign y334 = ~n2007 ;
  assign y335 = ~n2013 ;
  assign y336 = ~n2019 ;
  assign y337 = ~n2023 ;
  assign y338 = ~n2027 ;
  assign y339 = ~n2030 ;
  assign y340 = ~n2039 ;
  assign y341 = n2045 ;
  assign y342 = ~n2053 ;
  assign y343 = ~n2058 ;
  assign y344 = n2071 ;
  assign y345 = n2075 ;
  assign y346 = ~n2081 ;
  assign y347 = ~n2083 ;
  assign y348 = ~n2100 ;
  assign y349 = n2104 ;
  assign y350 = ~n2110 ;
  assign y351 = ~n2113 ;
  assign y352 = ~n2124 ;
  assign y353 = ~1'b0 ;
  assign y354 = n2143 ;
  assign y355 = ~n2152 ;
  assign y356 = n2153 ;
  assign y357 = ~n2154 ;
  assign y358 = n2164 ;
  assign y359 = n2168 ;
  assign y360 = n2169 ;
  assign y361 = ~n2179 ;
  assign y362 = n2182 ;
  assign y363 = ~n2195 ;
  assign y364 = ~n2198 ;
  assign y365 = ~n2202 ;
  assign y366 = ~n2205 ;
  assign y367 = ~n2208 ;
  assign y368 = n2225 ;
  assign y369 = ~n425 ;
  assign y370 = ~n2230 ;
  assign y371 = ~n2236 ;
  assign y372 = ~n2238 ;
  assign y373 = n2239 ;
  assign y374 = n2240 ;
  assign y375 = ~n2249 ;
  assign y376 = ~n2252 ;
  assign y377 = n2264 ;
  assign y378 = ~n2272 ;
  assign y379 = ~n2285 ;
  assign y380 = n2296 ;
  assign y381 = ~n2300 ;
  assign y382 = n2304 ;
  assign y383 = ~n2306 ;
  assign y384 = ~n2312 ;
  assign y385 = ~n2316 ;
  assign y386 = n2322 ;
  assign y387 = n2326 ;
  assign y388 = ~n2334 ;
  assign y389 = n2336 ;
  assign y390 = n2337 ;
  assign y391 = n2340 ;
  assign y392 = n2346 ;
  assign y393 = ~n2350 ;
  assign y394 = ~n2353 ;
  assign y395 = n2354 ;
  assign y396 = n2381 ;
  assign y397 = ~n2383 ;
  assign y398 = ~n2389 ;
  assign y399 = ~n2398 ;
  assign y400 = ~1'b0 ;
  assign y401 = n2408 ;
  assign y402 = n2415 ;
  assign y403 = n2421 ;
  assign y404 = ~n2429 ;
  assign y405 = n2431 ;
  assign y406 = n2433 ;
  assign y407 = ~n2439 ;
  assign y408 = n2446 ;
  assign y409 = n2449 ;
  assign y410 = n2457 ;
  assign y411 = n2471 ;
  assign y412 = ~n2472 ;
  assign y413 = ~n2479 ;
  assign y414 = n2482 ;
  assign y415 = ~n2484 ;
  assign y416 = ~n2486 ;
  assign y417 = n2517 ;
  assign y418 = ~1'b0 ;
  assign y419 = n2535 ;
  assign y420 = n2536 ;
  assign y421 = ~n2537 ;
  assign y422 = ~1'b0 ;
  assign y423 = n2561 ;
  assign y424 = ~1'b0 ;
  assign y425 = n2570 ;
  assign y426 = ~n2572 ;
  assign y427 = n2574 ;
  assign y428 = ~n2575 ;
  assign y429 = n2584 ;
  assign y430 = ~n2585 ;
  assign y431 = n2588 ;
  assign y432 = n2594 ;
  assign y433 = n2602 ;
  assign y434 = n2608 ;
  assign y435 = n2613 ;
  assign y436 = ~n2617 ;
  assign y437 = n2625 ;
  assign y438 = n2632 ;
  assign y439 = ~n2644 ;
  assign y440 = ~n2647 ;
  assign y441 = n2648 ;
  assign y442 = n2649 ;
  assign y443 = ~n2652 ;
  assign y444 = ~1'b0 ;
  assign y445 = ~n2668 ;
  assign y446 = ~n2696 ;
  assign y447 = n2700 ;
  assign y448 = ~n2701 ;
  assign y449 = ~n2735 ;
  assign y450 = ~n2740 ;
  assign y451 = ~n2743 ;
  assign y452 = ~n2745 ;
  assign y453 = n2747 ;
  assign y454 = n2748 ;
  assign y455 = n2753 ;
  assign y456 = ~n2755 ;
  assign y457 = ~n2760 ;
  assign y458 = ~n2771 ;
  assign y459 = ~n2777 ;
  assign y460 = n2801 ;
  assign y461 = n2804 ;
  assign y462 = ~n2808 ;
  assign y463 = 1'b0 ;
  assign y464 = n2818 ;
  assign y465 = n2828 ;
  assign y466 = n2829 ;
  assign y467 = ~n2836 ;
  assign y468 = n2847 ;
  assign y469 = ~n2850 ;
  assign y470 = n2861 ;
  assign y471 = ~1'b0 ;
  assign y472 = ~n2864 ;
  assign y473 = ~n2866 ;
  assign y474 = ~n2874 ;
  assign y475 = n2889 ;
  assign y476 = n2895 ;
  assign y477 = ~n2896 ;
  assign y478 = ~n2906 ;
  assign y479 = n2909 ;
  assign y480 = n2913 ;
  assign y481 = ~n2915 ;
  assign y482 = ~n2920 ;
  assign y483 = ~n2928 ;
  assign y484 = n2944 ;
  assign y485 = n2948 ;
  assign y486 = ~n2950 ;
  assign y487 = ~n2957 ;
  assign y488 = ~1'b0 ;
  assign y489 = n2966 ;
  assign y490 = ~1'b0 ;
  assign y491 = n2967 ;
  assign y492 = n2972 ;
  assign y493 = n2978 ;
  assign y494 = n2984 ;
  assign y495 = ~n2987 ;
  assign y496 = ~n2991 ;
  assign y497 = n2993 ;
  assign y498 = ~n2999 ;
  assign y499 = n3004 ;
  assign y500 = ~n3006 ;
  assign y501 = n3008 ;
  assign y502 = n3011 ;
  assign y503 = n3014 ;
  assign y504 = ~n3018 ;
  assign y505 = n3022 ;
  assign y506 = ~n3032 ;
  assign y507 = n3038 ;
  assign y508 = n3044 ;
  assign y509 = ~n3047 ;
  assign y510 = ~n3051 ;
  assign y511 = n3052 ;
  assign y512 = n3054 ;
  assign y513 = ~n3058 ;
  assign y514 = ~n3060 ;
  assign y515 = ~n3074 ;
  assign y516 = n3090 ;
  assign y517 = ~n3091 ;
  assign y518 = n3099 ;
  assign y519 = ~n3104 ;
  assign y520 = ~n3118 ;
  assign y521 = n3129 ;
  assign y522 = ~n3130 ;
  assign y523 = ~n3134 ;
  assign y524 = ~n3145 ;
  assign y525 = n3150 ;
  assign y526 = ~n3153 ;
  assign y527 = n3158 ;
  assign y528 = n3170 ;
  assign y529 = n3187 ;
  assign y530 = n3191 ;
  assign y531 = ~1'b0 ;
  assign y532 = n3205 ;
  assign y533 = ~n3209 ;
  assign y534 = ~n3216 ;
  assign y535 = n3232 ;
  assign y536 = ~n3246 ;
  assign y537 = n3247 ;
  assign y538 = n3250 ;
  assign y539 = ~n3252 ;
  assign y540 = ~n3253 ;
  assign y541 = ~n3255 ;
  assign y542 = n3262 ;
  assign y543 = ~n3275 ;
  assign y544 = n3278 ;
  assign y545 = n3289 ;
  assign y546 = ~1'b0 ;
  assign y547 = ~n3290 ;
  assign y548 = ~n3292 ;
  assign y549 = ~1'b0 ;
  assign y550 = n3295 ;
  assign y551 = ~n3299 ;
  assign y552 = n3303 ;
  assign y553 = ~n3314 ;
  assign y554 = ~n3321 ;
  assign y555 = n3323 ;
  assign y556 = n3324 ;
  assign y557 = n3328 ;
  assign y558 = n3329 ;
  assign y559 = n3346 ;
  assign y560 = ~n3348 ;
  assign y561 = ~1'b0 ;
  assign y562 = n3349 ;
  assign y563 = n3352 ;
  assign y564 = ~n3353 ;
  assign y565 = n3362 ;
  assign y566 = n3364 ;
  assign y567 = n3378 ;
  assign y568 = n3387 ;
  assign y569 = ~n3398 ;
  assign y570 = ~n3402 ;
  assign y571 = n3405 ;
  assign y572 = n3411 ;
  assign y573 = n3413 ;
  assign y574 = ~n3418 ;
  assign y575 = n3439 ;
  assign y576 = ~n3443 ;
  assign y577 = ~n3453 ;
  assign y578 = ~n3457 ;
  assign y579 = n3459 ;
  assign y580 = ~1'b0 ;
  assign y581 = n3462 ;
  assign y582 = ~n3464 ;
  assign y583 = ~n3469 ;
  assign y584 = ~n3475 ;
  assign y585 = ~n3479 ;
  assign y586 = ~n3481 ;
  assign y587 = n3493 ;
  assign y588 = ~n3494 ;
  assign y589 = ~1'b0 ;
  assign y590 = n3497 ;
  assign y591 = ~n3503 ;
  assign y592 = n3509 ;
  assign y593 = ~n3511 ;
  assign y594 = ~n3519 ;
  assign y595 = ~n3530 ;
  assign y596 = n3532 ;
  assign y597 = ~n3554 ;
  assign y598 = n3557 ;
  assign y599 = n3558 ;
  assign y600 = n3570 ;
  assign y601 = ~n3588 ;
  assign y602 = n3591 ;
  assign y603 = ~1'b0 ;
  assign y604 = ~n3599 ;
  assign y605 = n3602 ;
  assign y606 = n3608 ;
  assign y607 = n3615 ;
  assign y608 = ~n3625 ;
  assign y609 = ~n3629 ;
  assign y610 = ~n3634 ;
  assign y611 = n3637 ;
  assign y612 = ~n3656 ;
  assign y613 = ~n3659 ;
  assign y614 = ~1'b0 ;
  assign y615 = ~n3663 ;
  assign y616 = ~n3674 ;
  assign y617 = ~n3682 ;
  assign y618 = ~n3689 ;
  assign y619 = ~1'b0 ;
  assign y620 = ~1'b0 ;
  assign y621 = ~n3702 ;
  assign y622 = ~n3725 ;
  assign y623 = ~n3726 ;
  assign y624 = ~n3727 ;
  assign y625 = n3729 ;
  assign y626 = n3732 ;
  assign y627 = n3735 ;
  assign y628 = ~n3736 ;
  assign y629 = n3739 ;
  assign y630 = ~n3745 ;
  assign y631 = ~n3753 ;
  assign y632 = n3758 ;
  assign y633 = ~n3759 ;
  assign y634 = n3763 ;
  assign y635 = n3768 ;
  assign y636 = n3772 ;
  assign y637 = ~1'b0 ;
  assign y638 = ~1'b0 ;
  assign y639 = n3774 ;
  assign y640 = ~n3781 ;
  assign y641 = ~n3800 ;
  assign y642 = ~n3802 ;
  assign y643 = n3804 ;
  assign y644 = n3808 ;
  assign y645 = n3814 ;
  assign y646 = n3830 ;
  assign y647 = ~n3831 ;
  assign y648 = n3833 ;
  assign y649 = ~n3839 ;
  assign y650 = ~1'b0 ;
  assign y651 = ~n3848 ;
  assign y652 = ~n3857 ;
  assign y653 = n3862 ;
  assign y654 = ~1'b0 ;
  assign y655 = ~1'b0 ;
  assign y656 = ~n3879 ;
  assign y657 = ~1'b0 ;
  assign y658 = ~n3884 ;
  assign y659 = ~n3885 ;
  assign y660 = ~n3889 ;
  assign y661 = n3904 ;
  assign y662 = ~n3909 ;
  assign y663 = ~n3913 ;
  assign y664 = n3919 ;
  assign y665 = ~n3924 ;
  assign y666 = n3939 ;
  assign y667 = n3951 ;
  assign y668 = ~n3958 ;
  assign y669 = n3965 ;
  assign y670 = n3967 ;
  assign y671 = n3969 ;
  assign y672 = n3974 ;
  assign y673 = n3977 ;
  assign y674 = n3978 ;
  assign y675 = ~n3986 ;
  assign y676 = n3988 ;
  assign y677 = ~n3991 ;
  assign y678 = ~n3992 ;
  assign y679 = ~n4004 ;
  assign y680 = ~1'b0 ;
  assign y681 = n4017 ;
  assign y682 = n4018 ;
  assign y683 = n4019 ;
  assign y684 = ~n4021 ;
  assign y685 = n4028 ;
  assign y686 = ~n4034 ;
  assign y687 = ~n4041 ;
  assign y688 = ~n4048 ;
  assign y689 = ~n4050 ;
  assign y690 = ~n4052 ;
  assign y691 = n4055 ;
  assign y692 = ~n4063 ;
  assign y693 = ~n4066 ;
  assign y694 = n4083 ;
  assign y695 = n4090 ;
  assign y696 = n4104 ;
  assign y697 = n4106 ;
  assign y698 = ~1'b0 ;
  assign y699 = ~n4110 ;
  assign y700 = ~1'b0 ;
  assign y701 = n4111 ;
  assign y702 = ~n4113 ;
  assign y703 = n4143 ;
  assign y704 = n4147 ;
  assign y705 = ~n4151 ;
  assign y706 = n4153 ;
  assign y707 = n4155 ;
  assign y708 = ~n4159 ;
  assign y709 = n4172 ;
  assign y710 = n4180 ;
  assign y711 = n4186 ;
  assign y712 = ~n4188 ;
  assign y713 = n4193 ;
  assign y714 = n4205 ;
  assign y715 = ~n4214 ;
  assign y716 = n4216 ;
  assign y717 = ~n4219 ;
  assign y718 = ~n4221 ;
  assign y719 = n4223 ;
  assign y720 = n4228 ;
  assign y721 = ~n4230 ;
  assign y722 = ~n4239 ;
  assign y723 = ~n4242 ;
  assign y724 = n4252 ;
  assign y725 = n4255 ;
  assign y726 = ~1'b0 ;
  assign y727 = n4258 ;
  assign y728 = ~n4259 ;
  assign y729 = ~n4264 ;
  assign y730 = n4269 ;
  assign y731 = ~n4273 ;
  assign y732 = n4275 ;
  assign y733 = n4281 ;
  assign y734 = n4282 ;
  assign y735 = n4284 ;
  assign y736 = ~n4291 ;
  assign y737 = ~n4301 ;
  assign y738 = ~1'b0 ;
  assign y739 = ~1'b0 ;
  assign y740 = ~n4311 ;
  assign y741 = ~n4316 ;
  assign y742 = n4328 ;
  assign y743 = n4330 ;
  assign y744 = ~n4332 ;
  assign y745 = ~n4342 ;
  assign y746 = n4345 ;
  assign y747 = ~n4354 ;
  assign y748 = ~n4361 ;
  assign y749 = n4367 ;
  assign y750 = ~n4386 ;
  assign y751 = n4388 ;
  assign y752 = n4394 ;
  assign y753 = ~1'b0 ;
  assign y754 = n4405 ;
  assign y755 = n4415 ;
  assign y756 = n4432 ;
  assign y757 = ~n4442 ;
  assign y758 = n4443 ;
  assign y759 = n4446 ;
  assign y760 = ~n4448 ;
  assign y761 = n4460 ;
  assign y762 = ~1'b0 ;
  assign y763 = ~n4470 ;
  assign y764 = n4480 ;
  assign y765 = ~n4490 ;
  assign y766 = n4493 ;
  assign y767 = ~n4501 ;
  assign y768 = n4504 ;
  assign y769 = n4506 ;
  assign y770 = ~1'b0 ;
  assign y771 = ~n4516 ;
  assign y772 = ~n4521 ;
  assign y773 = ~n4522 ;
  assign y774 = ~n4528 ;
  assign y775 = n4534 ;
  assign y776 = ~n4538 ;
  assign y777 = ~n4540 ;
  assign y778 = ~n4281 ;
  assign y779 = n4543 ;
  assign y780 = ~n4545 ;
  assign y781 = n4552 ;
  assign y782 = ~n4557 ;
  assign y783 = ~1'b0 ;
  assign y784 = n4563 ;
  assign y785 = ~n4575 ;
  assign y786 = n4579 ;
  assign y787 = n4591 ;
  assign y788 = ~n4601 ;
  assign y789 = ~1'b0 ;
  assign y790 = ~n4608 ;
  assign y791 = ~1'b0 ;
  assign y792 = ~n4611 ;
  assign y793 = n4623 ;
  assign y794 = ~n4625 ;
  assign y795 = ~n4632 ;
  assign y796 = ~1'b0 ;
  assign y797 = n4643 ;
  assign y798 = ~n4658 ;
  assign y799 = ~n4659 ;
  assign y800 = n4678 ;
  assign y801 = ~n4682 ;
  assign y802 = n4683 ;
  assign y803 = ~n4710 ;
  assign y804 = ~n4720 ;
  assign y805 = ~1'b0 ;
  assign y806 = ~n4726 ;
  assign y807 = n4743 ;
  assign y808 = ~n4746 ;
  assign y809 = ~n4747 ;
  assign y810 = n4749 ;
  assign y811 = ~n4751 ;
  assign y812 = ~n4761 ;
  assign y813 = n4766 ;
  assign y814 = ~1'b0 ;
  assign y815 = n4771 ;
  assign y816 = n4775 ;
  assign y817 = n956 ;
  assign y818 = n4776 ;
  assign y819 = n4781 ;
  assign y820 = n4785 ;
  assign y821 = n4799 ;
  assign y822 = n4801 ;
  assign y823 = ~n4808 ;
  assign y824 = n4810 ;
  assign y825 = ~n4815 ;
  assign y826 = n4822 ;
  assign y827 = ~n4834 ;
  assign y828 = ~n4842 ;
  assign y829 = n4844 ;
  assign y830 = ~n4859 ;
  assign y831 = ~n4869 ;
  assign y832 = ~1'b0 ;
  assign y833 = ~n4872 ;
  assign y834 = ~n4874 ;
  assign y835 = ~n4881 ;
  assign y836 = ~n4889 ;
  assign y837 = ~n4903 ;
  assign y838 = n4911 ;
  assign y839 = ~n4917 ;
  assign y840 = ~n4925 ;
  assign y841 = ~n4927 ;
  assign y842 = n4935 ;
  assign y843 = ~n4937 ;
  assign y844 = ~n4949 ;
  assign y845 = ~n4954 ;
  assign y846 = n4955 ;
  assign y847 = ~1'b0 ;
  assign y848 = n4962 ;
  assign y849 = n4968 ;
  assign y850 = ~n4971 ;
  assign y851 = ~n4981 ;
  assign y852 = n4982 ;
  assign y853 = ~n4984 ;
  assign y854 = ~n4986 ;
  assign y855 = n4998 ;
  assign y856 = n5011 ;
  assign y857 = n5040 ;
  assign y858 = n5041 ;
  assign y859 = n5051 ;
  assign y860 = ~n5055 ;
  assign y861 = n5065 ;
  assign y862 = ~n5066 ;
  assign y863 = ~n5067 ;
  assign y864 = ~1'b0 ;
  assign y865 = ~n5071 ;
  assign y866 = n5078 ;
  assign y867 = ~1'b0 ;
  assign y868 = ~n5081 ;
  assign y869 = ~n5085 ;
  assign y870 = n5093 ;
  assign y871 = ~n5095 ;
  assign y872 = n5101 ;
  assign y873 = n5117 ;
  assign y874 = n5120 ;
  assign y875 = n5122 ;
  assign y876 = ~n5127 ;
  assign y877 = ~n5130 ;
  assign y878 = n5135 ;
  assign y879 = ~n5147 ;
  assign y880 = ~n5151 ;
  assign y881 = ~n5152 ;
  assign y882 = n5155 ;
  assign y883 = ~n5158 ;
  assign y884 = n5164 ;
  assign y885 = ~n5168 ;
  assign y886 = n5172 ;
  assign y887 = ~n5179 ;
  assign y888 = ~n5187 ;
  assign y889 = ~n5191 ;
  assign y890 = n5193 ;
  assign y891 = n5197 ;
  assign y892 = ~n5201 ;
  assign y893 = n5220 ;
  assign y894 = ~n5225 ;
  assign y895 = n5239 ;
  assign y896 = ~n5243 ;
  assign y897 = n5262 ;
  assign y898 = ~n5263 ;
  assign y899 = n5268 ;
  assign y900 = ~n5271 ;
  assign y901 = ~1'b0 ;
  assign y902 = ~1'b0 ;
  assign y903 = ~n5278 ;
  assign y904 = ~n5290 ;
  assign y905 = n5294 ;
  assign y906 = n5304 ;
  assign y907 = ~n5321 ;
  assign y908 = ~1'b0 ;
  assign y909 = ~n5322 ;
  assign y910 = ~n5334 ;
  assign y911 = n5338 ;
  assign y912 = n5339 ;
  assign y913 = n5342 ;
  assign y914 = n5343 ;
  assign y915 = n5345 ;
  assign y916 = n5347 ;
  assign y917 = ~1'b0 ;
  assign y918 = ~n5349 ;
  assign y919 = ~n5357 ;
  assign y920 = ~n5377 ;
  assign y921 = n5393 ;
  assign y922 = ~n5396 ;
  assign y923 = ~n5398 ;
  assign y924 = ~n5401 ;
  assign y925 = n5405 ;
  assign y926 = ~n5409 ;
  assign y927 = ~1'b0 ;
  assign y928 = ~n5411 ;
  assign y929 = ~1'b0 ;
  assign y930 = ~n5422 ;
  assign y931 = n5425 ;
  assign y932 = n5434 ;
  assign y933 = n5441 ;
  assign y934 = n5449 ;
  assign y935 = ~n5456 ;
  assign y936 = n5457 ;
  assign y937 = ~n5459 ;
  assign y938 = n5461 ;
  assign y939 = ~1'b0 ;
  assign y940 = ~n5464 ;
  assign y941 = ~1'b0 ;
  assign y942 = n5466 ;
  assign y943 = ~n5470 ;
  assign y944 = ~n5471 ;
  assign y945 = n5472 ;
  assign y946 = ~n5480 ;
  assign y947 = ~n5508 ;
  assign y948 = n5512 ;
  assign y949 = ~n5523 ;
  assign y950 = ~n5525 ;
  assign y951 = ~n5527 ;
  assign y952 = ~n5532 ;
  assign y953 = ~1'b0 ;
  assign y954 = ~n5537 ;
  assign y955 = ~n5539 ;
  assign y956 = ~n5541 ;
  assign y957 = n5545 ;
  assign y958 = n5550 ;
  assign y959 = n5557 ;
  assign y960 = ~n5564 ;
  assign y961 = ~n5568 ;
  assign y962 = ~n5569 ;
  assign y963 = n5575 ;
  assign y964 = n5577 ;
  assign y965 = n5591 ;
  assign y966 = n5596 ;
  assign y967 = ~n5605 ;
  assign y968 = n5607 ;
  assign y969 = n5616 ;
  assign y970 = n5621 ;
  assign y971 = n5627 ;
  assign y972 = n5628 ;
  assign y973 = n5629 ;
  assign y974 = ~n5635 ;
  assign y975 = ~n5637 ;
  assign y976 = ~n5647 ;
  assign y977 = n5654 ;
  assign y978 = n5656 ;
  assign y979 = n5664 ;
  assign y980 = n5666 ;
  assign y981 = n5677 ;
  assign y982 = ~n5698 ;
  assign y983 = ~n5718 ;
  assign y984 = ~n5723 ;
  assign y985 = n5724 ;
  assign y986 = ~n5735 ;
  assign y987 = ~n5745 ;
  assign y988 = ~n5750 ;
  assign y989 = ~n5751 ;
  assign y990 = ~n5762 ;
  assign y991 = n5765 ;
  assign y992 = ~n5766 ;
  assign y993 = ~n5768 ;
  assign y994 = ~n5772 ;
  assign y995 = ~n5775 ;
  assign y996 = ~n5777 ;
  assign y997 = ~n5780 ;
  assign y998 = ~n5781 ;
  assign y999 = ~n5787 ;
  assign y1000 = ~n5789 ;
  assign y1001 = ~n5792 ;
  assign y1002 = ~n5798 ;
  assign y1003 = n5807 ;
  assign y1004 = ~n5810 ;
  assign y1005 = ~n5811 ;
  assign y1006 = n5812 ;
  assign y1007 = ~n5815 ;
  assign y1008 = ~n5819 ;
  assign y1009 = ~n5820 ;
  assign y1010 = ~n5821 ;
  assign y1011 = n5826 ;
  assign y1012 = ~n5827 ;
  assign y1013 = n5833 ;
  assign y1014 = ~n5840 ;
  assign y1015 = n5846 ;
  assign y1016 = ~n5847 ;
  assign y1017 = ~n5849 ;
  assign y1018 = ~n5856 ;
  assign y1019 = n5860 ;
  assign y1020 = n5874 ;
  assign y1021 = ~n5877 ;
  assign y1022 = n5887 ;
  assign y1023 = ~n5889 ;
  assign y1024 = n5894 ;
  assign y1025 = n5895 ;
  assign y1026 = ~n5913 ;
  assign y1027 = ~n5923 ;
  assign y1028 = ~n5934 ;
  assign y1029 = ~1'b0 ;
  assign y1030 = ~n5938 ;
  assign y1031 = ~n5940 ;
  assign y1032 = ~n5948 ;
  assign y1033 = ~1'b0 ;
  assign y1034 = ~n5951 ;
  assign y1035 = ~1'b0 ;
  assign y1036 = n5970 ;
  assign y1037 = n5992 ;
  assign y1038 = ~n5995 ;
  assign y1039 = ~n5998 ;
  assign y1040 = ~n6001 ;
  assign y1041 = n6002 ;
  assign y1042 = n6011 ;
  assign y1043 = ~n6018 ;
  assign y1044 = ~n6019 ;
  assign y1045 = n6022 ;
  assign y1046 = ~n6035 ;
  assign y1047 = ~1'b0 ;
  assign y1048 = ~n6036 ;
  assign y1049 = ~n6039 ;
  assign y1050 = n6041 ;
  assign y1051 = n6042 ;
  assign y1052 = n6051 ;
  assign y1053 = ~n6054 ;
  assign y1054 = n6056 ;
  assign y1055 = n6063 ;
  assign y1056 = n6085 ;
  assign y1057 = ~n6086 ;
  assign y1058 = ~n6097 ;
  assign y1059 = n6109 ;
  assign y1060 = ~n6115 ;
  assign y1061 = n6144 ;
  assign y1062 = ~n6151 ;
  assign y1063 = n6153 ;
  assign y1064 = ~n6155 ;
  assign y1065 = ~n6181 ;
  assign y1066 = ~n6182 ;
  assign y1067 = ~n6192 ;
  assign y1068 = n6195 ;
  assign y1069 = ~n6200 ;
  assign y1070 = n6205 ;
  assign y1071 = ~n6207 ;
  assign y1072 = n6213 ;
  assign y1073 = ~n6222 ;
  assign y1074 = n6238 ;
  assign y1075 = n6240 ;
  assign y1076 = ~n6242 ;
  assign y1077 = ~1'b0 ;
  assign y1078 = n6248 ;
  assign y1079 = ~n6250 ;
  assign y1080 = n6257 ;
  assign y1081 = ~n6258 ;
  assign y1082 = n6272 ;
  assign y1083 = ~n6274 ;
  assign y1084 = n6288 ;
  assign y1085 = ~n6294 ;
  assign y1086 = ~n6295 ;
  assign y1087 = ~n6298 ;
  assign y1088 = n6316 ;
  assign y1089 = n6317 ;
  assign y1090 = ~n6318 ;
  assign y1091 = ~n6321 ;
  assign y1092 = n6332 ;
  assign y1093 = n6339 ;
  assign y1094 = n6346 ;
  assign y1095 = ~n6348 ;
  assign y1096 = n6352 ;
  assign y1097 = n6364 ;
  assign y1098 = ~1'b0 ;
  assign y1099 = ~n6375 ;
  assign y1100 = n6377 ;
  assign y1101 = n6380 ;
  assign y1102 = ~1'b0 ;
  assign y1103 = ~n6387 ;
  assign y1104 = n6392 ;
  assign y1105 = ~1'b0 ;
  assign y1106 = n6395 ;
  assign y1107 = n6398 ;
  assign y1108 = n6403 ;
  assign y1109 = n6404 ;
  assign y1110 = ~n6408 ;
  assign y1111 = n6410 ;
  assign y1112 = ~n6420 ;
  assign y1113 = ~n6424 ;
  assign y1114 = n6431 ;
  assign y1115 = ~n6432 ;
  assign y1116 = n6442 ;
  assign y1117 = n6444 ;
  assign y1118 = n6457 ;
  assign y1119 = ~n6462 ;
  assign y1120 = n6463 ;
  assign y1121 = n6468 ;
  assign y1122 = n6474 ;
  assign y1123 = n6476 ;
  assign y1124 = n6477 ;
  assign y1125 = n6483 ;
  assign y1126 = n6484 ;
  assign y1127 = n6488 ;
  assign y1128 = ~n6494 ;
  assign y1129 = ~n6497 ;
  assign y1130 = n6506 ;
  assign y1131 = ~n6509 ;
  assign y1132 = n6512 ;
  assign y1133 = n6520 ;
  assign y1134 = ~1'b0 ;
  assign y1135 = ~n6524 ;
  assign y1136 = ~n6533 ;
  assign y1137 = ~n6539 ;
  assign y1138 = ~n6543 ;
  assign y1139 = n6544 ;
  assign y1140 = ~n6547 ;
  assign y1141 = ~n6555 ;
  assign y1142 = n6561 ;
  assign y1143 = ~1'b0 ;
  assign y1144 = ~n6563 ;
  assign y1145 = n6564 ;
  assign y1146 = n6565 ;
  assign y1147 = n6578 ;
  assign y1148 = n6593 ;
  assign y1149 = ~n1927 ;
  assign y1150 = n6598 ;
  assign y1151 = ~n6604 ;
  assign y1152 = ~n6606 ;
  assign y1153 = n6610 ;
  assign y1154 = ~n6612 ;
  assign y1155 = ~n6620 ;
  assign y1156 = n6622 ;
  assign y1157 = ~n6628 ;
  assign y1158 = ~1'b0 ;
  assign y1159 = n6632 ;
  assign y1160 = ~n6633 ;
  assign y1161 = n6634 ;
  assign y1162 = ~n6643 ;
  assign y1163 = ~n6647 ;
  assign y1164 = n6652 ;
  assign y1165 = ~n6656 ;
  assign y1166 = n6663 ;
  assign y1167 = ~n6664 ;
  assign y1168 = n6669 ;
  assign y1169 = ~n6673 ;
  assign y1170 = n6674 ;
  assign y1171 = ~n6683 ;
  assign y1172 = ~n6684 ;
  assign y1173 = ~1'b0 ;
  assign y1174 = n6696 ;
  assign y1175 = ~n6702 ;
  assign y1176 = n6708 ;
  assign y1177 = n6718 ;
  assign y1178 = ~n6725 ;
  assign y1179 = n6731 ;
  assign y1180 = n6734 ;
  assign y1181 = ~n6735 ;
  assign y1182 = n6744 ;
  assign y1183 = ~n6757 ;
  assign y1184 = n6759 ;
  assign y1185 = ~n6766 ;
  assign y1186 = n6777 ;
  assign y1187 = ~n6784 ;
  assign y1188 = n6785 ;
  assign y1189 = ~n6786 ;
  assign y1190 = n6790 ;
  assign y1191 = n6795 ;
  assign y1192 = ~1'b0 ;
  assign y1193 = ~n6796 ;
  assign y1194 = ~1'b0 ;
  assign y1195 = ~n6813 ;
  assign y1196 = n6816 ;
  assign y1197 = n6826 ;
  assign y1198 = n6834 ;
  assign y1199 = ~n6838 ;
  assign y1200 = n6840 ;
  assign y1201 = n6846 ;
  assign y1202 = n6847 ;
  assign y1203 = n6853 ;
  assign y1204 = n6854 ;
  assign y1205 = n6856 ;
  assign y1206 = n6859 ;
  assign y1207 = ~1'b0 ;
  assign y1208 = n6866 ;
  assign y1209 = n6869 ;
  assign y1210 = ~n6882 ;
  assign y1211 = ~1'b0 ;
  assign y1212 = ~n6888 ;
  assign y1213 = ~n6892 ;
  assign y1214 = ~n6893 ;
  assign y1215 = ~1'b0 ;
  assign y1216 = ~n6901 ;
  assign y1217 = ~n6912 ;
  assign y1218 = n6913 ;
  assign y1219 = ~1'b0 ;
  assign y1220 = ~n6923 ;
  assign y1221 = ~n6942 ;
  assign y1222 = ~1'b0 ;
  assign y1223 = ~n6947 ;
  assign y1224 = ~n6952 ;
  assign y1225 = 1'b0 ;
  assign y1226 = n6954 ;
  assign y1227 = n6964 ;
  assign y1228 = ~n6969 ;
  assign y1229 = n6970 ;
  assign y1230 = ~n6975 ;
  assign y1231 = ~n6982 ;
  assign y1232 = ~n6984 ;
  assign y1233 = n6990 ;
  assign y1234 = ~n6993 ;
  assign y1235 = ~n6994 ;
  assign y1236 = n6998 ;
  assign y1237 = ~n7005 ;
  assign y1238 = n7014 ;
  assign y1239 = ~1'b0 ;
  assign y1240 = n7017 ;
  assign y1241 = n7019 ;
  assign y1242 = n7026 ;
  assign y1243 = ~n7033 ;
  assign y1244 = ~1'b0 ;
  assign y1245 = ~n7036 ;
  assign y1246 = n7038 ;
  assign y1247 = ~n7043 ;
  assign y1248 = n7046 ;
  assign y1249 = ~n7053 ;
  assign y1250 = n7055 ;
  assign y1251 = n7058 ;
  assign y1252 = n7063 ;
  assign y1253 = ~n7078 ;
  assign y1254 = ~n7082 ;
  assign y1255 = n7085 ;
  assign y1256 = ~n7087 ;
  assign y1257 = ~n7088 ;
  assign y1258 = n7092 ;
  assign y1259 = ~n7094 ;
  assign y1260 = ~n7099 ;
  assign y1261 = n7100 ;
  assign y1262 = n7102 ;
  assign y1263 = ~n7110 ;
  assign y1264 = n7122 ;
  assign y1265 = n7127 ;
  assign y1266 = n7139 ;
  assign y1267 = ~1'b0 ;
  assign y1268 = ~n7141 ;
  assign y1269 = ~n7152 ;
  assign y1270 = ~n7160 ;
  assign y1271 = n7163 ;
  assign y1272 = ~n7165 ;
  assign y1273 = n7167 ;
  assign y1274 = ~n7169 ;
  assign y1275 = n7172 ;
  assign y1276 = n7189 ;
  assign y1277 = n7194 ;
  assign y1278 = ~n7202 ;
  assign y1279 = ~n7206 ;
  assign y1280 = n7209 ;
  assign y1281 = n7211 ;
  assign y1282 = ~n7213 ;
  assign y1283 = ~n7235 ;
  assign y1284 = n7240 ;
  assign y1285 = ~n7244 ;
  assign y1286 = n7250 ;
  assign y1287 = ~n7259 ;
  assign y1288 = ~n7263 ;
  assign y1289 = ~n7279 ;
  assign y1290 = ~n7280 ;
  assign y1291 = ~n7283 ;
  assign y1292 = ~n7289 ;
  assign y1293 = n7292 ;
  assign y1294 = ~n7304 ;
  assign y1295 = ~n7313 ;
  assign y1296 = ~1'b0 ;
  assign y1297 = ~n7319 ;
  assign y1298 = ~1'b0 ;
  assign y1299 = ~n7321 ;
  assign y1300 = ~n7339 ;
  assign y1301 = ~n7346 ;
  assign y1302 = ~n7350 ;
  assign y1303 = ~n7356 ;
  assign y1304 = n7357 ;
  assign y1305 = ~1'b0 ;
  assign y1306 = n7358 ;
  assign y1307 = n7360 ;
  assign y1308 = ~n7362 ;
  assign y1309 = ~n7363 ;
  assign y1310 = n7368 ;
  assign y1311 = ~n7375 ;
  assign y1312 = ~n7377 ;
  assign y1313 = ~n7379 ;
  assign y1314 = n7391 ;
  assign y1315 = ~n7392 ;
  assign y1316 = ~n7400 ;
  assign y1317 = ~n7402 ;
  assign y1318 = n7412 ;
  assign y1319 = ~n7423 ;
  assign y1320 = ~n7435 ;
  assign y1321 = n7440 ;
  assign y1322 = ~n7441 ;
  assign y1323 = ~n7448 ;
  assign y1324 = n7454 ;
  assign y1325 = n7455 ;
  assign y1326 = ~1'b0 ;
  assign y1327 = n7473 ;
  assign y1328 = ~n7484 ;
  assign y1329 = ~n7486 ;
  assign y1330 = ~n7492 ;
  assign y1331 = ~n7495 ;
  assign y1332 = n7501 ;
  assign y1333 = n7502 ;
  assign y1334 = n7504 ;
  assign y1335 = ~n7505 ;
  assign y1336 = ~n7517 ;
  assign y1337 = ~n7520 ;
  assign y1338 = ~n7522 ;
  assign y1339 = n7524 ;
  assign y1340 = n7530 ;
  assign y1341 = ~n7535 ;
  assign y1342 = n7539 ;
  assign y1343 = ~n7550 ;
  assign y1344 = ~n7553 ;
  assign y1345 = n7568 ;
  assign y1346 = ~n7570 ;
  assign y1347 = ~n7584 ;
  assign y1348 = ~n7591 ;
  assign y1349 = n7593 ;
  assign y1350 = ~n7595 ;
  assign y1351 = ~n7602 ;
  assign y1352 = n7606 ;
  assign y1353 = ~n7611 ;
  assign y1354 = n7614 ;
  assign y1355 = ~n7625 ;
  assign y1356 = n7628 ;
  assign y1357 = ~n7629 ;
  assign y1358 = ~n7633 ;
  assign y1359 = n7648 ;
  assign y1360 = ~n7652 ;
  assign y1361 = n7658 ;
  assign y1362 = ~n7663 ;
  assign y1363 = ~n7664 ;
  assign y1364 = n7667 ;
  assign y1365 = n7670 ;
  assign y1366 = ~n7672 ;
  assign y1367 = n7673 ;
  assign y1368 = ~1'b0 ;
  assign y1369 = ~1'b0 ;
  assign y1370 = ~n7681 ;
  assign y1371 = n7684 ;
  assign y1372 = ~n7696 ;
  assign y1373 = ~n7700 ;
  assign y1374 = ~n7702 ;
  assign y1375 = ~n7703 ;
  assign y1376 = n7707 ;
  assign y1377 = ~n7712 ;
  assign y1378 = ~n7719 ;
  assign y1379 = n7722 ;
  assign y1380 = n7725 ;
  assign y1381 = n7732 ;
  assign y1382 = n7740 ;
  assign y1383 = n7743 ;
  assign y1384 = ~n7749 ;
  assign y1385 = n7750 ;
  assign y1386 = ~n7751 ;
  assign y1387 = n7764 ;
  assign y1388 = n7765 ;
  assign y1389 = ~1'b0 ;
  assign y1390 = ~n7767 ;
  assign y1391 = ~n7768 ;
  assign y1392 = ~n7774 ;
  assign y1393 = ~n7777 ;
  assign y1394 = ~1'b0 ;
  assign y1395 = ~1'b0 ;
  assign y1396 = n7783 ;
  assign y1397 = n7793 ;
  assign y1398 = ~n7800 ;
  assign y1399 = n7803 ;
  assign y1400 = ~n7805 ;
  assign y1401 = n7808 ;
  assign y1402 = ~n7815 ;
  assign y1403 = ~n7818 ;
  assign y1404 = ~n7823 ;
  assign y1405 = n7825 ;
  assign y1406 = n7834 ;
  assign y1407 = ~n7835 ;
  assign y1408 = ~n7836 ;
  assign y1409 = ~n7841 ;
  assign y1410 = ~n7844 ;
  assign y1411 = ~n7854 ;
  assign y1412 = ~n7861 ;
  assign y1413 = n7872 ;
  assign y1414 = ~n7879 ;
  assign y1415 = n7882 ;
  assign y1416 = ~n7892 ;
  assign y1417 = n7902 ;
  assign y1418 = n7907 ;
  assign y1419 = ~n7913 ;
  assign y1420 = n7921 ;
  assign y1421 = ~n7930 ;
  assign y1422 = ~n7935 ;
  assign y1423 = ~n7940 ;
  assign y1424 = n7945 ;
  assign y1425 = ~n7948 ;
  assign y1426 = n7954 ;
  assign y1427 = ~n7970 ;
  assign y1428 = ~n7978 ;
  assign y1429 = ~n7983 ;
  assign y1430 = ~n7989 ;
  assign y1431 = ~n7992 ;
  assign y1432 = n7997 ;
  assign y1433 = ~n8005 ;
  assign y1434 = n8007 ;
  assign y1435 = n8011 ;
  assign y1436 = n8013 ;
  assign y1437 = n8020 ;
  assign y1438 = n8025 ;
  assign y1439 = ~1'b0 ;
  assign y1440 = n8028 ;
  assign y1441 = ~n8045 ;
  assign y1442 = ~1'b0 ;
  assign y1443 = n8053 ;
  assign y1444 = n8061 ;
  assign y1445 = ~n8064 ;
  assign y1446 = n8068 ;
  assign y1447 = n8076 ;
  assign y1448 = ~n8079 ;
  assign y1449 = ~1'b0 ;
  assign y1450 = ~n8089 ;
  assign y1451 = ~n8090 ;
  assign y1452 = ~n8101 ;
  assign y1453 = ~n8102 ;
  assign y1454 = ~n8110 ;
  assign y1455 = n8111 ;
  assign y1456 = n8112 ;
  assign y1457 = n8115 ;
  assign y1458 = n8117 ;
  assign y1459 = ~n8150 ;
  assign y1460 = ~n8160 ;
  assign y1461 = ~n8163 ;
  assign y1462 = ~n8170 ;
  assign y1463 = n8171 ;
  assign y1464 = ~n8180 ;
  assign y1465 = ~n8181 ;
  assign y1466 = n8183 ;
  assign y1467 = n8191 ;
  assign y1468 = ~1'b0 ;
  assign y1469 = n8193 ;
  assign y1470 = n8196 ;
  assign y1471 = ~n8200 ;
  assign y1472 = ~n8203 ;
  assign y1473 = n8209 ;
  assign y1474 = ~n8216 ;
  assign y1475 = n8221 ;
  assign y1476 = ~n8226 ;
  assign y1477 = ~n8229 ;
  assign y1478 = n8241 ;
  assign y1479 = ~1'b0 ;
  assign y1480 = n8244 ;
  assign y1481 = ~n8245 ;
  assign y1482 = ~n8257 ;
  assign y1483 = n8258 ;
  assign y1484 = n8263 ;
  assign y1485 = n8266 ;
  assign y1486 = ~n8272 ;
  assign y1487 = ~n8274 ;
  assign y1488 = n8276 ;
  assign y1489 = ~n8280 ;
  assign y1490 = n8281 ;
  assign y1491 = n8283 ;
  assign y1492 = ~n8289 ;
  assign y1493 = ~n8290 ;
  assign y1494 = n8291 ;
  assign y1495 = n8299 ;
  assign y1496 = ~n8303 ;
  assign y1497 = ~n8304 ;
  assign y1498 = n8306 ;
  assign y1499 = ~n8312 ;
  assign y1500 = n8315 ;
  assign y1501 = ~n8327 ;
  assign y1502 = n8331 ;
  assign y1503 = ~n8347 ;
  assign y1504 = ~1'b0 ;
  assign y1505 = ~n8353 ;
  assign y1506 = n8366 ;
  assign y1507 = n8369 ;
  assign y1508 = ~n8378 ;
  assign y1509 = ~n8387 ;
  assign y1510 = n8390 ;
  assign y1511 = n8396 ;
  assign y1512 = n8408 ;
  assign y1513 = ~n8413 ;
  assign y1514 = n8421 ;
  assign y1515 = ~1'b0 ;
  assign y1516 = ~n8425 ;
  assign y1517 = ~1'b0 ;
  assign y1518 = n8426 ;
  assign y1519 = ~n8432 ;
  assign y1520 = n8436 ;
  assign y1521 = n8442 ;
  assign y1522 = ~1'b0 ;
  assign y1523 = ~n8443 ;
  assign y1524 = ~n8445 ;
  assign y1525 = ~n8450 ;
  assign y1526 = n8456 ;
  assign y1527 = ~n8458 ;
  assign y1528 = ~n8459 ;
  assign y1529 = ~1'b0 ;
  assign y1530 = n8472 ;
  assign y1531 = ~n8473 ;
  assign y1532 = n8476 ;
  assign y1533 = ~n8477 ;
  assign y1534 = n8486 ;
  assign y1535 = n8487 ;
  assign y1536 = n8490 ;
  assign y1537 = n8493 ;
  assign y1538 = n8494 ;
  assign y1539 = ~n8498 ;
  assign y1540 = ~n8501 ;
  assign y1541 = n8505 ;
  assign y1542 = n8515 ;
  assign y1543 = ~n8520 ;
  assign y1544 = ~n8521 ;
  assign y1545 = ~n8529 ;
  assign y1546 = ~n8536 ;
  assign y1547 = ~n8548 ;
  assign y1548 = ~n8549 ;
  assign y1549 = ~n8552 ;
  assign y1550 = ~1'b0 ;
  assign y1551 = ~1'b0 ;
  assign y1552 = n8561 ;
  assign y1553 = ~n8564 ;
  assign y1554 = ~n8566 ;
  assign y1555 = ~n8572 ;
  assign y1556 = n8573 ;
  assign y1557 = n8575 ;
  assign y1558 = ~n8576 ;
  assign y1559 = ~1'b0 ;
  assign y1560 = ~n8579 ;
  assign y1561 = ~n8581 ;
  assign y1562 = n8583 ;
  assign y1563 = ~n8585 ;
  assign y1564 = ~n8586 ;
  assign y1565 = ~n8587 ;
  assign y1566 = ~n8595 ;
  assign y1567 = ~n8601 ;
  assign y1568 = ~n8602 ;
  assign y1569 = ~n8608 ;
  assign y1570 = ~n8614 ;
  assign y1571 = ~n8617 ;
  assign y1572 = ~1'b0 ;
  assign y1573 = n8622 ;
  assign y1574 = ~n8625 ;
  assign y1575 = ~n8631 ;
  assign y1576 = n8633 ;
  assign y1577 = n8636 ;
  assign y1578 = ~n8642 ;
  assign y1579 = ~n8645 ;
  assign y1580 = ~n8655 ;
  assign y1581 = ~n8656 ;
  assign y1582 = ~n8660 ;
  assign y1583 = ~n8661 ;
  assign y1584 = n8671 ;
  assign y1585 = n8681 ;
  assign y1586 = n8686 ;
  assign y1587 = n8707 ;
  assign y1588 = n8714 ;
  assign y1589 = n8719 ;
  assign y1590 = n8727 ;
  assign y1591 = n8735 ;
  assign y1592 = ~n8739 ;
  assign y1593 = n8744 ;
  assign y1594 = n8747 ;
  assign y1595 = n8748 ;
  assign y1596 = ~1'b0 ;
  assign y1597 = ~n8749 ;
  assign y1598 = n8753 ;
  assign y1599 = ~1'b0 ;
  assign y1600 = n8754 ;
  assign y1601 = ~n8760 ;
  assign y1602 = n8767 ;
  assign y1603 = n8768 ;
  assign y1604 = n8771 ;
  assign y1605 = ~n8783 ;
  assign y1606 = n8790 ;
  assign y1607 = ~n8794 ;
  assign y1608 = n8800 ;
  assign y1609 = ~1'b0 ;
  assign y1610 = n8805 ;
  assign y1611 = ~n8807 ;
  assign y1612 = n8808 ;
  assign y1613 = n8813 ;
  assign y1614 = ~n8814 ;
  assign y1615 = n8815 ;
  assign y1616 = n8819 ;
  assign y1617 = n8824 ;
  assign y1618 = n8825 ;
  assign y1619 = ~n8826 ;
  assign y1620 = ~n8829 ;
  assign y1621 = ~n8831 ;
  assign y1622 = n8842 ;
  assign y1623 = n8851 ;
  assign y1624 = ~n8855 ;
  assign y1625 = n8859 ;
  assign y1626 = ~n8865 ;
  assign y1627 = ~n8867 ;
  assign y1628 = n8872 ;
  assign y1629 = n8873 ;
  assign y1630 = n8876 ;
  assign y1631 = ~n8877 ;
  assign y1632 = ~n8891 ;
  assign y1633 = ~n8901 ;
  assign y1634 = ~n8908 ;
  assign y1635 = ~n8912 ;
  assign y1636 = ~n8914 ;
  assign y1637 = ~n8915 ;
  assign y1638 = ~n8918 ;
  assign y1639 = n8919 ;
  assign y1640 = n8929 ;
  assign y1641 = n8933 ;
  assign y1642 = n8934 ;
  assign y1643 = n8936 ;
  assign y1644 = n8943 ;
  assign y1645 = ~n8945 ;
  assign y1646 = ~n8951 ;
  assign y1647 = ~n8952 ;
  assign y1648 = ~n8955 ;
  assign y1649 = n8968 ;
  assign y1650 = ~n8971 ;
  assign y1651 = n8979 ;
  assign y1652 = ~1'b0 ;
  assign y1653 = ~n8980 ;
  assign y1654 = n8989 ;
  assign y1655 = ~n8990 ;
  assign y1656 = ~n8994 ;
  assign y1657 = n8999 ;
  assign y1658 = ~n9013 ;
  assign y1659 = ~n9016 ;
  assign y1660 = n9019 ;
  assign y1661 = n9027 ;
  assign y1662 = ~n9029 ;
  assign y1663 = ~n9034 ;
  assign y1664 = n9040 ;
  assign y1665 = ~n9041 ;
  assign y1666 = n9049 ;
  assign y1667 = ~n9060 ;
  assign y1668 = n9065 ;
  assign y1669 = ~n9069 ;
  assign y1670 = ~n9070 ;
  assign y1671 = ~n9076 ;
  assign y1672 = ~n9086 ;
  assign y1673 = n9089 ;
  assign y1674 = ~n9096 ;
  assign y1675 = ~n9101 ;
  assign y1676 = ~n9103 ;
  assign y1677 = n9108 ;
  assign y1678 = ~n9110 ;
  assign y1679 = ~n9112 ;
  assign y1680 = ~n9116 ;
  assign y1681 = n9126 ;
  assign y1682 = n9142 ;
  assign y1683 = ~n9143 ;
  assign y1684 = ~n9147 ;
  assign y1685 = ~n9150 ;
  assign y1686 = n9152 ;
  assign y1687 = n9160 ;
  assign y1688 = n9161 ;
  assign y1689 = n9165 ;
  assign y1690 = ~n9168 ;
  assign y1691 = n9173 ;
  assign y1692 = n9182 ;
  assign y1693 = n9193 ;
  assign y1694 = n9208 ;
  assign y1695 = ~n9209 ;
  assign y1696 = ~n9213 ;
  assign y1697 = n9214 ;
  assign y1698 = ~n9220 ;
  assign y1699 = ~n9230 ;
  assign y1700 = ~n9233 ;
  assign y1701 = ~n9234 ;
  assign y1702 = ~n9238 ;
  assign y1703 = n9239 ;
  assign y1704 = n9240 ;
  assign y1705 = n9245 ;
  assign y1706 = ~n9250 ;
  assign y1707 = n9264 ;
  assign y1708 = ~n9268 ;
  assign y1709 = n4513 ;
  assign y1710 = ~n9274 ;
  assign y1711 = ~n9281 ;
  assign y1712 = n9282 ;
  assign y1713 = ~n9283 ;
  assign y1714 = ~n9284 ;
  assign y1715 = ~n9290 ;
  assign y1716 = n9294 ;
  assign y1717 = ~n9305 ;
  assign y1718 = ~n9323 ;
  assign y1719 = ~n9339 ;
  assign y1720 = ~n9343 ;
  assign y1721 = ~n9350 ;
  assign y1722 = n9357 ;
  assign y1723 = ~n9360 ;
  assign y1724 = ~n9361 ;
  assign y1725 = ~n9363 ;
  assign y1726 = ~n9367 ;
  assign y1727 = n9370 ;
  assign y1728 = ~n9376 ;
  assign y1729 = n9380 ;
  assign y1730 = ~1'b0 ;
  assign y1731 = ~n9385 ;
  assign y1732 = n9386 ;
  assign y1733 = n9388 ;
  assign y1734 = n9389 ;
  assign y1735 = n9394 ;
  assign y1736 = n9404 ;
  assign y1737 = n9406 ;
  assign y1738 = n9411 ;
  assign y1739 = n9420 ;
  assign y1740 = n9429 ;
  assign y1741 = n9440 ;
  assign y1742 = ~n9452 ;
  assign y1743 = ~n9461 ;
  assign y1744 = ~n9464 ;
  assign y1745 = ~n9465 ;
  assign y1746 = n9474 ;
  assign y1747 = ~n9477 ;
  assign y1748 = ~n9481 ;
  assign y1749 = ~n9486 ;
  assign y1750 = n9493 ;
  assign y1751 = ~1'b0 ;
  assign y1752 = ~n9494 ;
  assign y1753 = n9500 ;
  assign y1754 = n9502 ;
  assign y1755 = ~n9504 ;
  assign y1756 = n9507 ;
  assign y1757 = n9513 ;
  assign y1758 = n9515 ;
  assign y1759 = ~1'b0 ;
  assign y1760 = n9521 ;
  assign y1761 = ~n9523 ;
  assign y1762 = n9528 ;
  assign y1763 = n9539 ;
  assign y1764 = ~n9550 ;
  assign y1765 = ~1'b0 ;
  assign y1766 = ~n9557 ;
  assign y1767 = n9566 ;
  assign y1768 = ~n9570 ;
  assign y1769 = ~1'b0 ;
  assign y1770 = ~n9571 ;
  assign y1771 = n9573 ;
  assign y1772 = ~n9578 ;
  assign y1773 = n9583 ;
  assign y1774 = ~n9589 ;
  assign y1775 = n9592 ;
  assign y1776 = ~n9598 ;
  assign y1777 = ~n9600 ;
  assign y1778 = ~n9605 ;
  assign y1779 = n9607 ;
  assign y1780 = ~n9615 ;
  assign y1781 = ~n9616 ;
  assign y1782 = n9623 ;
  assign y1783 = n9625 ;
  assign y1784 = ~1'b0 ;
  assign y1785 = n9628 ;
  assign y1786 = n9631 ;
  assign y1787 = n9634 ;
  assign y1788 = ~1'b0 ;
  assign y1789 = ~1'b0 ;
  assign y1790 = n9643 ;
  assign y1791 = ~n9645 ;
  assign y1792 = ~n9647 ;
  assign y1793 = ~n9655 ;
  assign y1794 = n9661 ;
  assign y1795 = ~n9674 ;
  assign y1796 = ~1'b0 ;
  assign y1797 = ~n9684 ;
  assign y1798 = ~n9689 ;
  assign y1799 = n9690 ;
  assign y1800 = n9693 ;
  assign y1801 = n9696 ;
  assign y1802 = n9698 ;
  assign y1803 = ~n9704 ;
  assign y1804 = ~n9710 ;
  assign y1805 = n9728 ;
  assign y1806 = n9740 ;
  assign y1807 = n9746 ;
  assign y1808 = ~n9748 ;
  assign y1809 = ~n9761 ;
  assign y1810 = ~n9764 ;
  assign y1811 = n9780 ;
  assign y1812 = n9784 ;
  assign y1813 = ~n9786 ;
  assign y1814 = ~n9789 ;
  assign y1815 = ~n9791 ;
  assign y1816 = n9795 ;
  assign y1817 = n9798 ;
  assign y1818 = ~n9800 ;
  assign y1819 = ~n9802 ;
  assign y1820 = n9805 ;
  assign y1821 = ~1'b0 ;
  assign y1822 = n9809 ;
  assign y1823 = n9820 ;
  assign y1824 = ~n9826 ;
  assign y1825 = ~n9830 ;
  assign y1826 = ~n9833 ;
  assign y1827 = n9838 ;
  assign y1828 = n9842 ;
  assign y1829 = ~n9843 ;
  assign y1830 = ~1'b0 ;
  assign y1831 = n9844 ;
  assign y1832 = n9849 ;
  assign y1833 = ~n9853 ;
  assign y1834 = n9857 ;
  assign y1835 = ~n9858 ;
  assign y1836 = ~n9867 ;
  assign y1837 = ~n9870 ;
  assign y1838 = ~1'b0 ;
  assign y1839 = ~1'b0 ;
  assign y1840 = ~n9873 ;
  assign y1841 = n9874 ;
  assign y1842 = n9877 ;
  assign y1843 = ~n9886 ;
  assign y1844 = n9888 ;
  assign y1845 = n9890 ;
  assign y1846 = ~n9899 ;
  assign y1847 = n9900 ;
  assign y1848 = n9904 ;
  assign y1849 = ~n9909 ;
  assign y1850 = n9910 ;
  assign y1851 = n9914 ;
  assign y1852 = ~n9924 ;
  assign y1853 = n9949 ;
  assign y1854 = n9950 ;
  assign y1855 = ~n9953 ;
  assign y1856 = ~n6360 ;
  assign y1857 = n9954 ;
  assign y1858 = n9956 ;
  assign y1859 = n9970 ;
  assign y1860 = ~n9978 ;
  assign y1861 = n9983 ;
  assign y1862 = ~n9991 ;
  assign y1863 = n9993 ;
  assign y1864 = ~n10005 ;
  assign y1865 = ~n10006 ;
  assign y1866 = n10007 ;
  assign y1867 = ~n10014 ;
  assign y1868 = n10015 ;
  assign y1869 = ~n10018 ;
  assign y1870 = n10020 ;
  assign y1871 = ~1'b0 ;
  assign y1872 = ~n10021 ;
  assign y1873 = ~n10022 ;
  assign y1874 = ~n10023 ;
  assign y1875 = n10032 ;
  assign y1876 = ~1'b0 ;
  assign y1877 = ~n10034 ;
  assign y1878 = n10037 ;
  assign y1879 = ~n10038 ;
  assign y1880 = n10044 ;
  assign y1881 = n10050 ;
  assign y1882 = ~n10056 ;
  assign y1883 = ~n10061 ;
  assign y1884 = n10069 ;
  assign y1885 = ~n10070 ;
  assign y1886 = ~n10072 ;
  assign y1887 = ~n10076 ;
  assign y1888 = ~n10080 ;
  assign y1889 = ~n10087 ;
  assign y1890 = ~n10088 ;
  assign y1891 = ~n10094 ;
  assign y1892 = ~n10103 ;
  assign y1893 = ~n10107 ;
  assign y1894 = n10110 ;
  assign y1895 = n10113 ;
  assign y1896 = ~n10132 ;
  assign y1897 = ~n10135 ;
  assign y1898 = ~n10139 ;
  assign y1899 = ~n10141 ;
  assign y1900 = ~n10144 ;
  assign y1901 = ~n10156 ;
  assign y1902 = n10163 ;
  assign y1903 = ~n10168 ;
  assign y1904 = ~n10169 ;
  assign y1905 = ~n10174 ;
  assign y1906 = ~n10175 ;
  assign y1907 = ~n10180 ;
  assign y1908 = ~n10184 ;
  assign y1909 = ~n10193 ;
  assign y1910 = ~n10194 ;
  assign y1911 = ~n10196 ;
  assign y1912 = ~n10200 ;
  assign y1913 = n10203 ;
  assign y1914 = ~n10212 ;
  assign y1915 = ~n10214 ;
  assign y1916 = n10222 ;
  assign y1917 = ~1'b0 ;
  assign y1918 = ~n10228 ;
  assign y1919 = ~n10236 ;
  assign y1920 = ~n10244 ;
  assign y1921 = ~n10246 ;
  assign y1922 = ~1'b0 ;
  assign y1923 = n10255 ;
  assign y1924 = n10257 ;
  assign y1925 = n10258 ;
  assign y1926 = ~n10267 ;
  assign y1927 = n10271 ;
  assign y1928 = ~n10275 ;
  assign y1929 = n10277 ;
  assign y1930 = ~n10281 ;
  assign y1931 = n10285 ;
  assign y1932 = n10286 ;
  assign y1933 = ~1'b0 ;
  assign y1934 = ~n10297 ;
  assign y1935 = ~1'b0 ;
  assign y1936 = n10302 ;
  assign y1937 = n10304 ;
  assign y1938 = n10306 ;
  assign y1939 = ~n10308 ;
  assign y1940 = ~1'b0 ;
  assign y1941 = ~n10310 ;
  assign y1942 = n10321 ;
  assign y1943 = ~n10323 ;
  assign y1944 = ~n10325 ;
  assign y1945 = n10336 ;
  assign y1946 = n10341 ;
  assign y1947 = ~n10345 ;
  assign y1948 = ~n10349 ;
  assign y1949 = n10353 ;
  assign y1950 = n10356 ;
  assign y1951 = ~n10357 ;
  assign y1952 = n10360 ;
  assign y1953 = ~n10364 ;
  assign y1954 = n10367 ;
  assign y1955 = ~n10369 ;
  assign y1956 = n10372 ;
  assign y1957 = ~n10384 ;
  assign y1958 = ~n10387 ;
  assign y1959 = ~1'b0 ;
  assign y1960 = ~n10403 ;
  assign y1961 = ~n10405 ;
  assign y1962 = ~n10408 ;
  assign y1963 = n10413 ;
  assign y1964 = ~n10425 ;
  assign y1965 = n10431 ;
  assign y1966 = ~n10433 ;
  assign y1967 = ~n10436 ;
  assign y1968 = ~n10440 ;
  assign y1969 = n10445 ;
  assign y1970 = ~n10447 ;
  assign y1971 = n10448 ;
  assign y1972 = ~n10450 ;
  assign y1973 = ~n8642 ;
  assign y1974 = n10455 ;
  assign y1975 = ~n10457 ;
  assign y1976 = n10460 ;
  assign y1977 = n10461 ;
  assign y1978 = ~1'b0 ;
  assign y1979 = n10469 ;
  assign y1980 = n10470 ;
  assign y1981 = ~1'b0 ;
  assign y1982 = ~n10474 ;
  assign y1983 = ~n10478 ;
  assign y1984 = ~1'b0 ;
  assign y1985 = ~n10480 ;
  assign y1986 = ~n10487 ;
  assign y1987 = ~n10497 ;
  assign y1988 = ~n10500 ;
  assign y1989 = ~n10501 ;
  assign y1990 = ~n10509 ;
  assign y1991 = n10510 ;
  assign y1992 = n10525 ;
  assign y1993 = n10530 ;
  assign y1994 = n10531 ;
  assign y1995 = ~1'b0 ;
  assign y1996 = ~n10537 ;
  assign y1997 = ~1'b0 ;
  assign y1998 = n10538 ;
  assign y1999 = ~n10539 ;
  assign y2000 = ~n10545 ;
  assign y2001 = ~n10548 ;
  assign y2002 = ~1'b0 ;
  assign y2003 = n10555 ;
  assign y2004 = ~n10561 ;
  assign y2005 = n10567 ;
  assign y2006 = n10582 ;
  assign y2007 = n10585 ;
  assign y2008 = n10592 ;
  assign y2009 = ~n10600 ;
  assign y2010 = ~n10602 ;
  assign y2011 = n10608 ;
  assign y2012 = ~n10617 ;
  assign y2013 = n10619 ;
  assign y2014 = ~n10624 ;
  assign y2015 = ~n10631 ;
  assign y2016 = n10637 ;
  assign y2017 = n10642 ;
  assign y2018 = ~n10648 ;
  assign y2019 = ~n10659 ;
  assign y2020 = n10663 ;
  assign y2021 = n10666 ;
  assign y2022 = ~n10673 ;
  assign y2023 = n10678 ;
  assign y2024 = n10679 ;
  assign y2025 = n10689 ;
  assign y2026 = n10690 ;
  assign y2027 = n10697 ;
  assign y2028 = ~n10698 ;
  assign y2029 = ~n10707 ;
  assign y2030 = ~n10716 ;
  assign y2031 = ~n10717 ;
  assign y2032 = ~n10723 ;
  assign y2033 = ~n10724 ;
  assign y2034 = ~n10726 ;
  assign y2035 = ~n10732 ;
  assign y2036 = ~n10739 ;
  assign y2037 = n10745 ;
  assign y2038 = ~n10751 ;
  assign y2039 = ~n10754 ;
  assign y2040 = ~n10756 ;
  assign y2041 = n10763 ;
  assign y2042 = n10767 ;
  assign y2043 = ~n10768 ;
  assign y2044 = ~n10775 ;
  assign y2045 = n10784 ;
  assign y2046 = n10789 ;
  assign y2047 = ~1'b0 ;
  assign y2048 = ~n10801 ;
  assign y2049 = n10805 ;
  assign y2050 = ~n10806 ;
  assign y2051 = n10807 ;
  assign y2052 = n10812 ;
  assign y2053 = n10813 ;
  assign y2054 = ~n10822 ;
  assign y2055 = n10824 ;
  assign y2056 = n10835 ;
  assign y2057 = n10836 ;
  assign y2058 = ~n10847 ;
  assign y2059 = n10851 ;
  assign y2060 = n10853 ;
  assign y2061 = ~n10855 ;
  assign y2062 = ~n10857 ;
  assign y2063 = ~n10862 ;
  assign y2064 = ~n10865 ;
  assign y2065 = ~n10870 ;
  assign y2066 = n10874 ;
  assign y2067 = n10879 ;
  assign y2068 = ~n10882 ;
  assign y2069 = ~n10890 ;
  assign y2070 = n10893 ;
  assign y2071 = ~n10896 ;
  assign y2072 = ~n10897 ;
  assign y2073 = n10898 ;
  assign y2074 = ~n10902 ;
  assign y2075 = ~n10918 ;
  assign y2076 = ~n10921 ;
  assign y2077 = n10924 ;
  assign y2078 = ~n10925 ;
  assign y2079 = ~n10926 ;
  assign y2080 = ~n10930 ;
  assign y2081 = ~n10932 ;
  assign y2082 = n10940 ;
  assign y2083 = n10943 ;
  assign y2084 = n10949 ;
  assign y2085 = ~n10954 ;
  assign y2086 = ~n10956 ;
  assign y2087 = n10965 ;
  assign y2088 = ~n10967 ;
  assign y2089 = n10975 ;
  assign y2090 = n10978 ;
  assign y2091 = n10988 ;
  assign y2092 = ~n10991 ;
  assign y2093 = ~n10994 ;
  assign y2094 = ~n10995 ;
  assign y2095 = ~n10997 ;
  assign y2096 = ~n11008 ;
  assign y2097 = n11009 ;
  assign y2098 = ~1'b0 ;
  assign y2099 = n11014 ;
  assign y2100 = ~n11017 ;
  assign y2101 = ~n11025 ;
  assign y2102 = n11026 ;
  assign y2103 = ~n11027 ;
  assign y2104 = n11028 ;
  assign y2105 = ~n11040 ;
  assign y2106 = n11044 ;
  assign y2107 = ~n11050 ;
  assign y2108 = ~n11051 ;
  assign y2109 = ~n11053 ;
  assign y2110 = ~n11061 ;
  assign y2111 = ~n11062 ;
  assign y2112 = n2047 ;
  assign y2113 = ~n11065 ;
  assign y2114 = ~n11069 ;
  assign y2115 = n11072 ;
  assign y2116 = ~n11082 ;
  assign y2117 = ~n11086 ;
  assign y2118 = n11089 ;
  assign y2119 = ~1'b0 ;
  assign y2120 = n11091 ;
  assign y2121 = ~n11095 ;
  assign y2122 = ~1'b0 ;
  assign y2123 = ~n11097 ;
  assign y2124 = n11098 ;
  assign y2125 = ~1'b0 ;
  assign y2126 = n11102 ;
  assign y2127 = n11104 ;
  assign y2128 = ~n11111 ;
  assign y2129 = n11118 ;
  assign y2130 = ~n11135 ;
  assign y2131 = ~n11142 ;
  assign y2132 = n11146 ;
  assign y2133 = n11151 ;
  assign y2134 = n11154 ;
  assign y2135 = ~1'b0 ;
  assign y2136 = ~n11167 ;
  assign y2137 = ~n11171 ;
  assign y2138 = ~n11177 ;
  assign y2139 = ~n11184 ;
  assign y2140 = ~n11187 ;
  assign y2141 = ~n11192 ;
  assign y2142 = n11196 ;
  assign y2143 = ~n11203 ;
  assign y2144 = ~n11205 ;
  assign y2145 = ~n11206 ;
  assign y2146 = ~n2224 ;
  assign y2147 = n11208 ;
  assign y2148 = ~n11210 ;
  assign y2149 = n11218 ;
  assign y2150 = ~n11221 ;
  assign y2151 = ~n11223 ;
  assign y2152 = n11226 ;
  assign y2153 = n11235 ;
  assign y2154 = n11239 ;
  assign y2155 = n11242 ;
  assign y2156 = ~n11253 ;
  assign y2157 = n11256 ;
  assign y2158 = n11257 ;
  assign y2159 = ~n11261 ;
  assign y2160 = ~n11265 ;
  assign y2161 = n11272 ;
  assign y2162 = n11276 ;
  assign y2163 = n11277 ;
  assign y2164 = ~n11282 ;
  assign y2165 = ~n11287 ;
  assign y2166 = ~n11288 ;
  assign y2167 = ~n11295 ;
  assign y2168 = ~n11296 ;
  assign y2169 = ~1'b0 ;
  assign y2170 = n11298 ;
  assign y2171 = n11300 ;
  assign y2172 = ~1'b0 ;
  assign y2173 = ~n11308 ;
  assign y2174 = n11309 ;
  assign y2175 = ~n11310 ;
  assign y2176 = n1008 ;
  assign y2177 = n11313 ;
  assign y2178 = ~n11314 ;
  assign y2179 = ~n11317 ;
  assign y2180 = n11319 ;
  assign y2181 = ~n11323 ;
  assign y2182 = n11329 ;
  assign y2183 = n11336 ;
  assign y2184 = ~n11339 ;
  assign y2185 = ~n11340 ;
  assign y2186 = ~n11346 ;
  assign y2187 = ~n11348 ;
  assign y2188 = n11350 ;
  assign y2189 = ~n11351 ;
  assign y2190 = ~n11358 ;
  assign y2191 = ~n11385 ;
  assign y2192 = n11386 ;
  assign y2193 = ~n11390 ;
  assign y2194 = ~n11392 ;
  assign y2195 = n11393 ;
  assign y2196 = ~n11401 ;
  assign y2197 = ~n11403 ;
  assign y2198 = ~n11406 ;
  assign y2199 = n11408 ;
  assign y2200 = n11412 ;
  assign y2201 = n11421 ;
  assign y2202 = ~n11423 ;
  assign y2203 = ~n11434 ;
  assign y2204 = ~n11443 ;
  assign y2205 = n11449 ;
  assign y2206 = n11453 ;
  assign y2207 = ~n11454 ;
  assign y2208 = n11458 ;
  assign y2209 = n11463 ;
  assign y2210 = n11464 ;
  assign y2211 = ~n11468 ;
  assign y2212 = ~1'b0 ;
  assign y2213 = ~n11472 ;
  assign y2214 = n11476 ;
  assign y2215 = ~n11481 ;
  assign y2216 = n11482 ;
  assign y2217 = n11486 ;
  assign y2218 = ~n11495 ;
  assign y2219 = n11507 ;
  assign y2220 = ~n11512 ;
  assign y2221 = ~1'b0 ;
  assign y2222 = n11517 ;
  assign y2223 = n11521 ;
  assign y2224 = ~1'b0 ;
  assign y2225 = ~n11527 ;
  assign y2226 = ~n11529 ;
  assign y2227 = ~n11531 ;
  assign y2228 = n11537 ;
  assign y2229 = ~n11539 ;
  assign y2230 = n11541 ;
  assign y2231 = n11546 ;
  assign y2232 = ~n11556 ;
  assign y2233 = ~n11560 ;
  assign y2234 = n11574 ;
  assign y2235 = n11579 ;
  assign y2236 = n11580 ;
  assign y2237 = n11581 ;
  assign y2238 = ~n11582 ;
  assign y2239 = n11585 ;
  assign y2240 = ~n11586 ;
  assign y2241 = ~n11588 ;
  assign y2242 = ~n11590 ;
  assign y2243 = ~n11593 ;
  assign y2244 = n11598 ;
  assign y2245 = ~1'b0 ;
  assign y2246 = ~n11599 ;
  assign y2247 = ~1'b0 ;
  assign y2248 = ~n9884 ;
  assign y2249 = ~n11607 ;
  assign y2250 = ~n11608 ;
  assign y2251 = ~n11621 ;
  assign y2252 = ~n11622 ;
  assign y2253 = n11626 ;
  assign y2254 = ~n11635 ;
  assign y2255 = ~n11637 ;
  assign y2256 = ~n11649 ;
  assign y2257 = ~n11659 ;
  assign y2258 = n11665 ;
  assign y2259 = n11668 ;
  assign y2260 = ~n11673 ;
  assign y2261 = ~n11679 ;
  assign y2262 = ~n11683 ;
  assign y2263 = n11687 ;
  assign y2264 = n11689 ;
  assign y2265 = n11693 ;
  assign y2266 = ~n11697 ;
  assign y2267 = n11710 ;
  assign y2268 = n11711 ;
  assign y2269 = n11721 ;
  assign y2270 = n11730 ;
  assign y2271 = ~1'b0 ;
  assign y2272 = n11739 ;
  assign y2273 = n11747 ;
  assign y2274 = n11749 ;
  assign y2275 = ~1'b0 ;
  assign y2276 = ~n11753 ;
  assign y2277 = ~n11762 ;
  assign y2278 = n11763 ;
  assign y2279 = ~n11766 ;
  assign y2280 = ~n11775 ;
  assign y2281 = ~n11777 ;
  assign y2282 = ~n11783 ;
  assign y2283 = n11788 ;
  assign y2284 = n11789 ;
  assign y2285 = ~n11800 ;
  assign y2286 = n11804 ;
  assign y2287 = ~1'b0 ;
  assign y2288 = n11805 ;
  assign y2289 = ~n11812 ;
  assign y2290 = n11816 ;
  assign y2291 = ~n11831 ;
  assign y2292 = ~n11833 ;
  assign y2293 = n11837 ;
  assign y2294 = n11838 ;
  assign y2295 = n11839 ;
  assign y2296 = n11842 ;
  assign y2297 = ~n11847 ;
  assign y2298 = ~n11849 ;
  assign y2299 = ~n11851 ;
  assign y2300 = ~n11854 ;
  assign y2301 = ~n11867 ;
  assign y2302 = n11875 ;
  assign y2303 = n11876 ;
  assign y2304 = ~n11882 ;
  assign y2305 = ~n11887 ;
  assign y2306 = n11888 ;
  assign y2307 = ~n11889 ;
  assign y2308 = n11890 ;
  assign y2309 = n11899 ;
  assign y2310 = n11906 ;
  assign y2311 = ~n11908 ;
  assign y2312 = ~n11913 ;
  assign y2313 = ~n11915 ;
  assign y2314 = ~n11919 ;
  assign y2315 = n11924 ;
  assign y2316 = ~n11931 ;
  assign y2317 = n11934 ;
  assign y2318 = n11942 ;
  assign y2319 = n11947 ;
  assign y2320 = n11950 ;
  assign y2321 = ~1'b0 ;
  assign y2322 = ~n11953 ;
  assign y2323 = n11955 ;
  assign y2324 = n11972 ;
  assign y2325 = ~n11974 ;
  assign y2326 = ~n11977 ;
  assign y2327 = ~n11988 ;
  assign y2328 = n11989 ;
  assign y2329 = n11996 ;
  assign y2330 = n12008 ;
  assign y2331 = ~1'b0 ;
  assign y2332 = ~n12009 ;
  assign y2333 = n12010 ;
  assign y2334 = ~n12014 ;
  assign y2335 = ~n12021 ;
  assign y2336 = n12024 ;
  assign y2337 = n12032 ;
  assign y2338 = ~n12038 ;
  assign y2339 = ~n12041 ;
  assign y2340 = n12042 ;
  assign y2341 = n12043 ;
  assign y2342 = ~n12046 ;
  assign y2343 = n12057 ;
  assign y2344 = n12062 ;
  assign y2345 = n12066 ;
  assign y2346 = n12069 ;
  assign y2347 = n12071 ;
  assign y2348 = ~n12072 ;
  assign y2349 = ~1'b0 ;
  assign y2350 = ~n12073 ;
  assign y2351 = ~n12077 ;
  assign y2352 = n12090 ;
  assign y2353 = ~n12097 ;
  assign y2354 = n12100 ;
  assign y2355 = n12104 ;
  assign y2356 = ~n12108 ;
  assign y2357 = n12122 ;
  assign y2358 = n12124 ;
  assign y2359 = ~n12129 ;
  assign y2360 = n12131 ;
  assign y2361 = ~n12135 ;
  assign y2362 = ~n12140 ;
  assign y2363 = ~1'b0 ;
  assign y2364 = n12144 ;
  assign y2365 = ~n12154 ;
  assign y2366 = n12161 ;
  assign y2367 = n12165 ;
  assign y2368 = ~n12176 ;
  assign y2369 = n12179 ;
  assign y2370 = ~n12182 ;
  assign y2371 = n12183 ;
  assign y2372 = n12184 ;
  assign y2373 = ~n12190 ;
  assign y2374 = n12197 ;
  assign y2375 = ~n12199 ;
  assign y2376 = n12202 ;
  assign y2377 = n12203 ;
  assign y2378 = ~n12207 ;
  assign y2379 = ~n12209 ;
  assign y2380 = ~1'b0 ;
  assign y2381 = ~n12232 ;
  assign y2382 = ~n12234 ;
  assign y2383 = ~n12235 ;
  assign y2384 = n12244 ;
  assign y2385 = ~n12246 ;
  assign y2386 = n12254 ;
  assign y2387 = ~n12258 ;
  assign y2388 = ~n12259 ;
  assign y2389 = ~n12262 ;
  assign y2390 = n12271 ;
  assign y2391 = n12272 ;
  assign y2392 = n12281 ;
  assign y2393 = n12282 ;
  assign y2394 = ~n12285 ;
  assign y2395 = n12289 ;
  assign y2396 = ~n12291 ;
  assign y2397 = n12298 ;
  assign y2398 = ~n12302 ;
  assign y2399 = ~1'b0 ;
  assign y2400 = ~n12303 ;
  assign y2401 = ~n12304 ;
  assign y2402 = ~1'b0 ;
  assign y2403 = n12311 ;
  assign y2404 = ~n12317 ;
  assign y2405 = n12318 ;
  assign y2406 = ~n12321 ;
  assign y2407 = ~n12325 ;
  assign y2408 = n12327 ;
  assign y2409 = ~n12328 ;
  assign y2410 = n12330 ;
  assign y2411 = ~n12332 ;
  assign y2412 = n12335 ;
  assign y2413 = n12343 ;
  assign y2414 = ~n12349 ;
  assign y2415 = ~n12351 ;
  assign y2416 = ~n12356 ;
  assign y2417 = ~n12361 ;
  assign y2418 = n12363 ;
  assign y2419 = n12370 ;
  assign y2420 = n12376 ;
  assign y2421 = ~n12379 ;
  assign y2422 = ~1'b0 ;
  assign y2423 = n12381 ;
  assign y2424 = n12383 ;
  assign y2425 = ~n12392 ;
  assign y2426 = ~n12396 ;
  assign y2427 = ~n12397 ;
  assign y2428 = ~n12403 ;
  assign y2429 = ~n12405 ;
  assign y2430 = ~n12409 ;
  assign y2431 = ~1'b0 ;
  assign y2432 = n12412 ;
  assign y2433 = n12413 ;
  assign y2434 = ~n12418 ;
  assign y2435 = ~n12428 ;
  assign y2436 = ~n12431 ;
  assign y2437 = ~n12432 ;
  assign y2438 = n12433 ;
  assign y2439 = ~n12434 ;
  assign y2440 = ~n12445 ;
  assign y2441 = ~1'b0 ;
  assign y2442 = ~n12450 ;
  assign y2443 = n12451 ;
  assign y2444 = ~n12452 ;
  assign y2445 = ~n12459 ;
  assign y2446 = ~n12461 ;
  assign y2447 = n12465 ;
  assign y2448 = ~n12467 ;
  assign y2449 = ~n12476 ;
  assign y2450 = n12479 ;
  assign y2451 = n12487 ;
  assign y2452 = n12494 ;
  assign y2453 = n12495 ;
  assign y2454 = ~n12506 ;
  assign y2455 = n12507 ;
  assign y2456 = ~n12514 ;
  assign y2457 = n12516 ;
  assign y2458 = ~n12518 ;
  assign y2459 = n12525 ;
  assign y2460 = n12533 ;
  assign y2461 = ~n12540 ;
  assign y2462 = n12545 ;
  assign y2463 = ~n12549 ;
  assign y2464 = n12556 ;
  assign y2465 = n12558 ;
  assign y2466 = n12560 ;
  assign y2467 = n12564 ;
  assign y2468 = n12568 ;
  assign y2469 = n12569 ;
  assign y2470 = n12574 ;
  assign y2471 = n12582 ;
  assign y2472 = ~1'b0 ;
  assign y2473 = ~n12585 ;
  assign y2474 = ~n12587 ;
  assign y2475 = ~n12588 ;
  assign y2476 = ~n12590 ;
  assign y2477 = n12591 ;
  assign y2478 = n12593 ;
  assign y2479 = ~n12597 ;
  assign y2480 = ~n12601 ;
  assign y2481 = ~n12604 ;
  assign y2482 = n12612 ;
  assign y2483 = n12619 ;
  assign y2484 = ~n12628 ;
  assign y2485 = n12629 ;
  assign y2486 = ~n12634 ;
  assign y2487 = ~n12638 ;
  assign y2488 = n12639 ;
  assign y2489 = ~n12641 ;
  assign y2490 = ~n12644 ;
  assign y2491 = ~n12645 ;
  assign y2492 = ~n12652 ;
  assign y2493 = n12655 ;
  assign y2494 = n12668 ;
  assign y2495 = n12669 ;
  assign y2496 = n12671 ;
  assign y2497 = n12675 ;
  assign y2498 = n12676 ;
  assign y2499 = n12680 ;
  assign y2500 = n12685 ;
  assign y2501 = n12693 ;
  assign y2502 = n12701 ;
  assign y2503 = ~n12702 ;
  assign y2504 = n12706 ;
  assign y2505 = n12715 ;
  assign y2506 = n12721 ;
  assign y2507 = ~n12725 ;
  assign y2508 = n12727 ;
  assign y2509 = n12733 ;
  assign y2510 = n12736 ;
  assign y2511 = ~n12738 ;
  assign y2512 = ~n12747 ;
  assign y2513 = n12755 ;
  assign y2514 = n12756 ;
  assign y2515 = n12759 ;
  assign y2516 = n12765 ;
  assign y2517 = ~n12766 ;
  assign y2518 = ~n12768 ;
  assign y2519 = n12769 ;
  assign y2520 = n12772 ;
  assign y2521 = n12783 ;
  assign y2522 = ~n12787 ;
  assign y2523 = n12788 ;
  assign y2524 = ~n12792 ;
  assign y2525 = n12804 ;
  assign y2526 = ~n4281 ;
  assign y2527 = ~n12807 ;
  assign y2528 = ~n12810 ;
  assign y2529 = ~n12815 ;
  assign y2530 = n12823 ;
  assign y2531 = ~n12825 ;
  assign y2532 = n12834 ;
  assign y2533 = ~n12838 ;
  assign y2534 = ~n12840 ;
  assign y2535 = ~n12841 ;
  assign y2536 = ~1'b0 ;
  assign y2537 = n12845 ;
  assign y2538 = ~n12847 ;
  assign y2539 = n12855 ;
  assign y2540 = n12861 ;
  assign y2541 = n12870 ;
  assign y2542 = n12872 ;
  assign y2543 = n12876 ;
  assign y2544 = n12891 ;
  assign y2545 = ~n12899 ;
  assign y2546 = ~n12901 ;
  assign y2547 = ~n12904 ;
  assign y2548 = ~n12905 ;
  assign y2549 = n12906 ;
  assign y2550 = ~n12908 ;
  assign y2551 = ~n12912 ;
  assign y2552 = n12915 ;
  assign y2553 = ~1'b0 ;
  assign y2554 = n12917 ;
  assign y2555 = ~n12920 ;
  assign y2556 = ~n12926 ;
  assign y2557 = ~n12927 ;
  assign y2558 = ~n12931 ;
  assign y2559 = n12933 ;
  assign y2560 = ~1'b0 ;
  assign y2561 = ~n12935 ;
  assign y2562 = ~n12937 ;
  assign y2563 = n12944 ;
  assign y2564 = ~n12950 ;
  assign y2565 = n12952 ;
  assign y2566 = n12954 ;
  assign y2567 = ~n12960 ;
  assign y2568 = n12964 ;
  assign y2569 = ~n12969 ;
  assign y2570 = n12972 ;
  assign y2571 = ~n12978 ;
  assign y2572 = n12981 ;
  assign y2573 = ~n12982 ;
  assign y2574 = ~n12984 ;
  assign y2575 = ~1'b0 ;
  assign y2576 = n12989 ;
  assign y2577 = n12995 ;
  assign y2578 = ~n12998 ;
  assign y2579 = ~n13000 ;
  assign y2580 = n13008 ;
  assign y2581 = ~n13013 ;
  assign y2582 = ~n13016 ;
  assign y2583 = ~n13020 ;
  assign y2584 = n13023 ;
  assign y2585 = n13024 ;
  assign y2586 = n13029 ;
  assign y2587 = ~n13033 ;
  assign y2588 = n13037 ;
  assign y2589 = n13041 ;
  assign y2590 = n13057 ;
  assign y2591 = n13059 ;
  assign y2592 = n13060 ;
  assign y2593 = n13068 ;
  assign y2594 = n13070 ;
  assign y2595 = ~n13076 ;
  assign y2596 = ~n13078 ;
  assign y2597 = ~n13086 ;
  assign y2598 = ~n13089 ;
  assign y2599 = n13092 ;
  assign y2600 = n13099 ;
  assign y2601 = n13101 ;
  assign y2602 = ~n13111 ;
  assign y2603 = ~1'b0 ;
  assign y2604 = ~n13112 ;
  assign y2605 = ~n13118 ;
  assign y2606 = ~n13119 ;
  assign y2607 = ~n13121 ;
  assign y2608 = ~1'b0 ;
  assign y2609 = ~n13122 ;
  assign y2610 = n4057 ;
  assign y2611 = ~n13130 ;
  assign y2612 = ~n13132 ;
  assign y2613 = ~n13133 ;
  assign y2614 = n13137 ;
  assign y2615 = ~n13142 ;
  assign y2616 = ~n13145 ;
  assign y2617 = n13148 ;
  assign y2618 = ~n13151 ;
  assign y2619 = ~n13157 ;
  assign y2620 = n13161 ;
  assign y2621 = ~n13167 ;
  assign y2622 = n13178 ;
  assign y2623 = ~n13181 ;
  assign y2624 = n13198 ;
  assign y2625 = ~n13201 ;
  assign y2626 = ~n13202 ;
  assign y2627 = n13204 ;
  assign y2628 = ~n13208 ;
  assign y2629 = n13211 ;
  assign y2630 = ~n13212 ;
  assign y2631 = ~1'b0 ;
  assign y2632 = ~n13215 ;
  assign y2633 = n13196 ;
  assign y2634 = ~n13219 ;
  assign y2635 = ~n13224 ;
  assign y2636 = n13225 ;
  assign y2637 = ~n13228 ;
  assign y2638 = ~n13231 ;
  assign y2639 = n13233 ;
  assign y2640 = ~n13238 ;
  assign y2641 = n13240 ;
  assign y2642 = ~n13241 ;
  assign y2643 = ~n13244 ;
  assign y2644 = ~n13251 ;
  assign y2645 = ~1'b0 ;
  assign y2646 = n13255 ;
  assign y2647 = ~1'b0 ;
  assign y2648 = n13256 ;
  assign y2649 = ~n13257 ;
  assign y2650 = ~1'b0 ;
  assign y2651 = n13259 ;
  assign y2652 = ~n13260 ;
  assign y2653 = n13268 ;
  assign y2654 = n13269 ;
  assign y2655 = n13277 ;
  assign y2656 = n13280 ;
  assign y2657 = n13281 ;
  assign y2658 = n13284 ;
  assign y2659 = ~n13287 ;
  assign y2660 = n13290 ;
  assign y2661 = ~n13296 ;
  assign y2662 = ~n13297 ;
  assign y2663 = n13302 ;
  assign y2664 = ~1'b0 ;
  assign y2665 = ~n13311 ;
  assign y2666 = ~n13320 ;
  assign y2667 = n13323 ;
  assign y2668 = ~n13330 ;
  assign y2669 = ~n13331 ;
  assign y2670 = n13332 ;
  assign y2671 = ~n13335 ;
  assign y2672 = n13344 ;
  assign y2673 = n13348 ;
  assign y2674 = ~1'b0 ;
  assign y2675 = ~n13353 ;
  assign y2676 = ~n13355 ;
  assign y2677 = n13358 ;
  assign y2678 = ~n13361 ;
  assign y2679 = n13363 ;
  assign y2680 = ~n2703 ;
  assign y2681 = ~n13370 ;
  assign y2682 = ~n13377 ;
  assign y2683 = n13381 ;
  assign y2684 = n13392 ;
  assign y2685 = ~n13393 ;
  assign y2686 = ~n13398 ;
  assign y2687 = n13401 ;
  assign y2688 = n13404 ;
  assign y2689 = n13408 ;
  assign y2690 = ~n13411 ;
  assign y2691 = n13413 ;
  assign y2692 = ~n13414 ;
  assign y2693 = n13417 ;
  assign y2694 = ~n13419 ;
  assign y2695 = n13423 ;
  assign y2696 = ~n13425 ;
  assign y2697 = n13431 ;
  assign y2698 = n13441 ;
  assign y2699 = n13450 ;
  assign y2700 = ~n13452 ;
  assign y2701 = ~n13454 ;
  assign y2702 = ~n13455 ;
  assign y2703 = ~n13456 ;
  assign y2704 = ~1'b0 ;
  assign y2705 = ~n13457 ;
  assign y2706 = ~n13461 ;
  assign y2707 = ~n13464 ;
  assign y2708 = ~n13469 ;
  assign y2709 = n13470 ;
  assign y2710 = ~n13472 ;
  assign y2711 = ~n13473 ;
  assign y2712 = ~n13474 ;
  assign y2713 = ~n13479 ;
  assign y2714 = ~n13483 ;
  assign y2715 = n13497 ;
  assign y2716 = n13503 ;
  assign y2717 = ~n13506 ;
  assign y2718 = ~1'b0 ;
  assign y2719 = n13508 ;
  assign y2720 = n13512 ;
  assign y2721 = ~n13514 ;
  assign y2722 = n13529 ;
  assign y2723 = ~1'b0 ;
  assign y2724 = ~n13531 ;
  assign y2725 = ~n13539 ;
  assign y2726 = ~n13541 ;
  assign y2727 = n13543 ;
  assign y2728 = n13545 ;
  assign y2729 = ~n13554 ;
  assign y2730 = ~n13560 ;
  assign y2731 = n13561 ;
  assign y2732 = n13562 ;
  assign y2733 = n13563 ;
  assign y2734 = ~n13565 ;
  assign y2735 = ~n13567 ;
  assign y2736 = ~n13569 ;
  assign y2737 = ~n13574 ;
  assign y2738 = ~n13575 ;
  assign y2739 = ~n13578 ;
  assign y2740 = ~1'b0 ;
  assign y2741 = ~n13579 ;
  assign y2742 = ~n13580 ;
  assign y2743 = ~n13585 ;
  assign y2744 = n13589 ;
  assign y2745 = ~n13591 ;
  assign y2746 = n13595 ;
  assign y2747 = ~n13599 ;
  assign y2748 = ~n13601 ;
  assign y2749 = ~n13608 ;
  assign y2750 = ~n13631 ;
  assign y2751 = n13632 ;
  assign y2752 = ~n13639 ;
  assign y2753 = ~n13641 ;
  assign y2754 = n13642 ;
  assign y2755 = n13644 ;
  assign y2756 = n13656 ;
  assign y2757 = ~n13659 ;
  assign y2758 = ~n13668 ;
  assign y2759 = ~n13670 ;
  assign y2760 = n13675 ;
  assign y2761 = ~n13677 ;
  assign y2762 = n13679 ;
  assign y2763 = ~n13681 ;
  assign y2764 = n13686 ;
  assign y2765 = ~n13687 ;
  assign y2766 = n13688 ;
  assign y2767 = ~n13689 ;
  assign y2768 = n13693 ;
  assign y2769 = ~1'b0 ;
  assign y2770 = n13707 ;
  assign y2771 = n13714 ;
  assign y2772 = n13716 ;
  assign y2773 = ~n13718 ;
  assign y2774 = ~n13726 ;
  assign y2775 = n13732 ;
  assign y2776 = ~1'b0 ;
  assign y2777 = n13733 ;
  assign y2778 = ~n13738 ;
  assign y2779 = ~n13746 ;
  assign y2780 = n13747 ;
  assign y2781 = n13755 ;
  assign y2782 = n13759 ;
  assign y2783 = n13760 ;
  assign y2784 = ~n13765 ;
  assign y2785 = n13766 ;
  assign y2786 = n13773 ;
  assign y2787 = ~n13784 ;
  assign y2788 = n13785 ;
  assign y2789 = ~n13788 ;
  assign y2790 = n13793 ;
  assign y2791 = n13794 ;
  assign y2792 = ~n13803 ;
  assign y2793 = n13806 ;
  assign y2794 = ~n13812 ;
  assign y2795 = n13819 ;
  assign y2796 = n13821 ;
  assign y2797 = ~n13828 ;
  assign y2798 = ~n13829 ;
  assign y2799 = n13831 ;
  assign y2800 = ~1'b0 ;
  assign y2801 = n13837 ;
  assign y2802 = ~n13840 ;
  assign y2803 = ~n13842 ;
  assign y2804 = ~n13845 ;
  assign y2805 = n13848 ;
  assign y2806 = ~n13851 ;
  assign y2807 = n13860 ;
  assign y2808 = ~1'b0 ;
  assign y2809 = ~n13861 ;
  assign y2810 = n13863 ;
  assign y2811 = n13869 ;
  assign y2812 = ~n13871 ;
  assign y2813 = ~n13877 ;
  assign y2814 = ~n13878 ;
  assign y2815 = n13888 ;
  assign y2816 = ~n13889 ;
  assign y2817 = ~n13891 ;
  assign y2818 = ~n13894 ;
  assign y2819 = ~n13897 ;
  assign y2820 = ~n13899 ;
  assign y2821 = n13902 ;
  assign y2822 = ~n13904 ;
  assign y2823 = n13905 ;
  assign y2824 = n13906 ;
  assign y2825 = ~n13908 ;
  assign y2826 = ~n13911 ;
  assign y2827 = n13914 ;
  assign y2828 = n13923 ;
  assign y2829 = n13926 ;
  assign y2830 = ~n13928 ;
  assign y2831 = ~n13936 ;
  assign y2832 = ~n13941 ;
  assign y2833 = n13942 ;
  assign y2834 = n13951 ;
  assign y2835 = ~n13953 ;
  assign y2836 = ~n13955 ;
  assign y2837 = ~n13956 ;
  assign y2838 = ~n13958 ;
  assign y2839 = ~n13961 ;
  assign y2840 = n13963 ;
  assign y2841 = ~n13964 ;
  assign y2842 = ~n13968 ;
  assign y2843 = n13969 ;
  assign y2844 = ~1'b0 ;
  assign y2845 = ~1'b0 ;
  assign y2846 = n13970 ;
  assign y2847 = ~n13973 ;
  assign y2848 = ~n13977 ;
  assign y2849 = ~n13986 ;
  assign y2850 = ~n13987 ;
  assign y2851 = ~n13989 ;
  assign y2852 = n13993 ;
  assign y2853 = n13996 ;
  assign y2854 = n13998 ;
  assign y2855 = n14014 ;
  assign y2856 = ~n14025 ;
  assign y2857 = ~n14028 ;
  assign y2858 = ~n14029 ;
  assign y2859 = ~n14031 ;
  assign y2860 = ~1'b0 ;
  assign y2861 = n14036 ;
  assign y2862 = ~1'b0 ;
  assign y2863 = n14037 ;
  assign y2864 = n14043 ;
  assign y2865 = ~n14048 ;
  assign y2866 = ~n14049 ;
  assign y2867 = ~n14050 ;
  assign y2868 = n14052 ;
  assign y2869 = n14058 ;
  assign y2870 = ~n14060 ;
  assign y2871 = n14061 ;
  assign y2872 = n14063 ;
  assign y2873 = n14064 ;
  assign y2874 = ~n14067 ;
  assign y2875 = ~n14071 ;
  assign y2876 = ~n14074 ;
  assign y2877 = n14075 ;
  assign y2878 = ~n14077 ;
  assign y2879 = ~n14078 ;
  assign y2880 = n14081 ;
  assign y2881 = ~n14083 ;
  assign y2882 = n14084 ;
  assign y2883 = n14097 ;
  assign y2884 = ~n14099 ;
  assign y2885 = ~n14110 ;
  assign y2886 = n14119 ;
  assign y2887 = n14121 ;
  assign y2888 = n14123 ;
  assign y2889 = n14124 ;
  assign y2890 = ~1'b0 ;
  assign y2891 = ~n14128 ;
  assign y2892 = ~1'b0 ;
  assign y2893 = n14130 ;
  assign y2894 = n14131 ;
  assign y2895 = ~n14132 ;
  assign y2896 = ~n14135 ;
  assign y2897 = ~n14139 ;
  assign y2898 = ~n14142 ;
  assign y2899 = ~n14150 ;
  assign y2900 = n14157 ;
  assign y2901 = n14162 ;
  assign y2902 = ~n14164 ;
  assign y2903 = ~n14170 ;
  assign y2904 = ~n14172 ;
  assign y2905 = ~n14174 ;
  assign y2906 = n14175 ;
  assign y2907 = n14179 ;
  assign y2908 = n14180 ;
  assign y2909 = ~n14185 ;
  assign y2910 = ~n14190 ;
  assign y2911 = n14191 ;
  assign y2912 = ~n14194 ;
  assign y2913 = n14199 ;
  assign y2914 = ~n14203 ;
  assign y2915 = ~n14204 ;
  assign y2916 = ~n14208 ;
  assign y2917 = n14210 ;
  assign y2918 = n14215 ;
  assign y2919 = ~n14219 ;
  assign y2920 = ~n14224 ;
  assign y2921 = ~n14226 ;
  assign y2922 = n14230 ;
  assign y2923 = ~n14237 ;
  assign y2924 = ~1'b0 ;
  assign y2925 = ~n14238 ;
  assign y2926 = n14240 ;
  assign y2927 = n14242 ;
  assign y2928 = ~n14245 ;
  assign y2929 = n14248 ;
  assign y2930 = ~n14250 ;
  assign y2931 = ~1'b0 ;
  assign y2932 = ~n14253 ;
  assign y2933 = n14255 ;
  assign y2934 = n14256 ;
  assign y2935 = n14258 ;
  assign y2936 = ~n14260 ;
  assign y2937 = ~n14263 ;
  assign y2938 = n14273 ;
  assign y2939 = ~n14276 ;
  assign y2940 = n14280 ;
  assign y2941 = ~n14281 ;
  assign y2942 = ~n14282 ;
  assign y2943 = ~n14292 ;
  assign y2944 = ~n14294 ;
  assign y2945 = n14295 ;
  assign y2946 = n14298 ;
  assign y2947 = n14304 ;
  assign y2948 = ~n14312 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = n13683 ;
  assign y2951 = n14314 ;
  assign y2952 = ~n14319 ;
  assign y2953 = n14320 ;
  assign y2954 = ~n14324 ;
  assign y2955 = ~n14327 ;
  assign y2956 = n14340 ;
  assign y2957 = ~n14341 ;
  assign y2958 = n14346 ;
  assign y2959 = ~n14350 ;
  assign y2960 = n14351 ;
  assign y2961 = ~n14355 ;
  assign y2962 = n14356 ;
  assign y2963 = n14361 ;
  assign y2964 = ~n14365 ;
  assign y2965 = ~n14369 ;
  assign y2966 = n14371 ;
  assign y2967 = n14373 ;
  assign y2968 = ~n14379 ;
  assign y2969 = n14385 ;
  assign y2970 = ~n14389 ;
  assign y2971 = ~n14390 ;
  assign y2972 = ~n14393 ;
  assign y2973 = n14394 ;
  assign y2974 = n14396 ;
  assign y2975 = ~n14398 ;
  assign y2976 = n14399 ;
  assign y2977 = n14400 ;
  assign y2978 = n14405 ;
  assign y2979 = ~n14409 ;
  assign y2980 = ~n14416 ;
  assign y2981 = ~n14419 ;
  assign y2982 = ~n14425 ;
  assign y2983 = ~n14427 ;
  assign y2984 = n14430 ;
  assign y2985 = n14432 ;
  assign y2986 = ~n14438 ;
  assign y2987 = ~n14447 ;
  assign y2988 = n14452 ;
  assign y2989 = ~n14457 ;
  assign y2990 = n14462 ;
  assign y2991 = n14463 ;
  assign y2992 = n14465 ;
  assign y2993 = n14467 ;
  assign y2994 = ~n14469 ;
  assign y2995 = ~n14471 ;
  assign y2996 = n14472 ;
  assign y2997 = n14473 ;
  assign y2998 = n14476 ;
  assign y2999 = ~n14479 ;
  assign y3000 = n14480 ;
  assign y3001 = ~n14482 ;
  assign y3002 = ~n14486 ;
  assign y3003 = n14494 ;
  assign y3004 = n14497 ;
  assign y3005 = n14502 ;
  assign y3006 = n14508 ;
  assign y3007 = ~n14511 ;
  assign y3008 = n14513 ;
  assign y3009 = n14519 ;
  assign y3010 = n14521 ;
  assign y3011 = n14523 ;
  assign y3012 = n14527 ;
  assign y3013 = n14529 ;
  assign y3014 = n14531 ;
  assign y3015 = n14542 ;
  assign y3016 = n14544 ;
  assign y3017 = n14549 ;
  assign y3018 = ~n14556 ;
  assign y3019 = n14558 ;
  assign y3020 = ~1'b0 ;
  assign y3021 = ~1'b0 ;
  assign y3022 = n14566 ;
  assign y3023 = n14572 ;
  assign y3024 = n14573 ;
  assign y3025 = n14574 ;
  assign y3026 = ~1'b0 ;
  assign y3027 = n14576 ;
  assign y3028 = ~n14580 ;
  assign y3029 = ~n14582 ;
  assign y3030 = ~n14586 ;
  assign y3031 = n14588 ;
  assign y3032 = n14598 ;
  assign y3033 = ~n14600 ;
  assign y3034 = ~n14601 ;
  assign y3035 = ~n14604 ;
  assign y3036 = n14605 ;
  assign y3037 = ~n14613 ;
  assign y3038 = n14617 ;
  assign y3039 = ~n14618 ;
  assign y3040 = ~n14620 ;
  assign y3041 = ~n14622 ;
  assign y3042 = n14626 ;
  assign y3043 = n14629 ;
  assign y3044 = ~n14630 ;
  assign y3045 = ~n14632 ;
  assign y3046 = ~n14633 ;
  assign y3047 = ~n14635 ;
  assign y3048 = ~1'b0 ;
  assign y3049 = ~n14636 ;
  assign y3050 = ~n14648 ;
  assign y3051 = ~1'b0 ;
  assign y3052 = ~n14655 ;
  assign y3053 = ~n14657 ;
  assign y3054 = n14658 ;
  assign y3055 = n14663 ;
  assign y3056 = n14666 ;
  assign y3057 = ~n14667 ;
  assign y3058 = n14674 ;
  assign y3059 = n14681 ;
  assign y3060 = ~n14683 ;
  assign y3061 = ~n14684 ;
  assign y3062 = ~n14685 ;
  assign y3063 = n14689 ;
  assign y3064 = ~n14692 ;
  assign y3065 = ~n14697 ;
  assign y3066 = ~n14700 ;
  assign y3067 = ~n14705 ;
  assign y3068 = ~1'b0 ;
  assign y3069 = ~n14707 ;
  assign y3070 = n14710 ;
  assign y3071 = ~n14718 ;
  assign y3072 = n14719 ;
  assign y3073 = n14723 ;
  assign y3074 = n14724 ;
  assign y3075 = n14726 ;
  assign y3076 = n14727 ;
  assign y3077 = n14733 ;
  assign y3078 = ~n14737 ;
  assign y3079 = n14749 ;
  assign y3080 = ~n14756 ;
  assign y3081 = n14757 ;
  assign y3082 = ~n14758 ;
  assign y3083 = n14760 ;
  assign y3084 = n14764 ;
  assign y3085 = ~n14766 ;
  assign y3086 = ~n14767 ;
  assign y3087 = ~n14771 ;
  assign y3088 = ~n14772 ;
  assign y3089 = n14773 ;
  assign y3090 = ~1'b0 ;
  assign y3091 = n14778 ;
  assign y3092 = ~n14779 ;
  assign y3093 = n14781 ;
  assign y3094 = n14782 ;
  assign y3095 = n14783 ;
  assign y3096 = n14785 ;
  assign y3097 = ~n14790 ;
  assign y3098 = n14792 ;
  assign y3099 = ~1'b0 ;
  assign y3100 = n14797 ;
  assign y3101 = n14798 ;
  assign y3102 = ~n14799 ;
  assign y3103 = ~1'b0 ;
  assign y3104 = n14812 ;
  assign y3105 = n14813 ;
  assign y3106 = n14816 ;
  assign y3107 = n14823 ;
  assign y3108 = n14825 ;
  assign y3109 = ~n14828 ;
  assign y3110 = ~n14831 ;
  assign y3111 = ~1'b0 ;
  assign y3112 = ~n14835 ;
  assign y3113 = ~n14854 ;
  assign y3114 = ~n14858 ;
  assign y3115 = n14862 ;
  assign y3116 = ~n14866 ;
  assign y3117 = n14872 ;
  assign y3118 = ~1'b0 ;
  assign y3119 = ~n14882 ;
  assign y3120 = ~n14885 ;
  assign y3121 = n14889 ;
  assign y3122 = n14895 ;
  assign y3123 = n14899 ;
  assign y3124 = n14908 ;
  assign y3125 = ~n14916 ;
  assign y3126 = ~n14918 ;
  assign y3127 = ~n14922 ;
  assign y3128 = n14924 ;
  assign y3129 = n14928 ;
  assign y3130 = ~n14930 ;
  assign y3131 = n14936 ;
  assign y3132 = n14944 ;
  assign y3133 = ~n14946 ;
  assign y3134 = ~n14948 ;
  assign y3135 = n14949 ;
  assign y3136 = ~n14956 ;
  assign y3137 = ~1'b0 ;
  assign y3138 = n14961 ;
  assign y3139 = ~n14967 ;
  assign y3140 = ~n14969 ;
  assign y3141 = ~n14970 ;
  assign y3142 = n14972 ;
  assign y3143 = n14973 ;
  assign y3144 = n14975 ;
  assign y3145 = ~1'b0 ;
  assign y3146 = n14982 ;
  assign y3147 = ~n14986 ;
  assign y3148 = n14990 ;
  assign y3149 = n14999 ;
  assign y3150 = n15005 ;
  assign y3151 = ~n15009 ;
  assign y3152 = ~n15010 ;
  assign y3153 = n15017 ;
  assign y3154 = n15020 ;
  assign y3155 = ~n15021 ;
  assign y3156 = ~n15032 ;
  assign y3157 = n15034 ;
  assign y3158 = n15043 ;
  assign y3159 = n15046 ;
  assign y3160 = n15047 ;
  assign y3161 = n15050 ;
  assign y3162 = ~n15056 ;
  assign y3163 = ~n15061 ;
  assign y3164 = ~n15062 ;
  assign y3165 = ~n15068 ;
  assign y3166 = n15070 ;
  assign y3167 = ~n15074 ;
  assign y3168 = n15079 ;
  assign y3169 = n15083 ;
  assign y3170 = ~n15087 ;
  assign y3171 = n15089 ;
  assign y3172 = n15092 ;
  assign y3173 = ~n15093 ;
  assign y3174 = ~n15095 ;
  assign y3175 = ~1'b0 ;
  assign y3176 = ~n15111 ;
  assign y3177 = n15112 ;
  assign y3178 = n15117 ;
  assign y3179 = n15119 ;
  assign y3180 = n15122 ;
  assign y3181 = ~n15123 ;
  assign y3182 = n15126 ;
  assign y3183 = n15127 ;
  assign y3184 = n15129 ;
  assign y3185 = ~n15130 ;
  assign y3186 = ~1'b0 ;
  assign y3187 = ~n15138 ;
  assign y3188 = ~n15142 ;
  assign y3189 = ~n15145 ;
  assign y3190 = ~n15147 ;
  assign y3191 = ~n15153 ;
  assign y3192 = ~n15166 ;
  assign y3193 = ~n15171 ;
  assign y3194 = ~n15173 ;
  assign y3195 = ~n15181 ;
  assign y3196 = ~n15185 ;
  assign y3197 = ~n15186 ;
  assign y3198 = ~1'b0 ;
  assign y3199 = n15189 ;
  assign y3200 = n15192 ;
  assign y3201 = n15194 ;
  assign y3202 = ~n15198 ;
  assign y3203 = n15200 ;
  assign y3204 = ~n15202 ;
  assign y3205 = n15204 ;
  assign y3206 = ~n15207 ;
  assign y3207 = ~n15209 ;
  assign y3208 = ~n15210 ;
  assign y3209 = n15211 ;
  assign y3210 = n15212 ;
  assign y3211 = n15220 ;
  assign y3212 = ~n15222 ;
  assign y3213 = n15227 ;
  assign y3214 = n15232 ;
  assign y3215 = ~n15236 ;
  assign y3216 = ~n15237 ;
  assign y3217 = ~n15238 ;
  assign y3218 = ~n15241 ;
  assign y3219 = ~n15244 ;
  assign y3220 = ~n15246 ;
  assign y3221 = n15249 ;
  assign y3222 = ~1'b0 ;
  assign y3223 = ~n15252 ;
  assign y3224 = n15255 ;
  assign y3225 = 1'b0 ;
  assign y3226 = ~n15259 ;
  assign y3227 = n15270 ;
  assign y3228 = n15273 ;
  assign y3229 = n15279 ;
  assign y3230 = 1'b0 ;
  assign y3231 = n15280 ;
  assign y3232 = ~n15282 ;
  assign y3233 = ~n15284 ;
  assign y3234 = ~n15287 ;
  assign y3235 = ~n15288 ;
  assign y3236 = n15296 ;
  assign y3237 = ~n15297 ;
  assign y3238 = n15300 ;
  assign y3239 = n15304 ;
  assign y3240 = n15307 ;
  assign y3241 = ~1'b0 ;
  assign y3242 = n15308 ;
  assign y3243 = ~n15309 ;
  assign y3244 = n15313 ;
  assign y3245 = n15315 ;
  assign y3246 = ~n15318 ;
  assign y3247 = ~n15321 ;
  assign y3248 = n15327 ;
  assign y3249 = n15329 ;
  assign y3250 = ~n15331 ;
  assign y3251 = ~n15335 ;
  assign y3252 = n15336 ;
  assign y3253 = ~1'b0 ;
  assign y3254 = n15342 ;
  assign y3255 = n15343 ;
  assign y3256 = ~n15344 ;
  assign y3257 = ~1'b0 ;
  assign y3258 = n15346 ;
  assign y3259 = n15353 ;
  assign y3260 = n15362 ;
  assign y3261 = ~n15367 ;
  assign y3262 = ~n15372 ;
  assign y3263 = n15374 ;
  assign y3264 = ~1'b0 ;
  assign y3265 = ~n15375 ;
  assign y3266 = ~n15376 ;
  assign y3267 = n15378 ;
  assign y3268 = ~1'b0 ;
  assign y3269 = ~n15382 ;
  assign y3270 = ~n15387 ;
  assign y3271 = ~1'b0 ;
  assign y3272 = n15394 ;
  assign y3273 = ~1'b0 ;
  assign y3274 = ~n15397 ;
  assign y3275 = ~n15404 ;
  assign y3276 = ~n15410 ;
  assign y3277 = ~n15411 ;
  assign y3278 = ~n15413 ;
  assign y3279 = ~n15416 ;
  assign y3280 = ~n15418 ;
  assign y3281 = n15419 ;
  assign y3282 = n15421 ;
  assign y3283 = ~n15424 ;
  assign y3284 = ~n15426 ;
  assign y3285 = n15431 ;
  assign y3286 = n15432 ;
  assign y3287 = ~n15437 ;
  assign y3288 = n15438 ;
  assign y3289 = n15442 ;
  assign y3290 = ~n15446 ;
  assign y3291 = ~n15460 ;
  assign y3292 = n15461 ;
  assign y3293 = n15466 ;
  assign y3294 = n15470 ;
  assign y3295 = n15471 ;
  assign y3296 = n15477 ;
  assign y3297 = n15480 ;
  assign y3298 = ~n15490 ;
  assign y3299 = n15492 ;
  assign y3300 = n15493 ;
  assign y3301 = n15494 ;
  assign y3302 = n12614 ;
  assign y3303 = n15497 ;
  assign y3304 = n15500 ;
  assign y3305 = ~n15505 ;
  assign y3306 = ~n15515 ;
  assign y3307 = ~n15520 ;
  assign y3308 = ~n15522 ;
  assign y3309 = n15530 ;
  assign y3310 = ~n15539 ;
  assign y3311 = ~n15540 ;
  assign y3312 = n15541 ;
  assign y3313 = ~n15542 ;
  assign y3314 = n15544 ;
  assign y3315 = ~n15548 ;
  assign y3316 = ~n15551 ;
  assign y3317 = ~n15552 ;
  assign y3318 = ~n15554 ;
  assign y3319 = n15555 ;
  assign y3320 = n15556 ;
  assign y3321 = ~n15558 ;
  assign y3322 = n15564 ;
  assign y3323 = ~1'b0 ;
  assign y3324 = ~n15567 ;
  assign y3325 = n15573 ;
  assign y3326 = ~n15577 ;
  assign y3327 = ~n15585 ;
  assign y3328 = n15586 ;
  assign y3329 = ~n15588 ;
  assign y3330 = ~n15591 ;
  assign y3331 = ~n15595 ;
  assign y3332 = n15596 ;
  assign y3333 = ~n15598 ;
  assign y3334 = ~n15601 ;
  assign y3335 = n15605 ;
  assign y3336 = ~n15607 ;
  assign y3337 = n15608 ;
  assign y3338 = ~n15611 ;
  assign y3339 = n15621 ;
  assign y3340 = ~n15623 ;
  assign y3341 = ~n15624 ;
  assign y3342 = n15627 ;
  assign y3343 = ~n15628 ;
  assign y3344 = n15630 ;
  assign y3345 = ~n15631 ;
  assign y3346 = ~n15632 ;
  assign y3347 = n15640 ;
  assign y3348 = ~n15641 ;
  assign y3349 = n15645 ;
  assign y3350 = n15650 ;
  assign y3351 = ~1'b0 ;
  assign y3352 = n15653 ;
  assign y3353 = ~n15658 ;
  assign y3354 = ~n15662 ;
  assign y3355 = n15663 ;
  assign y3356 = n15669 ;
  assign y3357 = n15672 ;
  assign y3358 = n15680 ;
  assign y3359 = ~n15682 ;
  assign y3360 = n15686 ;
  assign y3361 = ~n15688 ;
  assign y3362 = n15692 ;
  assign y3363 = ~1'b0 ;
  assign y3364 = ~1'b0 ;
  assign y3365 = ~n15693 ;
  assign y3366 = ~n15698 ;
  assign y3367 = ~n15700 ;
  assign y3368 = n15705 ;
  assign y3369 = n15707 ;
  assign y3370 = ~n15711 ;
  assign y3371 = ~n15713 ;
  assign y3372 = n15716 ;
  assign y3373 = ~n15719 ;
  assign y3374 = ~n15725 ;
  assign y3375 = ~n15730 ;
  assign y3376 = ~n15731 ;
  assign y3377 = ~n15732 ;
  assign y3378 = n15734 ;
  assign y3379 = ~n15742 ;
  assign y3380 = n15743 ;
  assign y3381 = ~n15745 ;
  assign y3382 = ~1'b0 ;
  assign y3383 = ~n15749 ;
  assign y3384 = ~n15752 ;
  assign y3385 = n15755 ;
  assign y3386 = n15757 ;
  assign y3387 = ~n15763 ;
  assign y3388 = ~n15767 ;
  assign y3389 = ~n15768 ;
  assign y3390 = n15771 ;
  assign y3391 = ~n15773 ;
  assign y3392 = ~1'b0 ;
  assign y3393 = n15777 ;
  assign y3394 = n15782 ;
  assign y3395 = n15787 ;
  assign y3396 = n15789 ;
  assign y3397 = ~n15794 ;
  assign y3398 = ~n15798 ;
  assign y3399 = n15806 ;
  assign y3400 = n15810 ;
  assign y3401 = ~n15811 ;
  assign y3402 = n15817 ;
  assign y3403 = ~1'b0 ;
  assign y3404 = n15820 ;
  assign y3405 = n15824 ;
  assign y3406 = ~n15829 ;
  assign y3407 = n15830 ;
  assign y3408 = n15836 ;
  assign y3409 = ~n15841 ;
  assign y3410 = ~n15848 ;
  assign y3411 = n15855 ;
  assign y3412 = ~n15857 ;
  assign y3413 = ~n15858 ;
  assign y3414 = n15859 ;
  assign y3415 = ~n15863 ;
  assign y3416 = n15870 ;
  assign y3417 = ~n15871 ;
  assign y3418 = ~n15875 ;
  assign y3419 = ~n15877 ;
  assign y3420 = ~n15882 ;
  assign y3421 = n15883 ;
  assign y3422 = ~n15884 ;
  assign y3423 = n15886 ;
  assign y3424 = n15893 ;
  assign y3425 = ~n15894 ;
  assign y3426 = n15896 ;
  assign y3427 = n15904 ;
  assign y3428 = ~n15906 ;
  assign y3429 = ~n15907 ;
  assign y3430 = ~n15912 ;
  assign y3431 = ~n15917 ;
  assign y3432 = ~n15920 ;
  assign y3433 = n15923 ;
  assign y3434 = n15926 ;
  assign y3435 = n15929 ;
  assign y3436 = ~n15935 ;
  assign y3437 = n15939 ;
  assign y3438 = n15946 ;
  assign y3439 = n15947 ;
  assign y3440 = ~n15949 ;
  assign y3441 = n15950 ;
  assign y3442 = ~1'b0 ;
  assign y3443 = ~n15952 ;
  assign y3444 = ~n15954 ;
  assign y3445 = ~n15955 ;
  assign y3446 = n15961 ;
  assign y3447 = ~n15962 ;
  assign y3448 = n15963 ;
  assign y3449 = n15964 ;
  assign y3450 = n15966 ;
  assign y3451 = ~1'b0 ;
  assign y3452 = n15970 ;
  assign y3453 = n15972 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = n15980 ;
  assign y3456 = n15982 ;
  assign y3457 = n15983 ;
  assign y3458 = ~n15987 ;
  assign y3459 = n15990 ;
  assign y3460 = ~n15992 ;
  assign y3461 = n15994 ;
  assign y3462 = n15998 ;
  assign y3463 = ~n16003 ;
  assign y3464 = n16004 ;
  assign y3465 = n16005 ;
  assign y3466 = ~n16006 ;
  assign y3467 = ~n16009 ;
  assign y3468 = n16010 ;
  assign y3469 = n16021 ;
  assign y3470 = n16024 ;
  assign y3471 = n16028 ;
  assign y3472 = n16029 ;
  assign y3473 = ~n16036 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = ~n16039 ;
  assign y3476 = ~n16041 ;
  assign y3477 = n16042 ;
  assign y3478 = n16045 ;
  assign y3479 = n16048 ;
  assign y3480 = ~n16050 ;
  assign y3481 = ~n16053 ;
  assign y3482 = n16054 ;
  assign y3483 = n16055 ;
  assign y3484 = n16056 ;
  assign y3485 = n16062 ;
  assign y3486 = ~1'b0 ;
  assign y3487 = ~n16065 ;
  assign y3488 = ~n16068 ;
  assign y3489 = ~1'b0 ;
  assign y3490 = ~n16069 ;
  assign y3491 = n16078 ;
  assign y3492 = n16080 ;
  assign y3493 = ~n16081 ;
  assign y3494 = ~n16087 ;
  assign y3495 = ~n16088 ;
  assign y3496 = ~n16096 ;
  assign y3497 = n16103 ;
  assign y3498 = n16111 ;
  assign y3499 = ~n16112 ;
  assign y3500 = ~n16117 ;
  assign y3501 = ~n16122 ;
  assign y3502 = n16125 ;
  assign y3503 = n16128 ;
  assign y3504 = n16130 ;
  assign y3505 = n16131 ;
  assign y3506 = n16136 ;
  assign y3507 = ~n16137 ;
  assign y3508 = n16140 ;
  assign y3509 = ~n16143 ;
  assign y3510 = n16149 ;
  assign y3511 = ~n16153 ;
  assign y3512 = ~n16160 ;
  assign y3513 = ~n16161 ;
  assign y3514 = ~n16175 ;
  assign y3515 = n16177 ;
  assign y3516 = n16178 ;
  assign y3517 = ~1'b0 ;
  assign y3518 = n16179 ;
  assign y3519 = ~n16180 ;
  assign y3520 = ~n16188 ;
  assign y3521 = ~n16190 ;
  assign y3522 = n16198 ;
  assign y3523 = ~n16200 ;
  assign y3524 = n16201 ;
  assign y3525 = ~n16203 ;
  assign y3526 = n16205 ;
  assign y3527 = n16208 ;
  assign y3528 = ~n16211 ;
  assign y3529 = n16219 ;
  assign y3530 = n16220 ;
  assign y3531 = ~n16221 ;
  assign y3532 = ~n16223 ;
  assign y3533 = n16225 ;
  assign y3534 = n16231 ;
  assign y3535 = ~n16240 ;
  assign y3536 = ~n16242 ;
  assign y3537 = ~n16244 ;
  assign y3538 = ~n16246 ;
  assign y3539 = ~n16253 ;
  assign y3540 = n16255 ;
  assign y3541 = n16257 ;
  assign y3542 = ~n16259 ;
  assign y3543 = ~n16262 ;
  assign y3544 = n16264 ;
  assign y3545 = ~n16268 ;
  assign y3546 = ~n16272 ;
  assign y3547 = n16274 ;
  assign y3548 = n16276 ;
  assign y3549 = ~1'b0 ;
  assign y3550 = ~n16279 ;
  assign y3551 = n16292 ;
  assign y3552 = ~1'b0 ;
  assign y3553 = ~1'b0 ;
  assign y3554 = ~n16298 ;
  assign y3555 = n16304 ;
  assign y3556 = n16311 ;
  assign y3557 = ~n16315 ;
  assign y3558 = n16317 ;
  assign y3559 = ~n16323 ;
  assign y3560 = ~n15612 ;
  assign y3561 = n16324 ;
  assign y3562 = n16331 ;
  assign y3563 = ~n16333 ;
  assign y3564 = ~n16337 ;
  assign y3565 = n16339 ;
  assign y3566 = n16343 ;
  assign y3567 = ~n16345 ;
  assign y3568 = ~n16351 ;
  assign y3569 = n16366 ;
  assign y3570 = ~n16370 ;
  assign y3571 = n16372 ;
  assign y3572 = ~n16376 ;
  assign y3573 = ~n16379 ;
  assign y3574 = ~n16385 ;
  assign y3575 = ~n16396 ;
  assign y3576 = n16401 ;
  assign y3577 = n16403 ;
  assign y3578 = ~1'b0 ;
  assign y3579 = ~n16406 ;
  assign y3580 = ~n16407 ;
  assign y3581 = ~n16412 ;
  assign y3582 = n16413 ;
  assign y3583 = ~n16418 ;
  assign y3584 = ~n16421 ;
  assign y3585 = n16430 ;
  assign y3586 = ~1'b0 ;
  assign y3587 = ~n16433 ;
  assign y3588 = n16437 ;
  assign y3589 = n16438 ;
  assign y3590 = n12331 ;
  assign y3591 = ~n16448 ;
  assign y3592 = ~n16453 ;
  assign y3593 = ~1'b0 ;
  assign y3594 = ~n16457 ;
  assign y3595 = n16465 ;
  assign y3596 = n16468 ;
  assign y3597 = n16469 ;
  assign y3598 = ~n16480 ;
  assign y3599 = ~n16484 ;
  assign y3600 = n16487 ;
  assign y3601 = ~n16488 ;
  assign y3602 = n16489 ;
  assign y3603 = ~n16490 ;
  assign y3604 = n16491 ;
  assign y3605 = ~n16494 ;
  assign y3606 = ~n16496 ;
  assign y3607 = ~n16498 ;
  assign y3608 = n16503 ;
  assign y3609 = ~n16504 ;
  assign y3610 = n16510 ;
  assign y3611 = n16515 ;
  assign y3612 = ~n16519 ;
  assign y3613 = ~n16522 ;
  assign y3614 = ~n16523 ;
  assign y3615 = ~1'b0 ;
  assign y3616 = n16528 ;
  assign y3617 = n16529 ;
  assign y3618 = ~n16533 ;
  assign y3619 = n16539 ;
  assign y3620 = ~n16543 ;
  assign y3621 = n16546 ;
  assign y3622 = n16547 ;
  assign y3623 = ~n16556 ;
  assign y3624 = ~n16562 ;
  assign y3625 = ~n16568 ;
  assign y3626 = n16572 ;
  assign y3627 = n16577 ;
  assign y3628 = ~n16579 ;
  assign y3629 = n16590 ;
  assign y3630 = n16594 ;
  assign y3631 = ~n16600 ;
  assign y3632 = n16604 ;
  assign y3633 = n16612 ;
  assign y3634 = ~1'b0 ;
  assign y3635 = ~1'b0 ;
  assign y3636 = n16615 ;
  assign y3637 = n16616 ;
  assign y3638 = ~n16621 ;
  assign y3639 = n16622 ;
  assign y3640 = ~1'b0 ;
  assign y3641 = ~n16624 ;
  assign y3642 = n16625 ;
  assign y3643 = n16629 ;
  assign y3644 = n16633 ;
  assign y3645 = n16637 ;
  assign y3646 = n16639 ;
  assign y3647 = n16641 ;
  assign y3648 = ~n16643 ;
  assign y3649 = n16646 ;
  assign y3650 = n16650 ;
  assign y3651 = ~n16653 ;
  assign y3652 = ~n16658 ;
  assign y3653 = ~n16662 ;
  assign y3654 = n16667 ;
  assign y3655 = n16673 ;
  assign y3656 = ~n16677 ;
  assign y3657 = n16678 ;
  assign y3658 = ~n16681 ;
  assign y3659 = n16687 ;
  assign y3660 = ~n16690 ;
  assign y3661 = ~1'b0 ;
  assign y3662 = n16695 ;
  assign y3663 = ~n16698 ;
  assign y3664 = ~n16699 ;
  assign y3665 = n16700 ;
  assign y3666 = n16703 ;
  assign y3667 = ~1'b0 ;
  assign y3668 = n16705 ;
  assign y3669 = n16707 ;
  assign y3670 = n16716 ;
  assign y3671 = ~n16718 ;
  assign y3672 = ~n16720 ;
  assign y3673 = ~n16725 ;
  assign y3674 = ~n16728 ;
  assign y3675 = n16731 ;
  assign y3676 = n16734 ;
  assign y3677 = n16735 ;
  assign y3678 = ~n16740 ;
  assign y3679 = ~1'b0 ;
  assign y3680 = n16744 ;
  assign y3681 = ~n16750 ;
  assign y3682 = ~n16753 ;
  assign y3683 = ~n16755 ;
  assign y3684 = n16756 ;
  assign y3685 = ~n16757 ;
  assign y3686 = n16759 ;
  assign y3687 = ~n16761 ;
  assign y3688 = ~n16764 ;
  assign y3689 = ~n16769 ;
  assign y3690 = n16773 ;
  assign y3691 = n16774 ;
  assign y3692 = n16781 ;
  assign y3693 = ~n16789 ;
  assign y3694 = ~n16794 ;
  assign y3695 = n16797 ;
  assign y3696 = n16809 ;
  assign y3697 = ~n16812 ;
  assign y3698 = ~n16815 ;
  assign y3699 = ~n16825 ;
  assign y3700 = n16829 ;
  assign y3701 = n16832 ;
  assign y3702 = n16837 ;
  assign y3703 = n16845 ;
  assign y3704 = ~n16846 ;
  assign y3705 = n16848 ;
  assign y3706 = n16850 ;
  assign y3707 = n16851 ;
  assign y3708 = n16854 ;
  assign y3709 = ~n16856 ;
  assign y3710 = n16861 ;
  assign y3711 = n16864 ;
  assign y3712 = ~1'b0 ;
  assign y3713 = n16866 ;
  assign y3714 = n16869 ;
  assign y3715 = ~n16877 ;
  assign y3716 = ~n16878 ;
  assign y3717 = ~1'b0 ;
  assign y3718 = n16879 ;
  assign y3719 = n16880 ;
  assign y3720 = ~n16882 ;
  assign y3721 = n16887 ;
  assign y3722 = ~n16890 ;
  assign y3723 = n16891 ;
  assign y3724 = ~n16894 ;
  assign y3725 = n16895 ;
  assign y3726 = ~n16901 ;
  assign y3727 = n16905 ;
  assign y3728 = n16907 ;
  assign y3729 = n16908 ;
  assign y3730 = ~n16918 ;
  assign y3731 = n16920 ;
  assign y3732 = ~n16922 ;
  assign y3733 = ~n16925 ;
  assign y3734 = ~n16929 ;
  assign y3735 = ~n16932 ;
  assign y3736 = ~1'b0 ;
  assign y3737 = ~n16933 ;
  assign y3738 = ~n16934 ;
  assign y3739 = ~n16940 ;
  assign y3740 = n16946 ;
  assign y3741 = n16950 ;
  assign y3742 = n16957 ;
  assign y3743 = ~n16960 ;
  assign y3744 = n16964 ;
  assign y3745 = ~n16968 ;
  assign y3746 = n16972 ;
  assign y3747 = ~n16973 ;
  assign y3748 = n16974 ;
  assign y3749 = ~n16978 ;
  assign y3750 = n16981 ;
  assign y3751 = n16984 ;
  assign y3752 = n16986 ;
  assign y3753 = ~n16989 ;
  assign y3754 = ~n16992 ;
  assign y3755 = ~n16996 ;
  assign y3756 = ~n17001 ;
  assign y3757 = ~n17003 ;
  assign y3758 = n17004 ;
  assign y3759 = ~n17008 ;
  assign y3760 = n17009 ;
  assign y3761 = ~n17014 ;
  assign y3762 = ~n17018 ;
  assign y3763 = ~n17019 ;
  assign y3764 = n17021 ;
  assign y3765 = ~1'b0 ;
  assign y3766 = ~n17030 ;
  assign y3767 = n17033 ;
  assign y3768 = ~n17035 ;
  assign y3769 = n17037 ;
  assign y3770 = n17040 ;
  assign y3771 = ~n17043 ;
  assign y3772 = ~1'b0 ;
  assign y3773 = n17045 ;
  assign y3774 = ~n17053 ;
  assign y3775 = n17055 ;
  assign y3776 = n17056 ;
  assign y3777 = ~n17062 ;
  assign y3778 = ~n17064 ;
  assign y3779 = ~n17066 ;
  assign y3780 = n17067 ;
  assign y3781 = n17073 ;
  assign y3782 = ~n17076 ;
  assign y3783 = ~n17079 ;
  assign y3784 = n17083 ;
  assign y3785 = ~1'b0 ;
  assign y3786 = ~1'b0 ;
  assign y3787 = ~1'b0 ;
  assign y3788 = n17087 ;
  assign y3789 = n17088 ;
  assign y3790 = ~n17089 ;
  assign y3791 = n17092 ;
  assign y3792 = ~1'b0 ;
  assign y3793 = ~1'b0 ;
  assign y3794 = n17097 ;
  assign y3795 = ~n17102 ;
  assign y3796 = ~n17103 ;
  assign y3797 = ~n17104 ;
  assign y3798 = n17106 ;
  assign y3799 = ~n17111 ;
  assign y3800 = ~n17113 ;
  assign y3801 = n17117 ;
  assign y3802 = n17119 ;
  assign y3803 = n17124 ;
  assign y3804 = ~n17125 ;
  assign y3805 = ~n17135 ;
  assign y3806 = ~n17146 ;
  assign y3807 = ~n17151 ;
  assign y3808 = ~n17155 ;
  assign y3809 = ~1'b0 ;
  assign y3810 = ~n17160 ;
  assign y3811 = ~1'b0 ;
  assign y3812 = n17161 ;
  assign y3813 = ~n17170 ;
  assign y3814 = n17172 ;
  assign y3815 = ~n17179 ;
  assign y3816 = ~n17183 ;
  assign y3817 = ~n17185 ;
  assign y3818 = n17188 ;
  assign y3819 = ~1'b0 ;
  assign y3820 = n17192 ;
  assign y3821 = ~n17196 ;
  assign y3822 = n17203 ;
  assign y3823 = ~n17205 ;
  assign y3824 = n17223 ;
  assign y3825 = n17225 ;
  assign y3826 = ~n17228 ;
  assign y3827 = ~n17239 ;
  assign y3828 = ~n17241 ;
  assign y3829 = n17247 ;
  assign y3830 = n17251 ;
  assign y3831 = n17253 ;
  assign y3832 = ~1'b0 ;
  assign y3833 = ~n17255 ;
  assign y3834 = ~1'b0 ;
  assign y3835 = n17257 ;
  assign y3836 = n17258 ;
  assign y3837 = ~n17266 ;
  assign y3838 = ~n17268 ;
  assign y3839 = ~n17269 ;
  assign y3840 = ~n17274 ;
  assign y3841 = n17276 ;
  assign y3842 = ~n17280 ;
  assign y3843 = n17282 ;
  assign y3844 = ~n17283 ;
  assign y3845 = ~n17285 ;
  assign y3846 = ~1'b0 ;
  assign y3847 = ~n17289 ;
  assign y3848 = ~n17290 ;
  assign y3849 = ~n17293 ;
  assign y3850 = ~n17299 ;
  assign y3851 = n17304 ;
  assign y3852 = n17307 ;
  assign y3853 = ~n17315 ;
  assign y3854 = ~n17320 ;
  assign y3855 = ~n17324 ;
  assign y3856 = ~n17327 ;
  assign y3857 = n17331 ;
  assign y3858 = n17335 ;
  assign y3859 = ~n17339 ;
  assign y3860 = ~n17340 ;
  assign y3861 = n17342 ;
  assign y3862 = ~n17343 ;
  assign y3863 = ~n17344 ;
  assign y3864 = ~n17346 ;
  assign y3865 = ~n17348 ;
  assign y3866 = ~n17356 ;
  assign y3867 = n17358 ;
  assign y3868 = n17360 ;
  assign y3869 = n17369 ;
  assign y3870 = n17370 ;
  assign y3871 = n17380 ;
  assign y3872 = ~n17381 ;
  assign y3873 = ~n17384 ;
  assign y3874 = n17385 ;
  assign y3875 = n17394 ;
  assign y3876 = ~n17399 ;
  assign y3877 = ~n17402 ;
  assign y3878 = n17421 ;
  assign y3879 = ~1'b0 ;
  assign y3880 = ~1'b0 ;
  assign y3881 = ~n17425 ;
  assign y3882 = ~n17426 ;
  assign y3883 = n17429 ;
  assign y3884 = ~n17436 ;
  assign y3885 = ~n17440 ;
  assign y3886 = ~n17441 ;
  assign y3887 = n17445 ;
  assign y3888 = n17449 ;
  assign y3889 = ~n17453 ;
  assign y3890 = n17456 ;
  assign y3891 = n17458 ;
  assign y3892 = ~1'b0 ;
  assign y3893 = ~n17464 ;
  assign y3894 = ~n17466 ;
  assign y3895 = ~n17472 ;
  assign y3896 = ~n17475 ;
  assign y3897 = ~n17476 ;
  assign y3898 = n17477 ;
  assign y3899 = ~n17482 ;
  assign y3900 = n17484 ;
  assign y3901 = ~n17490 ;
  assign y3902 = ~1'b0 ;
  assign y3903 = ~n17493 ;
  assign y3904 = ~n17497 ;
  assign y3905 = n17501 ;
  assign y3906 = n17502 ;
  assign y3907 = ~n17507 ;
  assign y3908 = n17510 ;
  assign y3909 = n17514 ;
  assign y3910 = ~n17516 ;
  assign y3911 = ~n17518 ;
  assign y3912 = n17521 ;
  assign y3913 = ~n17522 ;
  assign y3914 = n17523 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = n17531 ;
  assign y3917 = ~n17536 ;
  assign y3918 = ~n17538 ;
  assign y3919 = ~n17542 ;
  assign y3920 = ~n17543 ;
  assign y3921 = ~n17545 ;
  assign y3922 = ~n17547 ;
  assign y3923 = n17550 ;
  assign y3924 = n17552 ;
  assign y3925 = ~n17555 ;
  assign y3926 = n17559 ;
  assign y3927 = ~n17562 ;
  assign y3928 = ~1'b0 ;
  assign y3929 = n17564 ;
  assign y3930 = n17565 ;
  assign y3931 = ~n17566 ;
  assign y3932 = n17567 ;
  assign y3933 = ~n17568 ;
  assign y3934 = n17571 ;
  assign y3935 = n17573 ;
  assign y3936 = n17575 ;
  assign y3937 = ~n17578 ;
  assign y3938 = n17583 ;
  assign y3939 = ~n17584 ;
  assign y3940 = ~n17585 ;
  assign y3941 = n17590 ;
  assign y3942 = n17596 ;
  assign y3943 = n17597 ;
  assign y3944 = n17602 ;
  assign y3945 = n17606 ;
  assign y3946 = n17607 ;
  assign y3947 = n17610 ;
  assign y3948 = n17614 ;
  assign y3949 = n17617 ;
  assign y3950 = n17619 ;
  assign y3951 = n17620 ;
  assign y3952 = ~n17623 ;
  assign y3953 = n17624 ;
  assign y3954 = n17625 ;
  assign y3955 = ~n17627 ;
  assign y3956 = n17629 ;
  assign y3957 = ~n17633 ;
  assign y3958 = n17637 ;
  assign y3959 = ~1'b0 ;
  assign y3960 = n17638 ;
  assign y3961 = ~n17643 ;
  assign y3962 = ~n17649 ;
  assign y3963 = n17656 ;
  assign y3964 = n17658 ;
  assign y3965 = n17664 ;
  assign y3966 = ~n17665 ;
  assign y3967 = n17666 ;
  assign y3968 = n17671 ;
  assign y3969 = ~n17673 ;
  assign y3970 = n17679 ;
  assign y3971 = n17684 ;
  assign y3972 = ~n17685 ;
  assign y3973 = ~1'b0 ;
  assign y3974 = n17686 ;
  assign y3975 = ~n17689 ;
  assign y3976 = n17691 ;
  assign y3977 = n17692 ;
  assign y3978 = n17694 ;
  assign y3979 = ~n17697 ;
  assign y3980 = n17701 ;
  assign y3981 = n17707 ;
  assign y3982 = ~1'b0 ;
  assign y3983 = n17717 ;
  assign y3984 = ~n17718 ;
  assign y3985 = ~n17726 ;
  assign y3986 = ~1'b0 ;
  assign y3987 = n17727 ;
  assign y3988 = ~n17734 ;
  assign y3989 = ~n17737 ;
  assign y3990 = ~n17746 ;
  assign y3991 = ~n17750 ;
  assign y3992 = ~n17754 ;
  assign y3993 = ~n17760 ;
  assign y3994 = n17767 ;
  assign y3995 = n17768 ;
  assign y3996 = ~1'b0 ;
  assign y3997 = ~n17770 ;
  assign y3998 = ~1'b0 ;
  assign y3999 = n17773 ;
  assign y4000 = n17776 ;
  assign y4001 = ~n17783 ;
  assign y4002 = ~n17787 ;
  assign y4003 = n17794 ;
  assign y4004 = n17796 ;
  assign y4005 = ~n17798 ;
  assign y4006 = n17803 ;
  assign y4007 = ~1'b0 ;
  assign y4008 = n17808 ;
  assign y4009 = ~n17815 ;
  assign y4010 = n17823 ;
  assign y4011 = n17826 ;
  assign y4012 = ~n17829 ;
  assign y4013 = n17836 ;
  assign y4014 = n17839 ;
  assign y4015 = ~n17841 ;
  assign y4016 = n17842 ;
  assign y4017 = ~n17843 ;
  assign y4018 = ~n17856 ;
  assign y4019 = n17859 ;
  assign y4020 = ~1'b0 ;
  assign y4021 = ~n17860 ;
  assign y4022 = n17861 ;
  assign y4023 = n17863 ;
  assign y4024 = ~n17866 ;
  assign y4025 = ~1'b0 ;
  assign y4026 = ~n17868 ;
  assign y4027 = ~n17870 ;
  assign y4028 = ~n17871 ;
  assign y4029 = ~n17873 ;
  assign y4030 = n17874 ;
  assign y4031 = n17881 ;
  assign y4032 = n17882 ;
  assign y4033 = ~n17893 ;
  assign y4034 = ~n17895 ;
  assign y4035 = n17902 ;
  assign y4036 = n17903 ;
  assign y4037 = n17905 ;
  assign y4038 = ~1'b0 ;
  assign y4039 = n17907 ;
  assign y4040 = ~n17910 ;
  assign y4041 = ~n17919 ;
  assign y4042 = n15456 ;
  assign y4043 = ~n17925 ;
  assign y4044 = ~n17926 ;
  assign y4045 = ~n17929 ;
  assign y4046 = ~n17931 ;
  assign y4047 = ~1'b0 ;
  assign y4048 = n17932 ;
  assign y4049 = ~n17935 ;
  assign y4050 = ~n17939 ;
  assign y4051 = n17940 ;
  assign y4052 = n17942 ;
  assign y4053 = n17946 ;
  assign y4054 = ~n17949 ;
  assign y4055 = n17952 ;
  assign y4056 = ~n17959 ;
  assign y4057 = n17962 ;
  assign y4058 = ~n17964 ;
  assign y4059 = ~n17968 ;
  assign y4060 = ~n17970 ;
  assign y4061 = ~n17971 ;
  assign y4062 = ~n17972 ;
  assign y4063 = ~n17974 ;
  assign y4064 = n17975 ;
  assign y4065 = n17977 ;
  assign y4066 = n17979 ;
  assign y4067 = ~n17983 ;
  assign y4068 = n17985 ;
  assign y4069 = n17987 ;
  assign y4070 = ~n17990 ;
  assign y4071 = n17996 ;
  assign y4072 = ~n17997 ;
  assign y4073 = ~n18004 ;
  assign y4074 = n18010 ;
  assign y4075 = ~n18011 ;
  assign y4076 = ~n18012 ;
  assign y4077 = n18016 ;
  assign y4078 = n18017 ;
  assign y4079 = n18025 ;
  assign y4080 = n18026 ;
  assign y4081 = n18028 ;
  assign y4082 = n18029 ;
  assign y4083 = ~n18035 ;
  assign y4084 = ~n18038 ;
  assign y4085 = ~n18042 ;
  assign y4086 = n18047 ;
  assign y4087 = ~n18049 ;
  assign y4088 = n18051 ;
  assign y4089 = n18055 ;
  assign y4090 = ~1'b0 ;
  assign y4091 = n18059 ;
  assign y4092 = ~n18060 ;
  assign y4093 = ~n14468 ;
  assign y4094 = ~1'b0 ;
  assign y4095 = n18061 ;
  assign y4096 = ~n18073 ;
  assign y4097 = ~n18081 ;
  assign y4098 = ~n18088 ;
  assign y4099 = ~n18089 ;
  assign y4100 = ~1'b0 ;
  assign y4101 = ~n18091 ;
  assign y4102 = ~n18093 ;
  assign y4103 = ~n18101 ;
  assign y4104 = n18104 ;
  assign y4105 = n18110 ;
  assign y4106 = n18112 ;
  assign y4107 = ~n18113 ;
  assign y4108 = n18114 ;
  assign y4109 = ~n18115 ;
  assign y4110 = ~n18120 ;
  assign y4111 = ~n18122 ;
  assign y4112 = n18131 ;
  assign y4113 = n18133 ;
  assign y4114 = n18137 ;
  assign y4115 = n18141 ;
  assign y4116 = n18143 ;
  assign y4117 = ~n18145 ;
  assign y4118 = ~n18146 ;
  assign y4119 = n18150 ;
  assign y4120 = ~n18156 ;
  assign y4121 = n18161 ;
  assign y4122 = n18162 ;
  assign y4123 = ~1'b0 ;
  assign y4124 = ~n18170 ;
  assign y4125 = n18175 ;
  assign y4126 = n18176 ;
  assign y4127 = n18180 ;
  assign y4128 = n18182 ;
  assign y4129 = ~n18187 ;
  assign y4130 = ~n18188 ;
  assign y4131 = ~n18189 ;
  assign y4132 = ~n18191 ;
  assign y4133 = ~n18193 ;
  assign y4134 = n18201 ;
  assign y4135 = ~1'b0 ;
  assign y4136 = ~n18202 ;
  assign y4137 = ~n18215 ;
  assign y4138 = n18226 ;
  assign y4139 = n18227 ;
  assign y4140 = n18228 ;
  assign y4141 = ~n18233 ;
  assign y4142 = ~1'b0 ;
  assign y4143 = n18237 ;
  assign y4144 = ~n18241 ;
  assign y4145 = ~n18242 ;
  assign y4146 = n18245 ;
  assign y4147 = n18246 ;
  assign y4148 = ~1'b0 ;
  assign y4149 = ~n18251 ;
  assign y4150 = n18257 ;
  assign y4151 = ~n18261 ;
  assign y4152 = n18265 ;
  assign y4153 = n18269 ;
  assign y4154 = ~1'b0 ;
  assign y4155 = n18277 ;
  assign y4156 = ~n18284 ;
  assign y4157 = ~n18285 ;
  assign y4158 = ~n18286 ;
  assign y4159 = ~n18287 ;
  assign y4160 = n18289 ;
  assign y4161 = n18291 ;
  assign y4162 = ~n18294 ;
  assign y4163 = 1'b0 ;
  assign y4164 = ~1'b0 ;
  assign y4165 = n18300 ;
  assign y4166 = n18302 ;
  assign y4167 = n18305 ;
  assign y4168 = ~n18309 ;
  assign y4169 = ~n18313 ;
  assign y4170 = ~n18315 ;
  assign y4171 = n18320 ;
  assign y4172 = n18321 ;
  assign y4173 = n18322 ;
  assign y4174 = ~n18324 ;
  assign y4175 = ~n18332 ;
  assign y4176 = n18333 ;
  assign y4177 = n18341 ;
  assign y4178 = ~n18343 ;
  assign y4179 = n18356 ;
  assign y4180 = ~n18360 ;
  assign y4181 = n18361 ;
  assign y4182 = ~n18364 ;
  assign y4183 = ~n18369 ;
  assign y4184 = n18378 ;
  assign y4185 = n18382 ;
  assign y4186 = ~n5953 ;
  assign y4187 = n18385 ;
  assign y4188 = ~n18389 ;
  assign y4189 = n18392 ;
  assign y4190 = n18395 ;
  assign y4191 = ~n18409 ;
  assign y4192 = ~n18410 ;
  assign y4193 = ~n18415 ;
  assign y4194 = ~n18417 ;
  assign y4195 = n18420 ;
  assign y4196 = n18421 ;
  assign y4197 = n18428 ;
  assign y4198 = n18430 ;
  assign y4199 = n18431 ;
  assign y4200 = n18434 ;
  assign y4201 = n18439 ;
  assign y4202 = ~1'b0 ;
  assign y4203 = ~n18441 ;
  assign y4204 = n18442 ;
  assign y4205 = n18445 ;
  assign y4206 = n18453 ;
  assign y4207 = ~n18457 ;
  assign y4208 = n18461 ;
  assign y4209 = n18465 ;
  assign y4210 = n18471 ;
  assign y4211 = n18473 ;
  assign y4212 = ~n18474 ;
  assign y4213 = n18476 ;
  assign y4214 = n18477 ;
  assign y4215 = n18478 ;
  assign y4216 = ~n18481 ;
  assign y4217 = ~n18488 ;
  assign y4218 = ~n18493 ;
  assign y4219 = ~n18496 ;
  assign y4220 = ~n18498 ;
  assign y4221 = ~n18504 ;
  assign y4222 = n18505 ;
  assign y4223 = ~n18508 ;
  assign y4224 = ~n18512 ;
  assign y4225 = ~n18516 ;
  assign y4226 = n18518 ;
  assign y4227 = ~n18519 ;
  assign y4228 = ~n18520 ;
  assign y4229 = n18522 ;
  assign y4230 = ~n18524 ;
  assign y4231 = n18525 ;
  assign y4232 = n18532 ;
  assign y4233 = n18533 ;
  assign y4234 = ~1'b0 ;
  assign y4235 = n18538 ;
  assign y4236 = n18542 ;
  assign y4237 = ~n18543 ;
  assign y4238 = n18551 ;
  assign y4239 = n18552 ;
  assign y4240 = ~n18562 ;
  assign y4241 = ~n18565 ;
  assign y4242 = ~n18567 ;
  assign y4243 = ~n18570 ;
  assign y4244 = n18575 ;
  assign y4245 = ~n18578 ;
  assign y4246 = ~n18580 ;
  assign y4247 = n18583 ;
  assign y4248 = n18592 ;
  assign y4249 = n18593 ;
  assign y4250 = ~n18594 ;
  assign y4251 = ~n18598 ;
  assign y4252 = ~n18604 ;
  assign y4253 = n18605 ;
  assign y4254 = n18615 ;
  assign y4255 = n18620 ;
  assign y4256 = ~1'b0 ;
  assign y4257 = ~1'b0 ;
  assign y4258 = ~1'b0 ;
  assign y4259 = n18627 ;
  assign y4260 = ~n18630 ;
  assign y4261 = n18632 ;
  assign y4262 = ~n18635 ;
  assign y4263 = ~n18639 ;
  assign y4264 = ~1'b0 ;
  assign y4265 = n18640 ;
  assign y4266 = ~n18644 ;
  assign y4267 = ~n18647 ;
  assign y4268 = n18648 ;
  assign y4269 = n18650 ;
  assign y4270 = n18651 ;
  assign y4271 = ~n18655 ;
  assign y4272 = n18658 ;
  assign y4273 = n18661 ;
  assign y4274 = n18662 ;
  assign y4275 = ~n18668 ;
  assign y4276 = n18679 ;
  assign y4277 = ~n18684 ;
  assign y4278 = n18687 ;
  assign y4279 = ~n18690 ;
  assign y4280 = n18692 ;
  assign y4281 = ~n18697 ;
  assign y4282 = ~n18699 ;
  assign y4283 = ~n18706 ;
  assign y4284 = n18709 ;
  assign y4285 = ~n18713 ;
  assign y4286 = n18716 ;
  assign y4287 = n18719 ;
  assign y4288 = n18725 ;
  assign y4289 = n18727 ;
  assign y4290 = ~n18731 ;
  assign y4291 = n18735 ;
  assign y4292 = ~n18738 ;
  assign y4293 = ~n18742 ;
  assign y4294 = n18745 ;
  assign y4295 = n18747 ;
  assign y4296 = n18749 ;
  assign y4297 = ~n18750 ;
  assign y4298 = n18753 ;
  assign y4299 = ~n18757 ;
  assign y4300 = ~1'b0 ;
  assign y4301 = ~n18761 ;
  assign y4302 = n18764 ;
  assign y4303 = n18767 ;
  assign y4304 = n18768 ;
  assign y4305 = n18775 ;
  assign y4306 = ~1'b0 ;
  assign y4307 = n18778 ;
  assign y4308 = ~n18780 ;
  assign y4309 = ~n18784 ;
  assign y4310 = ~n18788 ;
  assign y4311 = ~n18791 ;
  assign y4312 = n18793 ;
  assign y4313 = n18796 ;
  assign y4314 = n18807 ;
  assign y4315 = n18810 ;
  assign y4316 = n18812 ;
  assign y4317 = ~n18814 ;
  assign y4318 = ~n18820 ;
  assign y4319 = n18827 ;
  assign y4320 = n18831 ;
  assign y4321 = n18835 ;
  assign y4322 = n18841 ;
  assign y4323 = ~n18852 ;
  assign y4324 = ~n18856 ;
  assign y4325 = ~n18858 ;
  assign y4326 = ~n18862 ;
  assign y4327 = ~n18869 ;
  assign y4328 = ~n18872 ;
  assign y4329 = n18873 ;
  assign y4330 = n18874 ;
  assign y4331 = ~n18876 ;
  assign y4332 = ~n18880 ;
  assign y4333 = n18881 ;
  assign y4334 = n18883 ;
  assign y4335 = ~n18886 ;
  assign y4336 = ~n18891 ;
  assign y4337 = n18895 ;
  assign y4338 = ~n18899 ;
  assign y4339 = n18900 ;
  assign y4340 = n18908 ;
  assign y4341 = ~n18909 ;
  assign y4342 = ~n18910 ;
  assign y4343 = n18912 ;
  assign y4344 = n18913 ;
  assign y4345 = ~n18915 ;
  assign y4346 = ~n18918 ;
  assign y4347 = ~n18924 ;
  assign y4348 = ~n18925 ;
  assign y4349 = n18926 ;
  assign y4350 = ~n18931 ;
  assign y4351 = n18932 ;
  assign y4352 = n18933 ;
  assign y4353 = ~1'b0 ;
  assign y4354 = ~1'b0 ;
  assign y4355 = n18939 ;
  assign y4356 = ~n18942 ;
  assign y4357 = ~n18946 ;
  assign y4358 = n18947 ;
  assign y4359 = n18950 ;
  assign y4360 = n18952 ;
  assign y4361 = n18954 ;
  assign y4362 = ~n18957 ;
  assign y4363 = n18959 ;
  assign y4364 = ~n18961 ;
  assign y4365 = ~1'b0 ;
  assign y4366 = n18963 ;
  assign y4367 = n18964 ;
  assign y4368 = n18965 ;
  assign y4369 = ~n18966 ;
  assign y4370 = ~1'b0 ;
  assign y4371 = ~n18971 ;
  assign y4372 = n18974 ;
  assign y4373 = ~n18975 ;
  assign y4374 = n18980 ;
  assign y4375 = n18983 ;
  assign y4376 = ~n18985 ;
  assign y4377 = ~n18989 ;
  assign y4378 = n18991 ;
  assign y4379 = ~n18994 ;
  assign y4380 = ~n18996 ;
  assign y4381 = ~n19002 ;
  assign y4382 = n19004 ;
  assign y4383 = n19005 ;
  assign y4384 = ~n19006 ;
  assign y4385 = n19009 ;
  assign y4386 = n19011 ;
  assign y4387 = n19012 ;
  assign y4388 = n19023 ;
  assign y4389 = n19028 ;
  assign y4390 = n19031 ;
  assign y4391 = n19032 ;
  assign y4392 = ~n19033 ;
  assign y4393 = n19035 ;
  assign y4394 = n19037 ;
  assign y4395 = ~1'b0 ;
  assign y4396 = ~n19039 ;
  assign y4397 = ~n19041 ;
  assign y4398 = ~n19042 ;
  assign y4399 = n19043 ;
  assign y4400 = n19046 ;
  assign y4401 = ~1'b0 ;
  assign y4402 = ~n19049 ;
  assign y4403 = ~n19050 ;
  assign y4404 = ~n19053 ;
  assign y4405 = n19054 ;
  assign y4406 = n19057 ;
  assign y4407 = n19059 ;
  assign y4408 = ~n19071 ;
  assign y4409 = n19072 ;
  assign y4410 = ~n19076 ;
  assign y4411 = ~n19080 ;
  assign y4412 = n19082 ;
  assign y4413 = ~1'b0 ;
  assign y4414 = ~n19086 ;
  assign y4415 = n19089 ;
  assign y4416 = ~n19094 ;
  assign y4417 = n19096 ;
  assign y4418 = ~n19101 ;
  assign y4419 = n19103 ;
  assign y4420 = n19107 ;
  assign y4421 = ~n19110 ;
  assign y4422 = n19111 ;
  assign y4423 = n19113 ;
  assign y4424 = ~n19114 ;
  assign y4425 = ~n19115 ;
  assign y4426 = ~n19117 ;
  assign y4427 = n19119 ;
  assign y4428 = n19124 ;
  assign y4429 = n19129 ;
  assign y4430 = ~n19130 ;
  assign y4431 = n19131 ;
  assign y4432 = ~1'b0 ;
  assign y4433 = ~n19132 ;
  assign y4434 = ~n19135 ;
  assign y4435 = ~n19137 ;
  assign y4436 = n19139 ;
  assign y4437 = ~n19144 ;
  assign y4438 = ~n19148 ;
  assign y4439 = n19151 ;
  assign y4440 = ~n19153 ;
  assign y4441 = n19156 ;
  assign y4442 = ~n19169 ;
  assign y4443 = n19174 ;
  assign y4444 = ~n19176 ;
  assign y4445 = ~n19179 ;
  assign y4446 = ~n19185 ;
  assign y4447 = ~n19188 ;
  assign y4448 = ~n19191 ;
  assign y4449 = ~n19192 ;
  assign y4450 = ~1'b0 ;
  assign y4451 = ~n19196 ;
  assign y4452 = ~n19197 ;
  assign y4453 = n19203 ;
  assign y4454 = n19210 ;
  assign y4455 = ~1'b0 ;
  assign y4456 = ~1'b0 ;
  assign y4457 = ~1'b0 ;
  assign y4458 = n19219 ;
  assign y4459 = n19222 ;
  assign y4460 = n19224 ;
  assign y4461 = ~1'b0 ;
  assign y4462 = ~n19229 ;
  assign y4463 = n19233 ;
  assign y4464 = ~n19235 ;
  assign y4465 = ~n19242 ;
  assign y4466 = n19246 ;
  assign y4467 = n19257 ;
  assign y4468 = ~n19260 ;
  assign y4469 = ~n19261 ;
  assign y4470 = n19262 ;
  assign y4471 = ~n19268 ;
  assign y4472 = ~n19269 ;
  assign y4473 = n19272 ;
  assign y4474 = n19274 ;
  assign y4475 = n19280 ;
  assign y4476 = ~n19288 ;
  assign y4477 = n19291 ;
  assign y4478 = ~n19297 ;
  assign y4479 = ~n19299 ;
  assign y4480 = n19301 ;
  assign y4481 = ~n19303 ;
  assign y4482 = ~n19305 ;
  assign y4483 = n19306 ;
  assign y4484 = ~n19308 ;
  assign y4485 = ~n19309 ;
  assign y4486 = n19313 ;
  assign y4487 = ~n19315 ;
  assign y4488 = ~n19320 ;
  assign y4489 = n19327 ;
  assign y4490 = n19328 ;
  assign y4491 = 1'b0 ;
  assign y4492 = ~n19334 ;
  assign y4493 = n19335 ;
  assign y4494 = n19343 ;
  assign y4495 = ~1'b0 ;
  assign y4496 = n19345 ;
  assign y4497 = n19349 ;
  assign y4498 = ~n19350 ;
  assign y4499 = n19351 ;
  assign y4500 = ~n19358 ;
  assign y4501 = ~n19360 ;
  assign y4502 = ~n19362 ;
  assign y4503 = ~n19368 ;
  assign y4504 = ~1'b0 ;
  assign y4505 = ~n19372 ;
  assign y4506 = ~n19373 ;
  assign y4507 = n19378 ;
  assign y4508 = ~n19381 ;
  assign y4509 = n19384 ;
  assign y4510 = n19388 ;
  assign y4511 = ~n19395 ;
  assign y4512 = ~n19396 ;
  assign y4513 = n19398 ;
  assign y4514 = n19399 ;
  assign y4515 = ~n19404 ;
  assign y4516 = ~n19409 ;
  assign y4517 = n19414 ;
  assign y4518 = ~1'b0 ;
  assign y4519 = n19415 ;
  assign y4520 = n19419 ;
  assign y4521 = n19420 ;
  assign y4522 = ~n19422 ;
  assign y4523 = n19428 ;
  assign y4524 = n19431 ;
  assign y4525 = n19436 ;
  assign y4526 = ~n19438 ;
  assign y4527 = n19441 ;
  assign y4528 = ~n19445 ;
  assign y4529 = ~n19446 ;
  assign y4530 = ~n19447 ;
  assign y4531 = n19454 ;
  assign y4532 = n19462 ;
  assign y4533 = ~n19467 ;
  assign y4534 = ~n19469 ;
  assign y4535 = ~n19472 ;
  assign y4536 = n19473 ;
  assign y4537 = ~n19475 ;
  assign y4538 = ~n19479 ;
  assign y4539 = n19480 ;
  assign y4540 = n19483 ;
  assign y4541 = n19488 ;
  assign y4542 = n19489 ;
  assign y4543 = n19498 ;
  assign y4544 = ~n19500 ;
  assign y4545 = n19502 ;
  assign y4546 = ~n19503 ;
  assign y4547 = n19506 ;
  assign y4548 = ~n19509 ;
  assign y4549 = n19511 ;
  assign y4550 = ~1'b0 ;
  assign y4551 = n19514 ;
  assign y4552 = n19516 ;
  assign y4553 = n19520 ;
  assign y4554 = n19523 ;
  assign y4555 = ~n19528 ;
  assign y4556 = ~1'b0 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = n19529 ;
  assign y4559 = n19533 ;
  assign y4560 = ~n19534 ;
  assign y4561 = ~n19536 ;
  assign y4562 = n19538 ;
  assign y4563 = ~n19541 ;
  assign y4564 = ~n19543 ;
  assign y4565 = ~n19548 ;
  assign y4566 = ~n19550 ;
  assign y4567 = ~1'b0 ;
  assign y4568 = ~1'b0 ;
  assign y4569 = ~n19551 ;
  assign y4570 = ~n19558 ;
  assign y4571 = ~n19560 ;
  assign y4572 = ~n19564 ;
  assign y4573 = ~n19573 ;
  assign y4574 = ~n19575 ;
  assign y4575 = n19578 ;
  assign y4576 = ~n19579 ;
  assign y4577 = n19581 ;
  assign y4578 = n19585 ;
  assign y4579 = n19588 ;
  assign y4580 = ~n19589 ;
  assign y4581 = ~n8281 ;
  assign y4582 = ~n19592 ;
  assign y4583 = n19593 ;
  assign y4584 = ~n19594 ;
  assign y4585 = ~n19601 ;
  assign y4586 = ~n19602 ;
  assign y4587 = n19606 ;
  assign y4588 = n19607 ;
  assign y4589 = ~n19614 ;
  assign y4590 = n19617 ;
  assign y4591 = ~n19620 ;
  assign y4592 = n19626 ;
  assign y4593 = ~n19628 ;
  assign y4594 = ~n19630 ;
  assign y4595 = n19632 ;
  assign y4596 = ~n19633 ;
  assign y4597 = ~n19637 ;
  assign y4598 = n19640 ;
  assign y4599 = ~n19643 ;
  assign y4600 = ~1'b0 ;
  assign y4601 = n19644 ;
  assign y4602 = ~n19649 ;
  assign y4603 = ~n19652 ;
  assign y4604 = n19653 ;
  assign y4605 = ~n19663 ;
  assign y4606 = n19667 ;
  assign y4607 = ~n19669 ;
  assign y4608 = ~1'b0 ;
  assign y4609 = ~n19670 ;
  assign y4610 = n19673 ;
  assign y4611 = n19678 ;
  assign y4612 = n19679 ;
  assign y4613 = n19682 ;
  assign y4614 = ~1'b0 ;
  assign y4615 = ~n19687 ;
  assign y4616 = ~n19692 ;
  assign y4617 = ~n19696 ;
  assign y4618 = ~n19697 ;
  assign y4619 = ~n19710 ;
  assign y4620 = ~n19712 ;
  assign y4621 = ~n19716 ;
  assign y4622 = ~n19717 ;
  assign y4623 = ~n19720 ;
  assign y4624 = n19725 ;
  assign y4625 = n19730 ;
  assign y4626 = ~n19734 ;
  assign y4627 = ~n19741 ;
  assign y4628 = n19745 ;
  assign y4629 = n19746 ;
  assign y4630 = n19752 ;
  assign y4631 = n19753 ;
  assign y4632 = ~n19764 ;
  assign y4633 = ~n19765 ;
  assign y4634 = n19769 ;
  assign y4635 = ~n19772 ;
  assign y4636 = ~1'b0 ;
  assign y4637 = ~n19775 ;
  assign y4638 = n19781 ;
  assign y4639 = n19786 ;
  assign y4640 = ~n19791 ;
  assign y4641 = n19793 ;
  assign y4642 = ~n19802 ;
  assign y4643 = ~n19804 ;
  assign y4644 = n19807 ;
  assign y4645 = ~n19809 ;
  assign y4646 = ~n19810 ;
  assign y4647 = n19814 ;
  assign y4648 = ~n19815 ;
  assign y4649 = ~1'b0 ;
  assign y4650 = ~1'b0 ;
  assign y4651 = n19819 ;
  assign y4652 = n19821 ;
  assign y4653 = n19826 ;
  assign y4654 = n19827 ;
  assign y4655 = n19830 ;
  assign y4656 = ~n19833 ;
  assign y4657 = n19838 ;
  assign y4658 = ~1'b0 ;
  assign y4659 = ~1'b0 ;
  assign y4660 = n19840 ;
  assign y4661 = ~n19843 ;
  assign y4662 = n19844 ;
  assign y4663 = ~n19845 ;
  assign y4664 = ~n19847 ;
  assign y4665 = n19849 ;
  assign y4666 = n19856 ;
  assign y4667 = ~n19858 ;
  assign y4668 = n19864 ;
  assign y4669 = ~n19868 ;
  assign y4670 = n19871 ;
  assign y4671 = n19879 ;
  assign y4672 = n19880 ;
  assign y4673 = ~n19886 ;
  assign y4674 = ~n19892 ;
  assign y4675 = n19893 ;
  assign y4676 = ~n19905 ;
  assign y4677 = ~n19907 ;
  assign y4678 = ~1'b0 ;
  assign y4679 = n19909 ;
  assign y4680 = n19913 ;
  assign y4681 = ~n19914 ;
  assign y4682 = n19921 ;
  assign y4683 = ~n19927 ;
  assign y4684 = n19928 ;
  assign y4685 = ~n19929 ;
  assign y4686 = ~n19932 ;
  assign y4687 = n19934 ;
  assign y4688 = ~n19938 ;
  assign y4689 = n19942 ;
  assign y4690 = ~n19943 ;
  assign y4691 = n19944 ;
  assign y4692 = ~n19948 ;
  assign y4693 = n19950 ;
  assign y4694 = n19952 ;
  assign y4695 = n19955 ;
  assign y4696 = ~n19960 ;
  assign y4697 = n19961 ;
  assign y4698 = n19963 ;
  assign y4699 = n19967 ;
  assign y4700 = n19970 ;
  assign y4701 = ~n19971 ;
  assign y4702 = n19978 ;
  assign y4703 = n19979 ;
  assign y4704 = n19983 ;
  assign y4705 = ~n19988 ;
  assign y4706 = ~n19996 ;
  assign y4707 = n20000 ;
  assign y4708 = n20003 ;
  assign y4709 = n20005 ;
  assign y4710 = ~n20007 ;
  assign y4711 = n20009 ;
  assign y4712 = n20011 ;
  assign y4713 = n20012 ;
  assign y4714 = ~n20015 ;
  assign y4715 = n20019 ;
  assign y4716 = ~n20020 ;
  assign y4717 = n20022 ;
  assign y4718 = ~n20025 ;
  assign y4719 = n20026 ;
  assign y4720 = n20027 ;
  assign y4721 = n20032 ;
  assign y4722 = n20035 ;
  assign y4723 = n20038 ;
  assign y4724 = ~n20043 ;
  assign y4725 = ~n20047 ;
  assign y4726 = ~n20052 ;
  assign y4727 = n20059 ;
  assign y4728 = ~n20062 ;
  assign y4729 = n20063 ;
  assign y4730 = ~n20065 ;
  assign y4731 = ~n20071 ;
  assign y4732 = n20073 ;
  assign y4733 = ~n20077 ;
  assign y4734 = n20081 ;
  assign y4735 = ~n20083 ;
  assign y4736 = ~n20097 ;
  assign y4737 = n20100 ;
  assign y4738 = n20103 ;
  assign y4739 = ~n20106 ;
  assign y4740 = n20107 ;
  assign y4741 = n20109 ;
  assign y4742 = n20110 ;
  assign y4743 = ~n20114 ;
  assign y4744 = ~n20116 ;
  assign y4745 = n20119 ;
  assign y4746 = n20125 ;
  assign y4747 = ~n20129 ;
  assign y4748 = ~n20131 ;
  assign y4749 = n20133 ;
  assign y4750 = ~n20134 ;
  assign y4751 = ~n20137 ;
  assign y4752 = n20138 ;
  assign y4753 = n20139 ;
  assign y4754 = ~1'b0 ;
  assign y4755 = n20145 ;
  assign y4756 = ~n20146 ;
  assign y4757 = ~n20149 ;
  assign y4758 = ~n20151 ;
  assign y4759 = n20152 ;
  assign y4760 = ~n20153 ;
  assign y4761 = n20154 ;
  assign y4762 = n20156 ;
  assign y4763 = n20158 ;
  assign y4764 = n20161 ;
  assign y4765 = ~n20164 ;
  assign y4766 = ~n20168 ;
  assign y4767 = ~n20172 ;
  assign y4768 = n20181 ;
  assign y4769 = ~n20182 ;
  assign y4770 = n20183 ;
  assign y4771 = ~n20185 ;
  assign y4772 = ~n20190 ;
  assign y4773 = ~1'b0 ;
  assign y4774 = n20193 ;
  assign y4775 = ~n20199 ;
  assign y4776 = n20203 ;
  assign y4777 = n20206 ;
  assign y4778 = ~n20208 ;
  assign y4779 = n20213 ;
  assign y4780 = ~n20218 ;
  assign y4781 = ~n20222 ;
  assign y4782 = n20223 ;
  assign y4783 = ~1'b0 ;
  assign y4784 = n20229 ;
  assign y4785 = ~n20230 ;
  assign y4786 = ~n20232 ;
  assign y4787 = n20235 ;
  assign y4788 = n20240 ;
  assign y4789 = n20242 ;
  assign y4790 = n20247 ;
  assign y4791 = ~n20249 ;
  assign y4792 = ~n20254 ;
  assign y4793 = ~n20256 ;
  assign y4794 = n20259 ;
  assign y4795 = n20271 ;
  assign y4796 = ~n20276 ;
  assign y4797 = ~n20277 ;
  assign y4798 = n20281 ;
  assign y4799 = n20286 ;
  assign y4800 = n20288 ;
  assign y4801 = n20289 ;
  assign y4802 = ~n20290 ;
  assign y4803 = n20296 ;
  assign y4804 = n20298 ;
  assign y4805 = ~n20303 ;
  assign y4806 = ~n20305 ;
  assign y4807 = n20309 ;
  assign y4808 = n20310 ;
  assign y4809 = 1'b0 ;
  assign y4810 = n20315 ;
  assign y4811 = ~n20316 ;
  assign y4812 = n20317 ;
  assign y4813 = n20318 ;
  assign y4814 = n20320 ;
  assign y4815 = n20323 ;
  assign y4816 = n20324 ;
  assign y4817 = n20329 ;
  assign y4818 = ~n20331 ;
  assign y4819 = n20332 ;
  assign y4820 = ~n20334 ;
  assign y4821 = ~n20337 ;
  assign y4822 = n20339 ;
  assign y4823 = n20342 ;
  assign y4824 = n20347 ;
  assign y4825 = ~n20349 ;
  assign y4826 = n20354 ;
  assign y4827 = n20355 ;
  assign y4828 = n20357 ;
  assign y4829 = ~1'b0 ;
  assign y4830 = ~n20360 ;
  assign y4831 = n20362 ;
  assign y4832 = n20364 ;
  assign y4833 = n20367 ;
  assign y4834 = ~n20369 ;
  assign y4835 = n20370 ;
  assign y4836 = n20374 ;
  assign y4837 = ~n20377 ;
  assign y4838 = n20378 ;
  assign y4839 = n20382 ;
  assign y4840 = n20388 ;
  assign y4841 = n20390 ;
  assign y4842 = ~n20391 ;
  assign y4843 = ~n20395 ;
  assign y4844 = ~n20397 ;
  assign y4845 = ~n20398 ;
  assign y4846 = n20399 ;
  assign y4847 = ~n20403 ;
  assign y4848 = ~n20404 ;
  assign y4849 = ~1'b0 ;
  assign y4850 = n20407 ;
  assign y4851 = n20410 ;
  assign y4852 = n20412 ;
  assign y4853 = n20413 ;
  assign y4854 = ~n20421 ;
  assign y4855 = n20426 ;
  assign y4856 = ~n20427 ;
  assign y4857 = ~n20429 ;
  assign y4858 = n20431 ;
  assign y4859 = ~n20436 ;
  assign y4860 = ~n20439 ;
  assign y4861 = ~n20441 ;
  assign y4862 = n20447 ;
  assign y4863 = ~n20448 ;
  assign y4864 = n20450 ;
  assign y4865 = ~n20453 ;
  assign y4866 = n20454 ;
  assign y4867 = n20457 ;
  assign y4868 = n20458 ;
  assign y4869 = ~n20463 ;
  assign y4870 = ~1'b0 ;
  assign y4871 = ~n20464 ;
  assign y4872 = ~n20465 ;
  assign y4873 = ~1'b0 ;
  assign y4874 = n20471 ;
  assign y4875 = ~n20472 ;
  assign y4876 = ~n20474 ;
  assign y4877 = ~n20476 ;
  assign y4878 = ~n20479 ;
  assign y4879 = ~n20480 ;
  assign y4880 = n20482 ;
  assign y4881 = ~n20483 ;
  assign y4882 = ~n20486 ;
  assign y4883 = ~n20487 ;
  assign y4884 = ~1'b0 ;
  assign y4885 = ~n20489 ;
  assign y4886 = ~n20492 ;
  assign y4887 = ~n20495 ;
  assign y4888 = ~n20498 ;
  assign y4889 = ~n20501 ;
  assign y4890 = n20503 ;
  assign y4891 = n20513 ;
  assign y4892 = n20515 ;
  assign y4893 = n20521 ;
  assign y4894 = n20522 ;
  assign y4895 = ~n20525 ;
  assign y4896 = n20526 ;
  assign y4897 = n20528 ;
  assign y4898 = ~n20531 ;
  assign y4899 = n20533 ;
  assign y4900 = ~n20537 ;
  assign y4901 = n20538 ;
  assign y4902 = ~n20543 ;
  assign y4903 = ~n20544 ;
  assign y4904 = ~n20546 ;
  assign y4905 = ~n20551 ;
  assign y4906 = ~n20552 ;
  assign y4907 = n20556 ;
  assign y4908 = n20561 ;
  assign y4909 = ~n20563 ;
  assign y4910 = n20566 ;
  assign y4911 = ~n20570 ;
  assign y4912 = n20575 ;
  assign y4913 = n20577 ;
  assign y4914 = ~n20582 ;
  assign y4915 = ~n20586 ;
  assign y4916 = n20596 ;
  assign y4917 = ~1'b0 ;
  assign y4918 = ~n20600 ;
  assign y4919 = ~n20601 ;
  assign y4920 = ~n20604 ;
  assign y4921 = n20608 ;
  assign y4922 = ~n20610 ;
  assign y4923 = ~n20611 ;
  assign y4924 = ~n20613 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = n20618 ;
  assign y4927 = ~n20623 ;
  assign y4928 = n20628 ;
  assign y4929 = ~n20629 ;
  assign y4930 = ~1'b0 ;
  assign y4931 = ~n20634 ;
  assign y4932 = ~n20639 ;
  assign y4933 = n20640 ;
  assign y4934 = ~n20642 ;
  assign y4935 = ~n20645 ;
  assign y4936 = n20649 ;
  assign y4937 = ~1'b0 ;
  assign y4938 = n20650 ;
  assign y4939 = ~n20653 ;
  assign y4940 = n20658 ;
  assign y4941 = n20660 ;
  assign y4942 = ~n20661 ;
  assign y4943 = ~n20663 ;
  assign y4944 = n20664 ;
  assign y4945 = n20668 ;
  assign y4946 = ~n20670 ;
  assign y4947 = ~n20671 ;
  assign y4948 = ~n20675 ;
  assign y4949 = ~n20678 ;
  assign y4950 = ~n20679 ;
  assign y4951 = n20684 ;
  assign y4952 = ~n20686 ;
  assign y4953 = n20691 ;
  assign y4954 = n20694 ;
  assign y4955 = ~n20700 ;
  assign y4956 = n6544 ;
  assign y4957 = ~n20701 ;
  assign y4958 = n20702 ;
  assign y4959 = n20704 ;
  assign y4960 = ~n20709 ;
  assign y4961 = n20714 ;
  assign y4962 = ~n20723 ;
  assign y4963 = ~n20725 ;
  assign y4964 = ~n20727 ;
  assign y4965 = ~n20730 ;
  assign y4966 = ~n20734 ;
  assign y4967 = ~n20735 ;
  assign y4968 = n20737 ;
  assign y4969 = n20741 ;
  assign y4970 = n20748 ;
  assign y4971 = ~1'b0 ;
  assign y4972 = n20750 ;
  assign y4973 = ~n20752 ;
  assign y4974 = ~n20755 ;
  assign y4975 = n20757 ;
  assign y4976 = n20758 ;
  assign y4977 = n20761 ;
  assign y4978 = n20763 ;
  assign y4979 = ~n20765 ;
  assign y4980 = n20766 ;
  assign y4981 = ~n20771 ;
  assign y4982 = n20773 ;
  assign y4983 = n20778 ;
  assign y4984 = n20782 ;
  assign y4985 = n20791 ;
  assign y4986 = ~1'b0 ;
  assign y4987 = ~n20793 ;
  assign y4988 = ~n20799 ;
  assign y4989 = n20800 ;
  assign y4990 = n20801 ;
  assign y4991 = n20803 ;
  assign y4992 = ~n20806 ;
  assign y4993 = n20808 ;
  assign y4994 = n20811 ;
  assign y4995 = ~n20816 ;
  assign y4996 = n20819 ;
  assign y4997 = ~n20821 ;
  assign y4998 = n20824 ;
  assign y4999 = ~n20825 ;
  assign y5000 = ~n20830 ;
  assign y5001 = ~n20831 ;
  assign y5002 = n20832 ;
  assign y5003 = n20836 ;
  assign y5004 = ~n20837 ;
  assign y5005 = ~n20841 ;
  assign y5006 = n20842 ;
  assign y5007 = ~n20845 ;
  assign y5008 = ~1'b0 ;
  assign y5009 = ~n20847 ;
  assign y5010 = n20848 ;
  assign y5011 = n20851 ;
  assign y5012 = ~n20852 ;
  assign y5013 = ~1'b0 ;
  assign y5014 = ~n20854 ;
  assign y5015 = n20856 ;
  assign y5016 = ~n20857 ;
  assign y5017 = ~n20860 ;
  assign y5018 = n20867 ;
  assign y5019 = n20872 ;
  assign y5020 = ~n20877 ;
  assign y5021 = ~n20879 ;
  assign y5022 = ~n20881 ;
  assign y5023 = n20884 ;
  assign y5024 = ~n20886 ;
  assign y5025 = ~n20889 ;
  assign y5026 = ~n20891 ;
  assign y5027 = ~n20892 ;
  assign y5028 = n20895 ;
  assign y5029 = n20899 ;
  assign y5030 = ~n20901 ;
  assign y5031 = n20905 ;
  assign y5032 = ~n20908 ;
  assign y5033 = ~n20909 ;
  assign y5034 = ~n20914 ;
  assign y5035 = n20919 ;
  assign y5036 = n20920 ;
  assign y5037 = ~n20926 ;
  assign y5038 = n20928 ;
  assign y5039 = n20932 ;
  assign y5040 = n20939 ;
  assign y5041 = ~n20941 ;
  assign y5042 = ~n20942 ;
  assign y5043 = ~1'b0 ;
  assign y5044 = n20943 ;
  assign y5045 = ~n20953 ;
  assign y5046 = ~n20955 ;
  assign y5047 = n20960 ;
  assign y5048 = n20961 ;
  assign y5049 = n20966 ;
  assign y5050 = ~1'b0 ;
  assign y5051 = n20968 ;
  assign y5052 = ~n20970 ;
  assign y5053 = ~n20974 ;
  assign y5054 = n20975 ;
  assign y5055 = n20976 ;
  assign y5056 = ~n20978 ;
  assign y5057 = ~n20982 ;
  assign y5058 = ~n20992 ;
  assign y5059 = ~n20999 ;
  assign y5060 = n21006 ;
  assign y5061 = ~n21007 ;
  assign y5062 = ~n21010 ;
  assign y5063 = n21011 ;
  assign y5064 = n21013 ;
  assign y5065 = ~n21014 ;
  assign y5066 = ~n21015 ;
  assign y5067 = ~n21017 ;
  assign y5068 = ~n21027 ;
  assign y5069 = ~1'b0 ;
  assign y5070 = n21030 ;
  assign y5071 = n21032 ;
  assign y5072 = n21034 ;
  assign y5073 = n21038 ;
  assign y5074 = n21040 ;
  assign y5075 = n21042 ;
  assign y5076 = ~1'b0 ;
  assign y5077 = ~n21044 ;
  assign y5078 = ~n21045 ;
  assign y5079 = ~n21046 ;
  assign y5080 = ~n21047 ;
  assign y5081 = ~n21051 ;
  assign y5082 = n21061 ;
  assign y5083 = ~n21062 ;
  assign y5084 = ~n21066 ;
  assign y5085 = ~n21068 ;
  assign y5086 = ~n21071 ;
  assign y5087 = ~1'b0 ;
  assign y5088 = n21073 ;
  assign y5089 = n21074 ;
  assign y5090 = ~n21075 ;
  assign y5091 = ~n21081 ;
  assign y5092 = ~1'b0 ;
  assign y5093 = ~n21085 ;
  assign y5094 = ~n21088 ;
  assign y5095 = ~n21090 ;
  assign y5096 = ~n21094 ;
  assign y5097 = ~n21098 ;
  assign y5098 = ~n21101 ;
  assign y5099 = ~1'b0 ;
  assign y5100 = ~n21102 ;
  assign y5101 = n21103 ;
  assign y5102 = n21105 ;
  assign y5103 = ~n21106 ;
  assign y5104 = ~n21107 ;
  assign y5105 = ~n21119 ;
  assign y5106 = ~1'b0 ;
  assign y5107 = ~n21123 ;
  assign y5108 = n21127 ;
  assign y5109 = n21130 ;
  assign y5110 = ~n21132 ;
  assign y5111 = n21137 ;
  assign y5112 = ~1'b0 ;
  assign y5113 = ~n21138 ;
  assign y5114 = n21145 ;
  assign y5115 = n21146 ;
  assign y5116 = ~n21147 ;
  assign y5117 = n21148 ;
  assign y5118 = n21153 ;
  assign y5119 = n21154 ;
  assign y5120 = n21156 ;
  assign y5121 = ~1'b0 ;
  assign y5122 = ~n21160 ;
  assign y5123 = ~n21162 ;
  assign y5124 = ~n21163 ;
  assign y5125 = n21165 ;
  assign y5126 = n21168 ;
  assign y5127 = ~n21169 ;
  assign y5128 = n21171 ;
  assign y5129 = ~n21172 ;
  assign y5130 = ~n21173 ;
  assign y5131 = ~n21184 ;
  assign y5132 = ~n21187 ;
  assign y5133 = ~n21189 ;
  assign y5134 = n21191 ;
  assign y5135 = ~n21193 ;
  assign y5136 = n21194 ;
  assign y5137 = ~n21195 ;
  assign y5138 = ~n21198 ;
  assign y5139 = ~n21202 ;
  assign y5140 = n21204 ;
  assign y5141 = n21207 ;
  assign y5142 = ~n21210 ;
  assign y5143 = ~n21212 ;
  assign y5144 = ~n21213 ;
  assign y5145 = n21214 ;
  assign y5146 = ~n21215 ;
  assign y5147 = ~n21217 ;
  assign y5148 = ~n21219 ;
  assign y5149 = ~n21221 ;
  assign y5150 = ~n21223 ;
  assign y5151 = ~n21229 ;
  assign y5152 = ~n21230 ;
  assign y5153 = n21233 ;
  assign y5154 = ~1'b0 ;
  assign y5155 = ~n21239 ;
  assign y5156 = ~n21240 ;
  assign y5157 = ~n21242 ;
  assign y5158 = n21244 ;
  assign y5159 = ~1'b0 ;
  assign y5160 = ~1'b0 ;
  assign y5161 = n21248 ;
  assign y5162 = n21249 ;
  assign y5163 = n21251 ;
  assign y5164 = ~n21253 ;
  assign y5165 = n21254 ;
  assign y5166 = n21256 ;
  assign y5167 = n21257 ;
  assign y5168 = ~n21261 ;
  assign y5169 = ~n21262 ;
  assign y5170 = ~n21266 ;
  assign y5171 = n21267 ;
  assign y5172 = ~n21271 ;
  assign y5173 = ~n21273 ;
  assign y5174 = ~n21274 ;
  assign y5175 = ~n21276 ;
  assign y5176 = ~n21277 ;
  assign y5177 = ~n21279 ;
  assign y5178 = ~1'b0 ;
  assign y5179 = ~n21284 ;
  assign y5180 = n21287 ;
  assign y5181 = n21290 ;
  assign y5182 = ~n21293 ;
  assign y5183 = ~n21294 ;
  assign y5184 = n21296 ;
  assign y5185 = ~n21298 ;
  assign y5186 = n21299 ;
  assign y5187 = n21300 ;
  assign y5188 = ~n21302 ;
  assign y5189 = ~n21308 ;
  assign y5190 = ~n21313 ;
  assign y5191 = ~n21315 ;
  assign y5192 = ~n21316 ;
  assign y5193 = n21317 ;
  assign y5194 = n21323 ;
  assign y5195 = n21324 ;
  assign y5196 = ~n21325 ;
  assign y5197 = n21329 ;
  assign y5198 = n21332 ;
  assign y5199 = ~n21333 ;
  assign y5200 = n21335 ;
  assign y5201 = n21337 ;
  assign y5202 = n21341 ;
  assign y5203 = ~1'b0 ;
  assign y5204 = ~n21345 ;
  assign y5205 = n21351 ;
  assign y5206 = ~n21357 ;
  assign y5207 = ~n21358 ;
  assign y5208 = ~n21359 ;
  assign y5209 = ~n21363 ;
  assign y5210 = n21366 ;
  assign y5211 = n21367 ;
  assign y5212 = ~n21369 ;
  assign y5213 = n21374 ;
  assign y5214 = ~1'b0 ;
  assign y5215 = n21377 ;
  assign y5216 = n21378 ;
  assign y5217 = n21381 ;
  assign y5218 = n21382 ;
  assign y5219 = ~n21384 ;
  assign y5220 = n21385 ;
  assign y5221 = n21386 ;
  assign y5222 = ~n21390 ;
  assign y5223 = n21391 ;
  assign y5224 = n21392 ;
  assign y5225 = n21394 ;
  assign y5226 = ~n21398 ;
  assign y5227 = n21399 ;
  assign y5228 = ~n21401 ;
  assign y5229 = ~1'b0 ;
  assign y5230 = ~n21404 ;
  assign y5231 = ~n21406 ;
  assign y5232 = ~n21409 ;
  assign y5233 = n21415 ;
  assign y5234 = ~n21418 ;
  assign y5235 = ~n21419 ;
  assign y5236 = n21423 ;
  assign y5237 = ~n21428 ;
  assign y5238 = ~1'b0 ;
  assign y5239 = n21430 ;
  assign y5240 = n21432 ;
  assign y5241 = ~n21434 ;
  assign y5242 = n21438 ;
  assign y5243 = ~n21439 ;
  assign y5244 = n21440 ;
  assign y5245 = ~1'b0 ;
  assign y5246 = ~n21442 ;
  assign y5247 = n21443 ;
  assign y5248 = n21444 ;
  assign y5249 = n21446 ;
  assign y5250 = n21451 ;
  assign y5251 = n21452 ;
  assign y5252 = ~n21454 ;
  assign y5253 = ~n21461 ;
  assign y5254 = n21473 ;
  assign y5255 = n21474 ;
  assign y5256 = ~n21476 ;
  assign y5257 = n21477 ;
  assign y5258 = ~n21478 ;
  assign y5259 = ~n21479 ;
  assign y5260 = n21481 ;
  assign y5261 = n21485 ;
  assign y5262 = ~n21494 ;
  assign y5263 = n21496 ;
  assign y5264 = ~n21498 ;
  assign y5265 = ~n21500 ;
  assign y5266 = ~1'b0 ;
  assign y5267 = n21501 ;
  assign y5268 = n21504 ;
  assign y5269 = ~n21505 ;
  assign y5270 = n21507 ;
  assign y5271 = ~n21512 ;
  assign y5272 = ~n21515 ;
  assign y5273 = ~1'b0 ;
  assign y5274 = n21518 ;
  assign y5275 = ~n21526 ;
  assign y5276 = n11031 ;
  assign y5277 = n21527 ;
  assign y5278 = n21529 ;
  assign y5279 = n21530 ;
  assign y5280 = n21533 ;
  assign y5281 = ~n21534 ;
  assign y5282 = n21537 ;
  assign y5283 = n21541 ;
  assign y5284 = ~n21544 ;
  assign y5285 = ~n21545 ;
  assign y5286 = ~n21546 ;
  assign y5287 = n21547 ;
  assign y5288 = n21549 ;
  assign y5289 = n21551 ;
  assign y5290 = n21554 ;
  assign y5291 = n21558 ;
  assign y5292 = ~n21562 ;
  assign y5293 = n21565 ;
  assign y5294 = ~n21566 ;
  assign y5295 = n21569 ;
  assign y5296 = ~n21571 ;
  assign y5297 = ~n21575 ;
  assign y5298 = ~n21576 ;
  assign y5299 = ~n21577 ;
  assign y5300 = n21578 ;
  assign y5301 = n21580 ;
  assign y5302 = ~n21586 ;
  assign y5303 = ~n21588 ;
  assign y5304 = n21602 ;
  assign y5305 = ~n21607 ;
  assign y5306 = n21608 ;
  assign y5307 = ~n21612 ;
  assign y5308 = ~n21613 ;
  assign y5309 = n21614 ;
  assign y5310 = n21616 ;
  assign y5311 = ~n21618 ;
  assign y5312 = n21620 ;
  assign y5313 = n21628 ;
  assign y5314 = n21630 ;
  assign y5315 = ~n21634 ;
  assign y5316 = ~n21638 ;
  assign y5317 = ~1'b0 ;
  assign y5318 = ~n21643 ;
  assign y5319 = ~n21650 ;
  assign y5320 = ~n21651 ;
  assign y5321 = ~n21652 ;
  assign y5322 = n21655 ;
  assign y5323 = n21662 ;
  assign y5324 = ~n21670 ;
  assign y5325 = ~n21672 ;
  assign y5326 = ~n21673 ;
  assign y5327 = n21678 ;
  assign y5328 = ~1'b0 ;
  assign y5329 = n21679 ;
  assign y5330 = n21687 ;
  assign y5331 = n21691 ;
  assign y5332 = n21696 ;
  assign y5333 = ~1'b0 ;
  assign y5334 = n21701 ;
  assign y5335 = n21703 ;
  assign y5336 = ~n21704 ;
  assign y5337 = ~n21707 ;
  assign y5338 = ~n21709 ;
  assign y5339 = ~n21710 ;
  assign y5340 = ~n21713 ;
  assign y5341 = ~1'b0 ;
  assign y5342 = ~n21714 ;
  assign y5343 = n21715 ;
  assign y5344 = ~n21717 ;
  assign y5345 = ~n21720 ;
  assign y5346 = ~n21724 ;
  assign y5347 = ~n21728 ;
  assign y5348 = n21729 ;
  assign y5349 = n21735 ;
  assign y5350 = n21742 ;
  assign y5351 = ~n21744 ;
  assign y5352 = n21749 ;
  assign y5353 = ~1'b0 ;
  assign y5354 = ~n21753 ;
  assign y5355 = ~n21755 ;
  assign y5356 = ~n21758 ;
  assign y5357 = ~n21763 ;
  assign y5358 = ~n21771 ;
  assign y5359 = ~n21772 ;
  assign y5360 = ~n21774 ;
  assign y5361 = ~1'b0 ;
  assign y5362 = n21777 ;
  assign y5363 = ~n21779 ;
  assign y5364 = ~n21780 ;
  assign y5365 = ~n21783 ;
  assign y5366 = n21786 ;
  assign y5367 = n21792 ;
  assign y5368 = n21798 ;
  assign y5369 = ~n21802 ;
  assign y5370 = ~n21806 ;
  assign y5371 = n21808 ;
  assign y5372 = n21810 ;
  assign y5373 = ~n21812 ;
  assign y5374 = n21815 ;
  assign y5375 = ~n21817 ;
  assign y5376 = ~n21820 ;
  assign y5377 = n21827 ;
  assign y5378 = ~n21830 ;
  assign y5379 = n21833 ;
  assign y5380 = ~n21838 ;
  assign y5381 = n21840 ;
  assign y5382 = n21841 ;
  assign y5383 = n21842 ;
  assign y5384 = ~n21847 ;
  assign y5385 = n21850 ;
  assign y5386 = n21855 ;
  assign y5387 = ~n21860 ;
  assign y5388 = n21862 ;
  assign y5389 = ~n21864 ;
  assign y5390 = ~n21870 ;
  assign y5391 = n21875 ;
  assign y5392 = ~n21876 ;
  assign y5393 = n21878 ;
  assign y5394 = ~n21881 ;
  assign y5395 = ~n21883 ;
  assign y5396 = n21884 ;
  assign y5397 = ~n21885 ;
  assign y5398 = ~n21890 ;
  assign y5399 = n21891 ;
  assign y5400 = n21893 ;
  assign y5401 = ~n21896 ;
  assign y5402 = ~n21898 ;
  assign y5403 = ~n21903 ;
  assign y5404 = ~n21905 ;
  assign y5405 = ~n21907 ;
  assign y5406 = n21909 ;
  assign y5407 = n21911 ;
  assign y5408 = n21913 ;
  assign y5409 = n21915 ;
  assign y5410 = n21916 ;
  assign y5411 = ~n21919 ;
  assign y5412 = n21922 ;
  assign y5413 = n21933 ;
  assign y5414 = ~n21934 ;
  assign y5415 = ~n21938 ;
  assign y5416 = ~n21941 ;
  assign y5417 = ~n21944 ;
  assign y5418 = n21946 ;
  assign y5419 = n21951 ;
  assign y5420 = ~n21953 ;
  assign y5421 = ~n21955 ;
  assign y5422 = ~n21973 ;
  assign y5423 = ~n21975 ;
  assign y5424 = n21977 ;
  assign y5425 = n21981 ;
  assign y5426 = ~n21985 ;
  assign y5427 = n21986 ;
  assign y5428 = ~n21987 ;
  assign y5429 = n21992 ;
  assign y5430 = n21994 ;
  assign y5431 = n21995 ;
  assign y5432 = ~n21997 ;
  assign y5433 = n21999 ;
  assign y5434 = n22003 ;
  assign y5435 = ~n22006 ;
  assign y5436 = n22009 ;
  assign y5437 = ~n22011 ;
  assign y5438 = ~1'b0 ;
  assign y5439 = ~n22015 ;
  assign y5440 = ~n22023 ;
  assign y5441 = ~n22026 ;
  assign y5442 = n22027 ;
  assign y5443 = ~n22030 ;
  assign y5444 = n22031 ;
  assign y5445 = n22033 ;
  assign y5446 = n22037 ;
  assign y5447 = n22038 ;
  assign y5448 = n22040 ;
  assign y5449 = ~n22041 ;
  assign y5450 = ~1'b0 ;
  assign y5451 = n22045 ;
  assign y5452 = ~n22047 ;
  assign y5453 = ~n22052 ;
  assign y5454 = n22058 ;
  assign y5455 = n22060 ;
  assign y5456 = ~n22065 ;
  assign y5457 = n22067 ;
  assign y5458 = n22068 ;
  assign y5459 = ~n22069 ;
  assign y5460 = n22074 ;
  assign y5461 = ~n22076 ;
  assign y5462 = n22079 ;
  assign y5463 = ~n22083 ;
  assign y5464 = ~1'b0 ;
  assign y5465 = n22086 ;
  assign y5466 = n22091 ;
  assign y5467 = n22093 ;
  assign y5468 = ~n22094 ;
  assign y5469 = ~n8481 ;
  assign y5470 = ~n22098 ;
  assign y5471 = n22104 ;
  assign y5472 = ~n22105 ;
  assign y5473 = n22106 ;
  assign y5474 = ~n22108 ;
  assign y5475 = ~n22113 ;
  assign y5476 = ~n22114 ;
  assign y5477 = n22115 ;
  assign y5478 = ~n22116 ;
  assign y5479 = n22120 ;
  assign y5480 = ~n22123 ;
  assign y5481 = ~n22128 ;
  assign y5482 = n22131 ;
  assign y5483 = n22133 ;
  assign y5484 = ~n22135 ;
  assign y5485 = ~n22147 ;
  assign y5486 = n22148 ;
  assign y5487 = n22150 ;
  assign y5488 = n22153 ;
  assign y5489 = ~n22154 ;
  assign y5490 = n22160 ;
  assign y5491 = ~n22163 ;
  assign y5492 = ~n22170 ;
  assign y5493 = ~n22174 ;
  assign y5494 = n22175 ;
  assign y5495 = n22176 ;
  assign y5496 = n22177 ;
  assign y5497 = ~n22181 ;
  assign y5498 = n22187 ;
  assign y5499 = ~n22191 ;
  assign y5500 = n22193 ;
  assign y5501 = n22194 ;
  assign y5502 = n22197 ;
  assign y5503 = ~n22202 ;
  assign y5504 = n22205 ;
  assign y5505 = n22211 ;
  assign y5506 = n22212 ;
  assign y5507 = n22225 ;
  assign y5508 = n22233 ;
  assign y5509 = ~n22235 ;
  assign y5510 = ~n22236 ;
  assign y5511 = n22237 ;
  assign y5512 = n22240 ;
  assign y5513 = n22247 ;
  assign y5514 = n22249 ;
  assign y5515 = ~n22252 ;
  assign y5516 = n22253 ;
  assign y5517 = ~n22254 ;
  assign y5518 = n22258 ;
  assign y5519 = ~n22261 ;
  assign y5520 = n22265 ;
  assign y5521 = n22266 ;
  assign y5522 = n22269 ;
  assign y5523 = n22270 ;
  assign y5524 = n22273 ;
  assign y5525 = n22280 ;
  assign y5526 = n22288 ;
  assign y5527 = ~n22291 ;
  assign y5528 = n22292 ;
  assign y5529 = n22297 ;
  assign y5530 = n22300 ;
  assign y5531 = ~n22303 ;
  assign y5532 = ~n22306 ;
  assign y5533 = ~n22308 ;
  assign y5534 = ~n22309 ;
  assign y5535 = ~n22311 ;
  assign y5536 = ~n22313 ;
  assign y5537 = ~n22314 ;
  assign y5538 = ~n22315 ;
  assign y5539 = ~n22316 ;
  assign y5540 = ~n22318 ;
  assign y5541 = n22321 ;
  assign y5542 = n22324 ;
  assign y5543 = n22325 ;
  assign y5544 = ~n22327 ;
  assign y5545 = n22333 ;
  assign y5546 = n22339 ;
  assign y5547 = n22342 ;
  assign y5548 = n22345 ;
  assign y5549 = ~n22353 ;
  assign y5550 = n22355 ;
  assign y5551 = n22362 ;
  assign y5552 = n22366 ;
  assign y5553 = ~n22367 ;
  assign y5554 = n22369 ;
  assign y5555 = n22374 ;
  assign y5556 = ~n22375 ;
  assign y5557 = ~n22380 ;
  assign y5558 = n22382 ;
  assign y5559 = ~n22383 ;
  assign y5560 = n22386 ;
  assign y5561 = n22390 ;
  assign y5562 = ~n22391 ;
  assign y5563 = ~n22393 ;
  assign y5564 = ~n22396 ;
  assign y5565 = n22397 ;
  assign y5566 = n22401 ;
  assign y5567 = ~n22415 ;
  assign y5568 = ~n22417 ;
  assign y5569 = ~n22418 ;
  assign y5570 = n22422 ;
  assign y5571 = n22423 ;
  assign y5572 = n22425 ;
  assign y5573 = ~n22427 ;
  assign y5574 = n22430 ;
  assign y5575 = ~1'b0 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~n22431 ;
  assign y5578 = n22434 ;
  assign y5579 = n22435 ;
  assign y5580 = n22438 ;
  assign y5581 = n22444 ;
  assign y5582 = ~1'b0 ;
  assign y5583 = n22446 ;
  assign y5584 = n22449 ;
  assign y5585 = n22451 ;
  assign y5586 = n22454 ;
  assign y5587 = n22457 ;
  assign y5588 = ~n22462 ;
  assign y5589 = n22464 ;
  assign y5590 = ~n22466 ;
  assign y5591 = ~n22471 ;
  assign y5592 = ~n22474 ;
  assign y5593 = n22477 ;
  assign y5594 = ~n22478 ;
  assign y5595 = ~n22482 ;
  assign y5596 = n22487 ;
  assign y5597 = n22488 ;
  assign y5598 = n22491 ;
  assign y5599 = ~n22493 ;
  assign y5600 = n22495 ;
  assign y5601 = ~n22497 ;
  assign y5602 = ~n22502 ;
  assign y5603 = n22503 ;
  assign y5604 = ~n22505 ;
  assign y5605 = ~n22506 ;
  assign y5606 = ~n22511 ;
  assign y5607 = ~n22514 ;
  assign y5608 = n22516 ;
  assign y5609 = ~1'b0 ;
  assign y5610 = ~n22517 ;
  assign y5611 = ~n22520 ;
  assign y5612 = n22523 ;
  assign y5613 = n22526 ;
  assign y5614 = ~n22530 ;
  assign y5615 = ~n22533 ;
  assign y5616 = n22534 ;
  assign y5617 = ~n22536 ;
  assign y5618 = n22537 ;
  assign y5619 = n22539 ;
  assign y5620 = ~n22540 ;
  assign y5621 = ~n22543 ;
  assign y5622 = ~n22545 ;
  assign y5623 = ~n22548 ;
  assign y5624 = ~n22549 ;
  assign y5625 = ~n22551 ;
  assign y5626 = ~n22555 ;
  assign y5627 = ~n22559 ;
  assign y5628 = n22560 ;
  assign y5629 = ~n22566 ;
  assign y5630 = ~n22572 ;
  assign y5631 = ~n22573 ;
  assign y5632 = n22574 ;
  assign y5633 = ~n22575 ;
  assign y5634 = n22577 ;
  assign y5635 = n22580 ;
  assign y5636 = n22581 ;
  assign y5637 = ~n22586 ;
  assign y5638 = ~n22587 ;
  assign y5639 = ~1'b0 ;
  assign y5640 = ~n22591 ;
  assign y5641 = ~1'b0 ;
  assign y5642 = n22592 ;
  assign y5643 = n22595 ;
  assign y5644 = n22605 ;
  assign y5645 = n22612 ;
  assign y5646 = ~n22615 ;
  assign y5647 = ~n22618 ;
  assign y5648 = ~n22619 ;
  assign y5649 = ~n22622 ;
  assign y5650 = n22623 ;
  assign y5651 = n22624 ;
  assign y5652 = ~n22625 ;
  assign y5653 = n22627 ;
  assign y5654 = ~n22630 ;
  assign y5655 = ~1'b0 ;
  assign y5656 = n22631 ;
  assign y5657 = ~n22632 ;
  assign y5658 = ~n22633 ;
  assign y5659 = ~n22635 ;
  assign y5660 = ~n22636 ;
  assign y5661 = n22640 ;
  assign y5662 = n22641 ;
  assign y5663 = ~n22643 ;
  assign y5664 = n22644 ;
  assign y5665 = n22649 ;
  assign y5666 = n22650 ;
  assign y5667 = ~n22651 ;
  assign y5668 = ~n22653 ;
  assign y5669 = ~1'b0 ;
  assign y5670 = n22655 ;
  assign y5671 = ~n22657 ;
  assign y5672 = ~n22660 ;
  assign y5673 = ~n22665 ;
  assign y5674 = n22666 ;
  assign y5675 = ~n22671 ;
  assign y5676 = ~1'b0 ;
  assign y5677 = n22672 ;
  assign y5678 = ~n22680 ;
  assign y5679 = n22681 ;
  assign y5680 = n22682 ;
  assign y5681 = ~n22683 ;
  assign y5682 = n22684 ;
  assign y5683 = n22687 ;
  assign y5684 = ~1'b0 ;
  assign y5685 = n22688 ;
  assign y5686 = ~n22691 ;
  assign y5687 = n22692 ;
  assign y5688 = n22699 ;
  assign y5689 = ~n22700 ;
  assign y5690 = ~n22702 ;
  assign y5691 = n22703 ;
  assign y5692 = n22713 ;
  assign y5693 = n22717 ;
  assign y5694 = ~1'b0 ;
  assign y5695 = n22722 ;
  assign y5696 = n22726 ;
  assign y5697 = ~n22729 ;
  assign y5698 = ~n22732 ;
  assign y5699 = ~n22735 ;
  assign y5700 = ~1'b0 ;
  assign y5701 = n22740 ;
  assign y5702 = ~n22744 ;
  assign y5703 = n22746 ;
  assign y5704 = n22747 ;
  assign y5705 = ~n22748 ;
  assign y5706 = n22751 ;
  assign y5707 = ~n22753 ;
  assign y5708 = n22754 ;
  assign y5709 = ~n22756 ;
  assign y5710 = ~n22759 ;
  assign y5711 = n22761 ;
  assign y5712 = ~n22762 ;
  assign y5713 = n22763 ;
  assign y5714 = n22764 ;
  assign y5715 = n22766 ;
  assign y5716 = n22769 ;
  assign y5717 = ~n22771 ;
  assign y5718 = n22776 ;
  assign y5719 = ~n22778 ;
  assign y5720 = n22781 ;
  assign y5721 = ~n22785 ;
  assign y5722 = ~n22787 ;
  assign y5723 = ~n22788 ;
  assign y5724 = ~n22797 ;
  assign y5725 = n22798 ;
  assign y5726 = ~n22800 ;
  assign y5727 = n22802 ;
  assign y5728 = ~1'b0 ;
  assign y5729 = ~1'b0 ;
  assign y5730 = ~n22804 ;
  assign y5731 = n22812 ;
  assign y5732 = ~n22813 ;
  assign y5733 = ~n22814 ;
  assign y5734 = ~n22815 ;
  assign y5735 = n22818 ;
  assign y5736 = ~n22819 ;
  assign y5737 = ~n22823 ;
  assign y5738 = n22825 ;
  assign y5739 = n22828 ;
  assign y5740 = n22829 ;
  assign y5741 = n22835 ;
  assign y5742 = ~n22836 ;
  assign y5743 = ~n22838 ;
  assign y5744 = ~n22843 ;
  assign y5745 = ~1'b0 ;
  assign y5746 = ~n22847 ;
  assign y5747 = n22854 ;
  assign y5748 = n22857 ;
  assign y5749 = ~n22858 ;
  assign y5750 = ~n22865 ;
  assign y5751 = ~n22866 ;
  assign y5752 = ~n22868 ;
  assign y5753 = n22870 ;
  assign y5754 = ~n22872 ;
  assign y5755 = ~n22880 ;
  assign y5756 = ~n22881 ;
  assign y5757 = ~n22882 ;
  assign y5758 = n22884 ;
  assign y5759 = ~1'b0 ;
  assign y5760 = ~n22891 ;
  assign y5761 = n22897 ;
  assign y5762 = ~n22899 ;
  assign y5763 = n22906 ;
  assign y5764 = n22917 ;
  assign y5765 = ~n22918 ;
  assign y5766 = ~n22919 ;
  assign y5767 = ~1'b0 ;
  assign y5768 = ~n22922 ;
  assign y5769 = ~n22924 ;
  assign y5770 = ~n22925 ;
  assign y5771 = n22926 ;
  assign y5772 = n22933 ;
  assign y5773 = ~n22935 ;
  assign y5774 = ~n22939 ;
  assign y5775 = ~n22943 ;
  assign y5776 = ~n22945 ;
  assign y5777 = n22946 ;
  assign y5778 = n22947 ;
  assign y5779 = ~1'b0 ;
  assign y5780 = ~n22950 ;
  assign y5781 = n22957 ;
  assign y5782 = ~n22959 ;
  assign y5783 = n22960 ;
  assign y5784 = ~n22961 ;
  assign y5785 = n22966 ;
  assign y5786 = n22969 ;
  assign y5787 = ~1'b0 ;
  assign y5788 = n22972 ;
  assign y5789 = n22979 ;
  assign y5790 = ~n22983 ;
  assign y5791 = ~n22985 ;
  assign y5792 = ~n22987 ;
  assign y5793 = n22992 ;
  assign y5794 = ~n22994 ;
  assign y5795 = ~n22996 ;
  assign y5796 = n22998 ;
  assign y5797 = n22999 ;
  assign y5798 = n23000 ;
  assign y5799 = n23004 ;
  assign y5800 = n23011 ;
  assign y5801 = ~n23014 ;
  assign y5802 = ~n23024 ;
  assign y5803 = n23026 ;
  assign y5804 = ~n23029 ;
  assign y5805 = n23033 ;
  assign y5806 = n23035 ;
  assign y5807 = n23038 ;
  assign y5808 = ~n23039 ;
  assign y5809 = ~1'b0 ;
  assign y5810 = ~1'b0 ;
  assign y5811 = n23042 ;
  assign y5812 = ~n23043 ;
  assign y5813 = ~n23044 ;
  assign y5814 = n23049 ;
  assign y5815 = n23053 ;
  assign y5816 = ~n23056 ;
  assign y5817 = ~n23062 ;
  assign y5818 = ~n23063 ;
  assign y5819 = n23064 ;
  assign y5820 = ~n23067 ;
  assign y5821 = n23068 ;
  assign y5822 = n23070 ;
  assign y5823 = n23072 ;
  assign y5824 = ~n23073 ;
  assign y5825 = ~n23074 ;
  assign y5826 = ~1'b0 ;
  assign y5827 = n23079 ;
  assign y5828 = ~n23081 ;
  assign y5829 = n23083 ;
  assign y5830 = ~n23087 ;
  assign y5831 = n23091 ;
  assign y5832 = ~n23095 ;
  assign y5833 = ~n23099 ;
  assign y5834 = ~n23102 ;
  assign y5835 = ~n23106 ;
  assign y5836 = n23112 ;
  assign y5837 = ~n23117 ;
  assign y5838 = ~n23120 ;
  assign y5839 = ~n23121 ;
  assign y5840 = n23122 ;
  assign y5841 = ~n23123 ;
  assign y5842 = n23125 ;
  assign y5843 = ~n23129 ;
  assign y5844 = n23131 ;
  assign y5845 = ~n23132 ;
  assign y5846 = ~n23133 ;
  assign y5847 = ~n23135 ;
  assign y5848 = n23139 ;
  assign y5849 = ~n23143 ;
  assign y5850 = n23145 ;
  assign y5851 = ~n23151 ;
  assign y5852 = ~n23160 ;
  assign y5853 = n23161 ;
  assign y5854 = ~n23163 ;
  assign y5855 = n23164 ;
  assign y5856 = ~n23166 ;
  assign y5857 = n23169 ;
  assign y5858 = n23171 ;
  assign y5859 = ~n23173 ;
  assign y5860 = n23175 ;
  assign y5861 = n23177 ;
  assign y5862 = ~n23182 ;
  assign y5863 = ~1'b0 ;
  assign y5864 = ~1'b0 ;
  assign y5865 = ~n23183 ;
  assign y5866 = n23188 ;
  assign y5867 = n23189 ;
  assign y5868 = ~n23191 ;
  assign y5869 = n23192 ;
  assign y5870 = n23196 ;
  assign y5871 = ~n23200 ;
  assign y5872 = ~n23203 ;
  assign y5873 = n23206 ;
  assign y5874 = n23210 ;
  assign y5875 = n23212 ;
  assign y5876 = n23213 ;
  assign y5877 = n23214 ;
  assign y5878 = ~1'b0 ;
  assign y5879 = ~1'b0 ;
  assign y5880 = n23216 ;
  assign y5881 = n23220 ;
  assign y5882 = n23222 ;
  assign y5883 = n23224 ;
  assign y5884 = n23225 ;
  assign y5885 = n23230 ;
  assign y5886 = n23231 ;
  assign y5887 = ~n23233 ;
  assign y5888 = n23236 ;
  assign y5889 = ~n23237 ;
  assign y5890 = ~n23239 ;
  assign y5891 = ~n23240 ;
  assign y5892 = ~n23243 ;
  assign y5893 = ~n23245 ;
  assign y5894 = n23247 ;
  assign y5895 = ~n23249 ;
  assign y5896 = ~1'b0 ;
  assign y5897 = ~n23251 ;
  assign y5898 = n23252 ;
  assign y5899 = ~n23255 ;
  assign y5900 = ~n23260 ;
  assign y5901 = n23261 ;
  assign y5902 = ~n23264 ;
  assign y5903 = ~n23267 ;
  assign y5904 = n23269 ;
  assign y5905 = ~n23277 ;
  assign y5906 = n23278 ;
  assign y5907 = n23280 ;
  assign y5908 = n23282 ;
  assign y5909 = ~n23286 ;
  assign y5910 = n23289 ;
  assign y5911 = n23296 ;
  assign y5912 = ~n23297 ;
  assign y5913 = ~n23299 ;
  assign y5914 = ~n23306 ;
  assign y5915 = n23309 ;
  assign y5916 = ~n23312 ;
  assign y5917 = n23319 ;
  assign y5918 = n23323 ;
  assign y5919 = ~n23329 ;
  assign y5920 = n23332 ;
  assign y5921 = n23334 ;
  assign y5922 = ~1'b0 ;
  assign y5923 = n23337 ;
  assign y5924 = ~n23339 ;
  assign y5925 = ~n23343 ;
  assign y5926 = ~n23344 ;
  assign y5927 = n23347 ;
  assign y5928 = n23349 ;
  assign y5929 = n23351 ;
  assign y5930 = ~1'b0 ;
  assign y5931 = n23352 ;
  assign y5932 = n23354 ;
  assign y5933 = ~n23360 ;
  assign y5934 = n23365 ;
  assign y5935 = ~n23368 ;
  assign y5936 = ~n23372 ;
  assign y5937 = n23373 ;
  assign y5938 = ~n23377 ;
  assign y5939 = n23378 ;
  assign y5940 = n23380 ;
  assign y5941 = ~n23385 ;
  assign y5942 = ~n23386 ;
  assign y5943 = n18681 ;
  assign y5944 = ~n23388 ;
  assign y5945 = ~n23393 ;
  assign y5946 = ~n23394 ;
  assign y5947 = n23396 ;
  assign y5948 = ~n23397 ;
  assign y5949 = n23399 ;
  assign y5950 = n23400 ;
  assign y5951 = ~n23402 ;
  assign y5952 = ~1'b0 ;
  assign y5953 = ~n23409 ;
  assign y5954 = n23411 ;
  assign y5955 = n23413 ;
  assign y5956 = ~n23415 ;
  assign y5957 = n23418 ;
  assign y5958 = n23422 ;
  assign y5959 = ~n23423 ;
  assign y5960 = n23425 ;
  assign y5961 = n23433 ;
  assign y5962 = ~n23435 ;
  assign y5963 = ~n23441 ;
  assign y5964 = ~1'b0 ;
  assign y5965 = n23442 ;
  assign y5966 = ~n23446 ;
  assign y5967 = n23449 ;
  assign y5968 = ~n23452 ;
  assign y5969 = n23457 ;
  assign y5970 = ~n23459 ;
  assign y5971 = n23465 ;
  assign y5972 = n23467 ;
  assign y5973 = ~n23468 ;
  assign y5974 = ~n23472 ;
  assign y5975 = n23474 ;
  assign y5976 = n23475 ;
  assign y5977 = n23476 ;
  assign y5978 = n23480 ;
  assign y5979 = ~1'b0 ;
  assign y5980 = ~n23487 ;
  assign y5981 = ~n23490 ;
  assign y5982 = ~n23499 ;
  assign y5983 = n23501 ;
  assign y5984 = n23502 ;
  assign y5985 = n23504 ;
  assign y5986 = n23505 ;
  assign y5987 = ~n23507 ;
  assign y5988 = ~n23509 ;
  assign y5989 = ~n23522 ;
  assign y5990 = ~n23526 ;
  assign y5991 = ~n23528 ;
  assign y5992 = ~n23531 ;
  assign y5993 = n23534 ;
  assign y5994 = n23537 ;
  assign y5995 = ~n23538 ;
  assign y5996 = n23543 ;
  assign y5997 = ~n23545 ;
  assign y5998 = n23546 ;
  assign y5999 = n23548 ;
  assign y6000 = ~1'b0 ;
  assign y6001 = n23550 ;
  assign y6002 = n23553 ;
  assign y6003 = n23556 ;
  assign y6004 = n23560 ;
  assign y6005 = n23566 ;
  assign y6006 = ~n23567 ;
  assign y6007 = n23568 ;
  assign y6008 = ~n23572 ;
  assign y6009 = n23574 ;
  assign y6010 = ~n23577 ;
  assign y6011 = ~n23579 ;
  assign y6012 = ~n23581 ;
  assign y6013 = n23582 ;
  assign y6014 = n23584 ;
  assign y6015 = n23588 ;
  assign y6016 = n23593 ;
  assign y6017 = ~n23594 ;
  assign y6018 = n23598 ;
  assign y6019 = ~n23602 ;
  assign y6020 = ~n23604 ;
  assign y6021 = n23611 ;
  assign y6022 = n23612 ;
  assign y6023 = ~n23615 ;
  assign y6024 = ~n23619 ;
  assign y6025 = n23621 ;
  assign y6026 = n23622 ;
  assign y6027 = ~n23624 ;
  assign y6028 = ~n23626 ;
  assign y6029 = ~1'b0 ;
  assign y6030 = ~n23631 ;
  assign y6031 = ~n23634 ;
  assign y6032 = n23639 ;
  assign y6033 = n23640 ;
  assign y6034 = n23643 ;
  assign y6035 = n23645 ;
  assign y6036 = ~n23647 ;
  assign y6037 = ~n23649 ;
  assign y6038 = n23659 ;
  assign y6039 = ~n23667 ;
  assign y6040 = n23674 ;
  assign y6041 = n23676 ;
  assign y6042 = ~1'b0 ;
  assign y6043 = n23678 ;
  assign y6044 = ~n23679 ;
  assign y6045 = n23680 ;
  assign y6046 = ~n23682 ;
  assign y6047 = ~n23683 ;
  assign y6048 = n23688 ;
  assign y6049 = ~n23691 ;
  assign y6050 = n23694 ;
  assign y6051 = n23697 ;
  assign y6052 = ~n23698 ;
  assign y6053 = n23700 ;
  assign y6054 = n23701 ;
  assign y6055 = ~n23703 ;
  assign y6056 = ~n23707 ;
  assign y6057 = n23710 ;
  assign y6058 = ~n23712 ;
  assign y6059 = n23713 ;
  assign y6060 = ~n23714 ;
  assign y6061 = n23715 ;
  assign y6062 = ~n23720 ;
  assign y6063 = ~1'b0 ;
  assign y6064 = ~n23727 ;
  assign y6065 = ~n23728 ;
  assign y6066 = ~n23733 ;
  assign y6067 = ~n23738 ;
  assign y6068 = ~n23741 ;
  assign y6069 = ~n23744 ;
  assign y6070 = n23747 ;
  assign y6071 = n23750 ;
  assign y6072 = ~n23752 ;
  assign y6073 = ~n23758 ;
  assign y6074 = ~n23762 ;
  assign y6075 = n23769 ;
  assign y6076 = ~n23780 ;
  assign y6077 = n23784 ;
  assign y6078 = ~n23787 ;
  assign y6079 = ~n23790 ;
  assign y6080 = n23792 ;
  assign y6081 = n23793 ;
  assign y6082 = ~n23794 ;
  assign y6083 = ~1'b0 ;
  assign y6084 = ~1'b0 ;
  assign y6085 = ~n23798 ;
  assign y6086 = n23806 ;
  assign y6087 = ~n23807 ;
  assign y6088 = ~n23809 ;
  assign y6089 = ~n23811 ;
  assign y6090 = ~n23813 ;
  assign y6091 = n23815 ;
  assign y6092 = ~n23828 ;
  assign y6093 = ~n23830 ;
  assign y6094 = n23839 ;
  assign y6095 = ~n23842 ;
  assign y6096 = ~n23844 ;
  assign y6097 = ~n23845 ;
  assign y6098 = ~n23848 ;
  assign y6099 = ~n23850 ;
  assign y6100 = n23854 ;
  assign y6101 = ~n23857 ;
  assign y6102 = ~n23863 ;
  assign y6103 = ~n23866 ;
  assign y6104 = ~n23867 ;
  assign y6105 = n23868 ;
  assign y6106 = ~1'b0 ;
  assign y6107 = ~n23872 ;
  assign y6108 = ~n23873 ;
  assign y6109 = ~n23874 ;
  assign y6110 = n23875 ;
  assign y6111 = n23877 ;
  assign y6112 = n23878 ;
  assign y6113 = n23882 ;
  assign y6114 = n23883 ;
  assign y6115 = ~1'b0 ;
  assign y6116 = n23884 ;
  assign y6117 = n23886 ;
  assign y6118 = ~n23890 ;
  assign y6119 = ~n23899 ;
  assign y6120 = ~n23900 ;
  assign y6121 = n23902 ;
  assign y6122 = n23907 ;
  assign y6123 = n23912 ;
  assign y6124 = ~n23913 ;
  assign y6125 = ~n23916 ;
  assign y6126 = n23923 ;
  assign y6127 = n23924 ;
  assign y6128 = ~n23925 ;
  assign y6129 = ~1'b0 ;
  assign y6130 = n23930 ;
  assign y6131 = n23933 ;
  assign y6132 = n23934 ;
  assign y6133 = n23941 ;
  assign y6134 = ~n23942 ;
  assign y6135 = n23944 ;
  assign y6136 = ~1'b0 ;
  assign y6137 = n23945 ;
  assign y6138 = n23946 ;
  assign y6139 = ~n23947 ;
  assign y6140 = ~n23954 ;
  assign y6141 = ~n23956 ;
  assign y6142 = ~1'b0 ;
  assign y6143 = ~1'b0 ;
  assign y6144 = n23959 ;
  assign y6145 = ~n23962 ;
  assign y6146 = n23963 ;
  assign y6147 = ~n23964 ;
  assign y6148 = ~n23966 ;
  assign y6149 = ~n23978 ;
  assign y6150 = ~1'b0 ;
  assign y6151 = ~n23982 ;
  assign y6152 = n23984 ;
  assign y6153 = n23985 ;
  assign y6154 = ~n23987 ;
  assign y6155 = n23988 ;
  assign y6156 = ~1'b0 ;
  assign y6157 = n23992 ;
  assign y6158 = ~n23998 ;
  assign y6159 = n24002 ;
  assign y6160 = n24005 ;
  assign y6161 = ~n24006 ;
  assign y6162 = n24007 ;
  assign y6163 = n24008 ;
  assign y6164 = n24011 ;
  assign y6165 = n24013 ;
  assign y6166 = ~n24015 ;
  assign y6167 = n24017 ;
  assign y6168 = n24019 ;
  assign y6169 = ~n24020 ;
  assign y6170 = n24022 ;
  assign y6171 = ~n24025 ;
  assign y6172 = n24027 ;
  assign y6173 = ~n24029 ;
  assign y6174 = ~n24031 ;
  assign y6175 = ~n24037 ;
  assign y6176 = n24040 ;
  assign y6177 = ~n24045 ;
  assign y6178 = n24046 ;
  assign y6179 = n24050 ;
  assign y6180 = ~n24056 ;
  assign y6181 = n24060 ;
  assign y6182 = ~n24061 ;
  assign y6183 = ~n24062 ;
  assign y6184 = ~n24064 ;
  assign y6185 = ~n24068 ;
  assign y6186 = n24071 ;
  assign y6187 = ~n24075 ;
  assign y6188 = n24077 ;
  assign y6189 = ~n24078 ;
  assign y6190 = ~n24082 ;
  assign y6191 = ~n24084 ;
  assign y6192 = n24091 ;
  assign y6193 = n24093 ;
  assign y6194 = ~n24094 ;
  assign y6195 = n24097 ;
  assign y6196 = ~n24098 ;
  assign y6197 = ~n24099 ;
  assign y6198 = n24102 ;
  assign y6199 = ~n24104 ;
  assign y6200 = ~1'b0 ;
  assign y6201 = ~n24105 ;
  assign y6202 = n24110 ;
  assign y6203 = n24114 ;
  assign y6204 = ~n24117 ;
  assign y6205 = ~1'b0 ;
  assign y6206 = ~1'b0 ;
  assign y6207 = ~n24120 ;
  assign y6208 = n24121 ;
  assign y6209 = n24126 ;
  assign y6210 = n24127 ;
  assign y6211 = n24133 ;
  assign y6212 = ~n24135 ;
  assign y6213 = n24136 ;
  assign y6214 = n24142 ;
  assign y6215 = ~n24154 ;
  assign y6216 = ~n24158 ;
  assign y6217 = ~n24170 ;
  assign y6218 = n24173 ;
  assign y6219 = ~n24176 ;
  assign y6220 = ~1'b0 ;
  assign y6221 = ~n24178 ;
  assign y6222 = n24189 ;
  assign y6223 = ~n24192 ;
  assign y6224 = n24194 ;
  assign y6225 = ~n24199 ;
  assign y6226 = n24200 ;
  assign y6227 = n24201 ;
  assign y6228 = ~n24202 ;
  assign y6229 = ~n24206 ;
  assign y6230 = ~n24207 ;
  assign y6231 = ~n24213 ;
  assign y6232 = ~n24216 ;
  assign y6233 = n24218 ;
  assign y6234 = ~1'b0 ;
  assign y6235 = ~n24219 ;
  assign y6236 = ~n24220 ;
  assign y6237 = n24225 ;
  assign y6238 = ~n24226 ;
  assign y6239 = n24229 ;
  assign y6240 = ~n24230 ;
  assign y6241 = ~n24231 ;
  assign y6242 = ~n24233 ;
  assign y6243 = ~n24234 ;
  assign y6244 = ~n24239 ;
  assign y6245 = n24241 ;
  assign y6246 = ~1'b0 ;
  assign y6247 = n24248 ;
  assign y6248 = n24249 ;
  assign y6249 = ~n24250 ;
  assign y6250 = n24251 ;
  assign y6251 = ~1'b0 ;
  assign y6252 = n24253 ;
  assign y6253 = ~n24258 ;
  assign y6254 = n24261 ;
  assign y6255 = ~n24264 ;
  assign y6256 = ~n24265 ;
  assign y6257 = ~n24271 ;
  assign y6258 = n24278 ;
  assign y6259 = ~n24284 ;
  assign y6260 = ~n24287 ;
  assign y6261 = ~n24289 ;
  assign y6262 = n24292 ;
  assign y6263 = n24296 ;
  assign y6264 = n24299 ;
  assign y6265 = n24302 ;
  assign y6266 = ~n24303 ;
  assign y6267 = n24305 ;
  assign y6268 = n24308 ;
  assign y6269 = n24309 ;
  assign y6270 = n24311 ;
  assign y6271 = ~n12729 ;
  assign y6272 = n24317 ;
  assign y6273 = n24321 ;
  assign y6274 = n24324 ;
  assign y6275 = ~n24325 ;
  assign y6276 = n24327 ;
  assign y6277 = ~n24330 ;
  assign y6278 = n24331 ;
  assign y6279 = n24332 ;
  assign y6280 = ~n24333 ;
  assign y6281 = n24335 ;
  assign y6282 = n24337 ;
  assign y6283 = ~1'b0 ;
  assign y6284 = ~1'b0 ;
  assign y6285 = ~n24340 ;
  assign y6286 = n24343 ;
  assign y6287 = ~n24347 ;
  assign y6288 = ~n24351 ;
  assign y6289 = ~n24355 ;
  assign y6290 = ~n24356 ;
  assign y6291 = n24357 ;
  assign y6292 = ~n24359 ;
  assign y6293 = n24363 ;
  assign y6294 = ~n24364 ;
  assign y6295 = ~n24366 ;
  assign y6296 = ~n24368 ;
  assign y6297 = ~n24369 ;
  assign y6298 = ~n24373 ;
  assign y6299 = ~n24375 ;
  assign y6300 = ~1'b0 ;
  assign y6301 = ~n24380 ;
  assign y6302 = n24383 ;
  assign y6303 = ~n24384 ;
  assign y6304 = ~n24385 ;
  assign y6305 = n24387 ;
  assign y6306 = n24391 ;
  assign y6307 = ~n24392 ;
  assign y6308 = ~n24396 ;
  assign y6309 = n24398 ;
  assign y6310 = n24401 ;
  assign y6311 = n24402 ;
  assign y6312 = ~n24404 ;
  assign y6313 = n24405 ;
  assign y6314 = n24406 ;
  assign y6315 = n24407 ;
  assign y6316 = n24412 ;
  assign y6317 = ~1'b0 ;
  assign y6318 = ~n24416 ;
  assign y6319 = n24421 ;
  assign y6320 = ~n24422 ;
  assign y6321 = ~n24427 ;
  assign y6322 = n24429 ;
  assign y6323 = ~1'b0 ;
  assign y6324 = ~n24430 ;
  assign y6325 = ~n24440 ;
  assign y6326 = n24445 ;
  assign y6327 = n24447 ;
  assign y6328 = n24451 ;
  assign y6329 = ~n24461 ;
  assign y6330 = ~n24466 ;
  assign y6331 = ~n24468 ;
  assign y6332 = ~n24469 ;
  assign y6333 = n24471 ;
  assign y6334 = n24472 ;
  assign y6335 = ~n24473 ;
  assign y6336 = ~n24474 ;
  assign y6337 = n24481 ;
  assign y6338 = ~n24484 ;
  assign y6339 = ~n24487 ;
  assign y6340 = n24488 ;
  assign y6341 = ~n24490 ;
  assign y6342 = ~n24493 ;
  assign y6343 = n24495 ;
  assign y6344 = n24496 ;
  assign y6345 = ~1'b0 ;
  assign y6346 = ~n24498 ;
  assign y6347 = ~1'b0 ;
  assign y6348 = n24507 ;
  assign y6349 = n24509 ;
  assign y6350 = n24513 ;
  assign y6351 = n24514 ;
  assign y6352 = n24516 ;
  assign y6353 = ~n24518 ;
  assign y6354 = n24521 ;
  assign y6355 = ~n24522 ;
  assign y6356 = n24524 ;
  assign y6357 = ~n24526 ;
  assign y6358 = n24531 ;
  assign y6359 = n24532 ;
  assign y6360 = n24533 ;
  assign y6361 = ~n24538 ;
  assign y6362 = n24541 ;
  assign y6363 = ~1'b0 ;
  assign y6364 = ~1'b0 ;
  assign y6365 = n24544 ;
  assign y6366 = ~n24549 ;
  assign y6367 = ~n24552 ;
  assign y6368 = n24555 ;
  assign y6369 = ~n24556 ;
  assign y6370 = ~n24557 ;
  assign y6371 = ~1'b0 ;
  assign y6372 = n24560 ;
  assign y6373 = ~1'b0 ;
  assign y6374 = ~n24561 ;
  assign y6375 = n24563 ;
  assign y6376 = ~n24564 ;
  assign y6377 = n24567 ;
  assign y6378 = n24568 ;
  assign y6379 = ~n24572 ;
  assign y6380 = ~n24578 ;
  assign y6381 = ~1'b0 ;
  assign y6382 = ~1'b0 ;
  assign y6383 = n24580 ;
  assign y6384 = ~n24584 ;
  assign y6385 = ~n24585 ;
  assign y6386 = ~n24587 ;
  assign y6387 = n24590 ;
  assign y6388 = n24592 ;
  assign y6389 = n24594 ;
  assign y6390 = ~n24596 ;
  assign y6391 = n15513 ;
  assign y6392 = n24599 ;
  assign y6393 = ~n24600 ;
  assign y6394 = n24606 ;
  assign y6395 = n24609 ;
  assign y6396 = n24611 ;
  assign y6397 = n24617 ;
  assign y6398 = n24618 ;
  assign y6399 = n24620 ;
  assign y6400 = n24622 ;
  assign y6401 = ~n24624 ;
  assign y6402 = ~n24636 ;
  assign y6403 = ~n4856 ;
  assign y6404 = n24638 ;
  assign y6405 = n24642 ;
  assign y6406 = ~n24644 ;
  assign y6407 = n24645 ;
  assign y6408 = ~n24647 ;
  assign y6409 = ~n24649 ;
  assign y6410 = ~n24652 ;
  assign y6411 = ~n24653 ;
  assign y6412 = n24655 ;
  assign y6413 = n24657 ;
  assign y6414 = ~1'b0 ;
  assign y6415 = ~n24658 ;
  assign y6416 = ~n24661 ;
  assign y6417 = ~n24664 ;
  assign y6418 = n24666 ;
  assign y6419 = ~n24675 ;
  assign y6420 = n24676 ;
  assign y6421 = ~n24678 ;
  assign y6422 = ~1'b0 ;
  assign y6423 = ~1'b0 ;
  assign y6424 = ~n24679 ;
  assign y6425 = n24680 ;
  assign y6426 = ~n24682 ;
  assign y6427 = ~n24684 ;
  assign y6428 = ~n24686 ;
  assign y6429 = n24688 ;
  assign y6430 = n24690 ;
  assign y6431 = n24692 ;
  assign y6432 = n24693 ;
  assign y6433 = n24694 ;
  assign y6434 = n24695 ;
  assign y6435 = ~n24696 ;
  assign y6436 = ~n24706 ;
  assign y6437 = n24709 ;
  assign y6438 = ~n24714 ;
  assign y6439 = ~1'b0 ;
  assign y6440 = ~1'b0 ;
  assign y6441 = ~1'b0 ;
  assign y6442 = ~n24719 ;
  assign y6443 = n24720 ;
  assign y6444 = n24721 ;
  assign y6445 = ~n24722 ;
  assign y6446 = ~n24723 ;
  assign y6447 = ~1'b0 ;
  assign y6448 = ~1'b0 ;
  assign y6449 = n24725 ;
  assign y6450 = ~n24726 ;
  assign y6451 = ~n24736 ;
  assign y6452 = n24737 ;
  assign y6453 = ~n24738 ;
  assign y6454 = ~n24740 ;
  assign y6455 = n24742 ;
  assign y6456 = n24744 ;
  assign y6457 = ~1'b0 ;
  assign y6458 = ~n24745 ;
  assign y6459 = n24748 ;
  assign y6460 = ~n24749 ;
  assign y6461 = n24750 ;
  assign y6462 = ~n24751 ;
  assign y6463 = ~1'b0 ;
  assign y6464 = ~n24753 ;
  assign y6465 = ~n24755 ;
  assign y6466 = ~n24756 ;
  assign y6467 = n24757 ;
  assign y6468 = n24759 ;
  assign y6469 = n24764 ;
  assign y6470 = ~1'b0 ;
  assign y6471 = ~1'b0 ;
  assign y6472 = ~n24767 ;
  assign y6473 = ~n24773 ;
  assign y6474 = n24776 ;
  assign y6475 = ~n24777 ;
  assign y6476 = n24781 ;
  assign y6477 = ~n24784 ;
  assign y6478 = ~n24786 ;
  assign y6479 = ~n24790 ;
  assign y6480 = ~1'b0 ;
  assign y6481 = n24792 ;
  assign y6482 = n24796 ;
  assign y6483 = n24799 ;
  assign y6484 = ~n24803 ;
  assign y6485 = n24804 ;
  assign y6486 = n24805 ;
  assign y6487 = ~n24807 ;
  assign y6488 = ~n24811 ;
  assign y6489 = n24813 ;
  assign y6490 = ~n24814 ;
  assign y6491 = ~n24815 ;
  assign y6492 = ~n24822 ;
  assign y6493 = n24826 ;
  assign y6494 = n24832 ;
  assign y6495 = n24834 ;
  assign y6496 = ~n24836 ;
  assign y6497 = ~n24839 ;
  assign y6498 = n24842 ;
  assign y6499 = ~n24845 ;
  assign y6500 = ~n24847 ;
  assign y6501 = n24855 ;
  assign y6502 = ~n24862 ;
  assign y6503 = n24863 ;
  assign y6504 = ~n24864 ;
  assign y6505 = n24870 ;
  assign y6506 = ~n24873 ;
  assign y6507 = ~n24875 ;
  assign y6508 = ~n24876 ;
  assign y6509 = ~n24878 ;
  assign y6510 = ~n24879 ;
  assign y6511 = ~1'b0 ;
  assign y6512 = ~1'b0 ;
  assign y6513 = ~n24884 ;
  assign y6514 = n24887 ;
  assign y6515 = n24898 ;
  assign y6516 = ~n24902 ;
  assign y6517 = n24905 ;
  assign y6518 = n24906 ;
  assign y6519 = n24910 ;
  assign y6520 = n24913 ;
  assign y6521 = n24919 ;
  assign y6522 = ~n24921 ;
  assign y6523 = ~n24923 ;
  assign y6524 = n24935 ;
  assign y6525 = n24938 ;
  assign y6526 = n24941 ;
  assign y6527 = n24947 ;
  assign y6528 = ~n24948 ;
  assign y6529 = ~n24949 ;
  assign y6530 = ~n24951 ;
  assign y6531 = ~n24953 ;
  assign y6532 = n12442 ;
  assign y6533 = n24955 ;
  assign y6534 = n24959 ;
  assign y6535 = ~n24968 ;
  assign y6536 = ~n24971 ;
  assign y6537 = ~n24972 ;
  assign y6538 = ~1'b0 ;
  assign y6539 = ~n24973 ;
  assign y6540 = n24977 ;
  assign y6541 = ~n24978 ;
  assign y6542 = n24980 ;
  assign y6543 = n24982 ;
  assign y6544 = ~n24986 ;
  assign y6545 = n24988 ;
  assign y6546 = n24990 ;
  assign y6547 = n24991 ;
  assign y6548 = ~n24994 ;
  assign y6549 = n24995 ;
  assign y6550 = n24996 ;
  assign y6551 = ~n25001 ;
  assign y6552 = n25002 ;
  assign y6553 = ~n25004 ;
  assign y6554 = n25006 ;
  assign y6555 = ~n25008 ;
  assign y6556 = n25009 ;
  assign y6557 = n25013 ;
  assign y6558 = ~n25016 ;
  assign y6559 = ~n25023 ;
  assign y6560 = ~n25024 ;
  assign y6561 = n25028 ;
  assign y6562 = ~n25030 ;
  assign y6563 = n25035 ;
  assign y6564 = n25036 ;
  assign y6565 = ~n25038 ;
  assign y6566 = n25040 ;
  assign y6567 = n25042 ;
  assign y6568 = n25048 ;
  assign y6569 = n25053 ;
  assign y6570 = ~n25058 ;
  assign y6571 = n25060 ;
  assign y6572 = n25063 ;
  assign y6573 = ~n25070 ;
  assign y6574 = ~1'b0 ;
  assign y6575 = ~n25071 ;
  assign y6576 = n25072 ;
  assign y6577 = ~n25076 ;
  assign y6578 = n25081 ;
  assign y6579 = ~n25085 ;
  assign y6580 = ~n25086 ;
  assign y6581 = ~n25088 ;
  assign y6582 = ~n25089 ;
  assign y6583 = ~n25092 ;
  assign y6584 = ~n25099 ;
  assign y6585 = n25101 ;
  assign y6586 = ~1'b0 ;
  assign y6587 = ~1'b0 ;
  assign y6588 = n25102 ;
  assign y6589 = ~n25103 ;
  assign y6590 = n25108 ;
  assign y6591 = n25110 ;
  assign y6592 = ~n25113 ;
  assign y6593 = n25118 ;
  assign y6594 = ~n25120 ;
  assign y6595 = ~1'b0 ;
  assign y6596 = ~1'b0 ;
  assign y6597 = n25128 ;
  assign y6598 = n25130 ;
  assign y6599 = n25131 ;
  assign y6600 = ~n25134 ;
  assign y6601 = ~n25136 ;
  assign y6602 = ~n25141 ;
  assign y6603 = n25142 ;
  assign y6604 = ~1'b0 ;
  assign y6605 = ~n25144 ;
  assign y6606 = n25145 ;
  assign y6607 = n25148 ;
  assign y6608 = ~n25151 ;
  assign y6609 = ~n25152 ;
  assign y6610 = ~n25154 ;
  assign y6611 = ~n25155 ;
  assign y6612 = ~n25156 ;
  assign y6613 = n25157 ;
  assign y6614 = ~n25158 ;
  assign y6615 = n25159 ;
  assign y6616 = ~n25164 ;
  assign y6617 = ~n25165 ;
  assign y6618 = ~n25166 ;
  assign y6619 = ~n25169 ;
  assign y6620 = n25170 ;
  assign y6621 = ~1'b0 ;
  assign y6622 = n25175 ;
  assign y6623 = ~n25177 ;
  assign y6624 = ~n24183 ;
  assign y6625 = ~n25183 ;
  assign y6626 = n25187 ;
  assign y6627 = n25188 ;
  assign y6628 = n25190 ;
  assign y6629 = n25192 ;
  assign y6630 = ~1'b0 ;
  assign y6631 = ~1'b0 ;
  assign y6632 = ~n25194 ;
  assign y6633 = ~n25195 ;
  assign y6634 = ~n25202 ;
  assign y6635 = n25204 ;
  assign y6636 = ~n25205 ;
  assign y6637 = ~n25207 ;
  assign y6638 = n25214 ;
  assign y6639 = ~n25218 ;
  assign y6640 = n25220 ;
  assign y6641 = n25225 ;
  assign y6642 = ~n25227 ;
  assign y6643 = ~n25229 ;
  assign y6644 = ~n25232 ;
  assign y6645 = n25233 ;
  assign y6646 = ~n25234 ;
  assign y6647 = ~n25236 ;
  assign y6648 = n25238 ;
  assign y6649 = ~n25250 ;
  assign y6650 = n25253 ;
  assign y6651 = ~1'b0 ;
  assign y6652 = ~n25257 ;
  assign y6653 = n25259 ;
  assign y6654 = ~n9961 ;
  assign y6655 = n25261 ;
  assign y6656 = ~n25262 ;
  assign y6657 = n25271 ;
  assign y6658 = ~n25274 ;
  assign y6659 = ~n25279 ;
  assign y6660 = ~n25281 ;
  assign y6661 = n25282 ;
  assign y6662 = ~n25284 ;
  assign y6663 = ~n25287 ;
  assign y6664 = ~n25289 ;
  assign y6665 = n25290 ;
  assign y6666 = ~1'b0 ;
  assign y6667 = ~n25291 ;
  assign y6668 = n25295 ;
  assign y6669 = ~n13770 ;
  assign y6670 = ~n25296 ;
  assign y6671 = ~n25299 ;
  assign y6672 = n25300 ;
  assign y6673 = n25301 ;
  assign y6674 = ~n25304 ;
  assign y6675 = ~1'b0 ;
  assign y6676 = n25308 ;
  assign y6677 = ~n25309 ;
  assign y6678 = ~n25314 ;
  assign y6679 = n25317 ;
  assign y6680 = n25319 ;
  assign y6681 = ~n25322 ;
  assign y6682 = ~n25324 ;
  assign y6683 = n25326 ;
  assign y6684 = n25330 ;
  assign y6685 = ~n25331 ;
  assign y6686 = n25332 ;
  assign y6687 = n25334 ;
  assign y6688 = ~n25337 ;
  assign y6689 = ~n25339 ;
  assign y6690 = n25345 ;
  assign y6691 = ~n25349 ;
  assign y6692 = n25351 ;
  assign y6693 = n25353 ;
  assign y6694 = ~n25354 ;
  assign y6695 = ~n25358 ;
  assign y6696 = n25365 ;
  assign y6697 = ~1'b0 ;
  assign y6698 = ~n25368 ;
  assign y6699 = n25369 ;
  assign y6700 = ~n25372 ;
  assign y6701 = n25375 ;
  assign y6702 = n25378 ;
  assign y6703 = n25379 ;
  assign y6704 = n25382 ;
  assign y6705 = n25383 ;
  assign y6706 = n25385 ;
  assign y6707 = ~n25387 ;
  assign y6708 = n25388 ;
  assign y6709 = n25391 ;
  assign y6710 = n25395 ;
  assign y6711 = n25400 ;
  assign y6712 = n25406 ;
  assign y6713 = ~1'b0 ;
  assign y6714 = ~n25407 ;
  assign y6715 = ~n25408 ;
  assign y6716 = ~n25413 ;
  assign y6717 = n25418 ;
  assign y6718 = ~n25420 ;
  assign y6719 = ~1'b0 ;
  assign y6720 = ~n25422 ;
  assign y6721 = n25424 ;
  assign y6722 = ~n25426 ;
  assign y6723 = ~n25432 ;
  assign y6724 = n25434 ;
  assign y6725 = n25437 ;
  assign y6726 = n25438 ;
  assign y6727 = ~n25444 ;
  assign y6728 = ~n25445 ;
  assign y6729 = ~1'b0 ;
  assign y6730 = n25448 ;
  assign y6731 = ~n25449 ;
  assign y6732 = n25450 ;
  assign y6733 = ~n25453 ;
  assign y6734 = n25455 ;
  assign y6735 = n25456 ;
  assign y6736 = ~1'b0 ;
  assign y6737 = ~n25460 ;
  assign y6738 = ~n25462 ;
  assign y6739 = ~n25463 ;
  assign y6740 = ~n25466 ;
  assign y6741 = ~n25467 ;
  assign y6742 = n25470 ;
  assign y6743 = n25472 ;
  assign y6744 = ~n25473 ;
  assign y6745 = ~1'b0 ;
  assign y6746 = ~n25475 ;
  assign y6747 = n25478 ;
  assign y6748 = n25485 ;
  assign y6749 = ~n25490 ;
  assign y6750 = n25491 ;
  assign y6751 = n25497 ;
  assign y6752 = n25501 ;
  assign y6753 = ~n25502 ;
  assign y6754 = n25504 ;
  assign y6755 = ~1'b0 ;
  assign y6756 = n25507 ;
  assign y6757 = n25515 ;
  assign y6758 = n25517 ;
  assign y6759 = ~n25520 ;
  assign y6760 = ~n25521 ;
  assign y6761 = ~n25523 ;
  assign y6762 = n25526 ;
  assign y6763 = n25535 ;
  assign y6764 = n25536 ;
  assign y6765 = ~1'b0 ;
  assign y6766 = ~1'b0 ;
  assign y6767 = ~n25542 ;
  assign y6768 = ~n25547 ;
  assign y6769 = n25548 ;
  assign y6770 = ~n25551 ;
  assign y6771 = n1596 ;
  assign y6772 = ~n25552 ;
  assign y6773 = ~n25554 ;
  assign y6774 = n25557 ;
  assign y6775 = ~n25560 ;
  assign y6776 = ~n25561 ;
  assign y6777 = n25563 ;
  assign y6778 = ~1'b0 ;
  assign y6779 = n25564 ;
  assign y6780 = ~n25565 ;
  assign y6781 = ~n25567 ;
  assign y6782 = n25568 ;
  assign y6783 = ~n25571 ;
  assign y6784 = ~n25577 ;
  assign y6785 = n25582 ;
  assign y6786 = ~n25585 ;
  assign y6787 = ~n25589 ;
  assign y6788 = ~n25591 ;
  assign y6789 = n25594 ;
  assign y6790 = n25596 ;
  assign y6791 = n25599 ;
  assign y6792 = ~n25600 ;
  assign y6793 = ~n25601 ;
  assign y6794 = ~n25603 ;
  assign y6795 = n25607 ;
  assign y6796 = n25614 ;
  assign y6797 = ~n25616 ;
  assign y6798 = ~n25620 ;
  assign y6799 = ~n25622 ;
  assign y6800 = n25624 ;
  assign y6801 = ~n25626 ;
  assign y6802 = n25628 ;
  assign y6803 = ~n25631 ;
  assign y6804 = n25632 ;
  assign y6805 = n25636 ;
  assign y6806 = ~n25638 ;
  assign y6807 = ~1'b0 ;
  assign y6808 = ~n25639 ;
  assign y6809 = ~n25642 ;
  assign y6810 = ~n25643 ;
  assign y6811 = ~n25648 ;
  assign y6812 = ~n25655 ;
  assign y6813 = n25656 ;
  assign y6814 = ~n25658 ;
  assign y6815 = n25660 ;
  assign y6816 = ~n25664 ;
  assign y6817 = n25668 ;
  assign y6818 = ~n25669 ;
  assign y6819 = n25671 ;
  assign y6820 = ~n25673 ;
  assign y6821 = ~n25680 ;
  assign y6822 = n25686 ;
  assign y6823 = n25691 ;
  assign y6824 = n25698 ;
  assign y6825 = n25700 ;
  assign y6826 = n25701 ;
  assign y6827 = ~n25702 ;
  assign y6828 = ~n25705 ;
  assign y6829 = ~n25709 ;
  assign y6830 = ~n25715 ;
  assign y6831 = n25716 ;
  assign y6832 = n25719 ;
  assign y6833 = ~n25724 ;
  assign y6834 = ~n25726 ;
  assign y6835 = ~n25729 ;
  assign y6836 = ~n25730 ;
  assign y6837 = n25731 ;
  assign y6838 = n25734 ;
  assign y6839 = ~n25737 ;
  assign y6840 = n25738 ;
  assign y6841 = ~n25741 ;
  assign y6842 = n25743 ;
  assign y6843 = ~n25745 ;
  assign y6844 = n25746 ;
  assign y6845 = n25750 ;
  assign y6846 = n25752 ;
  assign y6847 = n25753 ;
  assign y6848 = ~n25758 ;
  assign y6849 = ~n25762 ;
  assign y6850 = n25765 ;
  assign y6851 = n25768 ;
  assign y6852 = ~1'b0 ;
  assign y6853 = ~n25769 ;
  assign y6854 = n25770 ;
  assign y6855 = n25771 ;
  assign y6856 = ~n25775 ;
  assign y6857 = ~n25776 ;
  assign y6858 = n25778 ;
  assign y6859 = n25782 ;
  assign y6860 = n25788 ;
  assign y6861 = ~1'b0 ;
  assign y6862 = ~n25791 ;
  assign y6863 = ~n25796 ;
  assign y6864 = ~n25799 ;
  assign y6865 = ~n25800 ;
  assign y6866 = ~n25801 ;
  assign y6867 = n25804 ;
  assign y6868 = ~n25805 ;
  assign y6869 = ~n25807 ;
  assign y6870 = n25812 ;
  assign y6871 = ~n25815 ;
  assign y6872 = n25816 ;
  assign y6873 = ~n25821 ;
  assign y6874 = n25824 ;
  assign y6875 = ~n25827 ;
  assign y6876 = n25830 ;
  assign y6877 = ~n25832 ;
  assign y6878 = n25833 ;
  assign y6879 = n25842 ;
  assign y6880 = n25843 ;
  assign y6881 = n25844 ;
  assign y6882 = n25849 ;
  assign y6883 = ~n25851 ;
  assign y6884 = ~1'b0 ;
  assign y6885 = n25853 ;
  assign y6886 = ~n25855 ;
  assign y6887 = ~n25858 ;
  assign y6888 = ~n25859 ;
  assign y6889 = ~n25860 ;
  assign y6890 = n25861 ;
  assign y6891 = n25862 ;
  assign y6892 = n25864 ;
  assign y6893 = ~n25866 ;
  assign y6894 = ~n25874 ;
  assign y6895 = ~n25879 ;
  assign y6896 = n25880 ;
  assign y6897 = n25881 ;
  assign y6898 = ~n25883 ;
  assign y6899 = n25885 ;
  assign y6900 = ~n25893 ;
  assign y6901 = ~n25894 ;
  assign y6902 = ~1'b0 ;
  assign y6903 = ~1'b0 ;
  assign y6904 = n25896 ;
  assign y6905 = n25899 ;
  assign y6906 = ~1'b0 ;
  assign y6907 = ~n25900 ;
  assign y6908 = ~n25904 ;
  assign y6909 = ~n25907 ;
  assign y6910 = n25910 ;
  assign y6911 = ~n25912 ;
  assign y6912 = ~n25913 ;
  assign y6913 = n25915 ;
  assign y6914 = ~1'b0 ;
  assign y6915 = ~n25917 ;
  assign y6916 = n25918 ;
  assign y6917 = ~n25927 ;
  assign y6918 = ~n25932 ;
  assign y6919 = n25935 ;
  assign y6920 = ~n25937 ;
  assign y6921 = ~1'b0 ;
  assign y6922 = ~n25938 ;
  assign y6923 = ~n25944 ;
  assign y6924 = n25948 ;
  assign y6925 = ~n25949 ;
  assign y6926 = ~n25950 ;
  assign y6927 = ~n25952 ;
  assign y6928 = n25953 ;
  assign y6929 = ~n25955 ;
  assign y6930 = ~n25957 ;
  assign y6931 = ~n25959 ;
  assign y6932 = ~n25962 ;
  assign y6933 = ~n25963 ;
  assign y6934 = n25964 ;
  assign y6935 = ~n25969 ;
  assign y6936 = ~n25970 ;
  assign y6937 = n25973 ;
  assign y6938 = ~n25976 ;
  assign y6939 = ~n25977 ;
  assign y6940 = ~n25978 ;
  assign y6941 = n25981 ;
  assign y6942 = ~n25983 ;
  assign y6943 = ~n25986 ;
  assign y6944 = ~n25991 ;
  assign y6945 = ~n25995 ;
  assign y6946 = ~1'b0 ;
  assign y6947 = ~n26004 ;
  assign y6948 = ~n26005 ;
  assign y6949 = n26006 ;
  assign y6950 = ~n26007 ;
  assign y6951 = n26015 ;
  assign y6952 = n26019 ;
  assign y6953 = ~n26021 ;
  assign y6954 = ~n26024 ;
  assign y6955 = ~n26027 ;
  assign y6956 = n26029 ;
  assign y6957 = ~n26030 ;
  assign y6958 = ~n26034 ;
  assign y6959 = n26035 ;
  assign y6960 = n26038 ;
  assign y6961 = ~n26042 ;
  assign y6962 = n26044 ;
  assign y6963 = ~1'b0 ;
  assign y6964 = n26054 ;
  assign y6965 = n26063 ;
  assign y6966 = ~n26064 ;
  assign y6967 = n26065 ;
  assign y6968 = ~n26068 ;
  assign y6969 = ~n26069 ;
  assign y6970 = n26073 ;
  assign y6971 = n26076 ;
  assign y6972 = n17302 ;
  assign y6973 = n26077 ;
  assign y6974 = ~n26079 ;
  assign y6975 = ~n13476 ;
  assign y6976 = ~n26080 ;
  assign y6977 = n26083 ;
  assign y6978 = ~n26085 ;
  assign y6979 = ~n26088 ;
  assign y6980 = ~n26091 ;
  assign y6981 = ~n26094 ;
  assign y6982 = ~n26095 ;
  assign y6983 = n26097 ;
  assign y6984 = n26099 ;
  assign y6985 = n26104 ;
  assign y6986 = ~n26107 ;
  assign y6987 = ~n26110 ;
  assign y6988 = n26114 ;
  assign y6989 = ~n26121 ;
  assign y6990 = ~n26122 ;
  assign y6991 = ~n26125 ;
  assign y6992 = ~1'b0 ;
  assign y6993 = n26128 ;
  assign y6994 = n26131 ;
  assign y6995 = ~n26133 ;
  assign y6996 = n26135 ;
  assign y6997 = n26136 ;
  assign y6998 = n26137 ;
  assign y6999 = ~n26140 ;
  assign y7000 = ~n26142 ;
  assign y7001 = ~1'b0 ;
  assign y7002 = n26144 ;
  assign y7003 = n26145 ;
  assign y7004 = ~n26146 ;
  assign y7005 = ~n26150 ;
  assign y7006 = ~n26151 ;
  assign y7007 = ~n26152 ;
  assign y7008 = n26154 ;
  assign y7009 = n26158 ;
  assign y7010 = ~n26161 ;
  assign y7011 = ~n26166 ;
  assign y7012 = n26172 ;
  assign y7013 = ~n26174 ;
  assign y7014 = n26176 ;
  assign y7015 = n26177 ;
  assign y7016 = n26181 ;
  assign y7017 = ~n26183 ;
  assign y7018 = ~1'b0 ;
  assign y7019 = n26187 ;
  assign y7020 = n26188 ;
  assign y7021 = ~n26191 ;
  assign y7022 = n26193 ;
  assign y7023 = n26195 ;
  assign y7024 = ~1'b0 ;
  assign y7025 = ~n26199 ;
  assign y7026 = ~n26201 ;
  assign y7027 = n26204 ;
  assign y7028 = n26205 ;
  assign y7029 = n26209 ;
  assign y7030 = ~n26212 ;
  assign y7031 = ~n26214 ;
  assign y7032 = ~n26219 ;
  assign y7033 = n26223 ;
  assign y7034 = ~n26227 ;
  assign y7035 = n26229 ;
  assign y7036 = ~n26230 ;
  assign y7037 = n26232 ;
  assign y7038 = n26234 ;
  assign y7039 = ~n26238 ;
  assign y7040 = ~n26239 ;
  assign y7041 = ~n26241 ;
  assign y7042 = ~1'b0 ;
  assign y7043 = ~1'b0 ;
  assign y7044 = n26242 ;
  assign y7045 = ~n26245 ;
  assign y7046 = n26246 ;
  assign y7047 = n26248 ;
  assign y7048 = n26252 ;
  assign y7049 = n26253 ;
  assign y7050 = ~n26256 ;
  assign y7051 = n26261 ;
  assign y7052 = ~1'b0 ;
  assign y7053 = ~1'b0 ;
  assign y7054 = n26264 ;
  assign y7055 = ~n26266 ;
  assign y7056 = ~n26267 ;
  assign y7057 = ~n26268 ;
  assign y7058 = ~n26273 ;
  assign y7059 = ~n26274 ;
  assign y7060 = ~n26275 ;
  assign y7061 = ~n26278 ;
  assign y7062 = ~n26280 ;
  assign y7063 = n26281 ;
  assign y7064 = ~n26282 ;
  assign y7065 = n26283 ;
  assign y7066 = ~n26285 ;
  assign y7067 = ~n26289 ;
  assign y7068 = n26292 ;
  assign y7069 = n26295 ;
  assign y7070 = ~n26297 ;
  assign y7071 = ~n26301 ;
  assign y7072 = ~n26302 ;
  assign y7073 = ~n26303 ;
  assign y7074 = n26311 ;
  assign y7075 = n26314 ;
  assign y7076 = n26315 ;
  assign y7077 = ~n26319 ;
  assign y7078 = n26321 ;
  assign y7079 = n26323 ;
  assign y7080 = ~n26324 ;
  assign y7081 = ~n26326 ;
  assign y7082 = n26330 ;
  assign y7083 = n26332 ;
  assign y7084 = n26333 ;
  assign y7085 = n26341 ;
  assign y7086 = ~n26343 ;
  assign y7087 = n26346 ;
  assign y7088 = ~n26351 ;
  assign y7089 = ~n26352 ;
  assign y7090 = ~n26355 ;
  assign y7091 = ~n26357 ;
  assign y7092 = ~1'b0 ;
  assign y7093 = n26359 ;
  assign y7094 = ~n26360 ;
  assign y7095 = ~n26363 ;
  assign y7096 = ~n26366 ;
  assign y7097 = ~n26367 ;
  assign y7098 = n26368 ;
  assign y7099 = ~n26372 ;
  assign y7100 = ~1'b0 ;
  assign y7101 = n26374 ;
  assign y7102 = ~n26375 ;
  assign y7103 = n26376 ;
  assign y7104 = ~n26378 ;
  assign y7105 = ~n26379 ;
  assign y7106 = n26384 ;
  assign y7107 = ~n26386 ;
  assign y7108 = ~n26387 ;
  assign y7109 = n26398 ;
  assign y7110 = ~n26400 ;
  assign y7111 = n26407 ;
  assign y7112 = n26410 ;
  assign y7113 = ~n26413 ;
  assign y7114 = n26415 ;
  assign y7115 = ~n26416 ;
  assign y7116 = ~n26419 ;
  assign y7117 = ~n26421 ;
  assign y7118 = n26428 ;
  assign y7119 = n26429 ;
  assign y7120 = n26431 ;
  assign y7121 = n26435 ;
  assign y7122 = ~1'b0 ;
  assign y7123 = ~n26437 ;
  assign y7124 = ~n26439 ;
  assign y7125 = n26445 ;
  assign y7126 = n26452 ;
  assign y7127 = ~n26453 ;
  assign y7128 = ~n26455 ;
  assign y7129 = ~n26458 ;
  assign y7130 = ~n26459 ;
  assign y7131 = n26462 ;
  assign y7132 = ~n26464 ;
  assign y7133 = n26465 ;
  assign y7134 = n26468 ;
  assign y7135 = n26470 ;
  assign y7136 = ~n26471 ;
  assign y7137 = n26476 ;
  assign y7138 = ~n26482 ;
  assign y7139 = ~n26485 ;
  assign y7140 = ~1'b0 ;
  assign y7141 = n26487 ;
  assign y7142 = ~n26489 ;
  assign y7143 = ~n26492 ;
  assign y7144 = ~n26493 ;
  assign y7145 = n26499 ;
  assign y7146 = n26502 ;
  assign y7147 = ~n26503 ;
  assign y7148 = ~n26505 ;
  assign y7149 = ~n26506 ;
  assign y7150 = ~n26507 ;
  assign y7151 = n26510 ;
  assign y7152 = ~n26511 ;
  assign y7153 = n26514 ;
  assign y7154 = n26517 ;
  assign y7155 = n26518 ;
  assign y7156 = ~n26519 ;
  assign y7157 = ~n26520 ;
  assign y7158 = ~n26523 ;
  assign y7159 = ~1'b0 ;
  assign y7160 = ~1'b0 ;
  assign y7161 = n26524 ;
  assign y7162 = ~n26526 ;
  assign y7163 = n26532 ;
  assign y7164 = n26536 ;
  assign y7165 = n26541 ;
  assign y7166 = ~n26542 ;
  assign y7167 = ~n26545 ;
  assign y7168 = ~1'b0 ;
  assign y7169 = ~1'b0 ;
  assign y7170 = n26548 ;
  assign y7171 = ~n26549 ;
  assign y7172 = ~n26551 ;
  assign y7173 = ~1'b0 ;
  assign y7174 = ~n26552 ;
  assign y7175 = n26554 ;
  assign y7176 = ~n26555 ;
  assign y7177 = n26562 ;
  assign y7178 = ~n26566 ;
  assign y7179 = ~n26567 ;
  assign y7180 = ~n26570 ;
  assign y7181 = ~n26576 ;
  assign y7182 = n26578 ;
  assign y7183 = ~n26582 ;
  assign y7184 = ~n26589 ;
  assign y7185 = n26594 ;
  assign y7186 = n26596 ;
  assign y7187 = ~n26600 ;
  assign y7188 = ~n26604 ;
  assign y7189 = ~n26605 ;
  assign y7190 = n26606 ;
  assign y7191 = ~n26607 ;
  assign y7192 = n26611 ;
  assign y7193 = ~n26614 ;
  assign y7194 = ~n26617 ;
  assign y7195 = ~1'b0 ;
  assign y7196 = n26618 ;
  assign y7197 = ~n26622 ;
  assign y7198 = n26627 ;
  assign y7199 = ~n11034 ;
  assign y7200 = ~n26628 ;
  assign y7201 = ~n26632 ;
  assign y7202 = ~n26634 ;
  assign y7203 = n26637 ;
  assign y7204 = n26638 ;
  assign y7205 = ~n26641 ;
  assign y7206 = n26644 ;
  assign y7207 = ~n26648 ;
  assign y7208 = ~n26649 ;
  assign y7209 = ~n26653 ;
  assign y7210 = n26657 ;
  assign y7211 = ~n26660 ;
  assign y7212 = ~n26662 ;
  assign y7213 = ~n26664 ;
  assign y7214 = n26669 ;
  assign y7215 = n26671 ;
  assign y7216 = ~n26672 ;
  assign y7217 = ~n26673 ;
  assign y7218 = ~n26675 ;
  assign y7219 = ~1'b0 ;
  assign y7220 = ~n26677 ;
  assign y7221 = ~n26682 ;
  assign y7222 = n26684 ;
  assign y7223 = ~n26686 ;
  assign y7224 = ~n26691 ;
  assign y7225 = n26694 ;
  assign y7226 = ~n26697 ;
  assign y7227 = ~1'b0 ;
  assign y7228 = ~1'b0 ;
  assign y7229 = ~n26700 ;
  assign y7230 = ~n26701 ;
  assign y7231 = ~n26702 ;
  assign y7232 = n26704 ;
  assign y7233 = n26707 ;
  assign y7234 = n26712 ;
  assign y7235 = n26715 ;
  assign y7236 = ~1'b0 ;
  assign y7237 = ~n26717 ;
  assign y7238 = n26720 ;
  assign y7239 = n26722 ;
  assign y7240 = ~n26723 ;
  assign y7241 = n26725 ;
  assign y7242 = n26730 ;
  assign y7243 = ~n26735 ;
  assign y7244 = ~n26737 ;
  assign y7245 = n26738 ;
  assign y7246 = n26742 ;
  assign y7247 = ~n26744 ;
  assign y7248 = n26745 ;
  assign y7249 = ~n26749 ;
  assign y7250 = ~n26752 ;
  assign y7251 = ~n26755 ;
  assign y7252 = n26759 ;
  assign y7253 = ~n26763 ;
  assign y7254 = ~1'b0 ;
  assign y7255 = ~n26765 ;
  assign y7256 = n26766 ;
  assign y7257 = n26767 ;
  assign y7258 = n26768 ;
  assign y7259 = n26771 ;
  assign y7260 = n26774 ;
  assign y7261 = ~n26779 ;
  assign y7262 = n26780 ;
  assign y7263 = ~n26785 ;
  assign y7264 = ~n26788 ;
  assign y7265 = ~n26789 ;
  assign y7266 = ~n26791 ;
  assign y7267 = ~n26793 ;
  assign y7268 = n26794 ;
  assign y7269 = n26796 ;
  assign y7270 = ~n26800 ;
  assign y7271 = ~n26801 ;
  assign y7272 = n26806 ;
  assign y7273 = n26810 ;
  assign y7274 = n26813 ;
  assign y7275 = n26817 ;
  assign y7276 = n26819 ;
  assign y7277 = n26823 ;
  assign y7278 = ~n26826 ;
  assign y7279 = n26833 ;
  assign y7280 = n26834 ;
  assign y7281 = ~1'b0 ;
  assign y7282 = ~n26837 ;
  assign y7283 = ~n26838 ;
  assign y7284 = n26841 ;
  assign y7285 = n26842 ;
  assign y7286 = ~n26845 ;
  assign y7287 = ~n26846 ;
  assign y7288 = n26850 ;
  assign y7289 = ~n26852 ;
  assign y7290 = n26854 ;
  assign y7291 = n26857 ;
  assign y7292 = ~1'b0 ;
  assign y7293 = ~n26859 ;
  assign y7294 = ~n26861 ;
  assign y7295 = n26862 ;
  assign y7296 = ~n26866 ;
  assign y7297 = ~n26868 ;
  assign y7298 = n26869 ;
  assign y7299 = ~1'b0 ;
  assign y7300 = ~n26871 ;
  assign y7301 = n26872 ;
  assign y7302 = n26875 ;
  assign y7303 = ~n26878 ;
  assign y7304 = n26879 ;
  assign y7305 = n26880 ;
  assign y7306 = ~n26882 ;
  assign y7307 = n26884 ;
  assign y7308 = n26888 ;
  assign y7309 = ~1'b0 ;
  assign y7310 = n26889 ;
  assign y7311 = n26891 ;
  assign y7312 = ~n26892 ;
  assign y7313 = ~n26893 ;
  assign y7314 = ~n26896 ;
  assign y7315 = ~1'b0 ;
  assign y7316 = n26901 ;
  assign y7317 = n26904 ;
  assign y7318 = n26911 ;
  assign y7319 = n26915 ;
  assign y7320 = ~n26918 ;
  assign y7321 = ~n26919 ;
  assign y7322 = ~n26921 ;
  assign y7323 = ~n26925 ;
  assign y7324 = n26926 ;
  assign y7325 = n26928 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = ~n26931 ;
  assign y7328 = ~n26932 ;
  assign y7329 = ~n26934 ;
  assign y7330 = n26935 ;
  assign y7331 = ~n26939 ;
  assign y7332 = n26941 ;
  assign y7333 = ~n26942 ;
  assign y7334 = ~1'b0 ;
  assign y7335 = ~1'b0 ;
  assign y7336 = ~1'b0 ;
  assign y7337 = n26947 ;
  assign y7338 = ~n26950 ;
  assign y7339 = ~n26951 ;
  assign y7340 = ~n26952 ;
  assign y7341 = n26953 ;
  assign y7342 = ~n26956 ;
  assign y7343 = ~1'b0 ;
  assign y7344 = n26958 ;
  assign y7345 = n26959 ;
  assign y7346 = ~n26960 ;
  assign y7347 = ~n26962 ;
  assign y7348 = ~n26965 ;
  assign y7349 = n26966 ;
  assign y7350 = ~n26971 ;
  assign y7351 = n26974 ;
  assign y7352 = ~n26976 ;
  assign y7353 = n26980 ;
  assign y7354 = n26981 ;
  assign y7355 = n26983 ;
  assign y7356 = n26989 ;
  assign y7357 = ~n26992 ;
  assign y7358 = ~n26996 ;
  assign y7359 = n26998 ;
  assign y7360 = ~1'b0 ;
  assign y7361 = n27000 ;
  assign y7362 = n27005 ;
  assign y7363 = n27006 ;
  assign y7364 = ~n27009 ;
  assign y7365 = ~n27011 ;
  assign y7366 = ~n27012 ;
  assign y7367 = n27014 ;
  assign y7368 = ~n27015 ;
  assign y7369 = ~n27017 ;
  assign y7370 = ~n27020 ;
  assign y7371 = n27022 ;
  assign y7372 = n27029 ;
  assign y7373 = ~n27030 ;
  assign y7374 = ~n27031 ;
  assign y7375 = ~n27033 ;
  assign y7376 = n27034 ;
  assign y7377 = ~n27038 ;
  assign y7378 = n27039 ;
  assign y7379 = ~1'b0 ;
  assign y7380 = ~1'b0 ;
  assign y7381 = n27044 ;
  assign y7382 = ~n27049 ;
  assign y7383 = n27053 ;
  assign y7384 = n27058 ;
  assign y7385 = n27059 ;
  assign y7386 = ~n27062 ;
  assign y7387 = n27066 ;
  assign y7388 = n27067 ;
  assign y7389 = n27069 ;
  assign y7390 = ~1'b0 ;
  assign y7391 = ~1'b0 ;
  assign y7392 = ~n27072 ;
  assign y7393 = n27075 ;
  assign y7394 = ~n27076 ;
  assign y7395 = n27082 ;
  assign y7396 = n27084 ;
  assign y7397 = ~n27089 ;
  assign y7398 = n27091 ;
  assign y7399 = ~1'b0 ;
  assign y7400 = ~n27095 ;
  assign y7401 = n27096 ;
  assign y7402 = ~n27097 ;
  assign y7403 = n27098 ;
  assign y7404 = n27105 ;
  assign y7405 = n27108 ;
  assign y7406 = ~n27109 ;
  assign y7407 = n27111 ;
  assign y7408 = n27112 ;
  assign y7409 = ~n27113 ;
  assign y7410 = n27114 ;
  assign y7411 = ~n27115 ;
  assign y7412 = ~n27119 ;
  assign y7413 = ~n27120 ;
  assign y7414 = n27122 ;
  assign y7415 = n27125 ;
  assign y7416 = ~n27131 ;
  assign y7417 = n27134 ;
  assign y7418 = ~1'b0 ;
  assign y7419 = n27138 ;
  assign y7420 = n27140 ;
  assign y7421 = n27142 ;
  assign y7422 = ~n27144 ;
  assign y7423 = ~1'b0 ;
  assign y7424 = ~n27148 ;
  assign y7425 = ~1'b0 ;
  assign y7426 = n27151 ;
  assign y7427 = ~n27153 ;
  assign y7428 = n27158 ;
  assign y7429 = n27159 ;
  assign y7430 = n27161 ;
  assign y7431 = ~n27162 ;
  assign y7432 = n27163 ;
  assign y7433 = ~n27165 ;
  assign y7434 = ~n27166 ;
  assign y7435 = ~n27170 ;
  assign y7436 = n27174 ;
  assign y7437 = n27178 ;
  assign y7438 = n27180 ;
  assign y7439 = n27182 ;
  assign y7440 = n27183 ;
  assign y7441 = ~1'b0 ;
  assign y7442 = ~1'b0 ;
  assign y7443 = ~n27184 ;
  assign y7444 = n27186 ;
  assign y7445 = n27194 ;
  assign y7446 = n27197 ;
  assign y7447 = ~n27200 ;
  assign y7448 = ~n27203 ;
  assign y7449 = ~1'b0 ;
  assign y7450 = ~n27208 ;
  assign y7451 = ~n27209 ;
  assign y7452 = n27210 ;
  assign y7453 = ~n27211 ;
  assign y7454 = ~n20762 ;
  assign y7455 = n27215 ;
  assign y7456 = n27222 ;
  assign y7457 = n27224 ;
  assign y7458 = ~n27229 ;
  assign y7459 = ~n27231 ;
  assign y7460 = n27233 ;
  assign y7461 = ~1'b0 ;
  assign y7462 = n27236 ;
  assign y7463 = n27238 ;
  assign y7464 = n27240 ;
  assign y7465 = n27241 ;
  assign y7466 = n27242 ;
  assign y7467 = ~n27243 ;
  assign y7468 = ~n27247 ;
  assign y7469 = ~1'b0 ;
  assign y7470 = n27248 ;
  assign y7471 = n27249 ;
  assign y7472 = n27251 ;
  assign y7473 = n27252 ;
  assign y7474 = ~n27254 ;
  assign y7475 = n27256 ;
  assign y7476 = ~1'b0 ;
  assign y7477 = n27260 ;
  assign y7478 = n27262 ;
  assign y7479 = ~n27264 ;
  assign y7480 = n27265 ;
  assign y7481 = ~n27267 ;
  assign y7482 = n27269 ;
  assign y7483 = n27270 ;
  assign y7484 = ~n27272 ;
  assign y7485 = n27281 ;
  assign y7486 = ~1'b0 ;
  assign y7487 = n27286 ;
  assign y7488 = ~n27287 ;
  assign y7489 = ~1'b0 ;
  assign y7490 = n27288 ;
  assign y7491 = n27289 ;
  assign y7492 = n27295 ;
  assign y7493 = n27297 ;
  assign y7494 = n27298 ;
  assign y7495 = n27300 ;
  assign y7496 = ~1'b0 ;
  assign y7497 = ~n27301 ;
  assign y7498 = ~n27303 ;
  assign y7499 = n27304 ;
  assign y7500 = ~n27306 ;
  assign y7501 = n27309 ;
  assign y7502 = n27310 ;
  assign y7503 = ~n27315 ;
  assign y7504 = ~n27316 ;
  assign y7505 = n27319 ;
  assign y7506 = n27320 ;
  assign y7507 = ~n27325 ;
  assign y7508 = ~n27328 ;
  assign y7509 = n27335 ;
  assign y7510 = n27338 ;
  assign y7511 = n27339 ;
  assign y7512 = n27340 ;
  assign y7513 = n27344 ;
  assign y7514 = ~n27346 ;
  assign y7515 = n27350 ;
  assign y7516 = ~n27352 ;
  assign y7517 = ~n27357 ;
  assign y7518 = n27358 ;
  assign y7519 = ~n27362 ;
  assign y7520 = ~n27372 ;
  assign y7521 = ~n27377 ;
  assign y7522 = n27384 ;
  assign y7523 = n27385 ;
  assign y7524 = ~1'b0 ;
  assign y7525 = n27388 ;
  assign y7526 = n27393 ;
  assign y7527 = ~n27394 ;
  assign y7528 = ~n27395 ;
  assign y7529 = n27396 ;
  assign y7530 = n27398 ;
  assign y7531 = n27399 ;
  assign y7532 = ~n27404 ;
  assign y7533 = n27407 ;
  assign y7534 = ~n27408 ;
  assign y7535 = n27410 ;
  assign y7536 = ~n3429 ;
  assign y7537 = ~n27411 ;
  assign y7538 = ~n27414 ;
  assign y7539 = n27415 ;
  assign y7540 = n27420 ;
  assign y7541 = n27423 ;
  assign y7542 = n27425 ;
  assign y7543 = ~1'b0 ;
  assign y7544 = n27428 ;
  assign y7545 = n27430 ;
  assign y7546 = n27433 ;
  assign y7547 = n27435 ;
  assign y7548 = n27437 ;
  assign y7549 = ~n27439 ;
  assign y7550 = n27443 ;
  assign y7551 = n27454 ;
  assign y7552 = ~n27456 ;
  assign y7553 = ~n27457 ;
  assign y7554 = ~n27467 ;
  assign y7555 = ~n27469 ;
  assign y7556 = n27470 ;
  assign y7557 = ~n27471 ;
  assign y7558 = ~1'b0 ;
  assign y7559 = n27473 ;
  assign y7560 = ~n27475 ;
  assign y7561 = ~n27479 ;
  assign y7562 = ~n27481 ;
  assign y7563 = n27486 ;
  assign y7564 = n27497 ;
  assign y7565 = n27499 ;
  assign y7566 = n27503 ;
  assign y7567 = ~n27506 ;
  assign y7568 = n27510 ;
  assign y7569 = ~1'b0 ;
  assign y7570 = n27513 ;
  assign y7571 = ~n27514 ;
  assign y7572 = n27516 ;
  assign y7573 = ~n27518 ;
  assign y7574 = ~n27524 ;
  assign y7575 = n27525 ;
  assign y7576 = ~n27526 ;
  assign y7577 = ~n27528 ;
  assign y7578 = ~n27531 ;
  assign y7579 = ~n27533 ;
  assign y7580 = n27539 ;
  assign y7581 = ~n27543 ;
  assign y7582 = ~n27544 ;
  assign y7583 = ~n27545 ;
  assign y7584 = ~n27549 ;
  assign y7585 = ~n27550 ;
  assign y7586 = ~n27553 ;
  assign y7587 = ~n27556 ;
  assign y7588 = ~n27558 ;
  assign y7589 = ~n27561 ;
  assign y7590 = n27562 ;
  assign y7591 = ~n27566 ;
  assign y7592 = ~n27569 ;
  assign y7593 = n27570 ;
  assign y7594 = ~n27572 ;
  assign y7595 = ~n27573 ;
  assign y7596 = n27575 ;
  assign y7597 = ~1'b0 ;
  assign y7598 = ~n27576 ;
  assign y7599 = ~n27583 ;
  assign y7600 = n27584 ;
  assign y7601 = n27586 ;
  assign y7602 = ~n27587 ;
  assign y7603 = ~n27588 ;
  assign y7604 = ~n27593 ;
  assign y7605 = ~n27597 ;
  assign y7606 = ~n27598 ;
  assign y7607 = ~n27600 ;
  assign y7608 = ~n27603 ;
  assign y7609 = n27606 ;
  assign y7610 = n27607 ;
  assign y7611 = n27609 ;
  assign y7612 = n27612 ;
  assign y7613 = ~n27617 ;
  assign y7614 = ~n27619 ;
  assign y7615 = n27623 ;
  assign y7616 = n27626 ;
  assign y7617 = n27629 ;
  assign y7618 = ~n27632 ;
  assign y7619 = ~n27634 ;
  assign y7620 = n27636 ;
  assign y7621 = n27637 ;
  assign y7622 = n27638 ;
  assign y7623 = ~1'b0 ;
  assign y7624 = ~n27642 ;
  assign y7625 = n27646 ;
  assign y7626 = ~n27657 ;
  assign y7627 = n27660 ;
  assign y7628 = n27663 ;
  assign y7629 = ~n27665 ;
  assign y7630 = n816 ;
  assign y7631 = ~n27670 ;
  assign y7632 = ~1'b0 ;
  assign y7633 = ~n27673 ;
  assign y7634 = ~1'b0 ;
  assign y7635 = ~n27675 ;
  assign y7636 = ~n27677 ;
  assign y7637 = n27678 ;
  assign y7638 = n27680 ;
  assign y7639 = ~n27682 ;
  assign y7640 = n27687 ;
  assign y7641 = ~n27688 ;
  assign y7642 = ~n27692 ;
  assign y7643 = ~n27694 ;
  assign y7644 = ~1'b0 ;
  assign y7645 = n27695 ;
  assign y7646 = ~n27696 ;
  assign y7647 = n27697 ;
  assign y7648 = ~n27698 ;
  assign y7649 = ~n27701 ;
  assign y7650 = ~n27704 ;
  assign y7651 = n27707 ;
  assign y7652 = n27710 ;
  assign y7653 = n27719 ;
  assign y7654 = n27722 ;
  assign y7655 = ~n27723 ;
  assign y7656 = n27725 ;
  assign y7657 = ~n27726 ;
  assign y7658 = ~n27727 ;
  assign y7659 = n27731 ;
  assign y7660 = ~n27736 ;
  assign y7661 = ~n27739 ;
  assign y7662 = ~n27740 ;
  assign y7663 = ~1'b0 ;
  assign y7664 = ~n27746 ;
  assign y7665 = n27749 ;
  assign y7666 = ~n27750 ;
  assign y7667 = ~n27751 ;
  assign y7668 = n27752 ;
  assign y7669 = n27758 ;
  assign y7670 = n27761 ;
  assign y7671 = ~n27770 ;
  assign y7672 = n27772 ;
  assign y7673 = n27774 ;
  assign y7674 = ~n27777 ;
  assign y7675 = ~n27778 ;
  assign y7676 = n27780 ;
  assign y7677 = ~n27786 ;
  assign y7678 = n27789 ;
  assign y7679 = ~n27793 ;
  assign y7680 = n27796 ;
  assign y7681 = n27798 ;
  assign y7682 = n27800 ;
  assign y7683 = ~n27801 ;
  assign y7684 = n27803 ;
  assign y7685 = n27804 ;
  assign y7686 = n27807 ;
  assign y7687 = n27809 ;
  assign y7688 = ~n27812 ;
  assign y7689 = ~n27814 ;
  assign y7690 = n27824 ;
  assign y7691 = n27826 ;
  assign y7692 = n27828 ;
  assign y7693 = ~n27833 ;
  assign y7694 = ~n27834 ;
  assign y7695 = n27838 ;
  assign y7696 = n27839 ;
  assign y7697 = n27843 ;
  assign y7698 = ~n27845 ;
  assign y7699 = ~1'b0 ;
  assign y7700 = ~n27846 ;
  assign y7701 = n27847 ;
  assign y7702 = ~n27850 ;
  assign y7703 = ~n27851 ;
  assign y7704 = n27853 ;
  assign y7705 = n27854 ;
  assign y7706 = n27855 ;
  assign y7707 = ~n27859 ;
  assign y7708 = ~1'b0 ;
  assign y7709 = ~n27862 ;
  assign y7710 = n27864 ;
  assign y7711 = n27867 ;
  assign y7712 = n27870 ;
  assign y7713 = ~n27871 ;
  assign y7714 = n27872 ;
  assign y7715 = n27873 ;
  assign y7716 = ~n27876 ;
  assign y7717 = n27878 ;
  assign y7718 = n27882 ;
  assign y7719 = n27887 ;
  assign y7720 = ~n27888 ;
  assign y7721 = ~n27890 ;
  assign y7722 = n27891 ;
  assign y7723 = ~n27898 ;
  assign y7724 = ~n27899 ;
  assign y7725 = ~n27902 ;
  assign y7726 = n27905 ;
  assign y7727 = ~n27907 ;
  assign y7728 = ~n6517 ;
  assign y7729 = n27908 ;
  assign y7730 = n27911 ;
  assign y7731 = ~n27914 ;
  assign y7732 = n27915 ;
  assign y7733 = n27917 ;
  assign y7734 = ~n27918 ;
  assign y7735 = n27922 ;
  assign y7736 = ~1'b0 ;
  assign y7737 = ~n27923 ;
  assign y7738 = ~n27926 ;
  assign y7739 = ~n27929 ;
  assign y7740 = ~n27932 ;
  assign y7741 = ~n27933 ;
  assign y7742 = ~n27934 ;
  assign y7743 = ~1'b0 ;
  assign y7744 = n27935 ;
  assign y7745 = ~n27937 ;
  assign y7746 = ~n27939 ;
  assign y7747 = n19641 ;
  assign y7748 = ~n27940 ;
  assign y7749 = ~n27944 ;
  assign y7750 = ~n27945 ;
  assign y7751 = n27949 ;
  assign y7752 = n27952 ;
  assign y7753 = ~n27954 ;
  assign y7754 = n27957 ;
  assign y7755 = n27962 ;
  assign y7756 = ~n27964 ;
  assign y7757 = ~n27968 ;
  assign y7758 = n27969 ;
  assign y7759 = n27972 ;
  assign y7760 = n27974 ;
  assign y7761 = ~n27976 ;
  assign y7762 = ~n27981 ;
  assign y7763 = ~n27984 ;
  assign y7764 = n27989 ;
  assign y7765 = ~n27993 ;
  assign y7766 = ~n27995 ;
  assign y7767 = ~n27996 ;
  assign y7768 = ~1'b0 ;
  assign y7769 = n27998 ;
  assign y7770 = ~1'b0 ;
  assign y7771 = n28000 ;
  assign y7772 = ~n28004 ;
  assign y7773 = n28005 ;
  assign y7774 = n28006 ;
  assign y7775 = ~n28012 ;
  assign y7776 = ~n28014 ;
  assign y7777 = ~1'b0 ;
  assign y7778 = ~n28016 ;
  assign y7779 = n28017 ;
  assign y7780 = n28020 ;
  assign y7781 = n28023 ;
  assign y7782 = ~n28025 ;
  assign y7783 = n28026 ;
  assign y7784 = n28028 ;
  assign y7785 = n28029 ;
  assign y7786 = ~n28031 ;
  assign y7787 = ~n28039 ;
  assign y7788 = ~n28041 ;
  assign y7789 = ~n28042 ;
  assign y7790 = ~n28050 ;
  assign y7791 = n28052 ;
  assign y7792 = ~n28053 ;
  assign y7793 = n28056 ;
  assign y7794 = ~1'b0 ;
  assign y7795 = n28059 ;
  assign y7796 = n28061 ;
  assign y7797 = ~n28062 ;
  assign y7798 = ~n28063 ;
  assign y7799 = ~n28064 ;
  assign y7800 = ~n28067 ;
  assign y7801 = ~n28068 ;
  assign y7802 = n28071 ;
  assign y7803 = n28074 ;
  assign y7804 = n28077 ;
  assign y7805 = ~n28085 ;
  assign y7806 = ~n28087 ;
  assign y7807 = ~n28091 ;
  assign y7808 = ~n28096 ;
  assign y7809 = n28100 ;
  assign y7810 = n28102 ;
  assign y7811 = ~n28104 ;
  assign y7812 = ~n28106 ;
  assign y7813 = ~n28110 ;
  assign y7814 = ~n28113 ;
  assign y7815 = ~n28115 ;
  assign y7816 = n28118 ;
  assign y7817 = ~n28124 ;
  assign y7818 = n28126 ;
  assign y7819 = n28130 ;
  assign y7820 = ~n28131 ;
  assign y7821 = ~n28137 ;
  assign y7822 = ~1'b0 ;
  assign y7823 = ~n28141 ;
  assign y7824 = ~n28142 ;
  assign y7825 = ~n28146 ;
  assign y7826 = ~n28148 ;
  assign y7827 = n28149 ;
  assign y7828 = ~n28153 ;
  assign y7829 = n28154 ;
  assign y7830 = ~n28155 ;
  assign y7831 = ~n28157 ;
  assign y7832 = n28159 ;
  assign y7833 = n28162 ;
  assign y7834 = ~n28170 ;
  assign y7835 = n28174 ;
  assign y7836 = n28175 ;
  assign y7837 = ~n28177 ;
  assign y7838 = n28178 ;
  assign y7839 = n28179 ;
  assign y7840 = n28185 ;
  assign y7841 = n28187 ;
  assign y7842 = ~n28189 ;
  assign y7843 = ~n28194 ;
  assign y7844 = ~n28196 ;
  assign y7845 = ~n28197 ;
  assign y7846 = n28201 ;
  assign y7847 = ~n28206 ;
  assign y7848 = n28208 ;
  assign y7849 = ~1'b0 ;
  assign y7850 = n28210 ;
  assign y7851 = ~n28213 ;
  assign y7852 = ~n28214 ;
  assign y7853 = n28217 ;
  assign y7854 = ~n28221 ;
  assign y7855 = ~n28224 ;
  assign y7856 = n28228 ;
  assign y7857 = ~n28230 ;
  assign y7858 = n28232 ;
  assign y7859 = ~1'b0 ;
  assign y7860 = ~1'b0 ;
  assign y7861 = ~n28233 ;
  assign y7862 = ~n28234 ;
  assign y7863 = n28235 ;
  assign y7864 = ~n28236 ;
  assign y7865 = n28242 ;
  assign y7866 = ~n28243 ;
  assign y7867 = ~n28244 ;
  assign y7868 = n28251 ;
  assign y7869 = n15543 ;
  assign y7870 = n4392 ;
  assign y7871 = ~n28255 ;
  assign y7872 = ~n28258 ;
  assign y7873 = n28259 ;
  assign y7874 = n28262 ;
  assign y7875 = n28264 ;
  assign y7876 = ~1'b0 ;
  assign y7877 = ~n28266 ;
  assign y7878 = n28270 ;
  assign y7879 = ~n28274 ;
  assign y7880 = ~n28276 ;
  assign y7881 = ~n28281 ;
  assign y7882 = n28282 ;
  assign y7883 = n28283 ;
  assign y7884 = n28289 ;
  assign y7885 = n28292 ;
  assign y7886 = n28294 ;
  assign y7887 = ~n28298 ;
  assign y7888 = n28301 ;
  assign y7889 = ~n28303 ;
  assign y7890 = n28307 ;
  assign y7891 = ~n28311 ;
  assign y7892 = n28313 ;
  assign y7893 = n28315 ;
  assign y7894 = n28320 ;
  assign y7895 = ~n28322 ;
  assign y7896 = ~n28327 ;
  assign y7897 = n28328 ;
  assign y7898 = n28329 ;
  assign y7899 = n28333 ;
  assign y7900 = ~n28334 ;
  assign y7901 = n28339 ;
  assign y7902 = n28344 ;
  assign y7903 = n28345 ;
  assign y7904 = ~n28351 ;
  assign y7905 = ~n28352 ;
  assign y7906 = n28355 ;
  assign y7907 = n28356 ;
  assign y7908 = ~n28359 ;
  assign y7909 = ~n28362 ;
  assign y7910 = ~n28369 ;
  assign y7911 = n28370 ;
  assign y7912 = ~1'b0 ;
  assign y7913 = ~1'b0 ;
  assign y7914 = n28371 ;
  assign y7915 = n28372 ;
  assign y7916 = ~n28373 ;
  assign y7917 = ~n28374 ;
  assign y7918 = ~n28376 ;
  assign y7919 = ~n28378 ;
  assign y7920 = n28380 ;
  assign y7921 = n28381 ;
  assign y7922 = ~n28385 ;
  assign y7923 = ~n28388 ;
  assign y7924 = ~n28390 ;
  assign y7925 = n28391 ;
  assign y7926 = ~n28395 ;
  assign y7927 = ~n28399 ;
  assign y7928 = ~n28400 ;
  assign y7929 = n28401 ;
  assign y7930 = ~n28406 ;
  assign y7931 = ~n28409 ;
  assign y7932 = ~n28411 ;
  assign y7933 = n28417 ;
  assign y7934 = ~n28418 ;
  assign y7935 = n28420 ;
  assign y7936 = n28424 ;
  assign y7937 = n28430 ;
  assign y7938 = ~n28433 ;
  assign y7939 = ~n28436 ;
  assign y7940 = n28437 ;
  assign y7941 = n28440 ;
  assign y7942 = n28443 ;
  assign y7943 = n28447 ;
  assign y7944 = ~n28449 ;
  assign y7945 = n28450 ;
  assign y7946 = ~n28456 ;
  assign y7947 = ~n28458 ;
  assign y7948 = n28459 ;
  assign y7949 = ~n28462 ;
  assign y7950 = ~n28463 ;
  assign y7951 = n28465 ;
  assign y7952 = n28469 ;
  assign y7953 = ~n28472 ;
  assign y7954 = n28474 ;
  assign y7955 = ~n28475 ;
  assign y7956 = ~n28476 ;
  assign y7957 = ~n28478 ;
  assign y7958 = n28479 ;
  assign y7959 = n28480 ;
  assign y7960 = n28482 ;
  assign y7961 = ~1'b0 ;
  assign y7962 = n28483 ;
  assign y7963 = ~n28484 ;
  assign y7964 = ~n28486 ;
  assign y7965 = ~n28487 ;
  assign y7966 = n28488 ;
  assign y7967 = ~n28491 ;
  assign y7968 = ~n28498 ;
  assign y7969 = ~n28506 ;
  assign y7970 = ~1'b0 ;
  assign y7971 = ~n28510 ;
  assign y7972 = ~n28512 ;
  assign y7973 = n28514 ;
  assign y7974 = ~n28521 ;
  assign y7975 = ~n28522 ;
  assign y7976 = n28525 ;
  assign y7977 = ~1'b0 ;
  assign y7978 = ~1'b0 ;
  assign y7979 = n28527 ;
  assign y7980 = n28530 ;
  assign y7981 = n28532 ;
  assign y7982 = n28537 ;
  assign y7983 = n28538 ;
  assign y7984 = n28539 ;
  assign y7985 = ~n28542 ;
  assign y7986 = n28544 ;
  assign y7987 = n28546 ;
  assign y7988 = ~1'b0 ;
  assign y7989 = n28554 ;
  assign y7990 = n28555 ;
  assign y7991 = ~n28558 ;
  assign y7992 = ~n28560 ;
  assign y7993 = n28561 ;
  assign y7994 = ~n28563 ;
  assign y7995 = ~n28569 ;
  assign y7996 = ~n28570 ;
  assign y7997 = n28575 ;
  assign y7998 = ~1'b0 ;
  assign y7999 = ~1'b0 ;
  assign y8000 = n28581 ;
  assign y8001 = n28582 ;
  assign y8002 = n28583 ;
  assign y8003 = n28585 ;
  assign y8004 = ~n28586 ;
  assign y8005 = ~n28589 ;
  assign y8006 = ~n28597 ;
  assign y8007 = ~1'b0 ;
  assign y8008 = ~1'b0 ;
  assign y8009 = ~n28598 ;
  assign y8010 = n28599 ;
  assign y8011 = ~n28600 ;
  assign y8012 = n28601 ;
  assign y8013 = n28602 ;
  assign y8014 = n28605 ;
  assign y8015 = n28607 ;
  assign y8016 = n28609 ;
  assign y8017 = ~n28619 ;
  assign y8018 = n28620 ;
  assign y8019 = n28624 ;
  assign y8020 = ~n28626 ;
  assign y8021 = ~n28628 ;
  assign y8022 = ~n28631 ;
  assign y8023 = n28632 ;
  assign y8024 = ~n28633 ;
  assign y8025 = n28637 ;
  assign y8026 = ~n28641 ;
  assign y8027 = ~n28642 ;
  assign y8028 = ~n28650 ;
  assign y8029 = n28653 ;
  assign y8030 = ~n28655 ;
  assign y8031 = ~1'b0 ;
  assign y8032 = n28656 ;
  assign y8033 = n28659 ;
  assign y8034 = ~n28660 ;
  assign y8035 = ~n28661 ;
  assign y8036 = ~n28663 ;
  assign y8037 = n28667 ;
  assign y8038 = n28668 ;
  assign y8039 = ~1'b0 ;
  assign y8040 = n28672 ;
  assign y8041 = n28674 ;
  assign y8042 = ~n28676 ;
  assign y8043 = n28677 ;
  assign y8044 = n28678 ;
  assign y8045 = ~n28680 ;
  assign y8046 = ~n28688 ;
  assign y8047 = ~n28690 ;
  assign y8048 = ~n28694 ;
  assign y8049 = n28695 ;
  assign y8050 = ~n28698 ;
  assign y8051 = n28704 ;
  assign y8052 = ~n28708 ;
  assign y8053 = n28709 ;
  assign y8054 = n28711 ;
  assign y8055 = n28724 ;
  assign y8056 = ~1'b0 ;
  assign y8057 = ~n28726 ;
  assign y8058 = n28728 ;
  assign y8059 = ~n28731 ;
  assign y8060 = n28732 ;
  assign y8061 = n28734 ;
  assign y8062 = n28735 ;
  assign y8063 = n28736 ;
  assign y8064 = ~n28741 ;
  assign y8065 = ~n28744 ;
  assign y8066 = n28746 ;
  assign y8067 = n28748 ;
  assign y8068 = ~n28749 ;
  assign y8069 = n28750 ;
  assign y8070 = ~n28753 ;
  assign y8071 = ~n28754 ;
  assign y8072 = ~n28757 ;
  assign y8073 = ~n28759 ;
  assign y8074 = n28765 ;
  assign y8075 = ~n28767 ;
  assign y8076 = ~n28768 ;
  assign y8077 = n28769 ;
  assign y8078 = n28772 ;
  assign y8079 = n28777 ;
  assign y8080 = ~n28778 ;
  assign y8081 = ~n28779 ;
  assign y8082 = ~n28781 ;
  assign y8083 = n28787 ;
  assign y8084 = ~n11599 ;
  assign y8085 = n28793 ;
  assign y8086 = n28794 ;
  assign y8087 = ~n28799 ;
  assign y8088 = ~n28801 ;
  assign y8089 = n28802 ;
  assign y8090 = ~n28803 ;
  assign y8091 = n28804 ;
  assign y8092 = ~n28807 ;
  assign y8093 = ~n28810 ;
  assign y8094 = ~n28812 ;
  assign y8095 = n28813 ;
  assign y8096 = ~n28816 ;
  assign y8097 = ~n28817 ;
  assign y8098 = n28818 ;
  assign y8099 = n28819 ;
  assign y8100 = n28821 ;
  assign y8101 = ~n28823 ;
  assign y8102 = ~1'b0 ;
  assign y8103 = ~n28825 ;
  assign y8104 = ~n28828 ;
  assign y8105 = n28829 ;
  assign y8106 = n28830 ;
  assign y8107 = ~n28833 ;
  assign y8108 = ~n28836 ;
  assign y8109 = ~n28837 ;
  assign y8110 = ~1'b0 ;
  assign y8111 = ~1'b0 ;
  assign y8112 = n28840 ;
  assign y8113 = n28845 ;
  assign y8114 = ~n28849 ;
  assign y8115 = n28850 ;
  assign y8116 = ~n28852 ;
  assign y8117 = ~n28859 ;
  assign y8118 = n28861 ;
  assign y8119 = n28863 ;
  assign y8120 = n28866 ;
  assign y8121 = n28868 ;
  assign y8122 = ~n28870 ;
  assign y8123 = n28876 ;
  assign y8124 = ~n28880 ;
  assign y8125 = n28882 ;
  assign y8126 = n28884 ;
  assign y8127 = ~n28886 ;
  assign y8128 = n28887 ;
  assign y8129 = ~n28888 ;
  assign y8130 = ~n28891 ;
  assign y8131 = ~n28894 ;
  assign y8132 = ~1'b0 ;
  assign y8133 = n28896 ;
  assign y8134 = n28898 ;
  assign y8135 = ~n28902 ;
  assign y8136 = ~n28904 ;
  assign y8137 = n28906 ;
  assign y8138 = n28910 ;
  assign y8139 = ~n28911 ;
  assign y8140 = n28912 ;
  assign y8141 = n28916 ;
  assign y8142 = ~n28917 ;
  assign y8143 = ~n28919 ;
  assign y8144 = ~n28921 ;
  assign y8145 = ~n28926 ;
  assign y8146 = n28930 ;
  assign y8147 = ~n28931 ;
  assign y8148 = ~n28936 ;
  assign y8149 = ~n28940 ;
  assign y8150 = n28941 ;
  assign y8151 = ~1'b0 ;
  assign y8152 = ~n28943 ;
  assign y8153 = n28944 ;
  assign y8154 = ~n28948 ;
  assign y8155 = ~n28949 ;
  assign y8156 = ~n28951 ;
  assign y8157 = ~n28952 ;
  assign y8158 = ~n28954 ;
  assign y8159 = ~n28958 ;
  assign y8160 = ~n28962 ;
  assign y8161 = n28964 ;
  assign y8162 = n28968 ;
  assign y8163 = ~n28969 ;
  assign y8164 = ~n28972 ;
  assign y8165 = n28978 ;
  assign y8166 = ~n28982 ;
  assign y8167 = n28986 ;
  assign y8168 = ~n28990 ;
  assign y8169 = ~1'b0 ;
  assign y8170 = ~n28993 ;
  assign y8171 = ~1'b0 ;
  assign y8172 = ~n28996 ;
  assign y8173 = n28998 ;
  assign y8174 = n29001 ;
  assign y8175 = n29004 ;
  assign y8176 = n29006 ;
  assign y8177 = ~n29012 ;
  assign y8178 = n29013 ;
  assign y8179 = n29018 ;
  assign y8180 = ~1'b0 ;
  assign y8181 = n29022 ;
  assign y8182 = n29024 ;
  assign y8183 = ~n29028 ;
  assign y8184 = n29030 ;
  assign y8185 = ~n29036 ;
  assign y8186 = ~n29037 ;
  assign y8187 = ~n29042 ;
  assign y8188 = n29043 ;
  assign y8189 = n29047 ;
  assign y8190 = ~1'b0 ;
  assign y8191 = ~1'b0 ;
  assign y8192 = n29049 ;
  assign y8193 = n29050 ;
  assign y8194 = n29052 ;
  assign y8195 = ~n29053 ;
  assign y8196 = ~n29059 ;
  assign y8197 = n29065 ;
  assign y8198 = n29070 ;
  assign y8199 = n29072 ;
  assign y8200 = ~n29081 ;
  assign y8201 = ~n29087 ;
  assign y8202 = ~1'b0 ;
  assign y8203 = ~n29088 ;
  assign y8204 = ~n29089 ;
  assign y8205 = ~n29092 ;
  assign y8206 = ~n29095 ;
  assign y8207 = ~n29096 ;
  assign y8208 = ~n29097 ;
  assign y8209 = ~n29101 ;
  assign y8210 = n29103 ;
  assign y8211 = ~n29109 ;
  assign y8212 = n29110 ;
  assign y8213 = n29112 ;
  assign y8214 = ~n29114 ;
  assign y8215 = ~n29116 ;
  assign y8216 = ~n29127 ;
  assign y8217 = n29128 ;
  assign y8218 = ~n29130 ;
  assign y8219 = ~n29131 ;
  assign y8220 = ~1'b0 ;
  assign y8221 = ~n29133 ;
  assign y8222 = n29137 ;
  assign y8223 = n29140 ;
  assign y8224 = ~n29147 ;
  assign y8225 = n29149 ;
  assign y8226 = n29151 ;
  assign y8227 = n29154 ;
  assign y8228 = n29155 ;
  assign y8229 = n29160 ;
  assign y8230 = ~n29161 ;
  assign y8231 = ~n29162 ;
  assign y8232 = n29163 ;
  assign y8233 = n29164 ;
  assign y8234 = n29165 ;
  assign y8235 = n29167 ;
  assign y8236 = ~n29168 ;
  assign y8237 = n29171 ;
  assign y8238 = ~n29172 ;
  assign y8239 = ~1'b0 ;
  assign y8240 = ~n29174 ;
  assign y8241 = n29175 ;
  assign y8242 = n29176 ;
  assign y8243 = ~n29177 ;
  assign y8244 = ~n29178 ;
  assign y8245 = ~n29179 ;
  assign y8246 = ~n29181 ;
  assign y8247 = n29188 ;
  assign y8248 = n29189 ;
  assign y8249 = n29191 ;
  assign y8250 = ~n29193 ;
  assign y8251 = n29195 ;
  assign y8252 = ~n29201 ;
  assign y8253 = n29202 ;
  assign y8254 = n29206 ;
  assign y8255 = n29207 ;
  assign y8256 = n29210 ;
  assign y8257 = ~n29211 ;
  assign y8258 = n29212 ;
  assign y8259 = n29217 ;
  assign y8260 = n29224 ;
  assign y8261 = ~n29230 ;
  assign y8262 = ~n29235 ;
  assign y8263 = ~n29237 ;
  assign y8264 = n29240 ;
  assign y8265 = n29243 ;
  assign y8266 = n29245 ;
  assign y8267 = ~n29247 ;
  assign y8268 = ~1'b0 ;
  assign y8269 = ~n29250 ;
  assign y8270 = ~n29253 ;
  assign y8271 = n29255 ;
  assign y8272 = ~n29256 ;
  assign y8273 = ~n29259 ;
  assign y8274 = ~n29260 ;
  assign y8275 = n29261 ;
  assign y8276 = ~1'b0 ;
  assign y8277 = n29264 ;
  assign y8278 = ~n29268 ;
  assign y8279 = ~n29269 ;
  assign y8280 = ~n29273 ;
  assign y8281 = ~n29277 ;
  assign y8282 = ~n29280 ;
  assign y8283 = n29281 ;
  assign y8284 = ~n12435 ;
  assign y8285 = ~n29283 ;
  assign y8286 = n29284 ;
  assign y8287 = n29290 ;
  assign y8288 = ~1'b0 ;
  assign y8289 = ~1'b0 ;
  assign y8290 = n29291 ;
  assign y8291 = n29294 ;
  assign y8292 = n29297 ;
  assign y8293 = ~n29300 ;
  assign y8294 = n29305 ;
  assign y8295 = n29306 ;
  assign y8296 = ~n29307 ;
  assign y8297 = ~n29311 ;
  assign y8298 = n29314 ;
  assign y8299 = ~1'b0 ;
  assign y8300 = n29315 ;
  assign y8301 = n29317 ;
  assign y8302 = ~n29318 ;
  assign y8303 = ~n12382 ;
  assign y8304 = ~n29319 ;
  assign y8305 = n29323 ;
  assign y8306 = ~n29324 ;
  assign y8307 = ~n29326 ;
  assign y8308 = n29330 ;
  assign y8309 = n29332 ;
  assign y8310 = n29335 ;
  assign y8311 = n29337 ;
  assign y8312 = n29338 ;
  assign y8313 = ~n29339 ;
  assign y8314 = n29341 ;
  assign y8315 = ~n29342 ;
  assign y8316 = ~n29344 ;
  assign y8317 = ~n29346 ;
  assign y8318 = ~n29348 ;
  assign y8319 = ~n29349 ;
  assign y8320 = n29358 ;
  assign y8321 = n29360 ;
  assign y8322 = ~n29364 ;
  assign y8323 = ~n29372 ;
  assign y8324 = n29373 ;
  assign y8325 = ~n29374 ;
  assign y8326 = ~n29376 ;
  assign y8327 = ~n8216 ;
  assign y8328 = ~1'b0 ;
  assign y8329 = ~n29377 ;
  assign y8330 = ~n29381 ;
  assign y8331 = ~n29383 ;
  assign y8332 = ~n29385 ;
  assign y8333 = n29386 ;
  assign y8334 = n29388 ;
  assign y8335 = n29390 ;
  assign y8336 = n29393 ;
  assign y8337 = ~n29395 ;
  assign y8338 = n29397 ;
  assign y8339 = ~n29399 ;
  assign y8340 = n29400 ;
  assign y8341 = n29402 ;
  assign y8342 = n29404 ;
  assign y8343 = n29405 ;
  assign y8344 = ~n29406 ;
  assign y8345 = n29409 ;
  assign y8346 = ~1'b0 ;
  assign y8347 = ~n29411 ;
  assign y8348 = ~n29412 ;
  assign y8349 = ~n25739 ;
  assign y8350 = n2907 ;
  assign y8351 = ~n29417 ;
  assign y8352 = ~n29418 ;
  assign y8353 = ~n29422 ;
  assign y8354 = n27453 ;
  assign y8355 = ~n29424 ;
  assign y8356 = ~n29426 ;
  assign y8357 = ~n29428 ;
  assign y8358 = n29429 ;
  assign y8359 = n29434 ;
  assign y8360 = ~n29439 ;
  assign y8361 = ~n29441 ;
  assign y8362 = n29442 ;
  assign y8363 = n29444 ;
  assign y8364 = n29445 ;
  assign y8365 = n29446 ;
  assign y8366 = n29448 ;
  assign y8367 = n29451 ;
  assign y8368 = ~1'b0 ;
  assign y8369 = ~n29457 ;
  assign y8370 = n29460 ;
  assign y8371 = n29461 ;
  assign y8372 = ~n29462 ;
  assign y8373 = ~n29465 ;
  assign y8374 = ~n29468 ;
  assign y8375 = n29474 ;
  assign y8376 = ~1'b0 ;
  assign y8377 = n29479 ;
  assign y8378 = n29481 ;
  assign y8379 = ~n29483 ;
  assign y8380 = ~n29484 ;
  assign y8381 = ~n29486 ;
  assign y8382 = n29487 ;
  assign y8383 = n29491 ;
  assign y8384 = ~n29493 ;
  assign y8385 = n29496 ;
  assign y8386 = n29498 ;
  assign y8387 = n29505 ;
  assign y8388 = n29508 ;
  assign y8389 = n29514 ;
  assign y8390 = ~n29520 ;
  assign y8391 = n29523 ;
  assign y8392 = ~n29525 ;
  assign y8393 = ~n29531 ;
  assign y8394 = n29534 ;
  assign y8395 = n29535 ;
  assign y8396 = ~n29540 ;
  assign y8397 = n29541 ;
  assign y8398 = n29543 ;
  assign y8399 = ~n29547 ;
  assign y8400 = n29550 ;
  assign y8401 = n29552 ;
  assign y8402 = n29556 ;
  assign y8403 = ~n29558 ;
  assign y8404 = ~n29560 ;
  assign y8405 = ~1'b0 ;
  assign y8406 = n29562 ;
  assign y8407 = n29563 ;
  assign y8408 = n29566 ;
  assign y8409 = n29569 ;
  assign y8410 = ~n29571 ;
  assign y8411 = ~n29573 ;
  assign y8412 = ~n29574 ;
  assign y8413 = ~n29578 ;
  assign y8414 = ~n29579 ;
  assign y8415 = ~n29581 ;
  assign y8416 = ~1'b0 ;
  assign y8417 = ~1'b0 ;
  assign y8418 = ~n29582 ;
  assign y8419 = n29584 ;
  assign y8420 = n29586 ;
  assign y8421 = n29588 ;
  assign y8422 = n29589 ;
  assign y8423 = ~n29590 ;
  assign y8424 = ~n29593 ;
  assign y8425 = ~1'b0 ;
  assign y8426 = n29595 ;
  assign y8427 = n29600 ;
  assign y8428 = n29602 ;
  assign y8429 = n29603 ;
  assign y8430 = ~n29606 ;
  assign y8431 = n29608 ;
  assign y8432 = n29609 ;
  assign y8433 = n29610 ;
  assign y8434 = n29611 ;
  assign y8435 = ~1'b0 ;
  assign y8436 = ~1'b0 ;
  assign y8437 = ~1'b0 ;
  assign y8438 = n29612 ;
  assign y8439 = ~n29614 ;
  assign y8440 = ~n29617 ;
  assign y8441 = ~n29618 ;
  assign y8442 = n29619 ;
  assign y8443 = ~n29623 ;
  assign y8444 = ~1'b0 ;
  assign y8445 = ~n29626 ;
  assign y8446 = ~n29627 ;
  assign y8447 = n29631 ;
  assign y8448 = ~n29632 ;
  assign y8449 = n29634 ;
  assign y8450 = n29635 ;
  assign y8451 = ~n29638 ;
  assign y8452 = n29642 ;
  assign y8453 = ~n29176 ;
  assign y8454 = n29643 ;
  assign y8455 = ~n29645 ;
  assign y8456 = ~n29651 ;
  assign y8457 = n29656 ;
  assign y8458 = ~n29659 ;
  assign y8459 = ~n29660 ;
  assign y8460 = n29670 ;
  assign y8461 = ~n29675 ;
  assign y8462 = n29683 ;
  assign y8463 = n29685 ;
  assign y8464 = n29688 ;
  assign y8465 = ~n29691 ;
  assign y8466 = ~n29692 ;
  assign y8467 = ~n29693 ;
  assign y8468 = ~n29695 ;
  assign y8469 = ~n29696 ;
  assign y8470 = ~n29700 ;
  assign y8471 = n29704 ;
  assign y8472 = ~n29707 ;
  assign y8473 = n29712 ;
  assign y8474 = n29713 ;
  assign y8475 = n29715 ;
  assign y8476 = n29716 ;
  assign y8477 = n29717 ;
  assign y8478 = n29720 ;
  assign y8479 = ~n29721 ;
  assign y8480 = n29723 ;
  assign y8481 = ~n29729 ;
  assign y8482 = n29732 ;
  assign y8483 = ~n29735 ;
  assign y8484 = ~n29740 ;
  assign y8485 = n29741 ;
  assign y8486 = ~1'b0 ;
  assign y8487 = ~n29744 ;
  assign y8488 = ~n29745 ;
  assign y8489 = ~n29747 ;
  assign y8490 = n29749 ;
  assign y8491 = n29752 ;
  assign y8492 = n29754 ;
  assign y8493 = ~n29756 ;
  assign y8494 = ~n29758 ;
  assign y8495 = ~n29761 ;
  assign y8496 = n29765 ;
  assign y8497 = n29766 ;
  assign y8498 = ~1'b0 ;
  assign y8499 = n29767 ;
  assign y8500 = ~n29768 ;
  assign y8501 = ~n29774 ;
  assign y8502 = n29775 ;
  assign y8503 = ~n29778 ;
  assign y8504 = ~1'b0 ;
  assign y8505 = n29779 ;
  assign y8506 = n29780 ;
  assign y8507 = n29782 ;
  assign y8508 = ~n29787 ;
  assign y8509 = ~n29788 ;
  assign y8510 = n29789 ;
  assign y8511 = n29793 ;
  assign y8512 = ~n29797 ;
  assign y8513 = ~n29803 ;
  assign y8514 = ~1'b0 ;
  assign y8515 = ~1'b0 ;
  assign y8516 = ~n29809 ;
  assign y8517 = ~n29813 ;
  assign y8518 = n29824 ;
  assign y8519 = ~n29825 ;
  assign y8520 = ~n29826 ;
  assign y8521 = ~n29827 ;
  assign y8522 = n29829 ;
  assign y8523 = ~n29831 ;
  assign y8524 = n29837 ;
  assign y8525 = n29840 ;
  assign y8526 = ~n29843 ;
  assign y8527 = n29844 ;
  assign y8528 = n29845 ;
  assign y8529 = ~n29850 ;
  assign y8530 = n29851 ;
  assign y8531 = ~n29852 ;
  assign y8532 = n29855 ;
  assign y8533 = ~n29857 ;
  assign y8534 = ~1'b0 ;
  assign y8535 = ~n29859 ;
  assign y8536 = n29864 ;
  assign y8537 = n29868 ;
  assign y8538 = n29874 ;
  assign y8539 = ~n29878 ;
  assign y8540 = n29881 ;
  assign y8541 = n29882 ;
  assign y8542 = n29883 ;
  assign y8543 = ~n29888 ;
  assign y8544 = n29891 ;
  assign y8545 = n29894 ;
  assign y8546 = ~1'b0 ;
  assign y8547 = ~n29895 ;
  assign y8548 = n29897 ;
  assign y8549 = ~n29899 ;
  assign y8550 = ~n29901 ;
  assign y8551 = n29904 ;
  assign y8552 = ~n29905 ;
  assign y8553 = ~n29906 ;
  assign y8554 = ~n29907 ;
  assign y8555 = ~1'b0 ;
  assign y8556 = ~1'b0 ;
  assign y8557 = n29908 ;
  assign y8558 = ~n29909 ;
  assign y8559 = n29910 ;
  assign y8560 = ~n29911 ;
  assign y8561 = n29915 ;
  assign y8562 = n29919 ;
  assign y8563 = n29922 ;
  assign y8564 = ~n29924 ;
  assign y8565 = n29926 ;
  assign y8566 = ~n29929 ;
  assign y8567 = n29932 ;
  assign y8568 = n29933 ;
  assign y8569 = ~n29934 ;
  assign y8570 = ~n29938 ;
  assign y8571 = ~n29941 ;
  assign y8572 = n29944 ;
  assign y8573 = ~n29945 ;
  assign y8574 = ~n29947 ;
  assign y8575 = n29949 ;
  assign y8576 = ~n29953 ;
  assign y8577 = ~n29957 ;
  assign y8578 = n29972 ;
  assign y8579 = ~n29973 ;
  assign y8580 = n29975 ;
  assign y8581 = ~n29977 ;
  assign y8582 = ~n29981 ;
  assign y8583 = ~1'b0 ;
  assign y8584 = ~n29983 ;
  assign y8585 = n29985 ;
  assign y8586 = ~n29986 ;
  assign y8587 = n29988 ;
  assign y8588 = n29990 ;
  assign y8589 = ~n29996 ;
  assign y8590 = ~n29997 ;
  assign y8591 = n30000 ;
  assign y8592 = ~n30003 ;
  assign y8593 = ~n30006 ;
  assign y8594 = ~1'b0 ;
  assign y8595 = ~1'b0 ;
  assign y8596 = ~n30011 ;
  assign y8597 = ~n30012 ;
  assign y8598 = ~n30013 ;
  assign y8599 = n30017 ;
  assign y8600 = ~n30024 ;
  assign y8601 = n30028 ;
  assign y8602 = n30030 ;
  assign y8603 = ~n30037 ;
  assign y8604 = ~n30039 ;
  assign y8605 = ~n30041 ;
  assign y8606 = n30042 ;
  assign y8607 = ~n30044 ;
  assign y8608 = n30045 ;
  assign y8609 = n30046 ;
  assign y8610 = n30048 ;
  assign y8611 = ~n30050 ;
  assign y8612 = n30051 ;
  assign y8613 = n30052 ;
  assign y8614 = ~1'b0 ;
  assign y8615 = ~n30056 ;
  assign y8616 = ~n30058 ;
  assign y8617 = ~n30059 ;
  assign y8618 = ~n30062 ;
  assign y8619 = n30065 ;
  assign y8620 = n30067 ;
  assign y8621 = ~n30071 ;
  assign y8622 = ~n30075 ;
  assign y8623 = ~1'b0 ;
  assign y8624 = ~1'b0 ;
  assign y8625 = n30080 ;
  assign y8626 = n30084 ;
  assign y8627 = ~n30085 ;
  assign y8628 = ~n30086 ;
  assign y8629 = n30088 ;
  assign y8630 = ~n30092 ;
  assign y8631 = ~n30094 ;
  assign y8632 = ~n30099 ;
  assign y8633 = n30100 ;
  assign y8634 = n30103 ;
  assign y8635 = ~n30104 ;
  assign y8636 = n30106 ;
  assign y8637 = ~n30112 ;
  assign y8638 = n30114 ;
  assign y8639 = ~n30116 ;
  assign y8640 = n30117 ;
  assign y8641 = n30120 ;
  assign y8642 = ~n30121 ;
  assign y8643 = n30122 ;
  assign y8644 = n30127 ;
  assign y8645 = ~n30128 ;
  assign y8646 = ~n30129 ;
  assign y8647 = ~n30130 ;
  assign y8648 = n30133 ;
  assign y8649 = n30145 ;
  assign y8650 = ~n30153 ;
  assign y8651 = n30157 ;
  assign y8652 = n30162 ;
  assign y8653 = n30164 ;
  assign y8654 = ~1'b0 ;
  assign y8655 = ~1'b0 ;
  assign y8656 = ~n30165 ;
  assign y8657 = n30167 ;
  assign y8658 = n30168 ;
  assign y8659 = ~n30169 ;
  assign y8660 = n30171 ;
  assign y8661 = ~n30172 ;
  assign y8662 = n30179 ;
  assign y8663 = ~n30189 ;
  assign y8664 = ~n30192 ;
  assign y8665 = ~n30197 ;
  assign y8666 = ~n30202 ;
  assign y8667 = ~n30204 ;
  assign y8668 = ~n30205 ;
  assign y8669 = ~n30206 ;
  assign y8670 = ~n30209 ;
  assign y8671 = ~n30217 ;
  assign y8672 = n30219 ;
  assign y8673 = ~n30222 ;
  assign y8674 = ~1'b0 ;
  assign y8675 = n30224 ;
  assign y8676 = ~n30227 ;
  assign y8677 = ~n30229 ;
  assign y8678 = n30230 ;
  assign y8679 = n30231 ;
  assign y8680 = n30232 ;
  assign y8681 = n30234 ;
  assign y8682 = ~n30235 ;
  assign y8683 = ~n30236 ;
  assign y8684 = n30237 ;
  assign y8685 = ~1'b0 ;
  assign y8686 = ~1'b0 ;
  assign y8687 = ~n30239 ;
  assign y8688 = n30240 ;
  assign y8689 = ~n30243 ;
  assign y8690 = n30249 ;
  assign y8691 = n30250 ;
  assign y8692 = ~n30251 ;
  assign y8693 = ~n30252 ;
  assign y8694 = ~n30253 ;
  assign y8695 = ~n30255 ;
  assign y8696 = ~1'b0 ;
  assign y8697 = ~1'b0 ;
  assign y8698 = n30257 ;
  assign y8699 = n30258 ;
  assign y8700 = n30260 ;
  assign y8701 = ~n30263 ;
  assign y8702 = n30264 ;
  assign y8703 = ~n30265 ;
  assign y8704 = ~n30266 ;
  assign y8705 = ~n30271 ;
  assign y8706 = n14762 ;
  assign y8707 = n30274 ;
  assign y8708 = n30276 ;
  assign y8709 = n30278 ;
  assign y8710 = ~n30288 ;
  assign y8711 = n30294 ;
  assign y8712 = n30297 ;
  assign y8713 = ~n30298 ;
  assign y8714 = ~n30299 ;
  assign y8715 = n30301 ;
  assign y8716 = ~n30303 ;
  assign y8717 = ~n17300 ;
  assign y8718 = n30305 ;
  assign y8719 = n30307 ;
  assign y8720 = ~n30311 ;
  assign y8721 = n30312 ;
  assign y8722 = n30317 ;
  assign y8723 = n30318 ;
  assign y8724 = ~n30321 ;
  assign y8725 = n30322 ;
  assign y8726 = n30323 ;
  assign y8727 = ~n30328 ;
  assign y8728 = n30329 ;
  assign y8729 = n30331 ;
  assign y8730 = n30335 ;
  assign y8731 = n30338 ;
  assign y8732 = n30339 ;
  assign y8733 = n30343 ;
  assign y8734 = n30348 ;
  assign y8735 = ~n30349 ;
  assign y8736 = n30351 ;
  assign y8737 = ~n30352 ;
  assign y8738 = n30356 ;
  assign y8739 = n30360 ;
  assign y8740 = ~n30362 ;
  assign y8741 = ~n30366 ;
  assign y8742 = ~n30368 ;
  assign y8743 = n30369 ;
  assign y8744 = ~n30374 ;
  assign y8745 = ~n30375 ;
  assign y8746 = n30376 ;
  assign y8747 = n30379 ;
  assign y8748 = ~n30382 ;
  assign y8749 = n30386 ;
  assign y8750 = n30388 ;
  assign y8751 = ~n30393 ;
  assign y8752 = ~n30400 ;
  assign y8753 = ~n30401 ;
  assign y8754 = ~n30404 ;
  assign y8755 = n30406 ;
  assign y8756 = n30409 ;
  assign y8757 = ~n30411 ;
  assign y8758 = ~1'b0 ;
  assign y8759 = ~1'b0 ;
  assign y8760 = n30413 ;
  assign y8761 = ~n30414 ;
  assign y8762 = n30415 ;
  assign y8763 = ~n30417 ;
  assign y8764 = n30418 ;
  assign y8765 = ~n30419 ;
  assign y8766 = ~n30420 ;
  assign y8767 = ~n30425 ;
  assign y8768 = ~n30427 ;
  assign y8769 = ~n30435 ;
  assign y8770 = n30438 ;
  assign y8771 = ~n30443 ;
  assign y8772 = ~n30446 ;
  assign y8773 = n30447 ;
  assign y8774 = ~n30452 ;
  assign y8775 = ~n30453 ;
  assign y8776 = ~1'b0 ;
  assign y8777 = ~n30460 ;
  assign y8778 = ~n30462 ;
  assign y8779 = n30463 ;
  assign y8780 = n30466 ;
  assign y8781 = ~n30468 ;
  assign y8782 = n30474 ;
  assign y8783 = n30477 ;
  assign y8784 = n30479 ;
  assign y8785 = n30480 ;
  assign y8786 = ~n30483 ;
  assign y8787 = ~1'b0 ;
  assign y8788 = ~1'b0 ;
  assign y8789 = ~1'b0 ;
  assign y8790 = n30485 ;
  assign y8791 = ~n30486 ;
  assign y8792 = n30488 ;
  assign y8793 = ~n30490 ;
  assign y8794 = ~n30492 ;
  assign y8795 = n30499 ;
  assign y8796 = ~n30503 ;
  assign y8797 = ~n30507 ;
  assign y8798 = n30509 ;
  assign y8799 = ~n30514 ;
  assign y8800 = n30522 ;
  assign y8801 = ~n30524 ;
  assign y8802 = ~n30527 ;
  assign y8803 = n30528 ;
  assign y8804 = ~n30529 ;
  assign y8805 = n30531 ;
  assign y8806 = ~n30533 ;
  assign y8807 = n30534 ;
  assign y8808 = ~n30537 ;
  assign y8809 = n30544 ;
  assign y8810 = ~n30549 ;
  assign y8811 = ~1'b0 ;
  assign y8812 = n30552 ;
  assign y8813 = n30555 ;
  assign y8814 = n30559 ;
  assign y8815 = ~n30564 ;
  assign y8816 = n30565 ;
  assign y8817 = n30566 ;
  assign y8818 = n30572 ;
  assign y8819 = ~n30574 ;
  assign y8820 = ~n30576 ;
  assign y8821 = ~1'b0 ;
  assign y8822 = n30578 ;
  assign y8823 = n30583 ;
  assign y8824 = ~n30586 ;
  assign y8825 = n30588 ;
  assign y8826 = ~n30589 ;
  assign y8827 = ~n30591 ;
  assign y8828 = n30592 ;
  assign y8829 = n30594 ;
  assign y8830 = ~1'b0 ;
  assign y8831 = ~n30595 ;
  assign y8832 = ~n30598 ;
  assign y8833 = ~n30600 ;
  assign y8834 = n30601 ;
  assign y8835 = ~n30602 ;
  assign y8836 = ~n30603 ;
  assign y8837 = ~n30606 ;
  assign y8838 = n30610 ;
  assign y8839 = ~n30613 ;
  assign y8840 = ~n30616 ;
  assign y8841 = ~n30618 ;
  assign y8842 = ~n30620 ;
  assign y8843 = ~n30622 ;
  assign y8844 = n30623 ;
  assign y8845 = n30624 ;
  assign y8846 = ~n30625 ;
  assign y8847 = n30626 ;
  assign y8848 = ~n30628 ;
  assign y8849 = ~n30629 ;
  assign y8850 = ~1'b0 ;
  assign y8851 = ~1'b0 ;
  assign y8852 = ~1'b0 ;
  assign y8853 = ~n30630 ;
  assign y8854 = n30633 ;
  assign y8855 = n30634 ;
  assign y8856 = n30635 ;
  assign y8857 = n30636 ;
  assign y8858 = n30641 ;
  assign y8859 = n30642 ;
  assign y8860 = ~n30644 ;
  assign y8861 = n30646 ;
  assign y8862 = n30649 ;
  assign y8863 = ~n30650 ;
  assign y8864 = ~n30652 ;
  assign y8865 = n30653 ;
  assign y8866 = n30654 ;
  assign y8867 = ~n30656 ;
  assign y8868 = ~n30658 ;
  assign y8869 = n30659 ;
  assign y8870 = ~n30660 ;
  assign y8871 = n30663 ;
  assign y8872 = n30665 ;
  assign y8873 = n30667 ;
  assign y8874 = ~n30669 ;
  assign y8875 = n30672 ;
  assign y8876 = ~n30675 ;
  assign y8877 = n30676 ;
  assign y8878 = ~n30677 ;
  assign y8879 = n4760 ;
  assign y8880 = n30679 ;
  assign y8881 = n30681 ;
  assign y8882 = n30684 ;
  assign y8883 = ~1'b0 ;
  assign y8884 = n30685 ;
  assign y8885 = n30688 ;
  assign y8886 = ~n30694 ;
  assign y8887 = ~n30696 ;
  assign y8888 = n30697 ;
  assign y8889 = n30698 ;
  assign y8890 = n30702 ;
  assign y8891 = ~n30704 ;
  assign y8892 = n30706 ;
  assign y8893 = ~n30709 ;
  assign y8894 = n30710 ;
  assign y8895 = n30712 ;
  assign y8896 = n30717 ;
  assign y8897 = n30719 ;
  assign y8898 = n30721 ;
  assign y8899 = ~n30723 ;
  assign y8900 = n30724 ;
  assign y8901 = ~n30732 ;
  assign y8902 = n30733 ;
  assign y8903 = n30736 ;
  assign y8904 = n30739 ;
  assign y8905 = ~n30741 ;
  assign y8906 = ~n30743 ;
  assign y8907 = n30744 ;
  assign y8908 = ~n30745 ;
  assign y8909 = n30747 ;
  assign y8910 = ~n30748 ;
  assign y8911 = ~n30749 ;
  assign y8912 = ~n30750 ;
  assign y8913 = ~n30751 ;
  assign y8914 = ~n30755 ;
  assign y8915 = n30758 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = n30763 ;
  assign y8918 = n30767 ;
  assign y8919 = ~n30770 ;
  assign y8920 = ~n30771 ;
  assign y8921 = n30773 ;
  assign y8922 = n30774 ;
  assign y8923 = n30778 ;
  assign y8924 = ~n30780 ;
  assign y8925 = ~n30781 ;
  assign y8926 = ~n30783 ;
  assign y8927 = ~n30785 ;
  assign y8928 = ~n30787 ;
  assign y8929 = ~n30789 ;
  assign y8930 = ~n30791 ;
  assign y8931 = ~n30792 ;
  assign y8932 = ~n30793 ;
  assign y8933 = n30794 ;
  assign y8934 = n30795 ;
  assign y8935 = n30796 ;
  assign y8936 = ~n30797 ;
  assign y8937 = ~1'b0 ;
  assign y8938 = n30800 ;
  assign y8939 = ~1'b0 ;
  assign y8940 = ~n30801 ;
  assign y8941 = n30803 ;
  assign y8942 = n30804 ;
  assign y8943 = ~n30805 ;
  assign y8944 = ~n30806 ;
  assign y8945 = ~n30810 ;
  assign y8946 = n30812 ;
  assign y8947 = ~n30813 ;
  assign y8948 = ~n30815 ;
  assign y8949 = ~n30817 ;
  assign y8950 = n30821 ;
  assign y8951 = n30822 ;
  assign y8952 = n30823 ;
  assign y8953 = n30825 ;
  assign y8954 = n30827 ;
  assign y8955 = n30829 ;
  assign y8956 = n30830 ;
  assign y8957 = ~n30833 ;
  assign y8958 = ~1'b0 ;
  assign y8959 = ~n30834 ;
  assign y8960 = ~n30838 ;
  assign y8961 = ~n30840 ;
  assign y8962 = ~n30841 ;
  assign y8963 = n30850 ;
  assign y8964 = n30853 ;
  assign y8965 = ~n30855 ;
  assign y8966 = n30858 ;
  assign y8967 = n30860 ;
  assign y8968 = n30861 ;
  assign y8969 = n30862 ;
  assign y8970 = ~n30863 ;
  assign y8971 = ~n30864 ;
  assign y8972 = ~n30868 ;
  assign y8973 = ~n30872 ;
  assign y8974 = ~n30876 ;
  assign y8975 = n30878 ;
  assign y8976 = ~n30880 ;
  assign y8977 = ~n30882 ;
  assign y8978 = n30886 ;
  assign y8979 = n30887 ;
  assign y8980 = n30892 ;
  assign y8981 = n30894 ;
  assign y8982 = ~n23855 ;
  assign y8983 = n30895 ;
  assign y8984 = n30898 ;
  assign y8985 = n30904 ;
  assign y8986 = ~n30906 ;
  assign y8987 = ~1'b0 ;
  assign y8988 = ~n30910 ;
  assign y8989 = n30912 ;
  assign y8990 = n30914 ;
  assign y8991 = n30920 ;
  assign y8992 = n30921 ;
  assign y8993 = n30924 ;
  assign y8994 = n30925 ;
  assign y8995 = n30926 ;
  assign y8996 = ~n30928 ;
  assign y8997 = n30930 ;
  assign y8998 = ~n30935 ;
  assign y8999 = ~n30936 ;
  assign y9000 = ~n30940 ;
  assign y9001 = n30942 ;
  assign y9002 = ~n30943 ;
  assign y9003 = ~n30944 ;
  assign y9004 = ~n30945 ;
  assign y9005 = ~n30946 ;
  assign y9006 = n30952 ;
  assign y9007 = ~n30960 ;
  assign y9008 = ~1'b0 ;
  assign y9009 = ~n30961 ;
  assign y9010 = ~n30963 ;
  assign y9011 = ~n30965 ;
  assign y9012 = ~n30967 ;
  assign y9013 = n30968 ;
  assign y9014 = ~n30969 ;
  assign y9015 = n30971 ;
  assign y9016 = ~n30977 ;
  assign y9017 = ~n30982 ;
  assign y9018 = ~1'b0 ;
  assign y9019 = ~n30983 ;
  assign y9020 = n30989 ;
  assign y9021 = n30992 ;
  assign y9022 = n30995 ;
  assign y9023 = n30997 ;
  assign y9024 = ~n30998 ;
  assign y9025 = ~n31000 ;
  assign y9026 = ~n31004 ;
  assign y9027 = ~n31007 ;
  assign y9028 = ~n31008 ;
  assign y9029 = ~n31010 ;
  assign y9030 = ~n31012 ;
  assign y9031 = ~n31017 ;
  assign y9032 = n31021 ;
  assign y9033 = n31023 ;
  assign y9034 = n31024 ;
  assign y9035 = ~n31026 ;
  assign y9036 = ~n31030 ;
  assign y9037 = ~n31035 ;
  assign y9038 = n31038 ;
  assign y9039 = ~n31039 ;
  assign y9040 = n31042 ;
  assign y9041 = n31045 ;
  assign y9042 = n31047 ;
  assign y9043 = n31050 ;
  assign y9044 = n31052 ;
  assign y9045 = ~n31054 ;
  assign y9046 = ~n31056 ;
  assign y9047 = n31059 ;
  assign y9048 = n31060 ;
  assign y9049 = ~n31064 ;
  assign y9050 = n31065 ;
  assign y9051 = n31066 ;
  assign y9052 = n31070 ;
  assign y9053 = ~n31076 ;
  assign y9054 = n31078 ;
  assign y9055 = ~n31080 ;
  assign y9056 = n31081 ;
  assign y9057 = n31085 ;
  assign y9058 = n31089 ;
  assign y9059 = n31092 ;
  assign y9060 = n31093 ;
  assign y9061 = ~n31095 ;
  assign y9062 = ~n31098 ;
  assign y9063 = ~n31100 ;
  assign y9064 = ~1'b0 ;
  assign y9065 = ~1'b0 ;
  assign y9066 = n31103 ;
  assign y9067 = ~n31107 ;
  assign y9068 = ~n31112 ;
  assign y9069 = ~n31116 ;
  assign y9070 = ~n31119 ;
  assign y9071 = ~n31120 ;
  assign y9072 = ~n31123 ;
  assign y9073 = ~1'b0 ;
  assign y9074 = ~n31124 ;
  assign y9075 = ~n31126 ;
  assign y9076 = n31129 ;
  assign y9077 = n31132 ;
  assign y9078 = ~n31133 ;
  assign y9079 = n31137 ;
  assign y9080 = n31144 ;
  assign y9081 = ~n31145 ;
  assign y9082 = ~n31148 ;
  assign y9083 = n31151 ;
  assign y9084 = ~n31153 ;
  assign y9085 = n31158 ;
  assign y9086 = ~n31159 ;
  assign y9087 = ~n31160 ;
  assign y9088 = n31161 ;
  assign y9089 = n31163 ;
  assign y9090 = ~n31165 ;
  assign y9091 = n31170 ;
  assign y9092 = ~n31171 ;
  assign y9093 = n31176 ;
  assign y9094 = ~n31182 ;
  assign y9095 = ~n31184 ;
  assign y9096 = ~n31186 ;
  assign y9097 = ~1'b0 ;
  assign y9098 = ~n31187 ;
  assign y9099 = n31188 ;
  assign y9100 = ~n31191 ;
  assign y9101 = ~n31192 ;
  assign y9102 = n31193 ;
  assign y9103 = ~n31198 ;
  assign y9104 = n31200 ;
  assign y9105 = n31201 ;
  assign y9106 = ~n31204 ;
  assign y9107 = ~1'b0 ;
  assign y9108 = n31206 ;
  assign y9109 = ~n31208 ;
  assign y9110 = ~n31211 ;
  assign y9111 = ~n31214 ;
  assign y9112 = ~n31216 ;
  assign y9113 = n31217 ;
  assign y9114 = n31222 ;
  assign y9115 = n31225 ;
  assign y9116 = n31227 ;
  assign y9117 = ~n31231 ;
  assign y9118 = ~1'b0 ;
  assign y9119 = ~n31233 ;
  assign y9120 = n31234 ;
  assign y9121 = n31237 ;
  assign y9122 = ~n31238 ;
  assign y9123 = n31240 ;
  assign y9124 = n31243 ;
  assign y9125 = ~n31248 ;
  assign y9126 = n31252 ;
  assign y9127 = n31255 ;
  assign y9128 = ~1'b0 ;
  assign y9129 = ~1'b0 ;
  assign y9130 = ~1'b0 ;
  assign y9131 = ~n31260 ;
  assign y9132 = n31263 ;
  assign y9133 = ~n31265 ;
  assign y9134 = n31266 ;
  assign y9135 = ~n31267 ;
  assign y9136 = n31270 ;
  assign y9137 = ~n31271 ;
  assign y9138 = ~n31273 ;
  assign y9139 = ~1'b0 ;
  assign y9140 = ~1'b0 ;
  assign y9141 = ~n31275 ;
  assign y9142 = n31277 ;
  assign y9143 = ~n31280 ;
  assign y9144 = ~n31283 ;
  assign y9145 = ~n31284 ;
  assign y9146 = n31285 ;
  assign y9147 = ~n31295 ;
  assign y9148 = ~n31297 ;
  assign y9149 = n31299 ;
  assign y9150 = ~n31300 ;
  assign y9151 = n31301 ;
  assign y9152 = ~n31306 ;
  assign y9153 = n31309 ;
  assign y9154 = ~n31310 ;
  assign y9155 = ~n31312 ;
  assign y9156 = n31313 ;
  assign y9157 = ~n31316 ;
  assign y9158 = ~n31317 ;
  assign y9159 = ~n31318 ;
  assign y9160 = ~n31319 ;
  assign y9161 = n31322 ;
  assign y9162 = ~1'b0 ;
  assign y9163 = n31324 ;
  assign y9164 = ~n31325 ;
  assign y9165 = ~n31326 ;
  assign y9166 = n31328 ;
  assign y9167 = ~n31329 ;
  assign y9168 = ~n31331 ;
  assign y9169 = ~n31332 ;
  assign y9170 = n31333 ;
  assign y9171 = ~1'b0 ;
  assign y9172 = n31335 ;
  assign y9173 = ~1'b0 ;
  assign y9174 = ~n31345 ;
  assign y9175 = n31346 ;
  assign y9176 = ~n31347 ;
  assign y9177 = ~n31350 ;
  assign y9178 = ~n31351 ;
  assign y9179 = n31353 ;
  assign y9180 = ~n31354 ;
  assign y9181 = n31355 ;
  assign y9182 = ~1'b0 ;
  assign y9183 = n31359 ;
  assign y9184 = ~n31361 ;
  assign y9185 = ~n31363 ;
  assign y9186 = ~n31364 ;
  assign y9187 = ~n31365 ;
  assign y9188 = n31370 ;
  assign y9189 = ~n31371 ;
  assign y9190 = n31372 ;
  assign y9191 = n31374 ;
  assign y9192 = n31377 ;
  assign y9193 = n31380 ;
  assign y9194 = ~1'b0 ;
  assign y9195 = n31383 ;
  assign y9196 = n31390 ;
  assign y9197 = ~n31391 ;
  assign y9198 = n31392 ;
  assign y9199 = n31395 ;
  assign y9200 = ~n31398 ;
  assign y9201 = ~n31399 ;
  assign y9202 = ~n31400 ;
  assign y9203 = ~n31402 ;
  assign y9204 = ~n31404 ;
  assign y9205 = ~1'b0 ;
  assign y9206 = ~n31409 ;
  assign y9207 = n31410 ;
  assign y9208 = ~n31412 ;
  assign y9209 = n31413 ;
  assign y9210 = n31415 ;
  assign y9211 = ~n31417 ;
  assign y9212 = ~n31419 ;
  assign y9213 = n31421 ;
  assign y9214 = ~n31424 ;
  assign y9215 = ~1'b0 ;
  assign y9216 = ~n31426 ;
  assign y9217 = n31428 ;
  assign y9218 = n31432 ;
  assign y9219 = n31433 ;
  assign y9220 = ~n31435 ;
  assign y9221 = ~n31439 ;
  assign y9222 = ~n31440 ;
  assign y9223 = ~n31441 ;
  assign y9224 = ~n31442 ;
  assign y9225 = n31444 ;
  assign y9226 = ~n31448 ;
  assign y9227 = n31450 ;
  assign y9228 = n31452 ;
  assign y9229 = ~n31458 ;
  assign y9230 = ~n31460 ;
  assign y9231 = ~n31464 ;
  assign y9232 = n31466 ;
  assign y9233 = n31470 ;
  assign y9234 = ~n31474 ;
  assign y9235 = ~n31475 ;
  assign y9236 = n31477 ;
  assign y9237 = n31480 ;
  assign y9238 = ~1'b0 ;
  assign y9239 = n31483 ;
  assign y9240 = n31484 ;
  assign y9241 = n31486 ;
  assign y9242 = n31493 ;
  assign y9243 = ~n31496 ;
  assign y9244 = ~n31503 ;
  assign y9245 = n31510 ;
  assign y9246 = ~n31511 ;
  assign y9247 = n31513 ;
  assign y9248 = n31514 ;
  assign y9249 = ~n31515 ;
  assign y9250 = ~n31517 ;
  assign y9251 = n31519 ;
  assign y9252 = ~n31520 ;
  assign y9253 = ~n31521 ;
  assign y9254 = n31523 ;
  assign y9255 = ~1'b0 ;
  assign y9256 = n31525 ;
  assign y9257 = n31528 ;
  assign y9258 = n31529 ;
  assign y9259 = ~n31538 ;
  assign y9260 = ~n31539 ;
  assign y9261 = ~n31541 ;
  assign y9262 = n31542 ;
  assign y9263 = ~n31546 ;
  assign y9264 = ~n31550 ;
  assign y9265 = ~1'b0 ;
  assign y9266 = n31551 ;
  assign y9267 = ~n31553 ;
  assign y9268 = n31556 ;
  assign y9269 = n31563 ;
  assign y9270 = n31569 ;
  assign y9271 = ~n31570 ;
  assign y9272 = ~n31571 ;
  assign y9273 = n31572 ;
  assign y9274 = n31577 ;
  assign y9275 = ~n31579 ;
  assign y9276 = n31584 ;
  assign y9277 = n11664 ;
  assign y9278 = n31590 ;
  assign y9279 = n31591 ;
  assign y9280 = n31596 ;
  assign y9281 = n31597 ;
  assign y9282 = n31598 ;
  assign y9283 = n31604 ;
  assign y9284 = ~n31606 ;
  assign y9285 = ~n31607 ;
  assign y9286 = n31608 ;
  assign y9287 = n31610 ;
  assign y9288 = n31612 ;
  assign y9289 = n31614 ;
  assign y9290 = ~n31615 ;
  assign y9291 = n31616 ;
  assign y9292 = n31617 ;
  assign y9293 = ~n31620 ;
  assign y9294 = n31621 ;
  assign y9295 = n31624 ;
  assign y9296 = ~n31625 ;
  assign y9297 = ~n31627 ;
  assign y9298 = ~n31631 ;
  assign y9299 = ~1'b0 ;
  assign y9300 = 1'b0 ;
  assign y9301 = n31632 ;
  assign y9302 = n31633 ;
  assign y9303 = ~n31634 ;
  assign y9304 = n31635 ;
  assign y9305 = ~n31636 ;
  assign y9306 = ~n31638 ;
  assign y9307 = n31639 ;
  assign y9308 = ~n31647 ;
  assign y9309 = ~n31649 ;
  assign y9310 = n31652 ;
  assign y9311 = ~n31653 ;
  assign y9312 = ~n31654 ;
  assign y9313 = ~n31656 ;
  assign y9314 = ~n31660 ;
  assign y9315 = ~n31661 ;
  assign y9316 = ~n31662 ;
  assign y9317 = ~n31664 ;
  assign y9318 = n31665 ;
  assign y9319 = ~n31667 ;
  assign y9320 = ~n31669 ;
  assign y9321 = ~n31673 ;
  assign y9322 = ~n31676 ;
  assign y9323 = ~n31677 ;
  assign y9324 = ~n31679 ;
  assign y9325 = n31682 ;
  assign y9326 = ~n31685 ;
  assign y9327 = ~n31687 ;
  assign y9328 = n31689 ;
  assign y9329 = ~n31691 ;
  assign y9330 = n31695 ;
  assign y9331 = ~n31697 ;
  assign y9332 = ~n31702 ;
  assign y9333 = ~n31703 ;
  assign y9334 = ~n31706 ;
  assign y9335 = ~n31707 ;
  assign y9336 = ~n31709 ;
  assign y9337 = ~n31712 ;
  assign y9338 = n31714 ;
  assign y9339 = ~n31716 ;
  assign y9340 = n31720 ;
  assign y9341 = ~1'b0 ;
  assign y9342 = ~1'b0 ;
  assign y9343 = n31724 ;
  assign y9344 = n31725 ;
  assign y9345 = n31727 ;
  assign y9346 = ~n31729 ;
  assign y9347 = n31730 ;
  assign y9348 = ~1'b0 ;
  assign y9349 = ~n31731 ;
  assign y9350 = ~n31732 ;
  assign y9351 = ~n31738 ;
  assign y9352 = n31740 ;
  assign y9353 = ~n31743 ;
  assign y9354 = ~n31744 ;
  assign y9355 = n31746 ;
  assign y9356 = n31750 ;
  assign y9357 = ~n31754 ;
  assign y9358 = n31757 ;
  assign y9359 = ~n31758 ;
  assign y9360 = n31760 ;
  assign y9361 = ~n31762 ;
  assign y9362 = n31764 ;
  assign y9363 = n31766 ;
  assign y9364 = ~1'b0 ;
  assign y9365 = ~n31769 ;
  assign y9366 = n31770 ;
  assign y9367 = ~n31771 ;
  assign y9368 = n31772 ;
  assign y9369 = ~n31773 ;
  assign y9370 = ~n31779 ;
  assign y9371 = n31780 ;
  assign y9372 = n31783 ;
  assign y9373 = ~n31785 ;
  assign y9374 = ~n31790 ;
  assign y9375 = n31792 ;
  assign y9376 = n31793 ;
  assign y9377 = n31794 ;
  assign y9378 = n31795 ;
  assign y9379 = n31796 ;
  assign y9380 = n31803 ;
  assign y9381 = ~n31805 ;
  assign y9382 = n31806 ;
  assign y9383 = n31808 ;
  assign y9384 = ~n31810 ;
  assign y9385 = ~1'b0 ;
  assign y9386 = ~1'b0 ;
  assign y9387 = ~n31812 ;
  assign y9388 = ~n31814 ;
  assign y9389 = ~n31815 ;
  assign y9390 = n31818 ;
  assign y9391 = ~n31819 ;
  assign y9392 = ~n31822 ;
  assign y9393 = ~n31823 ;
  assign y9394 = n31829 ;
  assign y9395 = ~n31832 ;
  assign y9396 = ~n31835 ;
  assign y9397 = ~1'b0 ;
  assign y9398 = ~n31836 ;
  assign y9399 = n31841 ;
  assign y9400 = n31845 ;
  assign y9401 = ~n31847 ;
  assign y9402 = n31848 ;
  assign y9403 = ~n31850 ;
  assign y9404 = n31851 ;
  assign y9405 = n31854 ;
  assign y9406 = n31856 ;
  assign y9407 = n31858 ;
  assign y9408 = n31859 ;
  assign y9409 = ~n31861 ;
  assign y9410 = ~n31863 ;
  assign y9411 = n31864 ;
  assign y9412 = n31869 ;
  assign y9413 = n31870 ;
  assign y9414 = ~n31872 ;
  assign y9415 = ~n31873 ;
  assign y9416 = ~n31877 ;
  assign y9417 = n31880 ;
  assign y9418 = n31881 ;
  assign y9419 = ~n31883 ;
  assign y9420 = ~n31887 ;
  assign y9421 = ~n31889 ;
  assign y9422 = ~n31893 ;
  assign y9423 = ~n31897 ;
  assign y9424 = n31898 ;
  assign y9425 = n31899 ;
  assign y9426 = ~n31900 ;
  assign y9427 = ~1'b0 ;
  assign y9428 = n31902 ;
  assign y9429 = n31904 ;
  assign y9430 = n31908 ;
  assign y9431 = n31909 ;
  assign y9432 = n31911 ;
  assign y9433 = n31914 ;
  assign y9434 = ~n31918 ;
  assign y9435 = n31921 ;
  assign y9436 = ~n31924 ;
  assign y9437 = ~1'b0 ;
  assign y9438 = n31928 ;
  assign y9439 = n31929 ;
  assign y9440 = ~n31930 ;
  assign y9441 = n31931 ;
  assign y9442 = ~n31934 ;
  assign y9443 = ~n31938 ;
  assign y9444 = n31943 ;
  assign y9445 = ~n31947 ;
  assign y9446 = n31950 ;
  assign y9447 = n31952 ;
  assign y9448 = ~1'b0 ;
  assign y9449 = ~1'b0 ;
  assign y9450 = ~1'b0 ;
  assign y9451 = ~n31953 ;
  assign y9452 = ~n31956 ;
  assign y9453 = ~n31958 ;
  assign y9454 = ~n31961 ;
  assign y9455 = ~n31964 ;
  assign y9456 = ~n31965 ;
  assign y9457 = n31966 ;
  assign y9458 = n31968 ;
  assign y9459 = ~1'b0 ;
  assign y9460 = ~1'b0 ;
  assign y9461 = n31969 ;
  assign y9462 = n31970 ;
  assign y9463 = ~n31972 ;
  assign y9464 = ~n31973 ;
  assign y9465 = ~n31974 ;
  assign y9466 = n31975 ;
  assign y9467 = ~n31976 ;
  assign y9468 = ~n31978 ;
  assign y9469 = n31980 ;
  assign y9470 = ~n31982 ;
  assign y9471 = ~1'b0 ;
  assign y9472 = ~n31983 ;
  assign y9473 = ~n31984 ;
  assign y9474 = ~n31986 ;
  assign y9475 = n31988 ;
  assign y9476 = n31990 ;
  assign y9477 = ~n31996 ;
  assign y9478 = ~n31997 ;
  assign y9479 = ~n31999 ;
  assign y9480 = n32002 ;
  assign y9481 = ~n32004 ;
  assign y9482 = ~n32009 ;
  assign y9483 = ~n32010 ;
  assign y9484 = ~n32011 ;
  assign y9485 = n32013 ;
  assign y9486 = n32017 ;
  assign y9487 = n32020 ;
  assign y9488 = ~n32023 ;
  assign y9489 = n32025 ;
  assign y9490 = ~n32026 ;
  assign y9491 = ~1'b0 ;
  assign y9492 = ~1'b0 ;
  assign y9493 = n32030 ;
  assign y9494 = ~n32032 ;
  assign y9495 = n32035 ;
  assign y9496 = n32037 ;
  assign y9497 = n32041 ;
  assign y9498 = ~n32042 ;
  assign y9499 = ~n32045 ;
  assign y9500 = ~n32046 ;
  assign y9501 = n32047 ;
  assign y9502 = ~n32049 ;
  assign y9503 = ~n32053 ;
  assign y9504 = n32057 ;
  assign y9505 = n32058 ;
  assign y9506 = ~n32059 ;
  assign y9507 = ~n32063 ;
  assign y9508 = ~n32074 ;
  assign y9509 = ~n32078 ;
  assign y9510 = ~n32080 ;
  assign y9511 = n32081 ;
  assign y9512 = ~n32082 ;
  assign y9513 = ~n32088 ;
  assign y9514 = n32090 ;
  assign y9515 = n32093 ;
  assign y9516 = ~n32096 ;
  assign y9517 = ~n32097 ;
  assign y9518 = n32100 ;
  assign y9519 = ~n32101 ;
  assign y9520 = ~n32102 ;
  assign y9521 = ~n32105 ;
  assign y9522 = n32106 ;
  assign y9523 = ~n32110 ;
  assign y9524 = n32112 ;
  assign y9525 = ~1'b0 ;
  assign y9526 = n32114 ;
  assign y9527 = n32116 ;
  assign y9528 = ~n32121 ;
  assign y9529 = ~n32126 ;
  assign y9530 = ~n32127 ;
  assign y9531 = n32131 ;
  assign y9532 = n32133 ;
  assign y9533 = ~n32134 ;
  assign y9534 = n32136 ;
  assign y9535 = ~n32138 ;
  assign y9536 = n32140 ;
  assign y9537 = ~1'b0 ;
  assign y9538 = ~n32146 ;
  assign y9539 = n32147 ;
  assign y9540 = ~n32148 ;
  assign y9541 = n32149 ;
  assign y9542 = n32152 ;
  assign y9543 = ~n32154 ;
  assign y9544 = ~n32156 ;
  assign y9545 = n32163 ;
  assign y9546 = ~n32165 ;
  assign y9547 = ~1'b0 ;
  assign y9548 = n32167 ;
  assign y9549 = n32168 ;
  assign y9550 = n32170 ;
  assign y9551 = n32171 ;
  assign y9552 = n32174 ;
  assign y9553 = n32176 ;
  assign y9554 = n32177 ;
  assign y9555 = ~n32183 ;
  assign y9556 = n32184 ;
  assign y9557 = ~n32186 ;
  assign y9558 = n32188 ;
  assign y9559 = ~n32190 ;
  assign y9560 = n32196 ;
  assign y9561 = n32199 ;
  assign y9562 = ~n32202 ;
  assign y9563 = ~n32203 ;
  assign y9564 = n32204 ;
  assign y9565 = ~n32206 ;
  assign y9566 = ~n32207 ;
  assign y9567 = n32214 ;
  assign y9568 = ~n32216 ;
  assign y9569 = n32218 ;
  assign y9570 = ~n32221 ;
  assign y9571 = n32222 ;
  assign y9572 = n32223 ;
  assign y9573 = n32225 ;
  assign y9574 = n31197 ;
  assign y9575 = ~n32227 ;
  assign y9576 = ~n32230 ;
  assign y9577 = n32231 ;
  assign y9578 = ~n32232 ;
  assign y9579 = ~n32233 ;
  assign y9580 = n32236 ;
  assign y9581 = n32239 ;
  assign y9582 = ~n32240 ;
  assign y9583 = ~n32243 ;
  assign y9584 = n32244 ;
  assign y9585 = ~n32248 ;
  assign y9586 = ~n32251 ;
  assign y9587 = n32253 ;
  assign y9588 = n32254 ;
  assign y9589 = ~n32257 ;
  assign y9590 = ~n32260 ;
  assign y9591 = ~n32262 ;
  assign y9592 = ~n32264 ;
  assign y9593 = n32266 ;
  assign y9594 = ~n32267 ;
  assign y9595 = ~n32269 ;
  assign y9596 = ~n32271 ;
  assign y9597 = n32272 ;
  assign y9598 = n32276 ;
  assign y9599 = n32277 ;
  assign y9600 = n32279 ;
  assign y9601 = ~n32283 ;
  assign y9602 = ~n32285 ;
  assign y9603 = n32291 ;
  assign y9604 = ~n32292 ;
  assign y9605 = ~n32293 ;
  assign y9606 = ~n32294 ;
  assign y9607 = ~n32295 ;
  assign y9608 = n32297 ;
  assign y9609 = ~n32300 ;
  assign y9610 = n32301 ;
  assign y9611 = n32303 ;
  assign y9612 = n32305 ;
  assign y9613 = ~1'b0 ;
  assign y9614 = n32306 ;
  assign y9615 = n32309 ;
  assign y9616 = n32310 ;
  assign y9617 = n32311 ;
  assign y9618 = n32312 ;
  assign y9619 = n32314 ;
  assign y9620 = n32323 ;
  assign y9621 = ~n32324 ;
  assign y9622 = n32326 ;
  assign y9623 = ~n32328 ;
  assign y9624 = ~1'b0 ;
  assign y9625 = ~n32329 ;
  assign y9626 = n32330 ;
  assign y9627 = n32331 ;
  assign y9628 = ~n32335 ;
  assign y9629 = ~n32338 ;
  assign y9630 = n32340 ;
  assign y9631 = ~n32345 ;
  assign y9632 = ~n32346 ;
  assign y9633 = ~n32350 ;
  assign y9634 = ~1'b0 ;
  assign y9635 = n32352 ;
  assign y9636 = n32353 ;
  assign y9637 = n32355 ;
  assign y9638 = n32361 ;
  assign y9639 = ~n32364 ;
  assign y9640 = ~n32365 ;
  assign y9641 = ~n32367 ;
  assign y9642 = n32370 ;
  assign y9643 = ~n32371 ;
  assign y9644 = ~n32377 ;
  assign y9645 = n32379 ;
  assign y9646 = ~n32381 ;
  assign y9647 = n32383 ;
  assign y9648 = ~n32386 ;
  assign y9649 = ~n32388 ;
  assign y9650 = ~n32392 ;
  assign y9651 = ~n32396 ;
  assign y9652 = ~n32397 ;
  assign y9653 = ~n32404 ;
  assign y9654 = ~n32406 ;
  assign y9655 = n32409 ;
  assign y9656 = n32411 ;
  assign y9657 = ~1'b0 ;
endmodule
