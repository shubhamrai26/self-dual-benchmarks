module top( x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 , y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 );
  input x0 , x1 , x2 , x3 , x4 , x5 , x6 , x7 , x8 , x9 , x10 , x11 , x12 , x13 , x14 , x15 , x16 , x17 , x18 , x19 , x20 , x21 , x22 , x23 , x24 , x25 , x26 , x27 , x28 , x29 , x30 , x31 , x32 , x33 , x34 , x35 , x36 , x37 , x38 , x39 , x40 , x41 , x42 , x43 , x44 , x45 , x46 , x47 , x48 , x49 , x50 , x51 , x52 , x53 , x54 , x55 , x56 , x57 , x58 , x59 , x60 , x61 , x62 , x63 , x64 , x65 , x66 , x67 , x68 , x69 , x70 , x71 , x72 , x73 , x74 , x75 , x76 , x77 , x78 , x79 , x80 , x81 , x82 , x83 , x84 , x85 , x86 , x87 , x88 , x89 , x90 , x91 , x92 , x93 , x94 , x95 , x96 , x97 , x98 , x99 , x100 , x101 , x102 , x103 , x104 , x105 , x106 , x107 , x108 , x109 , x110 , x111 , x112 , x113 , x114 , x115 , x116 , x117 , x118 , x119 , x120 , x121 , x122 , x123 , x124 , x125 , x126 , x127 ;
  output y0 , y1 , y2 , y3 , y4 , y5 , y6 , y7 , y8 , y9 , y10 , y11 , y12 , y13 , y14 , y15 , y16 , y17 , y18 , y19 , y20 , y21 , y22 , y23 , y24 , y25 , y26 , y27 , y28 , y29 , y30 , y31 , y32 , y33 , y34 , y35 , y36 , y37 , y38 , y39 , y40 , y41 , y42 , y43 , y44 , y45 , y46 , y47 , y48 , y49 , y50 , y51 , y52 , y53 , y54 , y55 , y56 , y57 , y58 , y59 , y60 , y61 , y62 , y63 , y64 , y65 , y66 , y67 , y68 , y69 , y70 , y71 , y72 , y73 , y74 , y75 , y76 , y77 , y78 , y79 , y80 , y81 , y82 , y83 , y84 , y85 , y86 , y87 , y88 , y89 , y90 , y91 , y92 , y93 , y94 , y95 , y96 , y97 , y98 , y99 , y100 , y101 , y102 , y103 , y104 , y105 , y106 , y107 , y108 , y109 , y110 , y111 , y112 , y113 , y114 , y115 , y116 , y117 , y118 , y119 , y120 , y121 , y122 , y123 , y124 , y125 , y126 , y127 , y128 , y129 , y130 , y131 , y132 , y133 , y134 , y135 , y136 , y137 , y138 , y139 , y140 , y141 , y142 , y143 , y144 , y145 , y146 , y147 , y148 , y149 , y150 , y151 , y152 , y153 , y154 , y155 , y156 , y157 , y158 , y159 , y160 , y161 , y162 , y163 , y164 , y165 , y166 , y167 , y168 , y169 , y170 , y171 , y172 , y173 , y174 , y175 , y176 , y177 , y178 , y179 , y180 , y181 , y182 , y183 , y184 , y185 , y186 , y187 , y188 , y189 , y190 , y191 , y192 , y193 , y194 , y195 , y196 , y197 , y198 , y199 , y200 , y201 , y202 , y203 , y204 , y205 , y206 , y207 , y208 , y209 , y210 , y211 , y212 , y213 , y214 , y215 , y216 , y217 , y218 , y219 , y220 , y221 , y222 , y223 , y224 , y225 , y226 , y227 , y228 , y229 , y230 , y231 , y232 , y233 , y234 , y235 , y236 , y237 , y238 , y239 , y240 , y241 , y242 , y243 , y244 , y245 , y246 , y247 , y248 , y249 , y250 , y251 , y252 , y253 , y254 , y255 , y256 , y257 , y258 , y259 , y260 , y261 , y262 , y263 , y264 , y265 , y266 , y267 , y268 , y269 , y270 , y271 , y272 , y273 , y274 , y275 , y276 , y277 , y278 , y279 , y280 , y281 , y282 , y283 , y284 , y285 , y286 , y287 , y288 , y289 , y290 , y291 , y292 , y293 , y294 , y295 , y296 , y297 , y298 , y299 , y300 , y301 , y302 , y303 , y304 , y305 , y306 , y307 , y308 , y309 , y310 , y311 , y312 , y313 , y314 , y315 , y316 , y317 , y318 , y319 , y320 , y321 , y322 , y323 , y324 , y325 , y326 , y327 , y328 , y329 , y330 , y331 , y332 , y333 , y334 , y335 , y336 , y337 , y338 , y339 , y340 , y341 , y342 , y343 , y344 , y345 , y346 , y347 , y348 , y349 , y350 , y351 , y352 , y353 , y354 , y355 , y356 , y357 , y358 , y359 , y360 , y361 , y362 , y363 , y364 , y365 , y366 , y367 , y368 , y369 , y370 , y371 , y372 , y373 , y374 , y375 , y376 , y377 , y378 , y379 , y380 , y381 , y382 , y383 , y384 , y385 , y386 , y387 , y388 , y389 , y390 , y391 , y392 , y393 , y394 , y395 , y396 , y397 , y398 , y399 , y400 , y401 , y402 , y403 , y404 , y405 , y406 , y407 , y408 , y409 , y410 , y411 , y412 , y413 , y414 , y415 , y416 , y417 , y418 , y419 , y420 , y421 , y422 , y423 , y424 , y425 , y426 , y427 , y428 , y429 , y430 , y431 , y432 , y433 , y434 , y435 , y436 , y437 , y438 , y439 , y440 , y441 , y442 , y443 , y444 , y445 , y446 , y447 , y448 , y449 , y450 , y451 , y452 , y453 , y454 , y455 , y456 , y457 , y458 , y459 , y460 , y461 , y462 , y463 , y464 , y465 , y466 , y467 , y468 , y469 , y470 , y471 , y472 , y473 , y474 , y475 , y476 , y477 , y478 , y479 , y480 , y481 , y482 , y483 , y484 , y485 , y486 , y487 , y488 , y489 , y490 , y491 , y492 , y493 , y494 , y495 , y496 , y497 , y498 , y499 , y500 , y501 , y502 , y503 , y504 , y505 , y506 , y507 , y508 , y509 , y510 , y511 , y512 , y513 , y514 , y515 , y516 , y517 , y518 , y519 , y520 , y521 , y522 , y523 , y524 , y525 , y526 , y527 , y528 , y529 , y530 , y531 , y532 , y533 , y534 , y535 , y536 , y537 , y538 , y539 , y540 , y541 , y542 , y543 , y544 , y545 , y546 , y547 , y548 , y549 , y550 , y551 , y552 , y553 , y554 , y555 , y556 , y557 , y558 , y559 , y560 , y561 , y562 , y563 , y564 , y565 , y566 , y567 , y568 , y569 , y570 , y571 , y572 , y573 , y574 , y575 , y576 , y577 , y578 , y579 , y580 , y581 , y582 , y583 , y584 , y585 , y586 , y587 , y588 , y589 , y590 , y591 , y592 , y593 , y594 , y595 , y596 , y597 , y598 , y599 , y600 , y601 , y602 , y603 , y604 , y605 , y606 , y607 , y608 , y609 , y610 , y611 , y612 , y613 , y614 , y615 , y616 , y617 , y618 , y619 , y620 , y621 , y622 , y623 , y624 , y625 , y626 , y627 , y628 , y629 , y630 , y631 , y632 , y633 , y634 , y635 , y636 , y637 , y638 , y639 , y640 , y641 , y642 , y643 , y644 , y645 , y646 , y647 , y648 , y649 , y650 , y651 , y652 , y653 , y654 , y655 , y656 , y657 , y658 , y659 , y660 , y661 , y662 , y663 , y664 , y665 , y666 , y667 , y668 , y669 , y670 , y671 , y672 , y673 , y674 , y675 , y676 , y677 , y678 , y679 , y680 , y681 , y682 , y683 , y684 , y685 , y686 , y687 , y688 , y689 , y690 , y691 , y692 , y693 , y694 , y695 , y696 , y697 , y698 , y699 , y700 , y701 , y702 , y703 , y704 , y705 , y706 , y707 , y708 , y709 , y710 , y711 , y712 , y713 , y714 , y715 , y716 , y717 , y718 , y719 , y720 , y721 , y722 , y723 , y724 , y725 , y726 , y727 , y728 , y729 , y730 , y731 , y732 , y733 , y734 , y735 , y736 , y737 , y738 , y739 , y740 , y741 , y742 , y743 , y744 , y745 , y746 , y747 , y748 , y749 , y750 , y751 , y752 , y753 , y754 , y755 , y756 , y757 , y758 , y759 , y760 , y761 , y762 , y763 , y764 , y765 , y766 , y767 , y768 , y769 , y770 , y771 , y772 , y773 , y774 , y775 , y776 , y777 , y778 , y779 , y780 , y781 , y782 , y783 , y784 , y785 , y786 , y787 , y788 , y789 , y790 , y791 , y792 , y793 , y794 , y795 , y796 , y797 , y798 , y799 , y800 , y801 , y802 , y803 , y804 , y805 , y806 , y807 , y808 , y809 , y810 , y811 , y812 , y813 , y814 , y815 , y816 , y817 , y818 , y819 , y820 , y821 , y822 , y823 , y824 , y825 , y826 , y827 , y828 , y829 , y830 , y831 , y832 , y833 , y834 , y835 , y836 , y837 , y838 , y839 , y840 , y841 , y842 , y843 , y844 , y845 , y846 , y847 , y848 , y849 , y850 , y851 , y852 , y853 , y854 , y855 , y856 , y857 , y858 , y859 , y860 , y861 , y862 , y863 , y864 , y865 , y866 , y867 , y868 , y869 , y870 , y871 , y872 , y873 , y874 , y875 , y876 , y877 , y878 , y879 , y880 , y881 , y882 , y883 , y884 , y885 , y886 , y887 , y888 , y889 , y890 , y891 , y892 , y893 , y894 , y895 , y896 , y897 , y898 , y899 , y900 , y901 , y902 , y903 , y904 , y905 , y906 , y907 , y908 , y909 , y910 , y911 , y912 , y913 , y914 , y915 , y916 , y917 , y918 , y919 , y920 , y921 , y922 , y923 , y924 , y925 , y926 , y927 , y928 , y929 , y930 , y931 , y932 , y933 , y934 , y935 , y936 , y937 , y938 , y939 , y940 , y941 , y942 , y943 , y944 , y945 , y946 , y947 , y948 , y949 , y950 , y951 , y952 , y953 , y954 , y955 , y956 , y957 , y958 , y959 , y960 , y961 , y962 , y963 , y964 , y965 , y966 , y967 , y968 , y969 , y970 , y971 , y972 , y973 , y974 , y975 , y976 , y977 , y978 , y979 , y980 , y981 , y982 , y983 , y984 , y985 , y986 , y987 , y988 , y989 , y990 , y991 , y992 , y993 , y994 , y995 , y996 , y997 , y998 , y999 , y1000 , y1001 , y1002 , y1003 , y1004 , y1005 , y1006 , y1007 , y1008 , y1009 , y1010 , y1011 , y1012 , y1013 , y1014 , y1015 , y1016 , y1017 , y1018 , y1019 , y1020 , y1021 , y1022 , y1023 , y1024 , y1025 , y1026 , y1027 , y1028 , y1029 , y1030 , y1031 , y1032 , y1033 , y1034 , y1035 , y1036 , y1037 , y1038 , y1039 , y1040 , y1041 , y1042 , y1043 , y1044 , y1045 , y1046 , y1047 , y1048 , y1049 , y1050 , y1051 , y1052 , y1053 , y1054 , y1055 , y1056 , y1057 , y1058 , y1059 , y1060 , y1061 , y1062 , y1063 , y1064 , y1065 , y1066 , y1067 , y1068 , y1069 , y1070 , y1071 , y1072 , y1073 , y1074 , y1075 , y1076 , y1077 , y1078 , y1079 , y1080 , y1081 , y1082 , y1083 , y1084 , y1085 , y1086 , y1087 , y1088 , y1089 , y1090 , y1091 , y1092 , y1093 , y1094 , y1095 , y1096 , y1097 , y1098 , y1099 , y1100 , y1101 , y1102 , y1103 , y1104 , y1105 , y1106 , y1107 , y1108 , y1109 , y1110 , y1111 , y1112 , y1113 , y1114 , y1115 , y1116 , y1117 , y1118 , y1119 , y1120 , y1121 , y1122 , y1123 , y1124 , y1125 , y1126 , y1127 , y1128 , y1129 , y1130 , y1131 , y1132 , y1133 , y1134 , y1135 , y1136 , y1137 , y1138 , y1139 , y1140 , y1141 , y1142 , y1143 , y1144 , y1145 , y1146 , y1147 , y1148 , y1149 , y1150 , y1151 , y1152 , y1153 , y1154 , y1155 , y1156 , y1157 , y1158 , y1159 , y1160 , y1161 , y1162 , y1163 , y1164 , y1165 , y1166 , y1167 , y1168 , y1169 , y1170 , y1171 , y1172 , y1173 , y1174 , y1175 , y1176 , y1177 , y1178 , y1179 , y1180 , y1181 , y1182 , y1183 , y1184 , y1185 , y1186 , y1187 , y1188 , y1189 , y1190 , y1191 , y1192 , y1193 , y1194 , y1195 , y1196 , y1197 , y1198 , y1199 , y1200 , y1201 , y1202 , y1203 , y1204 , y1205 , y1206 , y1207 , y1208 , y1209 , y1210 , y1211 , y1212 , y1213 , y1214 , y1215 , y1216 , y1217 , y1218 , y1219 , y1220 , y1221 , y1222 , y1223 , y1224 , y1225 , y1226 , y1227 , y1228 , y1229 , y1230 , y1231 , y1232 , y1233 , y1234 , y1235 , y1236 , y1237 , y1238 , y1239 , y1240 , y1241 , y1242 , y1243 , y1244 , y1245 , y1246 , y1247 , y1248 , y1249 , y1250 , y1251 , y1252 , y1253 , y1254 , y1255 , y1256 , y1257 , y1258 , y1259 , y1260 , y1261 , y1262 , y1263 , y1264 , y1265 , y1266 , y1267 , y1268 , y1269 , y1270 , y1271 , y1272 , y1273 , y1274 , y1275 , y1276 , y1277 , y1278 , y1279 , y1280 , y1281 , y1282 , y1283 , y1284 , y1285 , y1286 , y1287 , y1288 , y1289 , y1290 , y1291 , y1292 , y1293 , y1294 , y1295 , y1296 , y1297 , y1298 , y1299 , y1300 , y1301 , y1302 , y1303 , y1304 , y1305 , y1306 , y1307 , y1308 , y1309 , y1310 , y1311 , y1312 , y1313 , y1314 , y1315 , y1316 , y1317 , y1318 , y1319 , y1320 , y1321 , y1322 , y1323 , y1324 , y1325 , y1326 , y1327 , y1328 , y1329 , y1330 , y1331 , y1332 , y1333 , y1334 , y1335 , y1336 , y1337 , y1338 , y1339 , y1340 , y1341 , y1342 , y1343 , y1344 , y1345 , y1346 , y1347 , y1348 , y1349 , y1350 , y1351 , y1352 , y1353 , y1354 , y1355 , y1356 , y1357 , y1358 , y1359 , y1360 , y1361 , y1362 , y1363 , y1364 , y1365 , y1366 , y1367 , y1368 , y1369 , y1370 , y1371 , y1372 , y1373 , y1374 , y1375 , y1376 , y1377 , y1378 , y1379 , y1380 , y1381 , y1382 , y1383 , y1384 , y1385 , y1386 , y1387 , y1388 , y1389 , y1390 , y1391 , y1392 , y1393 , y1394 , y1395 , y1396 , y1397 , y1398 , y1399 , y1400 , y1401 , y1402 , y1403 , y1404 , y1405 , y1406 , y1407 , y1408 , y1409 , y1410 , y1411 , y1412 , y1413 , y1414 , y1415 , y1416 , y1417 , y1418 , y1419 , y1420 , y1421 , y1422 , y1423 , y1424 , y1425 , y1426 , y1427 , y1428 , y1429 , y1430 , y1431 , y1432 , y1433 , y1434 , y1435 , y1436 , y1437 , y1438 , y1439 , y1440 , y1441 , y1442 , y1443 , y1444 , y1445 , y1446 , y1447 , y1448 , y1449 , y1450 , y1451 , y1452 , y1453 , y1454 , y1455 , y1456 , y1457 , y1458 , y1459 , y1460 , y1461 , y1462 , y1463 , y1464 , y1465 , y1466 , y1467 , y1468 , y1469 , y1470 , y1471 , y1472 , y1473 , y1474 , y1475 , y1476 , y1477 , y1478 , y1479 , y1480 , y1481 , y1482 , y1483 , y1484 , y1485 , y1486 , y1487 , y1488 , y1489 , y1490 , y1491 , y1492 , y1493 , y1494 , y1495 , y1496 , y1497 , y1498 , y1499 , y1500 , y1501 , y1502 , y1503 , y1504 , y1505 , y1506 , y1507 , y1508 , y1509 , y1510 , y1511 , y1512 , y1513 , y1514 , y1515 , y1516 , y1517 , y1518 , y1519 , y1520 , y1521 , y1522 , y1523 , y1524 , y1525 , y1526 , y1527 , y1528 , y1529 , y1530 , y1531 , y1532 , y1533 , y1534 , y1535 , y1536 , y1537 , y1538 , y1539 , y1540 , y1541 , y1542 , y1543 , y1544 , y1545 , y1546 , y1547 , y1548 , y1549 , y1550 , y1551 , y1552 , y1553 , y1554 , y1555 , y1556 , y1557 , y1558 , y1559 , y1560 , y1561 , y1562 , y1563 , y1564 , y1565 , y1566 , y1567 , y1568 , y1569 , y1570 , y1571 , y1572 , y1573 , y1574 , y1575 , y1576 , y1577 , y1578 , y1579 , y1580 , y1581 , y1582 , y1583 , y1584 , y1585 , y1586 , y1587 , y1588 , y1589 , y1590 , y1591 , y1592 , y1593 , y1594 , y1595 , y1596 , y1597 , y1598 , y1599 , y1600 , y1601 , y1602 , y1603 , y1604 , y1605 , y1606 , y1607 , y1608 , y1609 , y1610 , y1611 , y1612 , y1613 , y1614 , y1615 , y1616 , y1617 , y1618 , y1619 , y1620 , y1621 , y1622 , y1623 , y1624 , y1625 , y1626 , y1627 , y1628 , y1629 , y1630 , y1631 , y1632 , y1633 , y1634 , y1635 , y1636 , y1637 , y1638 , y1639 , y1640 , y1641 , y1642 , y1643 , y1644 , y1645 , y1646 , y1647 , y1648 , y1649 , y1650 , y1651 , y1652 , y1653 , y1654 , y1655 , y1656 , y1657 , y1658 , y1659 , y1660 , y1661 , y1662 , y1663 , y1664 , y1665 , y1666 , y1667 , y1668 , y1669 , y1670 , y1671 , y1672 , y1673 , y1674 , y1675 , y1676 , y1677 , y1678 , y1679 , y1680 , y1681 , y1682 , y1683 , y1684 , y1685 , y1686 , y1687 , y1688 , y1689 , y1690 , y1691 , y1692 , y1693 , y1694 , y1695 , y1696 , y1697 , y1698 , y1699 , y1700 , y1701 , y1702 , y1703 , y1704 , y1705 , y1706 , y1707 , y1708 , y1709 , y1710 , y1711 , y1712 , y1713 , y1714 , y1715 , y1716 , y1717 , y1718 , y1719 , y1720 , y1721 , y1722 , y1723 , y1724 , y1725 , y1726 , y1727 , y1728 , y1729 , y1730 , y1731 , y1732 , y1733 , y1734 , y1735 , y1736 , y1737 , y1738 , y1739 , y1740 , y1741 , y1742 , y1743 , y1744 , y1745 , y1746 , y1747 , y1748 , y1749 , y1750 , y1751 , y1752 , y1753 , y1754 , y1755 , y1756 , y1757 , y1758 , y1759 , y1760 , y1761 , y1762 , y1763 , y1764 , y1765 , y1766 , y1767 , y1768 , y1769 , y1770 , y1771 , y1772 , y1773 , y1774 , y1775 , y1776 , y1777 , y1778 , y1779 , y1780 , y1781 , y1782 , y1783 , y1784 , y1785 , y1786 , y1787 , y1788 , y1789 , y1790 , y1791 , y1792 , y1793 , y1794 , y1795 , y1796 , y1797 , y1798 , y1799 , y1800 , y1801 , y1802 , y1803 , y1804 , y1805 , y1806 , y1807 , y1808 , y1809 , y1810 , y1811 , y1812 , y1813 , y1814 , y1815 , y1816 , y1817 , y1818 , y1819 , y1820 , y1821 , y1822 , y1823 , y1824 , y1825 , y1826 , y1827 , y1828 , y1829 , y1830 , y1831 , y1832 , y1833 , y1834 , y1835 , y1836 , y1837 , y1838 , y1839 , y1840 , y1841 , y1842 , y1843 , y1844 , y1845 , y1846 , y1847 , y1848 , y1849 , y1850 , y1851 , y1852 , y1853 , y1854 , y1855 , y1856 , y1857 , y1858 , y1859 , y1860 , y1861 , y1862 , y1863 , y1864 , y1865 , y1866 , y1867 , y1868 , y1869 , y1870 , y1871 , y1872 , y1873 , y1874 , y1875 , y1876 , y1877 , y1878 , y1879 , y1880 , y1881 , y1882 , y1883 , y1884 , y1885 , y1886 , y1887 , y1888 , y1889 , y1890 , y1891 , y1892 , y1893 , y1894 , y1895 , y1896 , y1897 , y1898 , y1899 , y1900 , y1901 , y1902 , y1903 , y1904 , y1905 , y1906 , y1907 , y1908 , y1909 , y1910 , y1911 , y1912 , y1913 , y1914 , y1915 , y1916 , y1917 , y1918 , y1919 , y1920 , y1921 , y1922 , y1923 , y1924 , y1925 , y1926 , y1927 , y1928 , y1929 , y1930 , y1931 , y1932 , y1933 , y1934 , y1935 , y1936 , y1937 , y1938 , y1939 , y1940 , y1941 , y1942 , y1943 , y1944 , y1945 , y1946 , y1947 , y1948 , y1949 , y1950 , y1951 , y1952 , y1953 , y1954 , y1955 , y1956 , y1957 , y1958 , y1959 , y1960 , y1961 , y1962 , y1963 , y1964 , y1965 , y1966 , y1967 , y1968 , y1969 , y1970 , y1971 , y1972 , y1973 , y1974 , y1975 , y1976 , y1977 , y1978 , y1979 , y1980 , y1981 , y1982 , y1983 , y1984 , y1985 , y1986 , y1987 , y1988 , y1989 , y1990 , y1991 , y1992 , y1993 , y1994 , y1995 , y1996 , y1997 , y1998 , y1999 , y2000 , y2001 , y2002 , y2003 , y2004 , y2005 , y2006 , y2007 , y2008 , y2009 , y2010 , y2011 , y2012 , y2013 , y2014 , y2015 , y2016 , y2017 , y2018 , y2019 , y2020 , y2021 , y2022 , y2023 , y2024 , y2025 , y2026 , y2027 , y2028 , y2029 , y2030 , y2031 , y2032 , y2033 , y2034 , y2035 , y2036 , y2037 , y2038 , y2039 , y2040 , y2041 , y2042 , y2043 , y2044 , y2045 , y2046 , y2047 , y2048 , y2049 , y2050 , y2051 , y2052 , y2053 , y2054 , y2055 , y2056 , y2057 , y2058 , y2059 , y2060 , y2061 , y2062 , y2063 , y2064 , y2065 , y2066 , y2067 , y2068 , y2069 , y2070 , y2071 , y2072 , y2073 , y2074 , y2075 , y2076 , y2077 , y2078 , y2079 , y2080 , y2081 , y2082 , y2083 , y2084 , y2085 , y2086 , y2087 , y2088 , y2089 , y2090 , y2091 , y2092 , y2093 , y2094 , y2095 , y2096 , y2097 , y2098 , y2099 , y2100 , y2101 , y2102 , y2103 , y2104 , y2105 , y2106 , y2107 , y2108 , y2109 , y2110 , y2111 , y2112 , y2113 , y2114 , y2115 , y2116 , y2117 , y2118 , y2119 , y2120 , y2121 , y2122 , y2123 , y2124 , y2125 , y2126 , y2127 , y2128 , y2129 , y2130 , y2131 , y2132 , y2133 , y2134 , y2135 , y2136 , y2137 , y2138 , y2139 , y2140 , y2141 , y2142 , y2143 , y2144 , y2145 , y2146 , y2147 , y2148 , y2149 , y2150 , y2151 , y2152 , y2153 , y2154 , y2155 , y2156 , y2157 , y2158 , y2159 , y2160 , y2161 , y2162 , y2163 , y2164 , y2165 , y2166 , y2167 , y2168 , y2169 , y2170 , y2171 , y2172 , y2173 , y2174 , y2175 , y2176 , y2177 , y2178 , y2179 , y2180 , y2181 , y2182 , y2183 , y2184 , y2185 , y2186 , y2187 , y2188 , y2189 , y2190 , y2191 , y2192 , y2193 , y2194 , y2195 , y2196 , y2197 , y2198 , y2199 , y2200 , y2201 , y2202 , y2203 , y2204 , y2205 , y2206 , y2207 , y2208 , y2209 , y2210 , y2211 , y2212 , y2213 , y2214 , y2215 , y2216 , y2217 , y2218 , y2219 , y2220 , y2221 , y2222 , y2223 , y2224 , y2225 , y2226 , y2227 , y2228 , y2229 , y2230 , y2231 , y2232 , y2233 , y2234 , y2235 , y2236 , y2237 , y2238 , y2239 , y2240 , y2241 , y2242 , y2243 , y2244 , y2245 , y2246 , y2247 , y2248 , y2249 , y2250 , y2251 , y2252 , y2253 , y2254 , y2255 , y2256 , y2257 , y2258 , y2259 , y2260 , y2261 , y2262 , y2263 , y2264 , y2265 , y2266 , y2267 , y2268 , y2269 , y2270 , y2271 , y2272 , y2273 , y2274 , y2275 , y2276 , y2277 , y2278 , y2279 , y2280 , y2281 , y2282 , y2283 , y2284 , y2285 , y2286 , y2287 , y2288 , y2289 , y2290 , y2291 , y2292 , y2293 , y2294 , y2295 , y2296 , y2297 , y2298 , y2299 , y2300 , y2301 , y2302 , y2303 , y2304 , y2305 , y2306 , y2307 , y2308 , y2309 , y2310 , y2311 , y2312 , y2313 , y2314 , y2315 , y2316 , y2317 , y2318 , y2319 , y2320 , y2321 , y2322 , y2323 , y2324 , y2325 , y2326 , y2327 , y2328 , y2329 , y2330 , y2331 , y2332 , y2333 , y2334 , y2335 , y2336 , y2337 , y2338 , y2339 , y2340 , y2341 , y2342 , y2343 , y2344 , y2345 , y2346 , y2347 , y2348 , y2349 , y2350 , y2351 , y2352 , y2353 , y2354 , y2355 , y2356 , y2357 , y2358 , y2359 , y2360 , y2361 , y2362 , y2363 , y2364 , y2365 , y2366 , y2367 , y2368 , y2369 , y2370 , y2371 , y2372 , y2373 , y2374 , y2375 , y2376 , y2377 , y2378 , y2379 , y2380 , y2381 , y2382 , y2383 , y2384 , y2385 , y2386 , y2387 , y2388 , y2389 , y2390 , y2391 , y2392 , y2393 , y2394 , y2395 , y2396 , y2397 , y2398 , y2399 , y2400 , y2401 , y2402 , y2403 , y2404 , y2405 , y2406 , y2407 , y2408 , y2409 , y2410 , y2411 , y2412 , y2413 , y2414 , y2415 , y2416 , y2417 , y2418 , y2419 , y2420 , y2421 , y2422 , y2423 , y2424 , y2425 , y2426 , y2427 , y2428 , y2429 , y2430 , y2431 , y2432 , y2433 , y2434 , y2435 , y2436 , y2437 , y2438 , y2439 , y2440 , y2441 , y2442 , y2443 , y2444 , y2445 , y2446 , y2447 , y2448 , y2449 , y2450 , y2451 , y2452 , y2453 , y2454 , y2455 , y2456 , y2457 , y2458 , y2459 , y2460 , y2461 , y2462 , y2463 , y2464 , y2465 , y2466 , y2467 , y2468 , y2469 , y2470 , y2471 , y2472 , y2473 , y2474 , y2475 , y2476 , y2477 , y2478 , y2479 , y2480 , y2481 , y2482 , y2483 , y2484 , y2485 , y2486 , y2487 , y2488 , y2489 , y2490 , y2491 , y2492 , y2493 , y2494 , y2495 , y2496 , y2497 , y2498 , y2499 , y2500 , y2501 , y2502 , y2503 , y2504 , y2505 , y2506 , y2507 , y2508 , y2509 , y2510 , y2511 , y2512 , y2513 , y2514 , y2515 , y2516 , y2517 , y2518 , y2519 , y2520 , y2521 , y2522 , y2523 , y2524 , y2525 , y2526 , y2527 , y2528 , y2529 , y2530 , y2531 , y2532 , y2533 , y2534 , y2535 , y2536 , y2537 , y2538 , y2539 , y2540 , y2541 , y2542 , y2543 , y2544 , y2545 , y2546 , y2547 , y2548 , y2549 , y2550 , y2551 , y2552 , y2553 , y2554 , y2555 , y2556 , y2557 , y2558 , y2559 , y2560 , y2561 , y2562 , y2563 , y2564 , y2565 , y2566 , y2567 , y2568 , y2569 , y2570 , y2571 , y2572 , y2573 , y2574 , y2575 , y2576 , y2577 , y2578 , y2579 , y2580 , y2581 , y2582 , y2583 , y2584 , y2585 , y2586 , y2587 , y2588 , y2589 , y2590 , y2591 , y2592 , y2593 , y2594 , y2595 , y2596 , y2597 , y2598 , y2599 , y2600 , y2601 , y2602 , y2603 , y2604 , y2605 , y2606 , y2607 , y2608 , y2609 , y2610 , y2611 , y2612 , y2613 , y2614 , y2615 , y2616 , y2617 , y2618 , y2619 , y2620 , y2621 , y2622 , y2623 , y2624 , y2625 , y2626 , y2627 , y2628 , y2629 , y2630 , y2631 , y2632 , y2633 , y2634 , y2635 , y2636 , y2637 , y2638 , y2639 , y2640 , y2641 , y2642 , y2643 , y2644 , y2645 , y2646 , y2647 , y2648 , y2649 , y2650 , y2651 , y2652 , y2653 , y2654 , y2655 , y2656 , y2657 , y2658 , y2659 , y2660 , y2661 , y2662 , y2663 , y2664 , y2665 , y2666 , y2667 , y2668 , y2669 , y2670 , y2671 , y2672 , y2673 , y2674 , y2675 , y2676 , y2677 , y2678 , y2679 , y2680 , y2681 , y2682 , y2683 , y2684 , y2685 , y2686 , y2687 , y2688 , y2689 , y2690 , y2691 , y2692 , y2693 , y2694 , y2695 , y2696 , y2697 , y2698 , y2699 , y2700 , y2701 , y2702 , y2703 , y2704 , y2705 , y2706 , y2707 , y2708 , y2709 , y2710 , y2711 , y2712 , y2713 , y2714 , y2715 , y2716 , y2717 , y2718 , y2719 , y2720 , y2721 , y2722 , y2723 , y2724 , y2725 , y2726 , y2727 , y2728 , y2729 , y2730 , y2731 , y2732 , y2733 , y2734 , y2735 , y2736 , y2737 , y2738 , y2739 , y2740 , y2741 , y2742 , y2743 , y2744 , y2745 , y2746 , y2747 , y2748 , y2749 , y2750 , y2751 , y2752 , y2753 , y2754 , y2755 , y2756 , y2757 , y2758 , y2759 , y2760 , y2761 , y2762 , y2763 , y2764 , y2765 , y2766 , y2767 , y2768 , y2769 , y2770 , y2771 , y2772 , y2773 , y2774 , y2775 , y2776 , y2777 , y2778 , y2779 , y2780 , y2781 , y2782 , y2783 , y2784 , y2785 , y2786 , y2787 , y2788 , y2789 , y2790 , y2791 , y2792 , y2793 , y2794 , y2795 , y2796 , y2797 , y2798 , y2799 , y2800 , y2801 , y2802 , y2803 , y2804 , y2805 , y2806 , y2807 , y2808 , y2809 , y2810 , y2811 , y2812 , y2813 , y2814 , y2815 , y2816 , y2817 , y2818 , y2819 , y2820 , y2821 , y2822 , y2823 , y2824 , y2825 , y2826 , y2827 , y2828 , y2829 , y2830 , y2831 , y2832 , y2833 , y2834 , y2835 , y2836 , y2837 , y2838 , y2839 , y2840 , y2841 , y2842 , y2843 , y2844 , y2845 , y2846 , y2847 , y2848 , y2849 , y2850 , y2851 , y2852 , y2853 , y2854 , y2855 , y2856 , y2857 , y2858 , y2859 , y2860 , y2861 , y2862 , y2863 , y2864 , y2865 , y2866 , y2867 , y2868 , y2869 , y2870 , y2871 , y2872 , y2873 , y2874 , y2875 , y2876 , y2877 , y2878 , y2879 , y2880 , y2881 , y2882 , y2883 , y2884 , y2885 , y2886 , y2887 , y2888 , y2889 , y2890 , y2891 , y2892 , y2893 , y2894 , y2895 , y2896 , y2897 , y2898 , y2899 , y2900 , y2901 , y2902 , y2903 , y2904 , y2905 , y2906 , y2907 , y2908 , y2909 , y2910 , y2911 , y2912 , y2913 , y2914 , y2915 , y2916 , y2917 , y2918 , y2919 , y2920 , y2921 , y2922 , y2923 , y2924 , y2925 , y2926 , y2927 , y2928 , y2929 , y2930 , y2931 , y2932 , y2933 , y2934 , y2935 , y2936 , y2937 , y2938 , y2939 , y2940 , y2941 , y2942 , y2943 , y2944 , y2945 , y2946 , y2947 , y2948 , y2949 , y2950 , y2951 , y2952 , y2953 , y2954 , y2955 , y2956 , y2957 , y2958 , y2959 , y2960 , y2961 , y2962 , y2963 , y2964 , y2965 , y2966 , y2967 , y2968 , y2969 , y2970 , y2971 , y2972 , y2973 , y2974 , y2975 , y2976 , y2977 , y2978 , y2979 , y2980 , y2981 , y2982 , y2983 , y2984 , y2985 , y2986 , y2987 , y2988 , y2989 , y2990 , y2991 , y2992 , y2993 , y2994 , y2995 , y2996 , y2997 , y2998 , y2999 , y3000 , y3001 , y3002 , y3003 , y3004 , y3005 , y3006 , y3007 , y3008 , y3009 , y3010 , y3011 , y3012 , y3013 , y3014 , y3015 , y3016 , y3017 , y3018 , y3019 , y3020 , y3021 , y3022 , y3023 , y3024 , y3025 , y3026 , y3027 , y3028 , y3029 , y3030 , y3031 , y3032 , y3033 , y3034 , y3035 , y3036 , y3037 , y3038 , y3039 , y3040 , y3041 , y3042 , y3043 , y3044 , y3045 , y3046 , y3047 , y3048 , y3049 , y3050 , y3051 , y3052 , y3053 , y3054 , y3055 , y3056 , y3057 , y3058 , y3059 , y3060 , y3061 , y3062 , y3063 , y3064 , y3065 , y3066 , y3067 , y3068 , y3069 , y3070 , y3071 , y3072 , y3073 , y3074 , y3075 , y3076 , y3077 , y3078 , y3079 , y3080 , y3081 , y3082 , y3083 , y3084 , y3085 , y3086 , y3087 , y3088 , y3089 , y3090 , y3091 , y3092 , y3093 , y3094 , y3095 , y3096 , y3097 , y3098 , y3099 , y3100 , y3101 , y3102 , y3103 , y3104 , y3105 , y3106 , y3107 , y3108 , y3109 , y3110 , y3111 , y3112 , y3113 , y3114 , y3115 , y3116 , y3117 , y3118 , y3119 , y3120 , y3121 , y3122 , y3123 , y3124 , y3125 , y3126 , y3127 , y3128 , y3129 , y3130 , y3131 , y3132 , y3133 , y3134 , y3135 , y3136 , y3137 , y3138 , y3139 , y3140 , y3141 , y3142 , y3143 , y3144 , y3145 , y3146 , y3147 , y3148 , y3149 , y3150 , y3151 , y3152 , y3153 , y3154 , y3155 , y3156 , y3157 , y3158 , y3159 , y3160 , y3161 , y3162 , y3163 , y3164 , y3165 , y3166 , y3167 , y3168 , y3169 , y3170 , y3171 , y3172 , y3173 , y3174 , y3175 , y3176 , y3177 , y3178 , y3179 , y3180 , y3181 , y3182 , y3183 , y3184 , y3185 , y3186 , y3187 , y3188 , y3189 , y3190 , y3191 , y3192 , y3193 , y3194 , y3195 , y3196 , y3197 , y3198 , y3199 , y3200 , y3201 , y3202 , y3203 , y3204 , y3205 , y3206 , y3207 , y3208 , y3209 , y3210 , y3211 , y3212 , y3213 , y3214 , y3215 , y3216 , y3217 , y3218 , y3219 , y3220 , y3221 , y3222 , y3223 , y3224 , y3225 , y3226 , y3227 , y3228 , y3229 , y3230 , y3231 , y3232 , y3233 , y3234 , y3235 , y3236 , y3237 , y3238 , y3239 , y3240 , y3241 , y3242 , y3243 , y3244 , y3245 , y3246 , y3247 , y3248 , y3249 , y3250 , y3251 , y3252 , y3253 , y3254 , y3255 , y3256 , y3257 , y3258 , y3259 , y3260 , y3261 , y3262 , y3263 , y3264 , y3265 , y3266 , y3267 , y3268 , y3269 , y3270 , y3271 , y3272 , y3273 , y3274 , y3275 , y3276 , y3277 , y3278 , y3279 , y3280 , y3281 , y3282 , y3283 , y3284 , y3285 , y3286 , y3287 , y3288 , y3289 , y3290 , y3291 , y3292 , y3293 , y3294 , y3295 , y3296 , y3297 , y3298 , y3299 , y3300 , y3301 , y3302 , y3303 , y3304 , y3305 , y3306 , y3307 , y3308 , y3309 , y3310 , y3311 , y3312 , y3313 , y3314 , y3315 , y3316 , y3317 , y3318 , y3319 , y3320 , y3321 , y3322 , y3323 , y3324 , y3325 , y3326 , y3327 , y3328 , y3329 , y3330 , y3331 , y3332 , y3333 , y3334 , y3335 , y3336 , y3337 , y3338 , y3339 , y3340 , y3341 , y3342 , y3343 , y3344 , y3345 , y3346 , y3347 , y3348 , y3349 , y3350 , y3351 , y3352 , y3353 , y3354 , y3355 , y3356 , y3357 , y3358 , y3359 , y3360 , y3361 , y3362 , y3363 , y3364 , y3365 , y3366 , y3367 , y3368 , y3369 , y3370 , y3371 , y3372 , y3373 , y3374 , y3375 , y3376 , y3377 , y3378 , y3379 , y3380 , y3381 , y3382 , y3383 , y3384 , y3385 , y3386 , y3387 , y3388 , y3389 , y3390 , y3391 , y3392 , y3393 , y3394 , y3395 , y3396 , y3397 , y3398 , y3399 , y3400 , y3401 , y3402 , y3403 , y3404 , y3405 , y3406 , y3407 , y3408 , y3409 , y3410 , y3411 , y3412 , y3413 , y3414 , y3415 , y3416 , y3417 , y3418 , y3419 , y3420 , y3421 , y3422 , y3423 , y3424 , y3425 , y3426 , y3427 , y3428 , y3429 , y3430 , y3431 , y3432 , y3433 , y3434 , y3435 , y3436 , y3437 , y3438 , y3439 , y3440 , y3441 , y3442 , y3443 , y3444 , y3445 , y3446 , y3447 , y3448 , y3449 , y3450 , y3451 , y3452 , y3453 , y3454 , y3455 , y3456 , y3457 , y3458 , y3459 , y3460 , y3461 , y3462 , y3463 , y3464 , y3465 , y3466 , y3467 , y3468 , y3469 , y3470 , y3471 , y3472 , y3473 , y3474 , y3475 , y3476 , y3477 , y3478 , y3479 , y3480 , y3481 , y3482 , y3483 , y3484 , y3485 , y3486 , y3487 , y3488 , y3489 , y3490 , y3491 , y3492 , y3493 , y3494 , y3495 , y3496 , y3497 , y3498 , y3499 , y3500 , y3501 , y3502 , y3503 , y3504 , y3505 , y3506 , y3507 , y3508 , y3509 , y3510 , y3511 , y3512 , y3513 , y3514 , y3515 , y3516 , y3517 , y3518 , y3519 , y3520 , y3521 , y3522 , y3523 , y3524 , y3525 , y3526 , y3527 , y3528 , y3529 , y3530 , y3531 , y3532 , y3533 , y3534 , y3535 , y3536 , y3537 , y3538 , y3539 , y3540 , y3541 , y3542 , y3543 , y3544 , y3545 , y3546 , y3547 , y3548 , y3549 , y3550 , y3551 , y3552 , y3553 , y3554 , y3555 , y3556 , y3557 , y3558 , y3559 , y3560 , y3561 , y3562 , y3563 , y3564 , y3565 , y3566 , y3567 , y3568 , y3569 , y3570 , y3571 , y3572 , y3573 , y3574 , y3575 , y3576 , y3577 , y3578 , y3579 , y3580 , y3581 , y3582 , y3583 , y3584 , y3585 , y3586 , y3587 , y3588 , y3589 , y3590 , y3591 , y3592 , y3593 , y3594 , y3595 , y3596 , y3597 , y3598 , y3599 , y3600 , y3601 , y3602 , y3603 , y3604 , y3605 , y3606 , y3607 , y3608 , y3609 , y3610 , y3611 , y3612 , y3613 , y3614 , y3615 , y3616 , y3617 , y3618 , y3619 , y3620 , y3621 , y3622 , y3623 , y3624 , y3625 , y3626 , y3627 , y3628 , y3629 , y3630 , y3631 , y3632 , y3633 , y3634 , y3635 , y3636 , y3637 , y3638 , y3639 , y3640 , y3641 , y3642 , y3643 , y3644 , y3645 , y3646 , y3647 , y3648 , y3649 , y3650 , y3651 , y3652 , y3653 , y3654 , y3655 , y3656 , y3657 , y3658 , y3659 , y3660 , y3661 , y3662 , y3663 , y3664 , y3665 , y3666 , y3667 , y3668 , y3669 , y3670 , y3671 , y3672 , y3673 , y3674 , y3675 , y3676 , y3677 , y3678 , y3679 , y3680 , y3681 , y3682 , y3683 , y3684 , y3685 , y3686 , y3687 , y3688 , y3689 , y3690 , y3691 , y3692 , y3693 , y3694 , y3695 , y3696 , y3697 , y3698 , y3699 , y3700 , y3701 , y3702 , y3703 , y3704 , y3705 , y3706 , y3707 , y3708 , y3709 , y3710 , y3711 , y3712 , y3713 , y3714 , y3715 , y3716 , y3717 , y3718 , y3719 , y3720 , y3721 , y3722 , y3723 , y3724 , y3725 , y3726 , y3727 , y3728 , y3729 , y3730 , y3731 , y3732 , y3733 , y3734 , y3735 , y3736 , y3737 , y3738 , y3739 , y3740 , y3741 , y3742 , y3743 , y3744 , y3745 , y3746 , y3747 , y3748 , y3749 , y3750 , y3751 , y3752 , y3753 , y3754 , y3755 , y3756 , y3757 , y3758 , y3759 , y3760 , y3761 , y3762 , y3763 , y3764 , y3765 , y3766 , y3767 , y3768 , y3769 , y3770 , y3771 , y3772 , y3773 , y3774 , y3775 , y3776 , y3777 , y3778 , y3779 , y3780 , y3781 , y3782 , y3783 , y3784 , y3785 , y3786 , y3787 , y3788 , y3789 , y3790 , y3791 , y3792 , y3793 , y3794 , y3795 , y3796 , y3797 , y3798 , y3799 , y3800 , y3801 , y3802 , y3803 , y3804 , y3805 , y3806 , y3807 , y3808 , y3809 , y3810 , y3811 , y3812 , y3813 , y3814 , y3815 , y3816 , y3817 , y3818 , y3819 , y3820 , y3821 , y3822 , y3823 , y3824 , y3825 , y3826 , y3827 , y3828 , y3829 , y3830 , y3831 , y3832 , y3833 , y3834 , y3835 , y3836 , y3837 , y3838 , y3839 , y3840 , y3841 , y3842 , y3843 , y3844 , y3845 , y3846 , y3847 , y3848 , y3849 , y3850 , y3851 , y3852 , y3853 , y3854 , y3855 , y3856 , y3857 , y3858 , y3859 , y3860 , y3861 , y3862 , y3863 , y3864 , y3865 , y3866 , y3867 , y3868 , y3869 , y3870 , y3871 , y3872 , y3873 , y3874 , y3875 , y3876 , y3877 , y3878 , y3879 , y3880 , y3881 , y3882 , y3883 , y3884 , y3885 , y3886 , y3887 , y3888 , y3889 , y3890 , y3891 , y3892 , y3893 , y3894 , y3895 , y3896 , y3897 , y3898 , y3899 , y3900 , y3901 , y3902 , y3903 , y3904 , y3905 , y3906 , y3907 , y3908 , y3909 , y3910 , y3911 , y3912 , y3913 , y3914 , y3915 , y3916 , y3917 , y3918 , y3919 , y3920 , y3921 , y3922 , y3923 , y3924 , y3925 , y3926 , y3927 , y3928 , y3929 , y3930 , y3931 , y3932 , y3933 , y3934 , y3935 , y3936 , y3937 , y3938 , y3939 , y3940 , y3941 , y3942 , y3943 , y3944 , y3945 , y3946 , y3947 , y3948 , y3949 , y3950 , y3951 , y3952 , y3953 , y3954 , y3955 , y3956 , y3957 , y3958 , y3959 , y3960 , y3961 , y3962 , y3963 , y3964 , y3965 , y3966 , y3967 , y3968 , y3969 , y3970 , y3971 , y3972 , y3973 , y3974 , y3975 , y3976 , y3977 , y3978 , y3979 , y3980 , y3981 , y3982 , y3983 , y3984 , y3985 , y3986 , y3987 , y3988 , y3989 , y3990 , y3991 , y3992 , y3993 , y3994 , y3995 , y3996 , y3997 , y3998 , y3999 , y4000 , y4001 , y4002 , y4003 , y4004 , y4005 , y4006 , y4007 , y4008 , y4009 , y4010 , y4011 , y4012 , y4013 , y4014 , y4015 , y4016 , y4017 , y4018 , y4019 , y4020 , y4021 , y4022 , y4023 , y4024 , y4025 , y4026 , y4027 , y4028 , y4029 , y4030 , y4031 , y4032 , y4033 , y4034 , y4035 , y4036 , y4037 , y4038 , y4039 , y4040 , y4041 , y4042 , y4043 , y4044 , y4045 , y4046 , y4047 , y4048 , y4049 , y4050 , y4051 , y4052 , y4053 , y4054 , y4055 , y4056 , y4057 , y4058 , y4059 , y4060 , y4061 , y4062 , y4063 , y4064 , y4065 , y4066 , y4067 , y4068 , y4069 , y4070 , y4071 , y4072 , y4073 , y4074 , y4075 , y4076 , y4077 , y4078 , y4079 , y4080 , y4081 , y4082 , y4083 , y4084 , y4085 , y4086 , y4087 , y4088 , y4089 , y4090 , y4091 , y4092 , y4093 , y4094 , y4095 , y4096 , y4097 , y4098 , y4099 , y4100 , y4101 , y4102 , y4103 , y4104 , y4105 , y4106 , y4107 , y4108 , y4109 , y4110 , y4111 , y4112 , y4113 , y4114 , y4115 , y4116 , y4117 , y4118 , y4119 , y4120 , y4121 , y4122 , y4123 , y4124 , y4125 , y4126 , y4127 , y4128 , y4129 , y4130 , y4131 , y4132 , y4133 , y4134 , y4135 , y4136 , y4137 , y4138 , y4139 , y4140 , y4141 , y4142 , y4143 , y4144 , y4145 , y4146 , y4147 , y4148 , y4149 , y4150 , y4151 , y4152 , y4153 , y4154 , y4155 , y4156 , y4157 , y4158 , y4159 , y4160 , y4161 , y4162 , y4163 , y4164 , y4165 , y4166 , y4167 , y4168 , y4169 , y4170 , y4171 , y4172 , y4173 , y4174 , y4175 , y4176 , y4177 , y4178 , y4179 , y4180 , y4181 , y4182 , y4183 , y4184 , y4185 , y4186 , y4187 , y4188 , y4189 , y4190 , y4191 , y4192 , y4193 , y4194 , y4195 , y4196 , y4197 , y4198 , y4199 , y4200 , y4201 , y4202 , y4203 , y4204 , y4205 , y4206 , y4207 , y4208 , y4209 , y4210 , y4211 , y4212 , y4213 , y4214 , y4215 , y4216 , y4217 , y4218 , y4219 , y4220 , y4221 , y4222 , y4223 , y4224 , y4225 , y4226 , y4227 , y4228 , y4229 , y4230 , y4231 , y4232 , y4233 , y4234 , y4235 , y4236 , y4237 , y4238 , y4239 , y4240 , y4241 , y4242 , y4243 , y4244 , y4245 , y4246 , y4247 , y4248 , y4249 , y4250 , y4251 , y4252 , y4253 , y4254 , y4255 , y4256 , y4257 , y4258 , y4259 , y4260 , y4261 , y4262 , y4263 , y4264 , y4265 , y4266 , y4267 , y4268 , y4269 , y4270 , y4271 , y4272 , y4273 , y4274 , y4275 , y4276 , y4277 , y4278 , y4279 , y4280 , y4281 , y4282 , y4283 , y4284 , y4285 , y4286 , y4287 , y4288 , y4289 , y4290 , y4291 , y4292 , y4293 , y4294 , y4295 , y4296 , y4297 , y4298 , y4299 , y4300 , y4301 , y4302 , y4303 , y4304 , y4305 , y4306 , y4307 , y4308 , y4309 , y4310 , y4311 , y4312 , y4313 , y4314 , y4315 , y4316 , y4317 , y4318 , y4319 , y4320 , y4321 , y4322 , y4323 , y4324 , y4325 , y4326 , y4327 , y4328 , y4329 , y4330 , y4331 , y4332 , y4333 , y4334 , y4335 , y4336 , y4337 , y4338 , y4339 , y4340 , y4341 , y4342 , y4343 , y4344 , y4345 , y4346 , y4347 , y4348 , y4349 , y4350 , y4351 , y4352 , y4353 , y4354 , y4355 , y4356 , y4357 , y4358 , y4359 , y4360 , y4361 , y4362 , y4363 , y4364 , y4365 , y4366 , y4367 , y4368 , y4369 , y4370 , y4371 , y4372 , y4373 , y4374 , y4375 , y4376 , y4377 , y4378 , y4379 , y4380 , y4381 , y4382 , y4383 , y4384 , y4385 , y4386 , y4387 , y4388 , y4389 , y4390 , y4391 , y4392 , y4393 , y4394 , y4395 , y4396 , y4397 , y4398 , y4399 , y4400 , y4401 , y4402 , y4403 , y4404 , y4405 , y4406 , y4407 , y4408 , y4409 , y4410 , y4411 , y4412 , y4413 , y4414 , y4415 , y4416 , y4417 , y4418 , y4419 , y4420 , y4421 , y4422 , y4423 , y4424 , y4425 , y4426 , y4427 , y4428 , y4429 , y4430 , y4431 , y4432 , y4433 , y4434 , y4435 , y4436 , y4437 , y4438 , y4439 , y4440 , y4441 , y4442 , y4443 , y4444 , y4445 , y4446 , y4447 , y4448 , y4449 , y4450 , y4451 , y4452 , y4453 , y4454 , y4455 , y4456 , y4457 , y4458 , y4459 , y4460 , y4461 , y4462 , y4463 , y4464 , y4465 , y4466 , y4467 , y4468 , y4469 , y4470 , y4471 , y4472 , y4473 , y4474 , y4475 , y4476 , y4477 , y4478 , y4479 , y4480 , y4481 , y4482 , y4483 , y4484 , y4485 , y4486 , y4487 , y4488 , y4489 , y4490 , y4491 , y4492 , y4493 , y4494 , y4495 , y4496 , y4497 , y4498 , y4499 , y4500 , y4501 , y4502 , y4503 , y4504 , y4505 , y4506 , y4507 , y4508 , y4509 , y4510 , y4511 , y4512 , y4513 , y4514 , y4515 , y4516 , y4517 , y4518 , y4519 , y4520 , y4521 , y4522 , y4523 , y4524 , y4525 , y4526 , y4527 , y4528 , y4529 , y4530 , y4531 , y4532 , y4533 , y4534 , y4535 , y4536 , y4537 , y4538 , y4539 , y4540 , y4541 , y4542 , y4543 , y4544 , y4545 , y4546 , y4547 , y4548 , y4549 , y4550 , y4551 , y4552 , y4553 , y4554 , y4555 , y4556 , y4557 , y4558 , y4559 , y4560 , y4561 , y4562 , y4563 , y4564 , y4565 , y4566 , y4567 , y4568 , y4569 , y4570 , y4571 , y4572 , y4573 , y4574 , y4575 , y4576 , y4577 , y4578 , y4579 , y4580 , y4581 , y4582 , y4583 , y4584 , y4585 , y4586 , y4587 , y4588 , y4589 , y4590 , y4591 , y4592 , y4593 , y4594 , y4595 , y4596 , y4597 , y4598 , y4599 , y4600 , y4601 , y4602 , y4603 , y4604 , y4605 , y4606 , y4607 , y4608 , y4609 , y4610 , y4611 , y4612 , y4613 , y4614 , y4615 , y4616 , y4617 , y4618 , y4619 , y4620 , y4621 , y4622 , y4623 , y4624 , y4625 , y4626 , y4627 , y4628 , y4629 , y4630 , y4631 , y4632 , y4633 , y4634 , y4635 , y4636 , y4637 , y4638 , y4639 , y4640 , y4641 , y4642 , y4643 , y4644 , y4645 , y4646 , y4647 , y4648 , y4649 , y4650 , y4651 , y4652 , y4653 , y4654 , y4655 , y4656 , y4657 , y4658 , y4659 , y4660 , y4661 , y4662 , y4663 , y4664 , y4665 , y4666 , y4667 , y4668 , y4669 , y4670 , y4671 , y4672 , y4673 , y4674 , y4675 , y4676 , y4677 , y4678 , y4679 , y4680 , y4681 , y4682 , y4683 , y4684 , y4685 , y4686 , y4687 , y4688 , y4689 , y4690 , y4691 , y4692 , y4693 , y4694 , y4695 , y4696 , y4697 , y4698 , y4699 , y4700 , y4701 , y4702 , y4703 , y4704 , y4705 , y4706 , y4707 , y4708 , y4709 , y4710 , y4711 , y4712 , y4713 , y4714 , y4715 , y4716 , y4717 , y4718 , y4719 , y4720 , y4721 , y4722 , y4723 , y4724 , y4725 , y4726 , y4727 , y4728 , y4729 , y4730 , y4731 , y4732 , y4733 , y4734 , y4735 , y4736 , y4737 , y4738 , y4739 , y4740 , y4741 , y4742 , y4743 , y4744 , y4745 , y4746 , y4747 , y4748 , y4749 , y4750 , y4751 , y4752 , y4753 , y4754 , y4755 , y4756 , y4757 , y4758 , y4759 , y4760 , y4761 , y4762 , y4763 , y4764 , y4765 , y4766 , y4767 , y4768 , y4769 , y4770 , y4771 , y4772 , y4773 , y4774 , y4775 , y4776 , y4777 , y4778 , y4779 , y4780 , y4781 , y4782 , y4783 , y4784 , y4785 , y4786 , y4787 , y4788 , y4789 , y4790 , y4791 , y4792 , y4793 , y4794 , y4795 , y4796 , y4797 , y4798 , y4799 , y4800 , y4801 , y4802 , y4803 , y4804 , y4805 , y4806 , y4807 , y4808 , y4809 , y4810 , y4811 , y4812 , y4813 , y4814 , y4815 , y4816 , y4817 , y4818 , y4819 , y4820 , y4821 , y4822 , y4823 , y4824 , y4825 , y4826 , y4827 , y4828 , y4829 , y4830 , y4831 , y4832 , y4833 , y4834 , y4835 , y4836 , y4837 , y4838 , y4839 , y4840 , y4841 , y4842 , y4843 , y4844 , y4845 , y4846 , y4847 , y4848 , y4849 , y4850 , y4851 , y4852 , y4853 , y4854 , y4855 , y4856 , y4857 , y4858 , y4859 , y4860 , y4861 , y4862 , y4863 , y4864 , y4865 , y4866 , y4867 , y4868 , y4869 , y4870 , y4871 , y4872 , y4873 , y4874 , y4875 , y4876 , y4877 , y4878 , y4879 , y4880 , y4881 , y4882 , y4883 , y4884 , y4885 , y4886 , y4887 , y4888 , y4889 , y4890 , y4891 , y4892 , y4893 , y4894 , y4895 , y4896 , y4897 , y4898 , y4899 , y4900 , y4901 , y4902 , y4903 , y4904 , y4905 , y4906 , y4907 , y4908 , y4909 , y4910 , y4911 , y4912 , y4913 , y4914 , y4915 , y4916 , y4917 , y4918 , y4919 , y4920 , y4921 , y4922 , y4923 , y4924 , y4925 , y4926 , y4927 , y4928 , y4929 , y4930 , y4931 , y4932 , y4933 , y4934 , y4935 , y4936 , y4937 , y4938 , y4939 , y4940 , y4941 , y4942 , y4943 , y4944 , y4945 , y4946 , y4947 , y4948 , y4949 , y4950 , y4951 , y4952 , y4953 , y4954 , y4955 , y4956 , y4957 , y4958 , y4959 , y4960 , y4961 , y4962 , y4963 , y4964 , y4965 , y4966 , y4967 , y4968 , y4969 , y4970 , y4971 , y4972 , y4973 , y4974 , y4975 , y4976 , y4977 , y4978 , y4979 , y4980 , y4981 , y4982 , y4983 , y4984 , y4985 , y4986 , y4987 , y4988 , y4989 , y4990 , y4991 , y4992 , y4993 , y4994 , y4995 , y4996 , y4997 , y4998 , y4999 , y5000 , y5001 , y5002 , y5003 , y5004 , y5005 , y5006 , y5007 , y5008 , y5009 , y5010 , y5011 , y5012 , y5013 , y5014 , y5015 , y5016 , y5017 , y5018 , y5019 , y5020 , y5021 , y5022 , y5023 , y5024 , y5025 , y5026 , y5027 , y5028 , y5029 , y5030 , y5031 , y5032 , y5033 , y5034 , y5035 , y5036 , y5037 , y5038 , y5039 , y5040 , y5041 , y5042 , y5043 , y5044 , y5045 , y5046 , y5047 , y5048 , y5049 , y5050 , y5051 , y5052 , y5053 , y5054 , y5055 , y5056 , y5057 , y5058 , y5059 , y5060 , y5061 , y5062 , y5063 , y5064 , y5065 , y5066 , y5067 , y5068 , y5069 , y5070 , y5071 , y5072 , y5073 , y5074 , y5075 , y5076 , y5077 , y5078 , y5079 , y5080 , y5081 , y5082 , y5083 , y5084 , y5085 , y5086 , y5087 , y5088 , y5089 , y5090 , y5091 , y5092 , y5093 , y5094 , y5095 , y5096 , y5097 , y5098 , y5099 , y5100 , y5101 , y5102 , y5103 , y5104 , y5105 , y5106 , y5107 , y5108 , y5109 , y5110 , y5111 , y5112 , y5113 , y5114 , y5115 , y5116 , y5117 , y5118 , y5119 , y5120 , y5121 , y5122 , y5123 , y5124 , y5125 , y5126 , y5127 , y5128 , y5129 , y5130 , y5131 , y5132 , y5133 , y5134 , y5135 , y5136 , y5137 , y5138 , y5139 , y5140 , y5141 , y5142 , y5143 , y5144 , y5145 , y5146 , y5147 , y5148 , y5149 , y5150 , y5151 , y5152 , y5153 , y5154 , y5155 , y5156 , y5157 , y5158 , y5159 , y5160 , y5161 , y5162 , y5163 , y5164 , y5165 , y5166 , y5167 , y5168 , y5169 , y5170 , y5171 , y5172 , y5173 , y5174 , y5175 , y5176 , y5177 , y5178 , y5179 , y5180 , y5181 , y5182 , y5183 , y5184 , y5185 , y5186 , y5187 , y5188 , y5189 , y5190 , y5191 , y5192 , y5193 , y5194 , y5195 , y5196 , y5197 , y5198 , y5199 , y5200 , y5201 , y5202 , y5203 , y5204 , y5205 , y5206 , y5207 , y5208 , y5209 , y5210 , y5211 , y5212 , y5213 , y5214 , y5215 , y5216 , y5217 , y5218 , y5219 , y5220 , y5221 , y5222 , y5223 , y5224 , y5225 , y5226 , y5227 , y5228 , y5229 , y5230 , y5231 , y5232 , y5233 , y5234 , y5235 , y5236 , y5237 , y5238 , y5239 , y5240 , y5241 , y5242 , y5243 , y5244 , y5245 , y5246 , y5247 , y5248 , y5249 , y5250 , y5251 , y5252 , y5253 , y5254 , y5255 , y5256 , y5257 , y5258 , y5259 , y5260 , y5261 , y5262 , y5263 , y5264 , y5265 , y5266 , y5267 , y5268 , y5269 , y5270 , y5271 , y5272 , y5273 , y5274 , y5275 , y5276 , y5277 , y5278 , y5279 , y5280 , y5281 , y5282 , y5283 , y5284 , y5285 , y5286 , y5287 , y5288 , y5289 , y5290 , y5291 , y5292 , y5293 , y5294 , y5295 , y5296 , y5297 , y5298 , y5299 , y5300 , y5301 , y5302 , y5303 , y5304 , y5305 , y5306 , y5307 , y5308 , y5309 , y5310 , y5311 , y5312 , y5313 , y5314 , y5315 , y5316 , y5317 , y5318 , y5319 , y5320 , y5321 , y5322 , y5323 , y5324 , y5325 , y5326 , y5327 , y5328 , y5329 , y5330 , y5331 , y5332 , y5333 , y5334 , y5335 , y5336 , y5337 , y5338 , y5339 , y5340 , y5341 , y5342 , y5343 , y5344 , y5345 , y5346 , y5347 , y5348 , y5349 , y5350 , y5351 , y5352 , y5353 , y5354 , y5355 , y5356 , y5357 , y5358 , y5359 , y5360 , y5361 , y5362 , y5363 , y5364 , y5365 , y5366 , y5367 , y5368 , y5369 , y5370 , y5371 , y5372 , y5373 , y5374 , y5375 , y5376 , y5377 , y5378 , y5379 , y5380 , y5381 , y5382 , y5383 , y5384 , y5385 , y5386 , y5387 , y5388 , y5389 , y5390 , y5391 , y5392 , y5393 , y5394 , y5395 , y5396 , y5397 , y5398 , y5399 , y5400 , y5401 , y5402 , y5403 , y5404 , y5405 , y5406 , y5407 , y5408 , y5409 , y5410 , y5411 , y5412 , y5413 , y5414 , y5415 , y5416 , y5417 , y5418 , y5419 , y5420 , y5421 , y5422 , y5423 , y5424 , y5425 , y5426 , y5427 , y5428 , y5429 , y5430 , y5431 , y5432 , y5433 , y5434 , y5435 , y5436 , y5437 , y5438 , y5439 , y5440 , y5441 , y5442 , y5443 , y5444 , y5445 , y5446 , y5447 , y5448 , y5449 , y5450 , y5451 , y5452 , y5453 , y5454 , y5455 , y5456 , y5457 , y5458 , y5459 , y5460 , y5461 , y5462 , y5463 , y5464 , y5465 , y5466 , y5467 , y5468 , y5469 , y5470 , y5471 , y5472 , y5473 , y5474 , y5475 , y5476 , y5477 , y5478 , y5479 , y5480 , y5481 , y5482 , y5483 , y5484 , y5485 , y5486 , y5487 , y5488 , y5489 , y5490 , y5491 , y5492 , y5493 , y5494 , y5495 , y5496 , y5497 , y5498 , y5499 , y5500 , y5501 , y5502 , y5503 , y5504 , y5505 , y5506 , y5507 , y5508 , y5509 , y5510 , y5511 , y5512 , y5513 , y5514 , y5515 , y5516 , y5517 , y5518 , y5519 , y5520 , y5521 , y5522 , y5523 , y5524 , y5525 , y5526 , y5527 , y5528 , y5529 , y5530 , y5531 , y5532 , y5533 , y5534 , y5535 , y5536 , y5537 , y5538 , y5539 , y5540 , y5541 , y5542 , y5543 , y5544 , y5545 , y5546 , y5547 , y5548 , y5549 , y5550 , y5551 , y5552 , y5553 , y5554 , y5555 , y5556 , y5557 , y5558 , y5559 , y5560 , y5561 , y5562 , y5563 , y5564 , y5565 , y5566 , y5567 , y5568 , y5569 , y5570 , y5571 , y5572 , y5573 , y5574 , y5575 , y5576 , y5577 , y5578 , y5579 , y5580 , y5581 , y5582 , y5583 , y5584 , y5585 , y5586 , y5587 , y5588 , y5589 , y5590 , y5591 , y5592 , y5593 , y5594 , y5595 , y5596 , y5597 , y5598 , y5599 , y5600 , y5601 , y5602 , y5603 , y5604 , y5605 , y5606 , y5607 , y5608 , y5609 , y5610 , y5611 , y5612 , y5613 , y5614 , y5615 , y5616 , y5617 , y5618 , y5619 , y5620 , y5621 , y5622 , y5623 , y5624 , y5625 , y5626 , y5627 , y5628 , y5629 , y5630 , y5631 , y5632 , y5633 , y5634 , y5635 , y5636 , y5637 , y5638 , y5639 , y5640 , y5641 , y5642 , y5643 , y5644 , y5645 , y5646 , y5647 , y5648 , y5649 , y5650 , y5651 , y5652 , y5653 , y5654 , y5655 , y5656 , y5657 , y5658 , y5659 , y5660 , y5661 , y5662 , y5663 , y5664 , y5665 , y5666 , y5667 , y5668 , y5669 , y5670 , y5671 , y5672 , y5673 , y5674 , y5675 , y5676 , y5677 , y5678 , y5679 , y5680 , y5681 , y5682 , y5683 , y5684 , y5685 , y5686 , y5687 , y5688 , y5689 , y5690 , y5691 , y5692 , y5693 , y5694 , y5695 , y5696 , y5697 , y5698 , y5699 , y5700 , y5701 , y5702 , y5703 , y5704 , y5705 , y5706 , y5707 , y5708 , y5709 , y5710 , y5711 , y5712 , y5713 , y5714 , y5715 , y5716 , y5717 , y5718 , y5719 , y5720 , y5721 , y5722 , y5723 , y5724 , y5725 , y5726 , y5727 , y5728 , y5729 , y5730 , y5731 , y5732 , y5733 , y5734 , y5735 , y5736 , y5737 , y5738 , y5739 , y5740 , y5741 , y5742 , y5743 , y5744 , y5745 , y5746 , y5747 , y5748 , y5749 , y5750 , y5751 , y5752 , y5753 , y5754 , y5755 , y5756 , y5757 , y5758 , y5759 , y5760 , y5761 , y5762 , y5763 , y5764 , y5765 , y5766 , y5767 , y5768 , y5769 , y5770 , y5771 , y5772 , y5773 , y5774 , y5775 , y5776 , y5777 , y5778 , y5779 , y5780 , y5781 , y5782 , y5783 , y5784 , y5785 , y5786 , y5787 , y5788 , y5789 , y5790 , y5791 , y5792 , y5793 , y5794 , y5795 , y5796 , y5797 , y5798 , y5799 , y5800 , y5801 , y5802 , y5803 , y5804 , y5805 , y5806 , y5807 , y5808 , y5809 , y5810 , y5811 , y5812 , y5813 , y5814 , y5815 , y5816 , y5817 , y5818 , y5819 , y5820 , y5821 , y5822 , y5823 , y5824 , y5825 , y5826 , y5827 , y5828 , y5829 , y5830 , y5831 , y5832 , y5833 , y5834 , y5835 , y5836 , y5837 , y5838 , y5839 , y5840 , y5841 , y5842 , y5843 , y5844 , y5845 , y5846 , y5847 , y5848 , y5849 , y5850 , y5851 , y5852 , y5853 , y5854 , y5855 , y5856 , y5857 , y5858 , y5859 , y5860 , y5861 , y5862 , y5863 , y5864 , y5865 , y5866 , y5867 , y5868 , y5869 , y5870 , y5871 , y5872 , y5873 , y5874 , y5875 , y5876 , y5877 , y5878 , y5879 , y5880 , y5881 , y5882 , y5883 , y5884 , y5885 , y5886 , y5887 , y5888 , y5889 , y5890 , y5891 , y5892 , y5893 , y5894 , y5895 , y5896 , y5897 , y5898 , y5899 , y5900 , y5901 , y5902 , y5903 , y5904 , y5905 , y5906 , y5907 , y5908 , y5909 , y5910 , y5911 , y5912 , y5913 , y5914 , y5915 , y5916 , y5917 , y5918 , y5919 , y5920 , y5921 , y5922 , y5923 , y5924 , y5925 , y5926 , y5927 , y5928 , y5929 , y5930 , y5931 , y5932 , y5933 , y5934 , y5935 , y5936 , y5937 , y5938 , y5939 , y5940 , y5941 , y5942 , y5943 , y5944 , y5945 , y5946 , y5947 , y5948 , y5949 , y5950 , y5951 , y5952 , y5953 , y5954 , y5955 , y5956 , y5957 , y5958 , y5959 , y5960 , y5961 , y5962 , y5963 , y5964 , y5965 , y5966 , y5967 , y5968 , y5969 , y5970 , y5971 , y5972 , y5973 , y5974 , y5975 , y5976 , y5977 , y5978 , y5979 , y5980 , y5981 , y5982 , y5983 , y5984 , y5985 , y5986 , y5987 , y5988 , y5989 , y5990 , y5991 , y5992 , y5993 , y5994 , y5995 , y5996 , y5997 , y5998 , y5999 , y6000 , y6001 , y6002 , y6003 , y6004 , y6005 , y6006 , y6007 , y6008 , y6009 , y6010 , y6011 , y6012 , y6013 , y6014 , y6015 , y6016 , y6017 , y6018 , y6019 , y6020 , y6021 , y6022 , y6023 , y6024 , y6025 , y6026 , y6027 , y6028 , y6029 , y6030 , y6031 , y6032 , y6033 , y6034 , y6035 , y6036 , y6037 , y6038 , y6039 , y6040 , y6041 , y6042 , y6043 , y6044 , y6045 , y6046 , y6047 , y6048 , y6049 , y6050 , y6051 , y6052 , y6053 , y6054 , y6055 , y6056 , y6057 , y6058 , y6059 , y6060 , y6061 , y6062 , y6063 , y6064 , y6065 , y6066 , y6067 , y6068 , y6069 , y6070 , y6071 , y6072 , y6073 , y6074 , y6075 , y6076 , y6077 , y6078 , y6079 , y6080 , y6081 , y6082 , y6083 , y6084 , y6085 , y6086 , y6087 , y6088 , y6089 , y6090 , y6091 , y6092 , y6093 , y6094 , y6095 , y6096 , y6097 , y6098 , y6099 , y6100 , y6101 , y6102 , y6103 , y6104 , y6105 , y6106 , y6107 , y6108 , y6109 , y6110 , y6111 , y6112 , y6113 , y6114 , y6115 , y6116 , y6117 , y6118 , y6119 , y6120 , y6121 , y6122 , y6123 , y6124 , y6125 , y6126 , y6127 , y6128 , y6129 , y6130 , y6131 , y6132 , y6133 , y6134 , y6135 , y6136 , y6137 , y6138 , y6139 , y6140 , y6141 , y6142 , y6143 , y6144 , y6145 , y6146 , y6147 , y6148 , y6149 , y6150 , y6151 , y6152 , y6153 , y6154 , y6155 , y6156 , y6157 , y6158 , y6159 , y6160 , y6161 , y6162 , y6163 , y6164 , y6165 , y6166 , y6167 , y6168 , y6169 , y6170 , y6171 , y6172 , y6173 , y6174 , y6175 , y6176 , y6177 , y6178 , y6179 , y6180 , y6181 , y6182 , y6183 , y6184 , y6185 , y6186 , y6187 , y6188 , y6189 , y6190 , y6191 , y6192 , y6193 , y6194 , y6195 , y6196 , y6197 , y6198 , y6199 , y6200 , y6201 , y6202 , y6203 , y6204 , y6205 , y6206 , y6207 , y6208 , y6209 , y6210 , y6211 , y6212 , y6213 , y6214 , y6215 , y6216 , y6217 , y6218 , y6219 , y6220 , y6221 , y6222 , y6223 , y6224 , y6225 , y6226 , y6227 , y6228 , y6229 , y6230 , y6231 , y6232 , y6233 , y6234 , y6235 , y6236 , y6237 , y6238 , y6239 , y6240 , y6241 , y6242 , y6243 , y6244 , y6245 , y6246 , y6247 , y6248 , y6249 , y6250 , y6251 , y6252 , y6253 , y6254 , y6255 , y6256 , y6257 , y6258 , y6259 , y6260 , y6261 , y6262 , y6263 , y6264 , y6265 , y6266 , y6267 , y6268 , y6269 , y6270 , y6271 , y6272 , y6273 , y6274 , y6275 , y6276 , y6277 , y6278 , y6279 , y6280 , y6281 , y6282 , y6283 , y6284 , y6285 , y6286 , y6287 , y6288 , y6289 , y6290 , y6291 , y6292 , y6293 , y6294 , y6295 , y6296 , y6297 , y6298 , y6299 , y6300 , y6301 , y6302 , y6303 , y6304 , y6305 , y6306 , y6307 , y6308 , y6309 , y6310 , y6311 , y6312 , y6313 , y6314 , y6315 , y6316 , y6317 , y6318 , y6319 , y6320 , y6321 , y6322 , y6323 , y6324 , y6325 , y6326 , y6327 , y6328 , y6329 , y6330 , y6331 , y6332 , y6333 , y6334 , y6335 , y6336 , y6337 , y6338 , y6339 , y6340 , y6341 , y6342 , y6343 , y6344 , y6345 , y6346 , y6347 , y6348 , y6349 , y6350 , y6351 , y6352 , y6353 , y6354 , y6355 , y6356 , y6357 , y6358 , y6359 , y6360 , y6361 , y6362 , y6363 , y6364 , y6365 , y6366 , y6367 , y6368 , y6369 , y6370 , y6371 , y6372 , y6373 , y6374 , y6375 , y6376 , y6377 , y6378 , y6379 , y6380 , y6381 , y6382 , y6383 , y6384 , y6385 , y6386 , y6387 , y6388 , y6389 , y6390 , y6391 , y6392 , y6393 , y6394 , y6395 , y6396 , y6397 , y6398 , y6399 , y6400 , y6401 , y6402 , y6403 , y6404 , y6405 , y6406 , y6407 , y6408 , y6409 , y6410 , y6411 , y6412 , y6413 , y6414 , y6415 , y6416 , y6417 , y6418 , y6419 , y6420 , y6421 , y6422 , y6423 , y6424 , y6425 , y6426 , y6427 , y6428 , y6429 , y6430 , y6431 , y6432 , y6433 , y6434 , y6435 , y6436 , y6437 , y6438 , y6439 , y6440 , y6441 , y6442 , y6443 , y6444 , y6445 , y6446 , y6447 , y6448 , y6449 , y6450 , y6451 , y6452 , y6453 , y6454 , y6455 , y6456 , y6457 , y6458 , y6459 , y6460 , y6461 , y6462 , y6463 , y6464 , y6465 , y6466 , y6467 , y6468 , y6469 , y6470 , y6471 , y6472 , y6473 , y6474 , y6475 , y6476 , y6477 , y6478 , y6479 , y6480 , y6481 , y6482 , y6483 , y6484 , y6485 , y6486 , y6487 , y6488 , y6489 , y6490 , y6491 , y6492 , y6493 , y6494 , y6495 , y6496 , y6497 , y6498 , y6499 , y6500 , y6501 , y6502 , y6503 , y6504 , y6505 , y6506 , y6507 , y6508 , y6509 , y6510 , y6511 , y6512 , y6513 , y6514 , y6515 , y6516 , y6517 , y6518 , y6519 , y6520 , y6521 , y6522 , y6523 , y6524 , y6525 , y6526 , y6527 , y6528 , y6529 , y6530 , y6531 , y6532 , y6533 , y6534 , y6535 , y6536 , y6537 , y6538 , y6539 , y6540 , y6541 , y6542 , y6543 , y6544 , y6545 , y6546 , y6547 , y6548 , y6549 , y6550 , y6551 , y6552 , y6553 , y6554 , y6555 , y6556 , y6557 , y6558 , y6559 , y6560 , y6561 , y6562 , y6563 , y6564 , y6565 , y6566 , y6567 , y6568 , y6569 , y6570 , y6571 , y6572 , y6573 , y6574 , y6575 , y6576 , y6577 , y6578 , y6579 , y6580 , y6581 , y6582 , y6583 , y6584 , y6585 , y6586 , y6587 , y6588 , y6589 , y6590 , y6591 , y6592 , y6593 , y6594 , y6595 , y6596 , y6597 , y6598 , y6599 , y6600 , y6601 , y6602 , y6603 , y6604 , y6605 , y6606 , y6607 , y6608 , y6609 , y6610 , y6611 , y6612 , y6613 , y6614 , y6615 , y6616 , y6617 , y6618 , y6619 , y6620 , y6621 , y6622 , y6623 , y6624 , y6625 , y6626 , y6627 , y6628 , y6629 , y6630 , y6631 , y6632 , y6633 , y6634 , y6635 , y6636 , y6637 , y6638 , y6639 , y6640 , y6641 , y6642 , y6643 , y6644 , y6645 , y6646 , y6647 , y6648 , y6649 , y6650 , y6651 , y6652 , y6653 , y6654 , y6655 , y6656 , y6657 , y6658 , y6659 , y6660 , y6661 , y6662 , y6663 , y6664 , y6665 , y6666 , y6667 , y6668 , y6669 , y6670 , y6671 , y6672 , y6673 , y6674 , y6675 , y6676 , y6677 , y6678 , y6679 , y6680 , y6681 , y6682 , y6683 , y6684 , y6685 , y6686 , y6687 , y6688 , y6689 , y6690 , y6691 , y6692 , y6693 , y6694 , y6695 , y6696 , y6697 , y6698 , y6699 , y6700 , y6701 , y6702 , y6703 , y6704 , y6705 , y6706 , y6707 , y6708 , y6709 , y6710 , y6711 , y6712 , y6713 , y6714 , y6715 , y6716 , y6717 , y6718 , y6719 , y6720 , y6721 , y6722 , y6723 , y6724 , y6725 , y6726 , y6727 , y6728 , y6729 , y6730 , y6731 , y6732 , y6733 , y6734 , y6735 , y6736 , y6737 , y6738 , y6739 , y6740 , y6741 , y6742 , y6743 , y6744 , y6745 , y6746 , y6747 , y6748 , y6749 , y6750 , y6751 , y6752 , y6753 , y6754 , y6755 , y6756 , y6757 , y6758 , y6759 , y6760 , y6761 , y6762 , y6763 , y6764 , y6765 , y6766 , y6767 , y6768 , y6769 , y6770 , y6771 , y6772 , y6773 , y6774 , y6775 , y6776 , y6777 , y6778 , y6779 , y6780 , y6781 , y6782 , y6783 , y6784 , y6785 , y6786 , y6787 , y6788 , y6789 , y6790 , y6791 , y6792 , y6793 , y6794 , y6795 , y6796 , y6797 , y6798 , y6799 , y6800 , y6801 , y6802 , y6803 , y6804 , y6805 , y6806 , y6807 , y6808 , y6809 , y6810 , y6811 , y6812 , y6813 , y6814 , y6815 , y6816 , y6817 , y6818 , y6819 , y6820 , y6821 , y6822 , y6823 , y6824 , y6825 , y6826 , y6827 , y6828 , y6829 , y6830 , y6831 , y6832 , y6833 , y6834 , y6835 , y6836 , y6837 , y6838 , y6839 , y6840 , y6841 , y6842 , y6843 , y6844 , y6845 , y6846 , y6847 , y6848 , y6849 , y6850 , y6851 , y6852 , y6853 , y6854 , y6855 , y6856 , y6857 , y6858 , y6859 , y6860 , y6861 , y6862 , y6863 , y6864 , y6865 , y6866 , y6867 , y6868 , y6869 , y6870 , y6871 , y6872 , y6873 , y6874 , y6875 , y6876 , y6877 , y6878 , y6879 , y6880 , y6881 , y6882 , y6883 , y6884 , y6885 , y6886 , y6887 , y6888 , y6889 , y6890 , y6891 , y6892 , y6893 , y6894 , y6895 , y6896 , y6897 , y6898 , y6899 , y6900 , y6901 , y6902 , y6903 , y6904 , y6905 , y6906 , y6907 , y6908 , y6909 , y6910 , y6911 , y6912 , y6913 , y6914 , y6915 , y6916 , y6917 , y6918 , y6919 , y6920 , y6921 , y6922 , y6923 , y6924 , y6925 , y6926 , y6927 , y6928 , y6929 , y6930 , y6931 , y6932 , y6933 , y6934 , y6935 , y6936 , y6937 , y6938 , y6939 , y6940 , y6941 , y6942 , y6943 , y6944 , y6945 , y6946 , y6947 , y6948 , y6949 , y6950 , y6951 , y6952 , y6953 , y6954 , y6955 , y6956 , y6957 , y6958 , y6959 , y6960 , y6961 , y6962 , y6963 , y6964 , y6965 , y6966 , y6967 , y6968 , y6969 , y6970 , y6971 , y6972 , y6973 , y6974 , y6975 , y6976 , y6977 , y6978 , y6979 , y6980 , y6981 , y6982 , y6983 , y6984 , y6985 , y6986 , y6987 , y6988 , y6989 , y6990 , y6991 , y6992 , y6993 , y6994 , y6995 , y6996 , y6997 , y6998 , y6999 , y7000 , y7001 , y7002 , y7003 , y7004 , y7005 , y7006 , y7007 , y7008 , y7009 , y7010 , y7011 , y7012 , y7013 , y7014 , y7015 , y7016 , y7017 , y7018 , y7019 , y7020 , y7021 , y7022 , y7023 , y7024 , y7025 , y7026 , y7027 , y7028 , y7029 , y7030 , y7031 , y7032 , y7033 , y7034 , y7035 , y7036 , y7037 , y7038 , y7039 , y7040 , y7041 , y7042 , y7043 , y7044 , y7045 , y7046 , y7047 , y7048 , y7049 , y7050 , y7051 , y7052 , y7053 , y7054 , y7055 , y7056 , y7057 , y7058 , y7059 , y7060 , y7061 , y7062 , y7063 , y7064 , y7065 , y7066 , y7067 , y7068 , y7069 , y7070 , y7071 , y7072 , y7073 , y7074 , y7075 , y7076 , y7077 , y7078 , y7079 , y7080 , y7081 , y7082 , y7083 , y7084 , y7085 , y7086 , y7087 , y7088 , y7089 , y7090 , y7091 , y7092 , y7093 , y7094 , y7095 , y7096 , y7097 , y7098 , y7099 , y7100 , y7101 , y7102 , y7103 , y7104 , y7105 , y7106 , y7107 , y7108 , y7109 , y7110 , y7111 , y7112 , y7113 , y7114 , y7115 , y7116 , y7117 , y7118 , y7119 , y7120 , y7121 , y7122 , y7123 , y7124 , y7125 , y7126 , y7127 , y7128 , y7129 , y7130 , y7131 , y7132 , y7133 , y7134 , y7135 , y7136 , y7137 , y7138 , y7139 , y7140 , y7141 , y7142 , y7143 , y7144 , y7145 , y7146 , y7147 , y7148 , y7149 , y7150 , y7151 , y7152 , y7153 , y7154 , y7155 , y7156 , y7157 , y7158 , y7159 , y7160 , y7161 , y7162 , y7163 , y7164 , y7165 , y7166 , y7167 , y7168 , y7169 , y7170 , y7171 , y7172 , y7173 , y7174 , y7175 , y7176 , y7177 , y7178 , y7179 , y7180 , y7181 , y7182 , y7183 , y7184 , y7185 , y7186 , y7187 , y7188 , y7189 , y7190 , y7191 , y7192 , y7193 , y7194 , y7195 , y7196 , y7197 , y7198 , y7199 , y7200 , y7201 , y7202 , y7203 , y7204 , y7205 , y7206 , y7207 , y7208 , y7209 , y7210 , y7211 , y7212 , y7213 , y7214 , y7215 , y7216 , y7217 , y7218 , y7219 , y7220 , y7221 , y7222 , y7223 , y7224 , y7225 , y7226 , y7227 , y7228 , y7229 , y7230 , y7231 , y7232 , y7233 , y7234 , y7235 , y7236 , y7237 , y7238 , y7239 , y7240 , y7241 , y7242 , y7243 , y7244 , y7245 , y7246 , y7247 , y7248 , y7249 , y7250 , y7251 , y7252 , y7253 , y7254 , y7255 , y7256 , y7257 , y7258 , y7259 , y7260 , y7261 , y7262 , y7263 , y7264 , y7265 , y7266 , y7267 , y7268 , y7269 , y7270 , y7271 , y7272 , y7273 , y7274 , y7275 , y7276 , y7277 , y7278 , y7279 , y7280 , y7281 , y7282 , y7283 , y7284 , y7285 , y7286 , y7287 , y7288 , y7289 , y7290 , y7291 , y7292 , y7293 , y7294 , y7295 , y7296 , y7297 , y7298 , y7299 , y7300 , y7301 , y7302 , y7303 , y7304 , y7305 , y7306 , y7307 , y7308 , y7309 , y7310 , y7311 , y7312 , y7313 , y7314 , y7315 , y7316 , y7317 , y7318 , y7319 , y7320 , y7321 , y7322 , y7323 , y7324 , y7325 , y7326 , y7327 , y7328 , y7329 , y7330 , y7331 , y7332 , y7333 , y7334 , y7335 , y7336 , y7337 , y7338 , y7339 , y7340 , y7341 , y7342 , y7343 , y7344 , y7345 , y7346 , y7347 , y7348 , y7349 , y7350 , y7351 , y7352 , y7353 , y7354 , y7355 , y7356 , y7357 , y7358 , y7359 , y7360 , y7361 , y7362 , y7363 , y7364 , y7365 , y7366 , y7367 , y7368 , y7369 , y7370 , y7371 , y7372 , y7373 , y7374 , y7375 , y7376 , y7377 , y7378 , y7379 , y7380 , y7381 , y7382 , y7383 , y7384 , y7385 , y7386 , y7387 , y7388 , y7389 , y7390 , y7391 , y7392 , y7393 , y7394 , y7395 , y7396 , y7397 , y7398 , y7399 , y7400 , y7401 , y7402 , y7403 , y7404 , y7405 , y7406 , y7407 , y7408 , y7409 , y7410 , y7411 , y7412 , y7413 , y7414 , y7415 , y7416 , y7417 , y7418 , y7419 , y7420 , y7421 , y7422 , y7423 , y7424 , y7425 , y7426 , y7427 , y7428 , y7429 , y7430 , y7431 , y7432 , y7433 , y7434 , y7435 , y7436 , y7437 , y7438 , y7439 , y7440 , y7441 , y7442 , y7443 , y7444 , y7445 , y7446 , y7447 , y7448 , y7449 , y7450 , y7451 , y7452 , y7453 , y7454 , y7455 , y7456 , y7457 , y7458 , y7459 , y7460 , y7461 , y7462 , y7463 , y7464 , y7465 , y7466 , y7467 , y7468 , y7469 , y7470 , y7471 , y7472 , y7473 , y7474 , y7475 , y7476 , y7477 , y7478 , y7479 , y7480 , y7481 , y7482 , y7483 , y7484 , y7485 , y7486 , y7487 , y7488 , y7489 , y7490 , y7491 , y7492 , y7493 , y7494 , y7495 , y7496 , y7497 , y7498 , y7499 , y7500 , y7501 , y7502 , y7503 , y7504 , y7505 , y7506 , y7507 , y7508 , y7509 , y7510 , y7511 , y7512 , y7513 , y7514 , y7515 , y7516 , y7517 , y7518 , y7519 , y7520 , y7521 , y7522 , y7523 , y7524 , y7525 , y7526 , y7527 , y7528 , y7529 , y7530 , y7531 , y7532 , y7533 , y7534 , y7535 , y7536 , y7537 , y7538 , y7539 , y7540 , y7541 , y7542 , y7543 , y7544 , y7545 , y7546 , y7547 , y7548 , y7549 , y7550 , y7551 , y7552 , y7553 , y7554 , y7555 , y7556 , y7557 , y7558 , y7559 , y7560 , y7561 , y7562 , y7563 , y7564 , y7565 , y7566 , y7567 , y7568 , y7569 , y7570 , y7571 , y7572 , y7573 , y7574 , y7575 , y7576 , y7577 , y7578 , y7579 , y7580 , y7581 , y7582 , y7583 , y7584 , y7585 , y7586 , y7587 , y7588 , y7589 , y7590 , y7591 , y7592 , y7593 , y7594 , y7595 , y7596 , y7597 , y7598 , y7599 , y7600 , y7601 , y7602 , y7603 , y7604 , y7605 , y7606 , y7607 , y7608 , y7609 , y7610 , y7611 , y7612 , y7613 , y7614 , y7615 , y7616 , y7617 , y7618 , y7619 , y7620 , y7621 , y7622 , y7623 , y7624 , y7625 , y7626 , y7627 , y7628 , y7629 , y7630 , y7631 , y7632 , y7633 , y7634 , y7635 , y7636 , y7637 , y7638 , y7639 , y7640 , y7641 , y7642 , y7643 , y7644 , y7645 , y7646 , y7647 , y7648 , y7649 , y7650 , y7651 , y7652 , y7653 , y7654 , y7655 , y7656 , y7657 , y7658 , y7659 , y7660 , y7661 , y7662 , y7663 , y7664 , y7665 , y7666 , y7667 , y7668 , y7669 , y7670 , y7671 , y7672 , y7673 , y7674 , y7675 , y7676 , y7677 , y7678 , y7679 , y7680 , y7681 , y7682 , y7683 , y7684 , y7685 , y7686 , y7687 , y7688 , y7689 , y7690 , y7691 , y7692 , y7693 , y7694 , y7695 , y7696 , y7697 , y7698 , y7699 , y7700 , y7701 , y7702 , y7703 , y7704 , y7705 , y7706 , y7707 , y7708 , y7709 , y7710 , y7711 , y7712 , y7713 , y7714 , y7715 , y7716 , y7717 , y7718 , y7719 , y7720 , y7721 , y7722 , y7723 , y7724 , y7725 , y7726 , y7727 , y7728 , y7729 , y7730 , y7731 , y7732 , y7733 , y7734 , y7735 , y7736 , y7737 , y7738 , y7739 , y7740 , y7741 , y7742 , y7743 , y7744 , y7745 , y7746 , y7747 , y7748 , y7749 , y7750 , y7751 , y7752 , y7753 , y7754 , y7755 , y7756 , y7757 , y7758 , y7759 , y7760 , y7761 , y7762 , y7763 , y7764 , y7765 , y7766 , y7767 , y7768 , y7769 , y7770 , y7771 , y7772 , y7773 , y7774 , y7775 , y7776 , y7777 , y7778 , y7779 , y7780 , y7781 , y7782 , y7783 , y7784 , y7785 , y7786 , y7787 , y7788 , y7789 , y7790 , y7791 , y7792 , y7793 , y7794 , y7795 , y7796 , y7797 , y7798 , y7799 , y7800 , y7801 , y7802 , y7803 , y7804 , y7805 , y7806 , y7807 , y7808 , y7809 , y7810 , y7811 , y7812 , y7813 , y7814 , y7815 , y7816 , y7817 , y7818 , y7819 , y7820 , y7821 , y7822 , y7823 , y7824 , y7825 , y7826 , y7827 , y7828 , y7829 , y7830 , y7831 , y7832 , y7833 , y7834 , y7835 , y7836 , y7837 , y7838 , y7839 , y7840 , y7841 , y7842 , y7843 , y7844 , y7845 , y7846 , y7847 , y7848 , y7849 , y7850 , y7851 , y7852 , y7853 , y7854 , y7855 , y7856 , y7857 , y7858 , y7859 , y7860 , y7861 , y7862 , y7863 , y7864 , y7865 , y7866 , y7867 , y7868 , y7869 , y7870 , y7871 , y7872 , y7873 , y7874 , y7875 , y7876 , y7877 , y7878 , y7879 , y7880 , y7881 , y7882 , y7883 , y7884 , y7885 , y7886 , y7887 , y7888 , y7889 , y7890 , y7891 , y7892 , y7893 , y7894 , y7895 , y7896 , y7897 , y7898 , y7899 , y7900 , y7901 , y7902 , y7903 , y7904 , y7905 , y7906 , y7907 , y7908 , y7909 , y7910 , y7911 , y7912 , y7913 , y7914 , y7915 , y7916 , y7917 , y7918 , y7919 , y7920 , y7921 , y7922 , y7923 , y7924 , y7925 , y7926 , y7927 , y7928 , y7929 , y7930 , y7931 , y7932 , y7933 , y7934 , y7935 , y7936 , y7937 , y7938 , y7939 , y7940 , y7941 , y7942 , y7943 , y7944 , y7945 , y7946 , y7947 , y7948 , y7949 , y7950 , y7951 , y7952 , y7953 , y7954 , y7955 , y7956 , y7957 , y7958 , y7959 , y7960 , y7961 , y7962 , y7963 , y7964 , y7965 , y7966 , y7967 , y7968 , y7969 , y7970 , y7971 , y7972 , y7973 , y7974 , y7975 , y7976 , y7977 , y7978 , y7979 , y7980 , y7981 , y7982 , y7983 , y7984 , y7985 , y7986 , y7987 , y7988 , y7989 , y7990 , y7991 , y7992 , y7993 , y7994 , y7995 , y7996 , y7997 , y7998 , y7999 , y8000 , y8001 , y8002 , y8003 , y8004 , y8005 , y8006 , y8007 , y8008 , y8009 , y8010 , y8011 , y8012 , y8013 , y8014 , y8015 , y8016 , y8017 , y8018 , y8019 , y8020 , y8021 , y8022 , y8023 , y8024 , y8025 , y8026 , y8027 , y8028 , y8029 , y8030 , y8031 , y8032 , y8033 , y8034 , y8035 , y8036 , y8037 , y8038 , y8039 , y8040 , y8041 , y8042 , y8043 , y8044 , y8045 , y8046 , y8047 , y8048 , y8049 , y8050 , y8051 , y8052 , y8053 , y8054 , y8055 , y8056 , y8057 , y8058 , y8059 , y8060 , y8061 , y8062 , y8063 , y8064 , y8065 , y8066 , y8067 , y8068 , y8069 , y8070 , y8071 , y8072 , y8073 , y8074 , y8075 , y8076 , y8077 , y8078 , y8079 , y8080 , y8081 , y8082 , y8083 , y8084 , y8085 , y8086 , y8087 , y8088 , y8089 , y8090 , y8091 , y8092 , y8093 , y8094 , y8095 , y8096 , y8097 , y8098 , y8099 , y8100 , y8101 , y8102 , y8103 , y8104 , y8105 , y8106 , y8107 , y8108 , y8109 , y8110 , y8111 , y8112 , y8113 , y8114 , y8115 , y8116 , y8117 , y8118 , y8119 , y8120 , y8121 , y8122 , y8123 , y8124 , y8125 , y8126 , y8127 , y8128 , y8129 , y8130 , y8131 , y8132 , y8133 , y8134 , y8135 , y8136 , y8137 , y8138 , y8139 , y8140 , y8141 , y8142 , y8143 , y8144 , y8145 , y8146 , y8147 , y8148 , y8149 , y8150 , y8151 , y8152 , y8153 , y8154 , y8155 , y8156 , y8157 , y8158 , y8159 , y8160 , y8161 , y8162 , y8163 , y8164 , y8165 , y8166 , y8167 , y8168 , y8169 , y8170 , y8171 , y8172 , y8173 , y8174 , y8175 , y8176 , y8177 , y8178 , y8179 , y8180 , y8181 , y8182 , y8183 , y8184 , y8185 , y8186 , y8187 , y8188 , y8189 , y8190 , y8191 , y8192 , y8193 , y8194 , y8195 , y8196 , y8197 , y8198 , y8199 , y8200 , y8201 , y8202 , y8203 , y8204 , y8205 , y8206 , y8207 , y8208 , y8209 , y8210 , y8211 , y8212 , y8213 , y8214 , y8215 , y8216 , y8217 , y8218 , y8219 , y8220 , y8221 , y8222 , y8223 , y8224 , y8225 , y8226 , y8227 , y8228 , y8229 , y8230 , y8231 , y8232 , y8233 , y8234 , y8235 , y8236 , y8237 , y8238 , y8239 , y8240 , y8241 , y8242 , y8243 , y8244 , y8245 , y8246 , y8247 , y8248 , y8249 , y8250 , y8251 , y8252 , y8253 , y8254 , y8255 , y8256 , y8257 , y8258 , y8259 , y8260 , y8261 , y8262 , y8263 , y8264 , y8265 , y8266 , y8267 , y8268 , y8269 , y8270 , y8271 , y8272 , y8273 , y8274 , y8275 , y8276 , y8277 , y8278 , y8279 , y8280 , y8281 , y8282 , y8283 , y8284 , y8285 , y8286 , y8287 , y8288 , y8289 , y8290 , y8291 , y8292 , y8293 , y8294 , y8295 , y8296 , y8297 , y8298 , y8299 , y8300 , y8301 , y8302 , y8303 , y8304 , y8305 , y8306 , y8307 , y8308 , y8309 , y8310 , y8311 , y8312 , y8313 , y8314 , y8315 , y8316 , y8317 , y8318 , y8319 , y8320 , y8321 , y8322 , y8323 , y8324 , y8325 , y8326 , y8327 , y8328 , y8329 , y8330 , y8331 , y8332 , y8333 , y8334 , y8335 , y8336 , y8337 , y8338 , y8339 , y8340 , y8341 , y8342 , y8343 , y8344 , y8345 , y8346 , y8347 , y8348 , y8349 , y8350 , y8351 , y8352 , y8353 , y8354 , y8355 , y8356 , y8357 , y8358 , y8359 , y8360 , y8361 , y8362 , y8363 , y8364 , y8365 , y8366 , y8367 , y8368 , y8369 , y8370 , y8371 , y8372 , y8373 , y8374 , y8375 , y8376 , y8377 , y8378 , y8379 , y8380 , y8381 , y8382 , y8383 , y8384 , y8385 , y8386 , y8387 , y8388 , y8389 , y8390 , y8391 , y8392 , y8393 , y8394 , y8395 , y8396 , y8397 , y8398 , y8399 , y8400 , y8401 , y8402 , y8403 , y8404 , y8405 , y8406 , y8407 , y8408 , y8409 , y8410 , y8411 , y8412 , y8413 , y8414 , y8415 , y8416 , y8417 , y8418 , y8419 , y8420 , y8421 , y8422 , y8423 , y8424 , y8425 , y8426 , y8427 , y8428 , y8429 , y8430 , y8431 , y8432 , y8433 , y8434 , y8435 , y8436 , y8437 , y8438 , y8439 , y8440 , y8441 , y8442 , y8443 , y8444 , y8445 , y8446 , y8447 , y8448 , y8449 , y8450 , y8451 , y8452 , y8453 , y8454 , y8455 , y8456 , y8457 , y8458 , y8459 , y8460 , y8461 , y8462 , y8463 , y8464 , y8465 , y8466 , y8467 , y8468 , y8469 , y8470 , y8471 , y8472 , y8473 , y8474 , y8475 , y8476 , y8477 , y8478 , y8479 , y8480 , y8481 , y8482 , y8483 , y8484 , y8485 , y8486 , y8487 , y8488 , y8489 , y8490 , y8491 , y8492 , y8493 , y8494 , y8495 , y8496 , y8497 , y8498 , y8499 , y8500 , y8501 , y8502 , y8503 , y8504 , y8505 , y8506 , y8507 , y8508 , y8509 , y8510 , y8511 , y8512 , y8513 , y8514 , y8515 , y8516 , y8517 , y8518 , y8519 , y8520 , y8521 , y8522 , y8523 , y8524 , y8525 , y8526 , y8527 , y8528 , y8529 , y8530 , y8531 , y8532 , y8533 , y8534 , y8535 , y8536 , y8537 , y8538 , y8539 , y8540 , y8541 , y8542 , y8543 , y8544 , y8545 , y8546 , y8547 , y8548 , y8549 , y8550 , y8551 , y8552 , y8553 , y8554 , y8555 , y8556 , y8557 , y8558 , y8559 , y8560 , y8561 , y8562 , y8563 , y8564 , y8565 , y8566 , y8567 , y8568 , y8569 , y8570 , y8571 , y8572 , y8573 , y8574 , y8575 , y8576 , y8577 , y8578 , y8579 , y8580 , y8581 , y8582 , y8583 , y8584 , y8585 , y8586 , y8587 , y8588 , y8589 , y8590 , y8591 , y8592 , y8593 , y8594 , y8595 , y8596 , y8597 , y8598 , y8599 , y8600 , y8601 , y8602 , y8603 , y8604 , y8605 , y8606 , y8607 , y8608 , y8609 , y8610 , y8611 , y8612 , y8613 , y8614 , y8615 , y8616 , y8617 , y8618 , y8619 , y8620 , y8621 , y8622 , y8623 , y8624 , y8625 , y8626 , y8627 , y8628 , y8629 , y8630 , y8631 , y8632 , y8633 , y8634 , y8635 , y8636 , y8637 , y8638 , y8639 , y8640 , y8641 , y8642 , y8643 , y8644 , y8645 , y8646 , y8647 , y8648 , y8649 , y8650 , y8651 , y8652 , y8653 , y8654 , y8655 , y8656 , y8657 , y8658 , y8659 , y8660 , y8661 , y8662 , y8663 , y8664 , y8665 , y8666 , y8667 , y8668 , y8669 , y8670 , y8671 , y8672 , y8673 , y8674 , y8675 , y8676 , y8677 , y8678 , y8679 , y8680 , y8681 , y8682 , y8683 , y8684 , y8685 , y8686 , y8687 , y8688 , y8689 , y8690 , y8691 , y8692 , y8693 , y8694 , y8695 , y8696 , y8697 , y8698 , y8699 , y8700 , y8701 , y8702 , y8703 , y8704 , y8705 , y8706 , y8707 , y8708 , y8709 , y8710 , y8711 , y8712 , y8713 , y8714 , y8715 , y8716 , y8717 , y8718 , y8719 , y8720 , y8721 , y8722 , y8723 , y8724 , y8725 , y8726 , y8727 , y8728 , y8729 , y8730 , y8731 , y8732 , y8733 , y8734 , y8735 , y8736 , y8737 , y8738 , y8739 , y8740 , y8741 , y8742 , y8743 , y8744 , y8745 , y8746 , y8747 , y8748 , y8749 , y8750 , y8751 , y8752 , y8753 , y8754 , y8755 , y8756 , y8757 , y8758 , y8759 , y8760 , y8761 , y8762 , y8763 , y8764 , y8765 , y8766 , y8767 , y8768 , y8769 , y8770 , y8771 , y8772 , y8773 , y8774 , y8775 , y8776 , y8777 , y8778 , y8779 , y8780 , y8781 , y8782 , y8783 , y8784 , y8785 , y8786 , y8787 , y8788 , y8789 , y8790 , y8791 , y8792 , y8793 , y8794 , y8795 , y8796 , y8797 , y8798 , y8799 , y8800 , y8801 , y8802 , y8803 , y8804 , y8805 , y8806 , y8807 , y8808 , y8809 , y8810 , y8811 , y8812 , y8813 , y8814 , y8815 , y8816 , y8817 , y8818 , y8819 , y8820 , y8821 , y8822 , y8823 , y8824 , y8825 , y8826 , y8827 , y8828 , y8829 , y8830 , y8831 , y8832 , y8833 , y8834 , y8835 , y8836 , y8837 , y8838 , y8839 , y8840 , y8841 , y8842 , y8843 , y8844 , y8845 , y8846 , y8847 , y8848 , y8849 , y8850 , y8851 , y8852 , y8853 , y8854 , y8855 , y8856 , y8857 , y8858 , y8859 , y8860 , y8861 , y8862 , y8863 , y8864 , y8865 , y8866 , y8867 , y8868 , y8869 , y8870 , y8871 , y8872 , y8873 , y8874 , y8875 , y8876 , y8877 , y8878 , y8879 , y8880 , y8881 , y8882 , y8883 , y8884 , y8885 , y8886 , y8887 , y8888 , y8889 , y8890 , y8891 , y8892 , y8893 , y8894 , y8895 , y8896 , y8897 , y8898 , y8899 , y8900 , y8901 , y8902 , y8903 , y8904 , y8905 , y8906 , y8907 , y8908 , y8909 , y8910 , y8911 , y8912 , y8913 , y8914 , y8915 , y8916 , y8917 , y8918 , y8919 , y8920 , y8921 , y8922 , y8923 , y8924 , y8925 , y8926 , y8927 , y8928 ;
  wire n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 ;
  assign n129 = ( ~x8 & x29 ) | ( ~x8 & x64 ) | ( x29 & x64 ) ;
  assign n130 = ( x71 & x86 ) | ( x71 & ~x89 ) | ( x86 & ~x89 ) ;
  assign n131 = ( ~x13 & x56 ) | ( ~x13 & x83 ) | ( x56 & x83 ) ;
  assign n132 = x111 ^ x42 ^ x15 ;
  assign n133 = x103 ^ x61 ^ x50 ;
  assign n134 = x118 ^ x78 ^ x34 ;
  assign n135 = n134 ^ x110 ^ x41 ;
  assign n136 = ( x4 & x35 ) | ( x4 & ~n135 ) | ( x35 & ~n135 ) ;
  assign n137 = x67 ^ x59 ^ x31 ;
  assign n138 = ~x63 & x123 ;
  assign n139 = ( x8 & x69 ) | ( x8 & ~x94 ) | ( x69 & ~x94 ) ;
  assign n140 = ( ~x48 & x85 ) | ( ~x48 & n139 ) | ( x85 & n139 ) ;
  assign n141 = x60 & x124 ;
  assign n142 = ~x58 & n141 ;
  assign n143 = ( x5 & ~x52 ) | ( x5 & n142 ) | ( ~x52 & n142 ) ;
  assign n144 = x113 ^ x74 ^ x26 ;
  assign n145 = x127 ^ x67 ^ x34 ;
  assign n152 = ( x65 & x70 ) | ( x65 & ~x73 ) | ( x70 & ~x73 ) ;
  assign n146 = x72 ^ x26 ^ x18 ;
  assign n147 = ( x32 & x86 ) | ( x32 & n146 ) | ( x86 & n146 ) ;
  assign n148 = ( x74 & n138 ) | ( x74 & n147 ) | ( n138 & n147 ) ;
  assign n149 = x91 ^ x16 ^ 1'b0 ;
  assign n150 = n148 & n149 ;
  assign n151 = ( ~x58 & x59 ) | ( ~x58 & n150 ) | ( x59 & n150 ) ;
  assign n153 = n152 ^ n151 ^ n144 ;
  assign n154 = x123 ^ x118 ^ x74 ;
  assign n155 = ( ~x72 & x100 ) | ( ~x72 & n154 ) | ( x100 & n154 ) ;
  assign n156 = n155 ^ x116 ^ 1'b0 ;
  assign n157 = x75 & ~n156 ;
  assign n158 = x106 ^ x105 ^ 1'b0 ;
  assign n159 = n157 & n158 ;
  assign n167 = n134 ^ x39 ^ x22 ;
  assign n165 = ( x93 & ~x98 ) | ( x93 & x103 ) | ( ~x98 & x103 ) ;
  assign n166 = ( ~x110 & x112 ) | ( ~x110 & n165 ) | ( x112 & n165 ) ;
  assign n160 = x94 ^ x88 ^ x24 ;
  assign n161 = n131 ^ x66 ^ x18 ;
  assign n162 = x96 & ~n161 ;
  assign n163 = ~x0 & n162 ;
  assign n164 = ( n144 & n160 ) | ( n144 & ~n163 ) | ( n160 & ~n163 ) ;
  assign n168 = n167 ^ n166 ^ n164 ;
  assign n169 = x110 ^ x90 ^ x21 ;
  assign n170 = n169 ^ x109 ^ x17 ;
  assign n175 = x90 ^ x2 ^ 1'b0 ;
  assign n171 = ( ~x0 & x40 ) | ( ~x0 & x44 ) | ( x40 & x44 ) ;
  assign n172 = x114 ^ x103 ^ x64 ;
  assign n173 = n172 ^ x41 ^ x1 ;
  assign n174 = ( n160 & ~n171 ) | ( n160 & n173 ) | ( ~n171 & n173 ) ;
  assign n176 = n175 ^ n174 ^ x39 ;
  assign n177 = x24 & x91 ;
  assign n178 = ~x110 & n177 ;
  assign n179 = n178 ^ x12 ^ 1'b0 ;
  assign n180 = x64 & ~n179 ;
  assign n181 = n180 ^ x97 ^ x95 ;
  assign n192 = x64 & x104 ;
  assign n188 = x71 ^ x55 ^ x41 ;
  assign n189 = n188 ^ x115 ^ x8 ;
  assign n190 = ( x50 & ~x113 ) | ( x50 & n189 ) | ( ~x113 & n189 ) ;
  assign n191 = ( x26 & x109 ) | ( x26 & ~n190 ) | ( x109 & ~n190 ) ;
  assign n182 = x22 & x124 ;
  assign n183 = ~x18 & n182 ;
  assign n184 = ( x15 & ~x28 ) | ( x15 & x80 ) | ( ~x28 & x80 ) ;
  assign n185 = ~n183 & n184 ;
  assign n186 = n185 ^ n171 ^ 1'b0 ;
  assign n187 = ( ~x3 & x78 ) | ( ~x3 & n186 ) | ( x78 & n186 ) ;
  assign n193 = n192 ^ n191 ^ n187 ;
  assign n194 = ( x66 & x96 ) | ( x66 & ~x124 ) | ( x96 & ~x124 ) ;
  assign n195 = n178 ^ x116 ^ x110 ;
  assign n196 = ( x32 & n154 ) | ( x32 & n195 ) | ( n154 & n195 ) ;
  assign n201 = n137 ^ x105 ^ x89 ;
  assign n199 = n148 ^ x54 ^ x52 ;
  assign n197 = n145 ^ x64 ^ x41 ;
  assign n198 = ( ~x36 & x60 ) | ( ~x36 & n197 ) | ( x60 & n197 ) ;
  assign n200 = n199 ^ n198 ^ n195 ;
  assign n202 = n201 ^ n200 ^ x30 ;
  assign n204 = ( x97 & x114 ) | ( x97 & ~n195 ) | ( x114 & ~n195 ) ;
  assign n203 = n130 ^ x45 ^ x1 ;
  assign n205 = n204 ^ n203 ^ x125 ;
  assign n206 = x86 & x97 ;
  assign n207 = ( x54 & ~n205 ) | ( x54 & n206 ) | ( ~n205 & n206 ) ;
  assign n208 = x43 ^ x37 ^ 1'b0 ;
  assign n209 = n129 & n208 ;
  assign n210 = ( x15 & ~x84 ) | ( x15 & n209 ) | ( ~x84 & n209 ) ;
  assign n211 = ( x80 & x103 ) | ( x80 & ~n210 ) | ( x103 & ~n210 ) ;
  assign n212 = ~x4 & x12 ;
  assign n213 = n212 ^ n195 ^ x28 ;
  assign n214 = n213 ^ x108 ^ x7 ;
  assign n215 = ( x57 & n130 ) | ( x57 & n178 ) | ( n130 & n178 ) ;
  assign n216 = n189 ^ x82 ^ x37 ;
  assign n217 = n216 ^ x73 ^ 1'b0 ;
  assign n218 = x76 & ~n217 ;
  assign n219 = ( n164 & ~n199 ) | ( n164 & n218 ) | ( ~n199 & n218 ) ;
  assign n220 = ( x14 & n215 ) | ( x14 & ~n219 ) | ( n215 & ~n219 ) ;
  assign n221 = x87 ^ x49 ^ x28 ;
  assign n222 = n221 ^ n192 ^ x102 ;
  assign n223 = ( ~x41 & x44 ) | ( ~x41 & n222 ) | ( x44 & n222 ) ;
  assign n224 = n223 ^ x115 ^ x41 ;
  assign n225 = x43 ^ x28 ^ x7 ;
  assign n226 = ( x19 & ~x36 ) | ( x19 & x88 ) | ( ~x36 & x88 ) ;
  assign n227 = ( x86 & ~x124 ) | ( x86 & n226 ) | ( ~x124 & n226 ) ;
  assign n228 = n227 ^ x70 ^ x13 ;
  assign n229 = ( x13 & x57 ) | ( x13 & ~x68 ) | ( x57 & ~x68 ) ;
  assign n230 = ( ~x99 & x118 ) | ( ~x99 & n229 ) | ( x118 & n229 ) ;
  assign n231 = x112 & n171 ;
  assign n232 = ~x64 & n231 ;
  assign n233 = n230 & n232 ;
  assign n234 = ( ~n147 & n228 ) | ( ~n147 & n233 ) | ( n228 & n233 ) ;
  assign n235 = n234 ^ n165 ^ x53 ;
  assign n236 = ~n225 & n235 ;
  assign n237 = n224 & n236 ;
  assign n241 = x111 ^ x87 ^ x42 ;
  assign n242 = n241 ^ x98 ^ x76 ;
  assign n243 = n242 ^ x50 ^ x36 ;
  assign n239 = ( x70 & ~n161 ) | ( x70 & n174 ) | ( ~n161 & n174 ) ;
  assign n240 = ( x70 & ~x119 ) | ( x70 & n239 ) | ( ~x119 & n239 ) ;
  assign n244 = n243 ^ n240 ^ x36 ;
  assign n238 = n215 ^ n209 ^ x85 ;
  assign n245 = n244 ^ n238 ^ x39 ;
  assign n246 = n243 ^ n242 ^ x94 ;
  assign n247 = ( x43 & ~x51 ) | ( x43 & n143 ) | ( ~x51 & n143 ) ;
  assign n248 = n246 | n247 ;
  assign n249 = ~x99 & n248 ;
  assign n250 = ( x29 & n245 ) | ( x29 & n249 ) | ( n245 & n249 ) ;
  assign n254 = n160 | n230 ;
  assign n251 = ( ~x17 & x54 ) | ( ~x17 & n131 ) | ( x54 & n131 ) ;
  assign n252 = n251 ^ x55 ^ x2 ;
  assign n253 = ( x82 & ~x91 ) | ( x82 & n252 ) | ( ~x91 & n252 ) ;
  assign n255 = n254 ^ n253 ^ n215 ;
  assign n260 = x62 ^ x57 ^ x22 ;
  assign n261 = n260 ^ x114 ^ x49 ;
  assign n262 = n261 ^ x11 ^ 1'b0 ;
  assign n263 = ~n164 & n262 ;
  assign n259 = ( ~x7 & x115 ) | ( ~x7 & n174 ) | ( x115 & n174 ) ;
  assign n256 = x2 & ~n225 ;
  assign n257 = ( x72 & x121 ) | ( x72 & ~n256 ) | ( x121 & ~n256 ) ;
  assign n258 = n257 ^ n191 ^ n146 ;
  assign n264 = n263 ^ n259 ^ n258 ;
  assign n265 = x117 ^ x97 ^ x22 ;
  assign n267 = n213 ^ x77 ^ 1'b0 ;
  assign n266 = ( n172 & n218 ) | ( n172 & ~n223 ) | ( n218 & ~n223 ) ;
  assign n268 = n267 ^ n266 ^ n234 ;
  assign n269 = ( n159 & n265 ) | ( n159 & n268 ) | ( n265 & n268 ) ;
  assign n270 = ( x29 & x88 ) | ( x29 & n133 ) | ( x88 & n133 ) ;
  assign n271 = x92 ^ x67 ^ x47 ;
  assign n272 = ( ~x19 & x80 ) | ( ~x19 & x97 ) | ( x80 & x97 ) ;
  assign n273 = n226 ^ x106 ^ x87 ;
  assign n274 = ( ~x12 & x25 ) | ( ~x12 & n273 ) | ( x25 & n273 ) ;
  assign n275 = x57 & ~n274 ;
  assign n276 = ~n272 & n275 ;
  assign n277 = n276 ^ n159 ^ x113 ;
  assign n278 = ( x42 & n271 ) | ( x42 & n277 ) | ( n271 & n277 ) ;
  assign n279 = ( x34 & n252 ) | ( x34 & n278 ) | ( n252 & n278 ) ;
  assign n285 = x105 ^ x68 ^ x52 ;
  assign n280 = ( x81 & n137 ) | ( x81 & n183 ) | ( n137 & n183 ) ;
  assign n281 = x74 & ~n137 ;
  assign n282 = x44 & ~n281 ;
  assign n283 = x122 & n282 ;
  assign n284 = ( x123 & n280 ) | ( x123 & n283 ) | ( n280 & n283 ) ;
  assign n286 = n285 ^ n284 ^ x92 ;
  assign n287 = n227 ^ n135 ^ x60 ;
  assign n288 = x77 ^ x32 ^ x13 ;
  assign n289 = n288 ^ x16 ^ x7 ;
  assign n290 = n289 ^ n151 ^ x111 ;
  assign n291 = n290 ^ n201 ^ n144 ;
  assign n292 = ( x28 & ~n246 ) | ( x28 & n291 ) | ( ~n246 & n291 ) ;
  assign n293 = ( ~x116 & n178 ) | ( ~x116 & n198 ) | ( n178 & n198 ) ;
  assign n294 = ( n180 & n202 ) | ( n180 & ~n293 ) | ( n202 & ~n293 ) ;
  assign n296 = ( x101 & ~n209 ) | ( x101 & n229 ) | ( ~n209 & n229 ) ;
  assign n295 = n263 ^ n146 ^ x91 ;
  assign n297 = n296 ^ n295 ^ 1'b0 ;
  assign n298 = n297 ^ x107 ^ x79 ;
  assign n299 = n294 & ~n298 ;
  assign n300 = n299 ^ n260 ^ 1'b0 ;
  assign n301 = n300 ^ n298 ^ n165 ;
  assign n302 = ( x27 & x59 ) | ( x27 & ~x125 ) | ( x59 & ~x125 ) ;
  assign n303 = ( x105 & x126 ) | ( x105 & ~n302 ) | ( x126 & ~n302 ) ;
  assign n304 = ( x106 & n172 ) | ( x106 & n303 ) | ( n172 & n303 ) ;
  assign n305 = x126 & n221 ;
  assign n306 = n227 ^ x41 ^ 1'b0 ;
  assign n307 = ~n188 & n306 ;
  assign n308 = x104 ^ x17 ^ 1'b0 ;
  assign n309 = ~n146 & n308 ;
  assign n310 = ( x3 & x78 ) | ( x3 & ~n309 ) | ( x78 & ~n309 ) ;
  assign n311 = ( n204 & ~n307 ) | ( n204 & n310 ) | ( ~n307 & n310 ) ;
  assign n322 = x96 ^ x43 ^ x23 ;
  assign n324 = x115 ^ x29 ^ x26 ;
  assign n325 = n225 ^ x106 ^ x1 ;
  assign n326 = n324 & n325 ;
  assign n323 = x113 ^ x76 ^ x74 ;
  assign n327 = n326 ^ n323 ^ 1'b0 ;
  assign n328 = x11 & n327 ;
  assign n329 = ( x120 & n322 ) | ( x120 & ~n328 ) | ( n322 & ~n328 ) ;
  assign n312 = n293 ^ x103 ^ x92 ;
  assign n313 = x46 ^ x19 ^ x11 ;
  assign n314 = ( x48 & x58 ) | ( x48 & n313 ) | ( x58 & n313 ) ;
  assign n315 = ( x60 & n160 ) | ( x60 & ~n314 ) | ( n160 & ~n314 ) ;
  assign n316 = x103 & ~n315 ;
  assign n317 = n316 ^ x52 ^ 1'b0 ;
  assign n318 = n317 ^ n145 ^ x111 ;
  assign n319 = n318 ^ n163 ^ x23 ;
  assign n320 = ( n225 & n312 ) | ( n225 & ~n319 ) | ( n312 & ~n319 ) ;
  assign n321 = n320 ^ n178 ^ x104 ;
  assign n330 = n329 ^ n321 ^ x100 ;
  assign n331 = ( ~x1 & x10 ) | ( ~x1 & n226 ) | ( x10 & n226 ) ;
  assign n332 = ( n145 & n170 ) | ( n145 & n331 ) | ( n170 & n331 ) ;
  assign n345 = ( x2 & ~n239 ) | ( x2 & n296 ) | ( ~n239 & n296 ) ;
  assign n346 = ( ~x38 & n183 ) | ( ~x38 & n345 ) | ( n183 & n345 ) ;
  assign n347 = n346 ^ x66 ^ x38 ;
  assign n348 = n347 ^ x116 ^ x98 ;
  assign n341 = x73 ^ x66 ^ 1'b0 ;
  assign n342 = n341 ^ x50 ^ 1'b0 ;
  assign n343 = ( n216 & ~n271 ) | ( n216 & n342 ) | ( ~n271 & n342 ) ;
  assign n340 = n246 ^ x73 ^ x42 ;
  assign n344 = n343 ^ n340 ^ n213 ;
  assign n333 = ( x27 & x33 ) | ( x27 & n322 ) | ( x33 & n322 ) ;
  assign n334 = ( x66 & ~n215 ) | ( x66 & n257 ) | ( ~n215 & n257 ) ;
  assign n335 = ( n312 & ~n333 ) | ( n312 & n334 ) | ( ~n333 & n334 ) ;
  assign n336 = n259 ^ n160 ^ x90 ;
  assign n337 = ( n168 & n202 ) | ( n168 & n336 ) | ( n202 & n336 ) ;
  assign n338 = n335 & ~n337 ;
  assign n339 = ~n165 & n338 ;
  assign n349 = n348 ^ n344 ^ n339 ;
  assign n351 = ( ~x36 & x99 ) | ( ~x36 & x124 ) | ( x99 & x124 ) ;
  assign n352 = ( x76 & n146 ) | ( x76 & ~n351 ) | ( n146 & ~n351 ) ;
  assign n353 = ( x10 & n132 ) | ( x10 & ~n352 ) | ( n132 & ~n352 ) ;
  assign n350 = n343 ^ n341 ^ 1'b0 ;
  assign n354 = n353 ^ n350 ^ n263 ;
  assign n355 = ~x106 & x116 ;
  assign n356 = n355 ^ n284 ^ x27 ;
  assign n357 = ( x92 & x121 ) | ( x92 & ~n356 ) | ( x121 & ~n356 ) ;
  assign n358 = ( x7 & ~x27 ) | ( x7 & n260 ) | ( ~x27 & n260 ) ;
  assign n359 = ( ~x10 & x27 ) | ( ~x10 & x91 ) | ( x27 & x91 ) ;
  assign n360 = ( ~x60 & x108 ) | ( ~x60 & n359 ) | ( x108 & n359 ) ;
  assign n361 = n360 ^ n353 ^ n147 ;
  assign n364 = n243 ^ n132 ^ x110 ;
  assign n365 = ( n154 & n188 ) | ( n154 & ~n364 ) | ( n188 & ~n364 ) ;
  assign n362 = n195 ^ x32 ^ x22 ;
  assign n363 = n362 ^ n315 ^ n190 ;
  assign n366 = n365 ^ n363 ^ n191 ;
  assign n367 = n199 ^ x79 ^ x38 ;
  assign n368 = ( ~x109 & n314 ) | ( ~x109 & n367 ) | ( n314 & n367 ) ;
  assign n369 = n368 ^ n267 ^ x18 ;
  assign n370 = ( x72 & n366 ) | ( x72 & n369 ) | ( n366 & n369 ) ;
  assign n371 = ( ~n358 & n361 ) | ( ~n358 & n370 ) | ( n361 & n370 ) ;
  assign n378 = x51 & x96 ;
  assign n379 = n378 ^ n131 ^ 1'b0 ;
  assign n380 = n226 ^ n169 ^ x41 ;
  assign n381 = ( ~x4 & n379 ) | ( ~x4 & n380 ) | ( n379 & n380 ) ;
  assign n376 = ( x81 & n152 ) | ( x81 & ~n281 ) | ( n152 & ~n281 ) ;
  assign n374 = n252 ^ x26 ^ x21 ;
  assign n375 = ( x88 & n186 ) | ( x88 & ~n374 ) | ( n186 & ~n374 ) ;
  assign n377 = n376 ^ n375 ^ x106 ;
  assign n372 = n140 ^ x44 ^ x32 ;
  assign n373 = ( x65 & n325 ) | ( x65 & n372 ) | ( n325 & n372 ) ;
  assign n382 = n381 ^ n377 ^ n373 ;
  assign n383 = ( x21 & n273 ) | ( x21 & n331 ) | ( n273 & n331 ) ;
  assign n384 = n383 ^ n178 ^ x64 ;
  assign n387 = ( ~x61 & n137 ) | ( ~x61 & n148 ) | ( n137 & n148 ) ;
  assign n388 = ( n140 & n326 ) | ( n140 & n387 ) | ( n326 & n387 ) ;
  assign n385 = x46 & x93 ;
  assign n386 = ( x4 & ~x85 ) | ( x4 & n385 ) | ( ~x85 & n385 ) ;
  assign n389 = n388 ^ n386 ^ x77 ;
  assign n390 = n247 & n389 ;
  assign n391 = n325 ^ n151 ^ x58 ;
  assign n392 = x16 & ~n291 ;
  assign n393 = ( n201 & n391 ) | ( n201 & n392 ) | ( n391 & n392 ) ;
  assign n394 = x40 & ~n365 ;
  assign n395 = n394 ^ n248 ^ 1'b0 ;
  assign n396 = n148 & n395 ;
  assign n397 = x37 & n396 ;
  assign n398 = n397 ^ n164 ^ 1'b0 ;
  assign n399 = ( n232 & n393 ) | ( n232 & n398 ) | ( n393 & n398 ) ;
  assign n412 = n391 ^ n353 ^ x121 ;
  assign n413 = x80 & n412 ;
  assign n414 = n322 & n413 ;
  assign n415 = x107 ^ x104 ^ x52 ;
  assign n416 = n415 ^ x53 ^ x18 ;
  assign n417 = ( ~n227 & n414 ) | ( ~n227 & n416 ) | ( n414 & n416 ) ;
  assign n418 = ( n280 & ~n282 ) | ( n280 & n417 ) | ( ~n282 & n417 ) ;
  assign n411 = ( ~x0 & n168 ) | ( ~x0 & n189 ) | ( n168 & n189 ) ;
  assign n405 = ( x59 & ~x116 ) | ( x59 & n221 ) | ( ~x116 & n221 ) ;
  assign n406 = ( ~x20 & x88 ) | ( ~x20 & x126 ) | ( x88 & x126 ) ;
  assign n407 = n406 ^ x88 ^ 1'b0 ;
  assign n408 = ~n405 & n407 ;
  assign n409 = n408 ^ x93 ^ x41 ;
  assign n400 = x27 & n143 ;
  assign n401 = x110 ^ x103 ^ x99 ;
  assign n402 = n296 & ~n401 ;
  assign n403 = n402 ^ x110 ^ 1'b0 ;
  assign n404 = ( n239 & n400 ) | ( n239 & n403 ) | ( n400 & n403 ) ;
  assign n410 = n409 ^ n404 ^ x47 ;
  assign n419 = n418 ^ n411 ^ n410 ;
  assign n420 = ( ~n166 & n201 ) | ( ~n166 & n277 ) | ( n201 & n277 ) ;
  assign n421 = n420 ^ n146 ^ x63 ;
  assign n422 = ( ~x62 & n197 ) | ( ~x62 & n421 ) | ( n197 & n421 ) ;
  assign n423 = ( n169 & ~n195 ) | ( n169 & n422 ) | ( ~n195 & n422 ) ;
  assign n424 = n181 ^ x36 ^ x28 ;
  assign n425 = ~n423 & n424 ;
  assign n426 = ~x37 & n425 ;
  assign n427 = n426 ^ n381 ^ 1'b0 ;
  assign n431 = x104 ^ x61 ^ x21 ;
  assign n432 = n431 ^ n129 ^ x32 ;
  assign n433 = n432 ^ n318 ^ x19 ;
  assign n434 = x3 & n433 ;
  assign n435 = n323 & n434 ;
  assign n428 = ( ~x2 & x115 ) | ( ~x2 & n365 ) | ( x115 & n365 ) ;
  assign n429 = n428 ^ x113 ^ x36 ;
  assign n430 = ( ~x1 & n178 ) | ( ~x1 & n429 ) | ( n178 & n429 ) ;
  assign n436 = n435 ^ n430 ^ n272 ;
  assign n448 = n345 ^ n335 ^ x86 ;
  assign n447 = ( x16 & ~n196 ) | ( x16 & n255 ) | ( ~n196 & n255 ) ;
  assign n437 = n142 ^ n139 ^ x111 ;
  assign n438 = ( n167 & n169 ) | ( n167 & n437 ) | ( n169 & n437 ) ;
  assign n439 = n438 ^ n257 ^ n175 ;
  assign n440 = ( ~n230 & n303 ) | ( ~n230 & n362 ) | ( n303 & n362 ) ;
  assign n441 = n438 ^ n163 ^ 1'b0 ;
  assign n442 = n440 | n441 ;
  assign n443 = n273 ^ n259 ^ x104 ;
  assign n444 = ( x120 & n418 ) | ( x120 & n443 ) | ( n418 & n443 ) ;
  assign n445 = ( n439 & n442 ) | ( n439 & ~n444 ) | ( n442 & ~n444 ) ;
  assign n446 = ( x126 & n154 ) | ( x126 & ~n445 ) | ( n154 & ~n445 ) ;
  assign n449 = n448 ^ n447 ^ n446 ;
  assign n457 = n256 ^ n188 ^ x5 ;
  assign n455 = n387 ^ x16 ^ x3 ;
  assign n454 = n388 ^ n246 ^ x92 ;
  assign n450 = ( x99 & ~n243 ) | ( x99 & n405 ) | ( ~n243 & n405 ) ;
  assign n451 = ( x42 & ~n331 ) | ( x42 & n450 ) | ( ~n331 & n450 ) ;
  assign n452 = ( n192 & n362 ) | ( n192 & ~n451 ) | ( n362 & ~n451 ) ;
  assign n453 = n452 ^ n283 ^ x67 ;
  assign n456 = n455 ^ n454 ^ n453 ;
  assign n458 = n457 ^ n456 ^ n160 ;
  assign n471 = ~x46 & n246 ;
  assign n469 = ( ~x42 & x105 ) | ( ~x42 & x107 ) | ( x105 & x107 ) ;
  assign n466 = n341 ^ x114 ^ x67 ;
  assign n467 = n466 ^ x105 ^ x91 ;
  assign n468 = n467 ^ n351 ^ n256 ;
  assign n470 = n469 ^ n468 ^ x20 ;
  assign n462 = ( ~x114 & n242 ) | ( ~x114 & n302 ) | ( n242 & n302 ) ;
  assign n463 = ( x10 & ~x120 ) | ( x10 & n462 ) | ( ~x120 & n462 ) ;
  assign n464 = ( n219 & ~n240 ) | ( n219 & n463 ) | ( ~n240 & n463 ) ;
  assign n459 = ( x52 & n155 ) | ( x52 & n366 ) | ( n155 & n366 ) ;
  assign n460 = n459 ^ x75 ^ x53 ;
  assign n461 = n460 ^ n347 ^ x71 ;
  assign n465 = n464 ^ n461 ^ n258 ;
  assign n472 = n471 ^ n470 ^ n465 ;
  assign n479 = ( x27 & x85 ) | ( x27 & ~x96 ) | ( x85 & ~x96 ) ;
  assign n480 = ( x67 & n212 ) | ( x67 & ~n479 ) | ( n212 & ~n479 ) ;
  assign n475 = ( x76 & ~n163 ) | ( x76 & n212 ) | ( ~n163 & n212 ) ;
  assign n476 = x75 ^ x53 ^ 1'b0 ;
  assign n477 = n475 & n476 ;
  assign n473 = n372 ^ n314 ^ x25 ;
  assign n474 = n473 ^ n313 ^ n164 ;
  assign n478 = n477 ^ n474 ^ n171 ;
  assign n481 = n480 ^ n478 ^ n375 ;
  assign n486 = n291 | n461 ;
  assign n482 = n392 ^ n260 ^ 1'b0 ;
  assign n483 = x69 & n157 ;
  assign n484 = ~x126 & n483 ;
  assign n485 = n482 | n484 ;
  assign n487 = n486 ^ n485 ^ 1'b0 ;
  assign n488 = ( n363 & ~n481 ) | ( n363 & n487 ) | ( ~n481 & n487 ) ;
  assign n491 = n405 ^ x41 ^ 1'b0 ;
  assign n492 = n491 ^ n261 ^ n221 ;
  assign n490 = n400 ^ n303 ^ n227 ;
  assign n493 = n492 ^ n490 ^ n282 ;
  assign n489 = n263 & ~n352 ;
  assign n494 = n493 ^ n489 ^ 1'b0 ;
  assign n495 = n494 ^ n237 ^ n206 ;
  assign n496 = n495 ^ n339 ^ n293 ;
  assign n501 = n131 & ~n132 ;
  assign n502 = ~x111 & n501 ;
  assign n497 = ( x19 & x44 ) | ( x19 & ~x70 ) | ( x44 & ~x70 ) ;
  assign n498 = ( x107 & n260 ) | ( x107 & ~n497 ) | ( n260 & ~n497 ) ;
  assign n499 = ( n184 & n440 ) | ( n184 & n498 ) | ( n440 & n498 ) ;
  assign n500 = ( n169 & ~n252 ) | ( n169 & n499 ) | ( ~n252 & n499 ) ;
  assign n503 = n502 ^ n500 ^ n401 ;
  assign n507 = ( x53 & n174 ) | ( x53 & n314 ) | ( n174 & n314 ) ;
  assign n506 = n439 ^ n194 ^ x68 ;
  assign n508 = n507 ^ n506 ^ x88 ;
  assign n509 = n508 ^ n160 ^ 1'b0 ;
  assign n510 = ~n400 & n509 ;
  assign n504 = ( x100 & n194 ) | ( x100 & ~n341 ) | ( n194 & ~n341 ) ;
  assign n505 = ~n155 & n504 ;
  assign n511 = n510 ^ n505 ^ 1'b0 ;
  assign n539 = n184 ^ n132 ^ 1'b0 ;
  assign n512 = ~n132 & n381 ;
  assign n513 = ( ~x27 & x48 ) | ( ~x27 & n507 ) | ( x48 & n507 ) ;
  assign n514 = ( x37 & n159 ) | ( x37 & ~n513 ) | ( n159 & ~n513 ) ;
  assign n515 = n514 ^ n130 ^ 1'b0 ;
  assign n516 = n512 & n515 ;
  assign n517 = n492 ^ n368 ^ x72 ;
  assign n518 = ( n445 & ~n516 ) | ( n445 & n517 ) | ( ~n516 & n517 ) ;
  assign n522 = n391 ^ n372 ^ x96 ;
  assign n523 = n522 ^ n391 ^ n258 ;
  assign n524 = n166 & n523 ;
  assign n519 = n138 ^ n133 ^ x47 ;
  assign n520 = x50 & n261 ;
  assign n521 = n519 & n520 ;
  assign n525 = n524 ^ n521 ^ n187 ;
  assign n533 = n219 & n437 ;
  assign n534 = ~n192 & n533 ;
  assign n530 = ( x34 & ~x107 ) | ( x34 & n462 ) | ( ~x107 & n462 ) ;
  assign n528 = ( x21 & n132 ) | ( x21 & n324 ) | ( n132 & n324 ) ;
  assign n529 = ( ~n319 & n475 ) | ( ~n319 & n528 ) | ( n475 & n528 ) ;
  assign n531 = n530 ^ n529 ^ 1'b0 ;
  assign n532 = ~n414 & n531 ;
  assign n526 = ( x23 & x117 ) | ( x23 & ~n197 ) | ( x117 & ~n197 ) ;
  assign n527 = n526 ^ n297 ^ x93 ;
  assign n535 = n534 ^ n532 ^ n527 ;
  assign n536 = ( x11 & ~n525 ) | ( x11 & n535 ) | ( ~n525 & n535 ) ;
  assign n537 = ( n421 & ~n518 ) | ( n421 & n536 ) | ( ~n518 & n536 ) ;
  assign n538 = n382 & n537 ;
  assign n540 = n539 ^ n538 ^ 1'b0 ;
  assign n541 = n473 ^ x68 ^ x36 ;
  assign n542 = n541 ^ n319 ^ n164 ;
  assign n543 = x48 ^ x36 ^ x23 ;
  assign n544 = ( n383 & n462 ) | ( n383 & n543 ) | ( n462 & n543 ) ;
  assign n545 = n544 ^ n491 ^ n396 ;
  assign n546 = ( x66 & n542 ) | ( x66 & ~n545 ) | ( n542 & ~n545 ) ;
  assign n547 = ( x2 & x16 ) | ( x2 & ~n421 ) | ( x16 & ~n421 ) ;
  assign n548 = x65 & n477 ;
  assign n549 = ~n547 & n548 ;
  assign n550 = ( ~n144 & n379 ) | ( ~n144 & n549 ) | ( n379 & n549 ) ;
  assign n552 = n406 ^ n138 ^ x95 ;
  assign n551 = n403 ^ n201 ^ x30 ;
  assign n553 = n552 ^ n551 ^ 1'b0 ;
  assign n554 = ~n502 & n553 ;
  assign n556 = n289 ^ n172 ^ x106 ;
  assign n557 = n556 ^ n507 ^ n480 ;
  assign n555 = ( n161 & n246 ) | ( n161 & ~n375 ) | ( n246 & ~n375 ) ;
  assign n558 = n557 ^ n555 ^ x7 ;
  assign n572 = n364 ^ x100 ^ x53 ;
  assign n559 = n329 ^ n245 ^ x11 ;
  assign n560 = x71 ^ x51 ^ x41 ;
  assign n561 = n193 & ~n560 ;
  assign n562 = ~n312 & n561 ;
  assign n563 = n562 ^ x111 ^ x2 ;
  assign n564 = ( n524 & ~n559 ) | ( n524 & n563 ) | ( ~n559 & n563 ) ;
  assign n565 = n172 ^ n155 ^ x26 ;
  assign n566 = ( ~n256 & n479 ) | ( ~n256 & n565 ) | ( n479 & n565 ) ;
  assign n567 = n457 ^ n130 ^ x126 ;
  assign n568 = ~n134 & n567 ;
  assign n569 = ( n564 & ~n566 ) | ( n564 & n568 ) | ( ~n566 & n568 ) ;
  assign n570 = n569 ^ x2 ^ 1'b0 ;
  assign n571 = n305 | n570 ;
  assign n573 = n572 ^ n571 ^ n477 ;
  assign n579 = ( x62 & ~x102 ) | ( x62 & n241 ) | ( ~x102 & n241 ) ;
  assign n574 = ( x120 & n190 ) | ( x120 & ~n245 ) | ( n190 & ~n245 ) ;
  assign n575 = ( x111 & n326 ) | ( x111 & n574 ) | ( n326 & n574 ) ;
  assign n576 = n575 ^ n526 ^ x59 ;
  assign n577 = n576 ^ n417 ^ n372 ;
  assign n578 = ( x20 & ~x47 ) | ( x20 & n577 ) | ( ~x47 & n577 ) ;
  assign n580 = n579 ^ n578 ^ 1'b0 ;
  assign n581 = n557 ^ x65 ^ x34 ;
  assign n582 = n581 ^ n432 ^ n258 ;
  assign n583 = n582 ^ x16 ^ 1'b0 ;
  assign n589 = n255 ^ n168 ^ n157 ;
  assign n586 = x103 ^ x53 ^ 1'b0 ;
  assign n587 = ( n195 & n232 ) | ( n195 & ~n586 ) | ( n232 & ~n586 ) ;
  assign n584 = n343 ^ n277 ^ x112 ;
  assign n585 = ( n300 & n323 ) | ( n300 & ~n584 ) | ( n323 & ~n584 ) ;
  assign n588 = n587 ^ n585 ^ n565 ;
  assign n590 = n589 ^ n588 ^ 1'b0 ;
  assign n591 = x92 & n590 ;
  assign n593 = n134 ^ x115 ^ 1'b0 ;
  assign n594 = x62 & ~n593 ;
  assign n595 = ( x112 & n560 ) | ( x112 & ~n594 ) | ( n560 & ~n594 ) ;
  assign n596 = x127 & ~n595 ;
  assign n592 = ( x50 & ~x81 ) | ( x50 & x88 ) | ( ~x81 & x88 ) ;
  assign n597 = n596 ^ n592 ^ n145 ;
  assign n598 = x85 & n200 ;
  assign n599 = ~n597 & n598 ;
  assign n600 = n439 | n599 ;
  assign n601 = n591 | n600 ;
  assign n606 = ( x42 & x43 ) | ( x42 & n285 ) | ( x43 & n285 ) ;
  assign n607 = ( x12 & ~n207 ) | ( x12 & n606 ) | ( ~n207 & n606 ) ;
  assign n608 = ( x37 & ~n245 ) | ( x37 & n607 ) | ( ~n245 & n607 ) ;
  assign n605 = n213 ^ x61 ^ x38 ;
  assign n602 = ( ~n143 & n529 ) | ( ~n143 & n539 ) | ( n529 & n539 ) ;
  assign n603 = ( ~n342 & n555 ) | ( ~n342 & n602 ) | ( n555 & n602 ) ;
  assign n604 = n303 & n603 ;
  assign n609 = n608 ^ n605 ^ n604 ;
  assign n616 = n253 & n582 ;
  assign n610 = n592 ^ n423 ^ n154 ;
  assign n611 = ( x63 & x91 ) | ( x63 & ~n173 ) | ( x91 & ~n173 ) ;
  assign n612 = n474 ^ n263 ^ x47 ;
  assign n613 = n611 & ~n612 ;
  assign n614 = n613 ^ n321 ^ 1'b0 ;
  assign n615 = n610 | n614 ;
  assign n617 = n616 ^ n615 ^ 1'b0 ;
  assign n618 = n251 ^ x97 ^ 1'b0 ;
  assign n619 = x117 & n618 ;
  assign n620 = n619 ^ x107 ^ x96 ;
  assign n621 = n597 ^ n540 ^ 1'b0 ;
  assign n622 = ( x9 & n256 ) | ( x9 & n337 ) | ( n256 & n337 ) ;
  assign n623 = n437 & ~n622 ;
  assign n624 = n623 ^ n416 ^ x78 ;
  assign n625 = ( n620 & ~n621 ) | ( n620 & n624 ) | ( ~n621 & n624 ) ;
  assign n636 = ( x79 & n133 ) | ( x79 & ~n165 ) | ( n133 & ~n165 ) ;
  assign n637 = ( n607 & n611 ) | ( n607 & n636 ) | ( n611 & n636 ) ;
  assign n638 = n637 ^ n313 ^ 1'b0 ;
  assign n634 = n312 ^ n289 ^ x67 ;
  assign n632 = ( x32 & n144 ) | ( x32 & ~n256 ) | ( n144 & ~n256 ) ;
  assign n633 = ( n544 & ~n567 ) | ( n544 & n632 ) | ( ~n567 & n632 ) ;
  assign n635 = n634 ^ n633 ^ x20 ;
  assign n630 = x64 ^ x55 ^ 1'b0 ;
  assign n626 = ( x80 & ~n204 ) | ( x80 & n346 ) | ( ~n204 & n346 ) ;
  assign n627 = ( n330 & n582 ) | ( n330 & n626 ) | ( n582 & n626 ) ;
  assign n628 = n356 & n627 ;
  assign n629 = ( ~n211 & n260 ) | ( ~n211 & n628 ) | ( n260 & n628 ) ;
  assign n631 = n630 ^ n629 ^ n210 ;
  assign n639 = n638 ^ n635 ^ n631 ;
  assign n640 = x82 ^ x56 ^ x1 ;
  assign n641 = n640 ^ n479 ^ x67 ;
  assign n642 = ( x107 & n322 ) | ( x107 & n484 ) | ( n322 & n484 ) ;
  assign n643 = ( ~x78 & n641 ) | ( ~x78 & n642 ) | ( n641 & n642 ) ;
  assign n646 = ( ~x75 & n135 ) | ( ~x75 & n457 ) | ( n135 & n457 ) ;
  assign n644 = n528 ^ n210 ^ x22 ;
  assign n645 = n644 ^ n290 ^ n268 ;
  assign n647 = n646 ^ n645 ^ n544 ;
  assign n648 = ( n202 & ~n596 ) | ( n202 & n646 ) | ( ~n596 & n646 ) ;
  assign n649 = ( ~n643 & n647 ) | ( ~n643 & n648 ) | ( n647 & n648 ) ;
  assign n656 = n592 ^ n206 ^ x111 ;
  assign n650 = n173 ^ n129 ^ 1'b0 ;
  assign n651 = n650 ^ n295 ^ n282 ;
  assign n652 = n278 ^ n235 ^ 1'b0 ;
  assign n653 = n651 & n652 ;
  assign n654 = x58 & n653 ;
  assign n655 = n654 ^ n248 ^ 1'b0 ;
  assign n657 = n656 ^ n655 ^ n512 ;
  assign n658 = n386 ^ n245 ^ x61 ;
  assign n659 = n658 ^ n575 ^ x110 ;
  assign n660 = n659 ^ n213 ^ n176 ;
  assign n661 = ( x102 & ~n446 ) | ( x102 & n660 ) | ( ~n446 & n660 ) ;
  assign n663 = n325 ^ n224 ^ 1'b0 ;
  assign n664 = n288 | n663 ;
  assign n662 = ( x56 & n318 ) | ( x56 & n383 ) | ( n318 & n383 ) ;
  assign n665 = n664 ^ n662 ^ n273 ;
  assign n666 = n665 ^ n637 ^ x32 ;
  assign n667 = n572 & n666 ;
  assign n668 = n667 ^ x113 ^ 1'b0 ;
  assign n669 = n530 ^ n209 ^ x123 ;
  assign n670 = ~n265 & n669 ;
  assign n673 = n498 ^ n462 ^ n318 ;
  assign n671 = n288 ^ n164 ^ x117 ;
  assign n672 = n502 | n671 ;
  assign n674 = n673 ^ n672 ^ 1'b0 ;
  assign n675 = n674 ^ n637 ^ 1'b0 ;
  assign n676 = n368 & ~n675 ;
  assign n677 = x80 & ~n676 ;
  assign n678 = ( n447 & n670 ) | ( n447 & n677 ) | ( n670 & n677 ) ;
  assign n679 = n474 ^ n437 ^ n161 ;
  assign n680 = ( n192 & n478 ) | ( n192 & n679 ) | ( n478 & n679 ) ;
  assign n681 = n680 ^ n525 ^ x57 ;
  assign n698 = x12 & ~n507 ;
  assign n686 = ( x96 & ~n201 ) | ( x96 & n534 ) | ( ~n201 & n534 ) ;
  assign n684 = ~x8 & n356 ;
  assign n682 = x106 & n646 ;
  assign n683 = n409 & n682 ;
  assign n685 = n684 ^ n683 ^ 1'b0 ;
  assign n687 = n686 ^ n685 ^ x12 ;
  assign n688 = n223 ^ x108 ^ 1'b0 ;
  assign n689 = ( ~n189 & n594 ) | ( ~n189 & n688 ) | ( n594 & n688 ) ;
  assign n691 = n463 ^ n391 ^ x85 ;
  assign n690 = ( x85 & ~n364 ) | ( x85 & n671 ) | ( ~n364 & n671 ) ;
  assign n692 = n691 ^ n690 ^ x116 ;
  assign n693 = n523 | n692 ;
  assign n694 = n581 & ~n693 ;
  assign n695 = n689 & ~n694 ;
  assign n696 = n587 & n695 ;
  assign n697 = ( n519 & n687 ) | ( n519 & ~n696 ) | ( n687 & ~n696 ) ;
  assign n699 = n698 ^ n697 ^ n444 ;
  assign n700 = n586 & n699 ;
  assign n701 = ( ~x15 & n191 ) | ( ~x15 & n291 ) | ( n191 & n291 ) ;
  assign n702 = n701 ^ n440 ^ x125 ;
  assign n705 = ( ~x42 & x56 ) | ( ~x42 & x107 ) | ( x56 & x107 ) ;
  assign n703 = n640 ^ n150 ^ x112 ;
  assign n704 = n703 ^ n459 ^ x123 ;
  assign n706 = n705 ^ n704 ^ n463 ;
  assign n707 = ( x31 & ~n312 ) | ( x31 & n436 ) | ( ~n312 & n436 ) ;
  assign n708 = ( n478 & n636 ) | ( n478 & n707 ) | ( n636 & n707 ) ;
  assign n709 = ~n232 & n258 ;
  assign n710 = n516 ^ n285 ^ x106 ;
  assign n727 = n196 ^ x121 ^ x117 ;
  assign n728 = ( ~x71 & n314 ) | ( ~x71 & n727 ) | ( n314 & n727 ) ;
  assign n723 = ( x3 & x87 ) | ( x3 & n388 ) | ( x87 & n388 ) ;
  assign n724 = n723 ^ n148 ^ 1'b0 ;
  assign n725 = ~n285 & n724 ;
  assign n719 = n227 ^ n213 ^ x42 ;
  assign n720 = n719 ^ n223 ^ n218 ;
  assign n721 = n720 ^ x70 ^ x0 ;
  assign n722 = n721 ^ n503 ^ n265 ;
  assign n726 = n725 ^ n722 ^ x87 ;
  assign n717 = ( x30 & ~x44 ) | ( x30 & n439 ) | ( ~x44 & n439 ) ;
  assign n716 = ( n210 & n352 ) | ( n210 & n486 ) | ( n352 & n486 ) ;
  assign n711 = x25 | n172 ;
  assign n712 = x64 & ~n482 ;
  assign n713 = n712 ^ x70 ^ 1'b0 ;
  assign n714 = ( x17 & n491 ) | ( x17 & n713 ) | ( n491 & n713 ) ;
  assign n715 = ( n641 & n711 ) | ( n641 & n714 ) | ( n711 & n714 ) ;
  assign n718 = n717 ^ n716 ^ n715 ;
  assign n729 = n728 ^ n726 ^ n718 ;
  assign n730 = ( ~n709 & n710 ) | ( ~n709 & n729 ) | ( n710 & n729 ) ;
  assign n734 = n482 ^ x113 ^ x30 ;
  assign n733 = n662 ^ n325 ^ 1'b0 ;
  assign n731 = ( x89 & n259 ) | ( x89 & ~n688 ) | ( n259 & ~n688 ) ;
  assign n732 = ( n206 & n245 ) | ( n206 & n731 ) | ( n245 & n731 ) ;
  assign n735 = n734 ^ n733 ^ n732 ;
  assign n736 = n335 & n428 ;
  assign n737 = n205 ^ n198 ^ n131 ;
  assign n738 = ( x24 & x87 ) | ( x24 & n266 ) | ( x87 & n266 ) ;
  assign n739 = n304 ^ x69 ^ 1'b0 ;
  assign n740 = n319 ^ n165 ^ x25 ;
  assign n741 = n740 ^ n470 ^ x17 ;
  assign n742 = ( n738 & n739 ) | ( n738 & n741 ) | ( n739 & n741 ) ;
  assign n743 = ( n364 & n737 ) | ( n364 & n742 ) | ( n737 & n742 ) ;
  assign n744 = n322 ^ n283 ^ x7 ;
  assign n745 = ( n438 & n581 ) | ( n438 & ~n744 ) | ( n581 & ~n744 ) ;
  assign n746 = ( n736 & ~n743 ) | ( n736 & n745 ) | ( ~n743 & n745 ) ;
  assign n747 = ( x32 & ~n280 ) | ( x32 & n713 ) | ( ~n280 & n713 ) ;
  assign n748 = ( n264 & ~n460 ) | ( n264 & n747 ) | ( ~n460 & n747 ) ;
  assign n749 = n611 ^ n146 ^ n134 ;
  assign n750 = ( n325 & n586 ) | ( n325 & n749 ) | ( n586 & n749 ) ;
  assign n751 = n750 ^ n504 ^ 1'b0 ;
  assign n752 = n500 ^ n284 ^ x121 ;
  assign n753 = ( n256 & n478 ) | ( n256 & ~n752 ) | ( n478 & ~n752 ) ;
  assign n754 = ( n154 & n734 ) | ( n154 & n753 ) | ( n734 & n753 ) ;
  assign n755 = ( x80 & n138 ) | ( x80 & n139 ) | ( n138 & n139 ) ;
  assign n756 = x3 & ~n755 ;
  assign n757 = ( n328 & ~n461 ) | ( n328 & n756 ) | ( ~n461 & n756 ) ;
  assign n758 = n757 ^ n666 ^ 1'b0 ;
  assign n779 = x112 & n252 ;
  assign n778 = n720 ^ n391 ^ x79 ;
  assign n780 = n779 ^ n778 ^ x57 ;
  assign n762 = ( x30 & n194 ) | ( x30 & n355 ) | ( n194 & n355 ) ;
  assign n763 = ~n288 & n530 ;
  assign n764 = n763 ^ n222 ^ 1'b0 ;
  assign n765 = n764 ^ n301 ^ x59 ;
  assign n766 = n762 & n765 ;
  assign n767 = n766 ^ x10 ^ 1'b0 ;
  assign n770 = x16 ^ x10 ^ 1'b0 ;
  assign n771 = n296 & n770 ;
  assign n768 = n644 ^ n288 ^ n280 ;
  assign n769 = n768 ^ n588 ^ n300 ;
  assign n772 = n771 ^ n769 ^ x38 ;
  assign n773 = n448 ^ n239 ^ 1'b0 ;
  assign n774 = n773 ^ n641 ^ n610 ;
  assign n775 = ( ~n767 & n772 ) | ( ~n767 & n774 ) | ( n772 & n774 ) ;
  assign n776 = ~n285 & n775 ;
  assign n777 = n776 ^ n355 ^ 1'b0 ;
  assign n759 = x87 & n479 ;
  assign n760 = n759 ^ n565 ^ n444 ;
  assign n761 = ( n303 & n596 ) | ( n303 & n760 ) | ( n596 & n760 ) ;
  assign n781 = n780 ^ n777 ^ n761 ;
  assign n782 = n556 ^ x23 ^ 1'b0 ;
  assign n784 = ( x105 & x110 ) | ( x105 & n660 ) | ( x110 & n660 ) ;
  assign n783 = n204 ^ n198 ^ 1'b0 ;
  assign n785 = n784 ^ n783 ^ n353 ;
  assign n786 = n785 ^ n722 ^ 1'b0 ;
  assign n787 = x21 & n786 ;
  assign n788 = ( n387 & n782 ) | ( n387 & n787 ) | ( n782 & n787 ) ;
  assign n789 = ( ~x15 & x43 ) | ( ~x15 & n637 ) | ( x43 & n637 ) ;
  assign n790 = ( ~x99 & x124 ) | ( ~x99 & n557 ) | ( x124 & n557 ) ;
  assign n791 = ( n211 & ~n353 ) | ( n211 & n736 ) | ( ~n353 & n736 ) ;
  assign n792 = n791 ^ n716 ^ n359 ;
  assign n793 = ( ~n684 & n790 ) | ( ~n684 & n792 ) | ( n790 & n792 ) ;
  assign n794 = ( x34 & n789 ) | ( x34 & ~n793 ) | ( n789 & ~n793 ) ;
  assign n795 = ~n453 & n689 ;
  assign n796 = n781 ^ n416 ^ n304 ;
  assign n797 = n606 ^ n369 ^ x0 ;
  assign n798 = ( x36 & n291 ) | ( x36 & ~n797 ) | ( n291 & ~n797 ) ;
  assign n799 = n739 ^ n620 ^ n139 ;
  assign n800 = ( n312 & n798 ) | ( n312 & ~n799 ) | ( n798 & ~n799 ) ;
  assign n801 = n504 ^ n421 ^ n312 ;
  assign n802 = n775 & ~n801 ;
  assign n803 = n800 & n802 ;
  assign n822 = n317 ^ x123 ^ x53 ;
  assign n823 = n822 ^ n168 ^ 1'b0 ;
  assign n824 = n823 ^ n272 ^ x9 ;
  assign n833 = n387 | n502 ;
  assign n825 = ( x47 & ~x49 ) | ( x47 & x50 ) | ( ~x49 & x50 ) ;
  assign n827 = ( ~n173 & n493 ) | ( ~n173 & n556 ) | ( n493 & n556 ) ;
  assign n828 = x97 & ~n827 ;
  assign n829 = n828 ^ n352 ^ 1'b0 ;
  assign n826 = ( x97 & ~x118 ) | ( x97 & n749 ) | ( ~x118 & n749 ) ;
  assign n830 = n829 ^ n826 ^ n771 ;
  assign n831 = n825 & n830 ;
  assign n832 = n831 ^ n178 ^ 1'b0 ;
  assign n834 = n833 ^ n832 ^ n243 ;
  assign n835 = ( n783 & n824 ) | ( n783 & n834 ) | ( n824 & n834 ) ;
  assign n818 = ( n228 & ~n292 ) | ( n228 & n484 ) | ( ~n292 & n484 ) ;
  assign n806 = ( x80 & x92 ) | ( x80 & ~n530 ) | ( x92 & ~n530 ) ;
  assign n812 = n148 ^ x38 ^ x23 ;
  assign n813 = x78 & ~n812 ;
  assign n814 = ~n806 & n813 ;
  assign n815 = ( ~x6 & n607 ) | ( ~x6 & n814 ) | ( n607 & n814 ) ;
  assign n810 = n688 ^ n560 ^ x70 ;
  assign n811 = n810 ^ n601 ^ n423 ;
  assign n816 = n815 ^ n811 ^ 1'b0 ;
  assign n807 = n806 ^ x63 ^ x54 ;
  assign n804 = ( n197 & ~n242 ) | ( n197 & n653 ) | ( ~n242 & n653 ) ;
  assign n805 = ( n307 & n784 ) | ( n307 & ~n804 ) | ( n784 & ~n804 ) ;
  assign n808 = n807 ^ n805 ^ 1'b0 ;
  assign n809 = n716 | n808 ;
  assign n817 = n816 ^ n809 ^ n390 ;
  assign n819 = n818 ^ n817 ^ n360 ;
  assign n820 = n819 ^ n399 ^ 1'b0 ;
  assign n821 = ~n673 & n820 ;
  assign n836 = n835 ^ n821 ^ x77 ;
  assign n837 = ( x15 & x23 ) | ( x15 & ~n175 ) | ( x23 & ~n175 ) ;
  assign n838 = n837 ^ n284 ^ x72 ;
  assign n839 = n838 ^ n419 ^ n132 ;
  assign n840 = n839 ^ n416 ^ n376 ;
  assign n845 = n688 ^ n499 ^ n341 ;
  assign n841 = n259 ^ n230 ^ n171 ;
  assign n842 = n220 ^ x24 ^ 1'b0 ;
  assign n843 = n841 & n842 ;
  assign n844 = n843 ^ n643 ^ n194 ;
  assign n846 = n845 ^ n844 ^ 1'b0 ;
  assign n847 = ~n840 & n846 ;
  assign n848 = n847 ^ n415 ^ n336 ;
  assign n850 = ( x12 & ~n343 ) | ( x12 & n469 ) | ( ~n343 & n469 ) ;
  assign n849 = n604 & n703 ;
  assign n851 = n850 ^ n849 ^ 1'b0 ;
  assign n853 = n329 ^ x66 ^ x45 ;
  assign n854 = n853 ^ n714 ^ n392 ;
  assign n855 = ( n223 & n691 ) | ( n223 & ~n854 ) | ( n691 & ~n854 ) ;
  assign n852 = n811 ^ n169 ^ 1'b0 ;
  assign n856 = n855 ^ n852 ^ x90 ;
  assign n857 = n830 ^ n599 ^ n372 ;
  assign n858 = n549 & ~n768 ;
  assign n859 = ( x9 & ~n857 ) | ( x9 & n858 ) | ( ~n857 & n858 ) ;
  assign n860 = ( n298 & ~n653 ) | ( n298 & n859 ) | ( ~n653 & n859 ) ;
  assign n861 = ( ~n238 & n474 ) | ( ~n238 & n860 ) | ( n474 & n860 ) ;
  assign n862 = x107 & ~n355 ;
  assign n863 = ~n201 & n862 ;
  assign n864 = ( x37 & n188 ) | ( x37 & ~n810 ) | ( n188 & ~n810 ) ;
  assign n865 = ( x7 & n863 ) | ( x7 & n864 ) | ( n863 & n864 ) ;
  assign n874 = ( x121 & n203 ) | ( x121 & ~n259 ) | ( n203 & ~n259 ) ;
  assign n878 = n619 ^ n480 ^ n240 ;
  assign n875 = n830 ^ n487 ^ 1'b0 ;
  assign n876 = n875 ^ n309 ^ x54 ;
  assign n877 = ( x88 & n372 ) | ( x88 & n876 ) | ( n372 & n876 ) ;
  assign n879 = n878 ^ n877 ^ x99 ;
  assign n880 = ( ~x94 & n589 ) | ( ~x94 & n759 ) | ( n589 & n759 ) ;
  assign n881 = ( n874 & n879 ) | ( n874 & n880 ) | ( n879 & n880 ) ;
  assign n866 = x43 & ~n199 ;
  assign n867 = n866 ^ n216 ^ 1'b0 ;
  assign n870 = n324 ^ n147 ^ x95 ;
  assign n868 = n559 ^ n254 ^ n250 ;
  assign n869 = n225 | n868 ;
  assign n871 = n870 ^ n869 ^ 1'b0 ;
  assign n872 = ( n292 & n867 ) | ( n292 & ~n871 ) | ( n867 & ~n871 ) ;
  assign n873 = ( x36 & ~n435 ) | ( x36 & n872 ) | ( ~n435 & n872 ) ;
  assign n882 = n881 ^ n873 ^ n521 ;
  assign n883 = n882 ^ n518 ^ 1'b0 ;
  assign n886 = n362 ^ n229 ^ 1'b0 ;
  assign n887 = n401 | n886 ;
  assign n888 = n887 ^ n198 ^ 1'b0 ;
  assign n889 = n888 ^ n359 ^ x64 ;
  assign n884 = n602 ^ n387 ^ n307 ;
  assign n885 = n439 | n884 ;
  assign n890 = n889 ^ n885 ^ x76 ;
  assign n891 = n479 ^ n206 ^ n154 ;
  assign n892 = n227 & n891 ;
  assign n893 = n892 ^ n771 ^ 1'b0 ;
  assign n894 = ~n645 & n893 ;
  assign n895 = ( ~n539 & n890 ) | ( ~n539 & n894 ) | ( n890 & n894 ) ;
  assign n896 = n895 ^ n804 ^ n704 ;
  assign n897 = n565 ^ n368 ^ 1'b0 ;
  assign n898 = n897 ^ n288 ^ x59 ;
  assign n899 = n898 ^ n375 ^ 1'b0 ;
  assign n900 = n896 & n899 ;
  assign n902 = x16 & n406 ;
  assign n903 = ~x74 & n902 ;
  assign n904 = ( ~x60 & x90 ) | ( ~x60 & n160 ) | ( x90 & n160 ) ;
  assign n905 = ( x120 & n373 ) | ( x120 & n904 ) | ( n373 & n904 ) ;
  assign n906 = ( n220 & n903 ) | ( n220 & ~n905 ) | ( n903 & ~n905 ) ;
  assign n901 = n879 ^ n709 ^ n218 ;
  assign n907 = n906 ^ n901 ^ n641 ;
  assign n908 = ( ~n452 & n692 ) | ( ~n452 & n762 ) | ( n692 & n762 ) ;
  assign n909 = ( n536 & n661 ) | ( n536 & n908 ) | ( n661 & n908 ) ;
  assign n920 = n894 ^ n722 ^ n267 ;
  assign n916 = n246 ^ x84 ^ 1'b0 ;
  assign n917 = x106 & n916 ;
  assign n918 = n917 ^ n574 ^ n257 ;
  assign n919 = n312 & ~n918 ;
  assign n921 = n920 ^ n919 ^ 1'b0 ;
  assign n913 = n186 ^ x18 ^ 1'b0 ;
  assign n914 = ( x20 & ~n841 ) | ( x20 & n913 ) | ( ~n841 & n913 ) ;
  assign n910 = ( x7 & ~n380 ) | ( x7 & n478 ) | ( ~n380 & n478 ) ;
  assign n911 = n321 & n910 ;
  assign n912 = ~n384 & n911 ;
  assign n915 = n914 ^ n912 ^ x96 ;
  assign n922 = n921 ^ n915 ^ n394 ;
  assign n928 = n572 ^ n250 ^ 1'b0 ;
  assign n929 = n281 & n928 ;
  assign n923 = ( x38 & n204 ) | ( x38 & n579 ) | ( n204 & n579 ) ;
  assign n924 = n438 ^ x28 ^ 1'b0 ;
  assign n925 = n555 & n924 ;
  assign n926 = ~n175 & n925 ;
  assign n927 = ( n139 & ~n923 ) | ( n139 & n926 ) | ( ~n923 & n926 ) ;
  assign n930 = n929 ^ n927 ^ n668 ;
  assign n939 = ( ~n460 & n762 ) | ( ~n460 & n887 ) | ( n762 & n887 ) ;
  assign n937 = ( ~n205 & n822 ) | ( ~n205 & n914 ) | ( n822 & n914 ) ;
  assign n932 = n471 ^ n188 ^ x41 ;
  assign n933 = n932 ^ n645 ^ n335 ;
  assign n934 = n737 ^ n438 ^ n401 ;
  assign n935 = n587 | n934 ;
  assign n936 = n933 & ~n935 ;
  assign n931 = n146 ^ x85 ^ 1'b0 ;
  assign n938 = n937 ^ n936 ^ n931 ;
  assign n940 = n939 ^ n938 ^ n734 ;
  assign n941 = n401 ^ n218 ^ x6 ;
  assign n961 = n825 ^ n309 ^ n201 ;
  assign n960 = n790 ^ n356 ^ n314 ;
  assign n962 = n961 ^ n960 ^ n196 ;
  assign n963 = ( x35 & ~n210 ) | ( x35 & n744 ) | ( ~n210 & n744 ) ;
  assign n964 = ( n454 & n962 ) | ( n454 & ~n963 ) | ( n962 & ~n963 ) ;
  assign n947 = n837 ^ x75 ^ x18 ;
  assign n944 = ( x34 & ~x85 ) | ( x34 & x95 ) | ( ~x85 & x95 ) ;
  assign n945 = n944 ^ n280 ^ n226 ;
  assign n946 = ( n151 & ~n662 ) | ( n151 & n945 ) | ( ~n662 & n945 ) ;
  assign n948 = n947 ^ n946 ^ n449 ;
  assign n953 = n606 ^ n560 ^ n302 ;
  assign n951 = n903 ^ n247 ^ x93 ;
  assign n952 = ( n218 & n692 ) | ( n218 & n951 ) | ( n692 & n951 ) ;
  assign n949 = n323 | n385 ;
  assign n950 = ( n727 & ~n945 ) | ( n727 & n949 ) | ( ~n945 & n949 ) ;
  assign n954 = n953 ^ n952 ^ n950 ;
  assign n955 = ( n201 & n391 ) | ( n201 & n574 ) | ( n391 & n574 ) ;
  assign n956 = ( x18 & ~x47 ) | ( x18 & n955 ) | ( ~x47 & n955 ) ;
  assign n957 = n956 ^ n490 ^ n376 ;
  assign n958 = ( n229 & n954 ) | ( n229 & ~n957 ) | ( n954 & ~n957 ) ;
  assign n959 = ( n648 & ~n948 ) | ( n648 & n958 ) | ( ~n948 & n958 ) ;
  assign n942 = n438 ^ n370 ^ x72 ;
  assign n943 = ( ~n242 & n934 ) | ( ~n242 & n942 ) | ( n934 & n942 ) ;
  assign n965 = n964 ^ n959 ^ n943 ;
  assign n966 = n400 ^ x32 ^ 1'b0 ;
  assign n977 = ( ~n212 & n274 ) | ( ~n212 & n646 ) | ( n274 & n646 ) ;
  assign n967 = n760 ^ n213 ^ n204 ;
  assign n968 = n967 ^ n614 ^ n336 ;
  assign n969 = n889 ^ n270 ^ n201 ;
  assign n970 = n713 | n913 ;
  assign n971 = n192 | n970 ;
  assign n972 = n971 ^ n305 ^ n221 ;
  assign n973 = n972 ^ n246 ^ 1'b0 ;
  assign n974 = ( ~n826 & n969 ) | ( ~n826 & n973 ) | ( n969 & n973 ) ;
  assign n975 = n974 ^ n954 ^ x72 ;
  assign n976 = n968 | n975 ;
  assign n978 = n977 ^ n976 ^ 1'b0 ;
  assign n989 = ( n210 & n214 ) | ( n210 & n565 ) | ( n214 & n565 ) ;
  assign n990 = x97 & n989 ;
  assign n986 = n971 ^ n740 ^ 1'b0 ;
  assign n985 = ( ~x49 & x120 ) | ( ~x49 & n674 ) | ( x120 & n674 ) ;
  assign n987 = n986 ^ n985 ^ 1'b0 ;
  assign n982 = ( n221 & n233 ) | ( n221 & ~n268 ) | ( n233 & ~n268 ) ;
  assign n983 = n982 ^ n680 ^ n479 ;
  assign n979 = n171 & ~n642 ;
  assign n980 = ~n296 & n979 ;
  assign n981 = n980 ^ n833 ^ n504 ;
  assign n984 = n983 ^ n981 ^ n474 ;
  assign n988 = n987 ^ n984 ^ n741 ;
  assign n991 = n990 ^ n988 ^ n683 ;
  assign n992 = ( x25 & n362 ) | ( x25 & n644 ) | ( n362 & n644 ) ;
  assign n993 = ( ~n630 & n917 ) | ( ~n630 & n992 ) | ( n917 & n992 ) ;
  assign n994 = n272 ^ x127 ^ x38 ;
  assign n995 = ( n642 & ~n727 ) | ( n642 & n994 ) | ( ~n727 & n994 ) ;
  assign n996 = ( n332 & ~n993 ) | ( n332 & n995 ) | ( ~n993 & n995 ) ;
  assign n997 = ( x92 & n351 ) | ( x92 & n996 ) | ( n351 & n996 ) ;
  assign n1005 = ~n260 & n494 ;
  assign n1006 = ~n377 & n1005 ;
  assign n1007 = n1006 ^ n197 ^ 1'b0 ;
  assign n1008 = n225 | n1007 ;
  assign n1009 = ( n277 & n674 ) | ( n277 & n1008 ) | ( n674 & n1008 ) ;
  assign n998 = n651 ^ n365 ^ 1'b0 ;
  assign n999 = n296 & ~n998 ;
  assign n1000 = n477 & n999 ;
  assign n1001 = ~n138 & n473 ;
  assign n1002 = n1001 ^ n487 ^ 1'b0 ;
  assign n1003 = ( n263 & n961 ) | ( n263 & ~n1002 ) | ( n961 & ~n1002 ) ;
  assign n1004 = ( ~n832 & n1000 ) | ( ~n832 & n1003 ) | ( n1000 & n1003 ) ;
  assign n1010 = n1009 ^ n1004 ^ n161 ;
  assign n1021 = n421 ^ x69 ^ x36 ;
  assign n1022 = n1021 ^ n187 ^ x125 ;
  assign n1011 = n260 ^ n165 ^ 1'b0 ;
  assign n1012 = n224 | n1011 ;
  assign n1013 = ( ~x108 & n129 ) | ( ~x108 & n528 ) | ( n129 & n528 ) ;
  assign n1014 = ( n579 & n992 ) | ( n579 & n1013 ) | ( n992 & n1013 ) ;
  assign n1015 = ( ~n792 & n1012 ) | ( ~n792 & n1014 ) | ( n1012 & n1014 ) ;
  assign n1016 = n1015 ^ n742 ^ n345 ;
  assign n1017 = ( ~x101 & n430 ) | ( ~x101 & n1016 ) | ( n430 & n1016 ) ;
  assign n1018 = ( ~x43 & n160 ) | ( ~x43 & n367 ) | ( n160 & n367 ) ;
  assign n1019 = n1018 ^ n437 ^ 1'b0 ;
  assign n1020 = n1017 | n1019 ;
  assign n1023 = n1022 ^ n1020 ^ 1'b0 ;
  assign n1024 = n994 ^ n209 ^ x35 ;
  assign n1029 = ( x88 & ~n302 ) | ( x88 & n381 ) | ( ~n302 & n381 ) ;
  assign n1030 = n1029 ^ n281 ^ x72 ;
  assign n1028 = ( n235 & ~n440 ) | ( n235 & n683 ) | ( ~n440 & n683 ) ;
  assign n1025 = x2 & ~n458 ;
  assign n1026 = n1025 ^ n969 ^ 1'b0 ;
  assign n1027 = n1026 ^ n616 ^ n492 ;
  assign n1031 = n1030 ^ n1028 ^ n1027 ;
  assign n1032 = ( n875 & ~n1024 ) | ( n875 & n1031 ) | ( ~n1024 & n1031 ) ;
  assign n1033 = x50 | n493 ;
  assign n1036 = ( n273 & ~n340 ) | ( n273 & n709 ) | ( ~n340 & n709 ) ;
  assign n1035 = n563 ^ n504 ^ n405 ;
  assign n1037 = n1036 ^ n1035 ^ n942 ;
  assign n1038 = n1037 ^ n755 ^ n736 ;
  assign n1034 = n894 ^ n287 ^ 1'b0 ;
  assign n1039 = n1038 ^ n1034 ^ n853 ;
  assign n1043 = ( x0 & ~n233 ) | ( x0 & n251 ) | ( ~n233 & n251 ) ;
  assign n1044 = ( x23 & ~n405 ) | ( x23 & n452 ) | ( ~n405 & n452 ) ;
  assign n1045 = n895 ^ n637 ^ n272 ;
  assign n1046 = ( ~n1043 & n1044 ) | ( ~n1043 & n1045 ) | ( n1044 & n1045 ) ;
  assign n1047 = ( n150 & n313 ) | ( n150 & n1046 ) | ( n313 & n1046 ) ;
  assign n1040 = ~n199 & n542 ;
  assign n1041 = n1040 ^ n634 ^ 1'b0 ;
  assign n1042 = n1041 ^ n537 ^ n536 ;
  assign n1048 = n1047 ^ n1042 ^ n189 ;
  assign n1049 = ( n1033 & n1039 ) | ( n1033 & ~n1048 ) | ( n1039 & ~n1048 ) ;
  assign n1050 = ( n225 & n289 ) | ( n225 & ~n549 ) | ( n289 & ~n549 ) ;
  assign n1051 = x76 & n1050 ;
  assign n1052 = n1051 ^ n715 ^ 1'b0 ;
  assign n1053 = ( n287 & n428 ) | ( n287 & ~n1052 ) | ( n428 & ~n1052 ) ;
  assign n1059 = ( n508 & n562 ) | ( n508 & ~n961 ) | ( n562 & ~n961 ) ;
  assign n1054 = ~n144 & n218 ;
  assign n1055 = n1054 ^ x88 ^ 1'b0 ;
  assign n1056 = n1055 ^ n502 ^ x5 ;
  assign n1057 = ( ~n423 & n962 ) | ( ~n423 & n1056 ) | ( n962 & n1056 ) ;
  assign n1058 = x108 & ~n1057 ;
  assign n1060 = n1059 ^ n1058 ^ 1'b0 ;
  assign n1061 = n469 ^ n347 ^ x18 ;
  assign n1062 = n690 ^ n344 ^ n170 ;
  assign n1063 = ( x113 & ~n1061 ) | ( x113 & n1062 ) | ( ~n1061 & n1062 ) ;
  assign n1065 = ( n190 & ~n242 ) | ( n190 & n341 ) | ( ~n242 & n341 ) ;
  assign n1066 = x56 & n1065 ;
  assign n1067 = n1066 ^ x113 ^ 1'b0 ;
  assign n1064 = n577 ^ n191 ^ x21 ;
  assign n1068 = n1067 ^ n1064 ^ n963 ;
  assign n1069 = n429 & ~n1068 ;
  assign n1070 = ( n857 & n1063 ) | ( n857 & n1069 ) | ( n1063 & n1069 ) ;
  assign n1075 = ( x124 & ~n392 ) | ( x124 & n401 ) | ( ~n392 & n401 ) ;
  assign n1073 = x5 & n335 ;
  assign n1074 = ~x124 & n1073 ;
  assign n1071 = n423 ^ n129 ^ 1'b0 ;
  assign n1072 = n563 & ~n1071 ;
  assign n1076 = n1075 ^ n1074 ^ n1072 ;
  assign n1085 = n980 ^ n312 ^ x118 ;
  assign n1081 = ( x57 & n265 ) | ( x57 & ~n673 ) | ( n265 & ~n673 ) ;
  assign n1082 = ~n484 & n1081 ;
  assign n1083 = n1082 ^ n797 ^ 1'b0 ;
  assign n1077 = n1018 ^ n698 ^ x1 ;
  assign n1078 = n875 | n1077 ;
  assign n1079 = n737 & ~n1078 ;
  assign n1080 = ( n475 & ~n559 ) | ( n475 & n1079 ) | ( ~n559 & n1079 ) ;
  assign n1084 = n1083 ^ n1080 ^ 1'b0 ;
  assign n1086 = n1085 ^ n1084 ^ n777 ;
  assign n1087 = ( n291 & ~n404 ) | ( n291 & n734 ) | ( ~n404 & n734 ) ;
  assign n1088 = ( n477 & ~n1044 ) | ( n477 & n1087 ) | ( ~n1044 & n1087 ) ;
  assign n1089 = ( n959 & ~n1081 ) | ( n959 & n1088 ) | ( ~n1081 & n1088 ) ;
  assign n1090 = n244 ^ x68 ^ x13 ;
  assign n1093 = ( x94 & n331 ) | ( x94 & ~n999 ) | ( n331 & ~n999 ) ;
  assign n1091 = n719 ^ n383 ^ x67 ;
  assign n1092 = ~n519 & n1091 ;
  assign n1094 = n1093 ^ n1092 ^ 1'b0 ;
  assign n1095 = n1094 ^ n224 ^ 1'b0 ;
  assign n1096 = ~n1090 & n1095 ;
  assign n1097 = n1096 ^ n404 ^ 1'b0 ;
  assign n1098 = n297 & n589 ;
  assign n1111 = x0 & x20 ;
  assign n1112 = n1111 ^ n142 ^ 1'b0 ;
  assign n1113 = n443 ^ n375 ^ n222 ;
  assign n1114 = n878 ^ n549 ^ n336 ;
  assign n1115 = ( n854 & ~n1113 ) | ( n854 & n1114 ) | ( ~n1113 & n1114 ) ;
  assign n1116 = ( n756 & ~n1112 ) | ( n756 & n1115 ) | ( ~n1112 & n1115 ) ;
  assign n1117 = n1116 ^ n933 ^ 1'b0 ;
  assign n1118 = ~n1003 & n1117 ;
  assign n1104 = ( x100 & ~n203 ) | ( x100 & n271 ) | ( ~n203 & n271 ) ;
  assign n1105 = n1104 ^ n585 ^ n226 ;
  assign n1106 = ( n138 & n193 ) | ( n138 & ~n715 ) | ( n193 & ~n715 ) ;
  assign n1107 = n321 & n449 ;
  assign n1108 = n1106 & n1107 ;
  assign n1109 = n1105 & ~n1108 ;
  assign n1099 = n315 ^ n291 ^ n272 ;
  assign n1100 = n1099 ^ n481 ^ n403 ;
  assign n1101 = ~n696 & n1100 ;
  assign n1102 = n1101 ^ n301 ^ 1'b0 ;
  assign n1103 = n1102 ^ n642 ^ n586 ;
  assign n1110 = n1109 ^ n1103 ^ n610 ;
  assign n1119 = n1118 ^ n1110 ^ n253 ;
  assign n1120 = ( ~n559 & n1098 ) | ( ~n559 & n1119 ) | ( n1098 & n1119 ) ;
  assign n1121 = n738 ^ n405 ^ n206 ;
  assign n1122 = ( n204 & n801 ) | ( n204 & n1121 ) | ( n801 & n1121 ) ;
  assign n1123 = ( n414 & n563 ) | ( n414 & ~n659 ) | ( n563 & ~n659 ) ;
  assign n1127 = n478 ^ n359 ^ 1'b0 ;
  assign n1128 = n334 & n1127 ;
  assign n1126 = ( ~n439 & n771 ) | ( ~n439 & n801 ) | ( n771 & n801 ) ;
  assign n1124 = ( ~n196 & n337 ) | ( ~n196 & n594 ) | ( n337 & n594 ) ;
  assign n1125 = n1124 ^ n823 ^ n494 ;
  assign n1129 = n1128 ^ n1126 ^ n1125 ;
  assign n1130 = ( n265 & n545 ) | ( n265 & n1129 ) | ( n545 & n1129 ) ;
  assign n1131 = ( n337 & ~n1123 ) | ( n337 & n1130 ) | ( ~n1123 & n1130 ) ;
  assign n1134 = n188 ^ x10 ^ x0 ;
  assign n1135 = n1134 ^ n452 ^ n260 ;
  assign n1136 = n321 & ~n1135 ;
  assign n1137 = n1136 ^ n207 ^ 1'b0 ;
  assign n1132 = n692 ^ n354 ^ 1'b0 ;
  assign n1133 = n229 & n1132 ;
  assign n1138 = n1137 ^ n1133 ^ n857 ;
  assign n1142 = n656 ^ n251 ^ 1'b0 ;
  assign n1143 = n609 & ~n1142 ;
  assign n1139 = n945 ^ n452 ^ n361 ;
  assign n1140 = n1139 ^ n658 ^ 1'b0 ;
  assign n1141 = ( n650 & n1123 ) | ( n650 & n1140 ) | ( n1123 & n1140 ) ;
  assign n1144 = n1143 ^ n1141 ^ n191 ;
  assign n1153 = n404 ^ n312 ^ n235 ;
  assign n1154 = ( x106 & ~n504 ) | ( x106 & n1153 ) | ( ~n504 & n1153 ) ;
  assign n1145 = n626 | n719 ;
  assign n1146 = n1145 ^ n405 ^ 1'b0 ;
  assign n1147 = n1146 ^ n242 ^ n210 ;
  assign n1148 = ( n186 & n364 ) | ( n186 & ~n969 ) | ( n364 & ~n969 ) ;
  assign n1149 = n1148 ^ n488 ^ 1'b0 ;
  assign n1150 = n325 & n1149 ;
  assign n1151 = ( n331 & n437 ) | ( n331 & ~n1150 ) | ( n437 & ~n1150 ) ;
  assign n1152 = ( x58 & ~n1147 ) | ( x58 & n1151 ) | ( ~n1147 & n1151 ) ;
  assign n1155 = n1154 ^ n1152 ^ n253 ;
  assign n1161 = n870 ^ x104 ^ x8 ;
  assign n1162 = n827 ^ n418 ^ x37 ;
  assign n1163 = ( x91 & n1161 ) | ( x91 & ~n1162 ) | ( n1161 & ~n1162 ) ;
  assign n1164 = n1163 ^ n994 ^ n814 ;
  assign n1156 = n197 & n1088 ;
  assign n1157 = n313 & n1156 ;
  assign n1158 = n824 ^ n195 ^ x9 ;
  assign n1159 = n1158 ^ n154 ^ 1'b0 ;
  assign n1160 = n1157 | n1159 ;
  assign n1165 = n1164 ^ n1160 ^ n192 ;
  assign n1166 = n1165 ^ n883 ^ n837 ;
  assign n1167 = ( x0 & ~n449 ) | ( x0 & n733 ) | ( ~n449 & n733 ) ;
  assign n1168 = n175 & n1167 ;
  assign n1169 = n1168 ^ n411 ^ 1'b0 ;
  assign n1179 = ( n273 & ~n363 ) | ( n273 & n466 ) | ( ~n363 & n466 ) ;
  assign n1175 = n727 ^ n529 ^ x117 ;
  assign n1176 = n1175 ^ n1099 ^ n388 ;
  assign n1171 = x120 ^ x97 ^ x40 ;
  assign n1172 = ( ~x97 & n529 ) | ( ~x97 & n1171 ) | ( n529 & n1171 ) ;
  assign n1173 = n1172 ^ n383 ^ x84 ;
  assign n1174 = ( n575 & ~n874 ) | ( n575 & n1173 ) | ( ~n874 & n1173 ) ;
  assign n1177 = n1176 ^ n1174 ^ 1'b0 ;
  assign n1178 = n1093 & ~n1177 ;
  assign n1170 = n875 ^ n507 ^ x58 ;
  assign n1180 = n1179 ^ n1178 ^ n1170 ;
  assign n1181 = ( x83 & ~n132 ) | ( x83 & n584 ) | ( ~n132 & n584 ) ;
  assign n1182 = n903 ^ n863 ^ n549 ;
  assign n1183 = ( n302 & n420 ) | ( n302 & n714 ) | ( n420 & n714 ) ;
  assign n1184 = ( n629 & ~n1182 ) | ( n629 & n1183 ) | ( ~n1182 & n1183 ) ;
  assign n1185 = ( n1069 & ~n1181 ) | ( n1069 & n1184 ) | ( ~n1181 & n1184 ) ;
  assign n1186 = n974 ^ n490 ^ 1'b0 ;
  assign n1187 = n1141 & ~n1186 ;
  assign n1188 = ( n264 & n1123 ) | ( n264 & n1187 ) | ( n1123 & n1187 ) ;
  assign n1191 = n444 ^ n375 ^ x113 ;
  assign n1192 = n1191 ^ n438 ^ n344 ;
  assign n1189 = n933 ^ n239 ^ 1'b0 ;
  assign n1190 = n1062 | n1189 ;
  assign n1193 = n1192 ^ n1190 ^ n1072 ;
  assign n1214 = n564 | n947 ;
  assign n1215 = n1214 ^ x67 ^ 1'b0 ;
  assign n1212 = ( ~n367 & n705 ) | ( ~n367 & n904 ) | ( n705 & n904 ) ;
  assign n1211 = n1173 ^ n737 ^ n582 ;
  assign n1213 = n1212 ^ n1211 ^ n981 ;
  assign n1207 = n713 ^ n463 ^ 1'b0 ;
  assign n1204 = n225 ^ n173 ^ x33 ;
  assign n1205 = ( n569 & ~n626 ) | ( n569 & n1204 ) | ( ~n626 & n1204 ) ;
  assign n1203 = n611 ^ n573 ^ 1'b0 ;
  assign n1206 = n1205 ^ n1203 ^ x102 ;
  assign n1195 = ( ~n138 & n252 ) | ( ~n138 & n1148 ) | ( n252 & n1148 ) ;
  assign n1197 = n914 ^ n891 ^ x81 ;
  assign n1196 = n263 & ~n610 ;
  assign n1198 = n1197 ^ n1196 ^ 1'b0 ;
  assign n1199 = ( ~x88 & n343 ) | ( ~x88 & n814 ) | ( n343 & n814 ) ;
  assign n1200 = n659 & ~n1199 ;
  assign n1201 = n1198 & n1200 ;
  assign n1202 = ( ~n634 & n1195 ) | ( ~n634 & n1201 ) | ( n1195 & n1201 ) ;
  assign n1208 = n1207 ^ n1206 ^ n1202 ;
  assign n1194 = n373 & n398 ;
  assign n1209 = n1208 ^ n1194 ^ 1'b0 ;
  assign n1210 = ( n167 & n710 ) | ( n167 & n1209 ) | ( n710 & n1209 ) ;
  assign n1216 = n1215 ^ n1213 ^ n1210 ;
  assign n1217 = n945 ^ n453 ^ x85 ;
  assign n1218 = ( x48 & ~n318 ) | ( x48 & n1217 ) | ( ~n318 & n1217 ) ;
  assign n1219 = n1218 ^ n1046 ^ n1022 ;
  assign n1220 = ~n752 & n1219 ;
  assign n1226 = n362 ^ n319 ^ n238 ;
  assign n1227 = n1226 ^ n416 ^ x101 ;
  assign n1225 = ( x40 & n138 ) | ( x40 & ~n549 ) | ( n138 & ~n549 ) ;
  assign n1222 = x107 & n597 ;
  assign n1223 = ~x85 & n1222 ;
  assign n1221 = n541 | n1032 ;
  assign n1224 = n1223 ^ n1221 ^ 1'b0 ;
  assign n1228 = n1227 ^ n1225 ^ n1224 ;
  assign n1229 = ~n774 & n782 ;
  assign n1230 = n491 & n1229 ;
  assign n1231 = n1230 ^ n680 ^ n195 ;
  assign n1232 = ( x44 & ~n599 ) | ( x44 & n791 ) | ( ~n599 & n791 ) ;
  assign n1233 = n1232 ^ n602 ^ 1'b0 ;
  assign n1234 = n992 ^ n645 ^ n295 ;
  assign n1235 = n1234 ^ n1131 ^ n154 ;
  assign n1236 = ~n355 & n680 ;
  assign n1237 = n1236 ^ n259 ^ 1'b0 ;
  assign n1239 = n258 ^ n161 ^ n148 ;
  assign n1240 = n1239 ^ n193 ^ x114 ;
  assign n1238 = ( x0 & ~x71 ) | ( x0 & n962 ) | ( ~x71 & n962 ) ;
  assign n1241 = n1240 ^ n1238 ^ 1'b0 ;
  assign n1242 = n1241 ^ n845 ^ 1'b0 ;
  assign n1243 = ( ~n1185 & n1237 ) | ( ~n1185 & n1242 ) | ( n1237 & n1242 ) ;
  assign n1247 = n502 ^ n406 ^ x52 ;
  assign n1249 = n358 ^ n201 ^ x26 ;
  assign n1250 = n205 ^ x87 ^ 1'b0 ;
  assign n1251 = n1249 & n1250 ;
  assign n1248 = n528 ^ n190 ^ 1'b0 ;
  assign n1252 = n1251 ^ n1248 ^ n722 ;
  assign n1253 = ( n334 & n532 ) | ( n334 & ~n784 ) | ( n532 & ~n784 ) ;
  assign n1254 = n1253 ^ n363 ^ n205 ;
  assign n1255 = ( x119 & n428 ) | ( x119 & ~n1254 ) | ( n428 & ~n1254 ) ;
  assign n1256 = ( n1247 & n1252 ) | ( n1247 & n1255 ) | ( n1252 & n1255 ) ;
  assign n1257 = n1256 ^ n601 ^ 1'b0 ;
  assign n1244 = n1012 ^ n414 ^ n210 ;
  assign n1245 = n690 & n1244 ;
  assign n1246 = ( ~n746 & n821 ) | ( ~n746 & n1245 ) | ( n821 & n1245 ) ;
  assign n1258 = n1257 ^ n1246 ^ n638 ;
  assign n1261 = n559 ^ x71 ^ 1'b0 ;
  assign n1259 = n987 ^ n877 ^ n703 ;
  assign n1260 = ( n388 & n499 ) | ( n388 & n1259 ) | ( n499 & n1259 ) ;
  assign n1262 = n1261 ^ n1260 ^ n701 ;
  assign n1263 = ( n302 & n315 ) | ( n302 & ~n468 ) | ( n315 & ~n468 ) ;
  assign n1264 = n1178 ^ n472 ^ 1'b0 ;
  assign n1265 = ~n1263 & n1264 ;
  assign n1266 = n419 ^ x121 ^ 1'b0 ;
  assign n1267 = n746 | n1266 ;
  assign n1269 = ( ~x116 & n471 ) | ( ~x116 & n771 ) | ( n471 & n771 ) ;
  assign n1270 = ( x100 & n388 ) | ( x100 & n1269 ) | ( n388 & n1269 ) ;
  assign n1271 = x96 | n471 ;
  assign n1272 = ~n1270 & n1271 ;
  assign n1273 = n1272 ^ n705 ^ 1'b0 ;
  assign n1274 = n1273 ^ n825 ^ n732 ;
  assign n1268 = ~n401 & n924 ;
  assign n1275 = n1274 ^ n1268 ^ 1'b0 ;
  assign n1276 = n1275 ^ n1273 ^ n233 ;
  assign n1277 = ( ~n163 & n1179 ) | ( ~n163 & n1276 ) | ( n1179 & n1276 ) ;
  assign n1278 = n1277 ^ n1003 ^ n775 ;
  assign n1279 = n433 ^ n251 ^ 1'b0 ;
  assign n1280 = ( n234 & ~n694 ) | ( n234 & n1238 ) | ( ~n694 & n1238 ) ;
  assign n1281 = n1280 ^ n229 ^ 1'b0 ;
  assign n1282 = ( n164 & n196 ) | ( n164 & n491 ) | ( n196 & n491 ) ;
  assign n1283 = n1282 ^ n510 ^ n490 ;
  assign n1284 = ( n137 & n344 ) | ( n137 & n1283 ) | ( n344 & n1283 ) ;
  assign n1285 = ( ~n191 & n1113 ) | ( ~n191 & n1284 ) | ( n1113 & n1284 ) ;
  assign n1286 = ( n463 & n1281 ) | ( n463 & ~n1285 ) | ( n1281 & ~n1285 ) ;
  assign n1287 = ~n1029 & n1045 ;
  assign n1288 = n1287 ^ n1153 ^ x46 ;
  assign n1289 = n1288 ^ n890 ^ n722 ;
  assign n1292 = n507 ^ n221 ^ n211 ;
  assign n1295 = n576 ^ n186 ^ n133 ;
  assign n1293 = n669 ^ n584 ^ n163 ;
  assign n1294 = n1293 ^ n1126 ^ n1099 ;
  assign n1296 = n1295 ^ n1294 ^ 1'b0 ;
  assign n1297 = n1292 & n1296 ;
  assign n1298 = n1297 ^ n1031 ^ n679 ;
  assign n1290 = n148 & ~n1102 ;
  assign n1291 = ( ~x115 & n410 ) | ( ~x115 & n1290 ) | ( n410 & n1290 ) ;
  assign n1299 = n1298 ^ n1291 ^ n155 ;
  assign n1300 = ~n416 & n830 ;
  assign n1301 = n1300 ^ n835 ^ n333 ;
  assign n1302 = n1301 ^ n1029 ^ n792 ;
  assign n1303 = n1302 ^ n717 ^ 1'b0 ;
  assign n1309 = n848 ^ n554 ^ n161 ;
  assign n1310 = n1309 ^ n756 ^ n630 ;
  assign n1304 = ( n172 & n512 ) | ( n172 & n566 ) | ( n512 & n566 ) ;
  assign n1305 = n1304 ^ n584 ^ n239 ;
  assign n1306 = n1305 ^ n542 ^ n285 ;
  assign n1307 = n858 | n974 ;
  assign n1308 = n1306 & ~n1307 ;
  assign n1311 = n1310 ^ n1308 ^ n277 ;
  assign n1312 = n569 | n1176 ;
  assign n1313 = x9 | n1312 ;
  assign n1314 = n1313 ^ n719 ^ x95 ;
  assign n1315 = ( n329 & ~n381 ) | ( n329 & n728 ) | ( ~n381 & n728 ) ;
  assign n1316 = ( n314 & ~n1102 ) | ( n314 & n1315 ) | ( ~n1102 & n1315 ) ;
  assign n1317 = n142 | n178 ;
  assign n1318 = n1317 ^ x73 ^ 1'b0 ;
  assign n1319 = ( x94 & n890 ) | ( x94 & n1318 ) | ( n890 & n1318 ) ;
  assign n1320 = n954 & n1319 ;
  assign n1321 = ( x114 & ~n341 ) | ( x114 & n710 ) | ( ~n341 & n710 ) ;
  assign n1322 = n1087 ^ n944 ^ n606 ;
  assign n1323 = n1322 ^ n298 ^ x125 ;
  assign n1324 = ( x1 & ~x37 ) | ( x1 & n989 ) | ( ~x37 & n989 ) ;
  assign n1325 = n537 & n602 ;
  assign n1326 = n1324 & n1325 ;
  assign n1327 = n1326 ^ n385 ^ n329 ;
  assign n1328 = ( n1321 & ~n1323 ) | ( n1321 & n1327 ) | ( ~n1323 & n1327 ) ;
  assign n1329 = ( ~n221 & n1320 ) | ( ~n221 & n1328 ) | ( n1320 & n1328 ) ;
  assign n1330 = ( n666 & n1114 ) | ( n666 & ~n1261 ) | ( n1114 & ~n1261 ) ;
  assign n1331 = ( n655 & n987 ) | ( n655 & n1330 ) | ( n987 & n1330 ) ;
  assign n1332 = n1331 ^ n513 ^ 1'b0 ;
  assign n1333 = x8 & ~n1332 ;
  assign n1334 = ( ~n370 & n855 ) | ( ~n370 & n1018 ) | ( n855 & n1018 ) ;
  assign n1335 = n1334 ^ n1018 ^ n282 ;
  assign n1336 = n790 & ~n1335 ;
  assign n1337 = n670 ^ n228 ^ x102 ;
  assign n1338 = n1337 ^ n555 ^ 1'b0 ;
  assign n1339 = ~n1105 & n1338 ;
  assign n1340 = ( ~n868 & n1112 ) | ( ~n868 & n1269 ) | ( n1112 & n1269 ) ;
  assign n1341 = ( n890 & ~n1339 ) | ( n890 & n1340 ) | ( ~n1339 & n1340 ) ;
  assign n1344 = x75 & ~n474 ;
  assign n1345 = n1344 ^ n336 ^ 1'b0 ;
  assign n1346 = ( x84 & n698 ) | ( x84 & ~n1345 ) | ( n698 & ~n1345 ) ;
  assign n1343 = n1213 ^ n969 ^ 1'b0 ;
  assign n1342 = n1197 ^ n793 ^ n490 ;
  assign n1347 = n1346 ^ n1343 ^ n1342 ;
  assign n1348 = n1081 ^ n450 ^ n424 ;
  assign n1349 = n263 | n1348 ;
  assign n1350 = ( n278 & n894 ) | ( n278 & ~n1349 ) | ( n894 & ~n1349 ) ;
  assign n1351 = ( ~n1085 & n1175 ) | ( ~n1085 & n1350 ) | ( n1175 & n1350 ) ;
  assign n1352 = n1178 ^ n768 ^ n430 ;
  assign n1353 = n1174 ^ n608 ^ x106 ;
  assign n1354 = n1353 ^ n1252 ^ n159 ;
  assign n1355 = ( n1085 & n1352 ) | ( n1085 & n1354 ) | ( n1352 & n1354 ) ;
  assign n1356 = n1351 & ~n1355 ;
  assign n1357 = n377 & ~n1292 ;
  assign n1358 = n1357 ^ n1106 ^ n586 ;
  assign n1359 = ( x54 & n340 ) | ( x54 & ~n1085 ) | ( n340 & ~n1085 ) ;
  assign n1360 = ( n894 & n1174 ) | ( n894 & n1175 ) | ( n1174 & n1175 ) ;
  assign n1361 = ( n1295 & n1359 ) | ( n1295 & n1360 ) | ( n1359 & n1360 ) ;
  assign n1362 = n1361 ^ n1287 ^ n991 ;
  assign n1374 = x100 & ~n210 ;
  assign n1375 = ( n474 & n1162 ) | ( n474 & n1374 ) | ( n1162 & n1374 ) ;
  assign n1376 = n1226 ^ n266 ^ n200 ;
  assign n1377 = ( n954 & n1375 ) | ( n954 & n1376 ) | ( n1375 & n1376 ) ;
  assign n1378 = ( n240 & ~n974 ) | ( n240 & n1377 ) | ( ~n974 & n1377 ) ;
  assign n1366 = ( x65 & n516 ) | ( x65 & n743 ) | ( n516 & n743 ) ;
  assign n1369 = ( x51 & n140 ) | ( x51 & n519 ) | ( n140 & n519 ) ;
  assign n1370 = n854 & n1369 ;
  assign n1367 = n1318 ^ n282 ^ x56 ;
  assign n1368 = n1367 ^ x30 ^ 1'b0 ;
  assign n1371 = n1370 ^ n1368 ^ n674 ;
  assign n1372 = ( n953 & n1366 ) | ( n953 & ~n1371 ) | ( n1366 & ~n1371 ) ;
  assign n1373 = n1372 ^ n952 ^ n212 ;
  assign n1363 = n814 ^ n285 ^ n136 ;
  assign n1364 = ( n252 & n691 ) | ( n252 & n1363 ) | ( n691 & n1363 ) ;
  assign n1365 = n1364 ^ n1045 ^ n503 ;
  assign n1379 = n1378 ^ n1373 ^ n1365 ;
  assign n1387 = n1173 ^ n581 ^ x28 ;
  assign n1386 = n1252 ^ n774 ^ n270 ;
  assign n1382 = n140 & ~n352 ;
  assign n1383 = n1382 ^ n1249 ^ 1'b0 ;
  assign n1381 = ( n258 & ~n609 ) | ( n258 & n881 ) | ( ~n609 & n881 ) ;
  assign n1380 = n858 ^ n640 ^ n517 ;
  assign n1384 = n1383 ^ n1381 ^ n1380 ;
  assign n1385 = ( n832 & n1255 ) | ( n832 & n1384 ) | ( n1255 & n1384 ) ;
  assign n1388 = n1387 ^ n1386 ^ n1385 ;
  assign n1389 = x8 & ~n282 ;
  assign n1390 = ~n325 & n1389 ;
  assign n1391 = n1390 ^ n643 ^ n331 ;
  assign n1392 = n1391 ^ n1226 ^ n1122 ;
  assign n1393 = x36 & ~n1008 ;
  assign n1416 = ~n232 & n889 ;
  assign n1417 = n1416 ^ x92 ^ 1'b0 ;
  assign n1418 = n1417 ^ n947 ^ n519 ;
  assign n1394 = ( x33 & ~n354 ) | ( x33 & n721 ) | ( ~n354 & n721 ) ;
  assign n1395 = ( x39 & ~x88 ) | ( x39 & n457 ) | ( ~x88 & n457 ) ;
  assign n1396 = x63 & n723 ;
  assign n1397 = ~n512 & n1396 ;
  assign n1398 = n1397 ^ n855 ^ 1'b0 ;
  assign n1399 = n189 & ~n1398 ;
  assign n1400 = ( x59 & ~x97 ) | ( x59 & n1399 ) | ( ~x97 & n1399 ) ;
  assign n1401 = ( n921 & n1395 ) | ( n921 & n1400 ) | ( n1395 & n1400 ) ;
  assign n1402 = n875 ^ n622 ^ 1'b0 ;
  assign n1403 = n282 | n1402 ;
  assign n1404 = n1403 ^ n569 ^ n495 ;
  assign n1405 = ( ~n1241 & n1401 ) | ( ~n1241 & n1404 ) | ( n1401 & n1404 ) ;
  assign n1406 = n1405 ^ n363 ^ n180 ;
  assign n1407 = ( n283 & n291 ) | ( n283 & n557 ) | ( n291 & n557 ) ;
  assign n1408 = ( x55 & n168 ) | ( x55 & ~n1407 ) | ( n168 & ~n1407 ) ;
  assign n1409 = ( x93 & ~n173 ) | ( x93 & n479 ) | ( ~n173 & n479 ) ;
  assign n1410 = n595 ^ n577 ^ n129 ;
  assign n1411 = ( ~x32 & x63 ) | ( ~x32 & n1410 ) | ( x63 & n1410 ) ;
  assign n1412 = n1411 ^ n336 ^ x102 ;
  assign n1413 = ( ~n1408 & n1409 ) | ( ~n1408 & n1412 ) | ( n1409 & n1412 ) ;
  assign n1414 = ( n1394 & ~n1406 ) | ( n1394 & n1413 ) | ( ~n1406 & n1413 ) ;
  assign n1415 = ( x87 & n1205 ) | ( x87 & ~n1414 ) | ( n1205 & ~n1414 ) ;
  assign n1419 = n1418 ^ n1415 ^ n1245 ;
  assign n1420 = ( n221 & n280 ) | ( n221 & n754 ) | ( n280 & n754 ) ;
  assign n1425 = ( n735 & n1084 ) | ( n735 & n1110 ) | ( n1084 & n1110 ) ;
  assign n1422 = n1270 ^ n426 ^ 1'b0 ;
  assign n1421 = n1178 ^ n805 ^ n611 ;
  assign n1423 = n1422 ^ n1421 ^ n195 ;
  assign n1424 = n1423 ^ n291 ^ n252 ;
  assign n1426 = n1425 ^ n1424 ^ n1404 ;
  assign n1427 = ( n859 & ~n1324 ) | ( n859 & n1426 ) | ( ~n1324 & n1426 ) ;
  assign n1431 = n908 ^ n632 ^ n370 ;
  assign n1428 = x42 & n1259 ;
  assign n1429 = n1428 ^ n710 ^ 1'b0 ;
  assign n1430 = ( x21 & n715 ) | ( x21 & n1429 ) | ( n715 & n1429 ) ;
  assign n1432 = n1431 ^ n1430 ^ n643 ;
  assign n1437 = n309 ^ n277 ^ n210 ;
  assign n1433 = n559 ^ n259 ^ n183 ;
  assign n1434 = n1433 ^ n992 ^ n365 ;
  assign n1435 = n1434 ^ n1140 ^ n555 ;
  assign n1436 = ( n250 & ~n566 ) | ( n250 & n1435 ) | ( ~n566 & n1435 ) ;
  assign n1438 = n1437 ^ n1436 ^ n1321 ;
  assign n1439 = ( n511 & ~n1432 ) | ( n511 & n1438 ) | ( ~n1432 & n1438 ) ;
  assign n1440 = n1439 ^ n835 ^ n460 ;
  assign n1450 = ( x50 & n390 ) | ( x50 & ~n1008 ) | ( n390 & ~n1008 ) ;
  assign n1451 = n1450 ^ n411 ^ n150 ;
  assign n1452 = n325 & n1451 ;
  assign n1442 = n1135 ^ n334 ^ x42 ;
  assign n1441 = n1036 ^ n326 ^ 1'b0 ;
  assign n1443 = n1442 ^ n1441 ^ x37 ;
  assign n1446 = n1239 ^ n513 ^ n460 ;
  assign n1447 = n1446 ^ n793 ^ n549 ;
  assign n1444 = x72 & n947 ;
  assign n1445 = n1444 ^ n643 ^ 1'b0 ;
  assign n1448 = n1447 ^ n1445 ^ x39 ;
  assign n1449 = ( n1094 & n1443 ) | ( n1094 & ~n1448 ) | ( n1443 & ~n1448 ) ;
  assign n1453 = n1452 ^ n1449 ^ 1'b0 ;
  assign n1454 = ~n792 & n1453 ;
  assign n1455 = n1009 ^ x112 ^ x5 ;
  assign n1456 = ( x70 & n1340 ) | ( x70 & ~n1455 ) | ( n1340 & ~n1455 ) ;
  assign n1457 = n1456 ^ n1100 ^ n843 ;
  assign n1458 = n1457 ^ n1399 ^ 1'b0 ;
  assign n1459 = n1357 | n1458 ;
  assign n1491 = n1340 ^ n1023 ^ n135 ;
  assign n1492 = n1399 & ~n1491 ;
  assign n1493 = n1409 ^ n400 ^ 1'b0 ;
  assign n1494 = n1492 & ~n1493 ;
  assign n1487 = x127 | n355 ;
  assign n1486 = n469 & n812 ;
  assign n1488 = n1487 ^ n1486 ^ n1359 ;
  assign n1489 = ( n798 & n995 ) | ( n798 & ~n1488 ) | ( n995 & ~n1488 ) ;
  assign n1476 = n701 ^ n507 ^ n432 ;
  assign n1479 = ( n152 & n324 ) | ( n152 & ~n1227 ) | ( n324 & ~n1227 ) ;
  assign n1480 = ( n271 & n474 ) | ( n271 & ~n1479 ) | ( n474 & ~n1479 ) ;
  assign n1481 = n334 & ~n1480 ;
  assign n1482 = n1481 ^ n574 ^ 1'b0 ;
  assign n1477 = ( ~x53 & n410 ) | ( ~x53 & n825 ) | ( n410 & n825 ) ;
  assign n1478 = ( n225 & n1043 ) | ( n225 & n1477 ) | ( n1043 & n1477 ) ;
  assign n1483 = n1482 ^ n1478 ^ n572 ;
  assign n1484 = n1483 ^ n727 ^ 1'b0 ;
  assign n1485 = n1476 & n1484 ;
  assign n1463 = ( ~x63 & x112 ) | ( ~x63 & n910 ) | ( x112 & n910 ) ;
  assign n1464 = x82 & n1463 ;
  assign n1465 = n1464 ^ n225 ^ 1'b0 ;
  assign n1460 = n229 ^ x80 ^ x65 ;
  assign n1461 = n1460 ^ n705 ^ x9 ;
  assign n1462 = n1461 ^ n676 ^ x96 ;
  assign n1466 = n1465 ^ n1462 ^ n727 ;
  assign n1467 = ( n261 & ~n1139 ) | ( n261 & n1383 ) | ( ~n1139 & n1383 ) ;
  assign n1468 = ( x17 & n567 ) | ( x17 & ~n603 ) | ( n567 & ~n603 ) ;
  assign n1469 = n609 & ~n1207 ;
  assign n1470 = n1469 ^ n1441 ^ 1'b0 ;
  assign n1471 = ~n1374 & n1470 ;
  assign n1472 = n1468 & n1471 ;
  assign n1473 = n1472 ^ n1036 ^ 1'b0 ;
  assign n1474 = ( n1466 & n1467 ) | ( n1466 & n1473 ) | ( n1467 & n1473 ) ;
  assign n1475 = ( n700 & n901 ) | ( n700 & n1474 ) | ( n901 & n1474 ) ;
  assign n1490 = n1489 ^ n1485 ^ n1475 ;
  assign n1495 = n1494 ^ n1490 ^ n983 ;
  assign n1496 = ( ~x22 & x41 ) | ( ~x22 & n500 ) | ( x41 & n500 ) ;
  assign n1497 = ( n352 & n374 ) | ( n352 & ~n1496 ) | ( n374 & ~n1496 ) ;
  assign n1498 = n1315 ^ n430 ^ 1'b0 ;
  assign n1499 = n1497 & n1498 ;
  assign n1500 = ( ~n797 & n1047 ) | ( ~n797 & n1148 ) | ( n1047 & n1148 ) ;
  assign n1501 = n1500 ^ n655 ^ n406 ;
  assign n1502 = n1501 ^ n1483 ^ x41 ;
  assign n1503 = ( ~n398 & n638 ) | ( ~n398 & n1274 ) | ( n638 & n1274 ) ;
  assign n1504 = n934 | n1503 ;
  assign n1505 = n1504 ^ n1349 ^ 1'b0 ;
  assign n1506 = n1331 ^ n949 ^ n418 ;
  assign n1507 = n1505 & ~n1506 ;
  assign n1508 = n734 & n1507 ;
  assign n1509 = n619 | n679 ;
  assign n1510 = ( n336 & n1043 ) | ( n336 & ~n1239 ) | ( n1043 & ~n1239 ) ;
  assign n1511 = n1510 ^ n170 ^ x54 ;
  assign n1512 = ( n364 & n630 ) | ( n364 & ~n1511 ) | ( n630 & ~n1511 ) ;
  assign n1513 = n1512 ^ x45 ^ 1'b0 ;
  assign n1514 = n1509 & n1513 ;
  assign n1524 = n994 ^ n261 ^ x70 ;
  assign n1519 = n1013 ^ n287 ^ x76 ;
  assign n1520 = ( ~n767 & n1056 ) | ( ~n767 & n1519 ) | ( n1056 & n1519 ) ;
  assign n1521 = ( x22 & n734 ) | ( x22 & n1520 ) | ( n734 & n1520 ) ;
  assign n1522 = n1521 ^ n1079 ^ n903 ;
  assign n1523 = n1522 ^ n157 ^ 1'b0 ;
  assign n1525 = n1524 ^ n1523 ^ n1123 ;
  assign n1515 = n513 ^ n465 ^ n283 ;
  assign n1516 = ( n867 & n949 ) | ( n867 & n1515 ) | ( n949 & n1515 ) ;
  assign n1517 = n1516 ^ n1423 ^ n512 ;
  assign n1518 = n713 | n1517 ;
  assign n1526 = n1525 ^ n1518 ^ 1'b0 ;
  assign n1528 = n1038 ^ n282 ^ x120 ;
  assign n1527 = ( n394 & n518 ) | ( n394 & ~n1052 ) | ( n518 & ~n1052 ) ;
  assign n1529 = n1528 ^ n1527 ^ n360 ;
  assign n1532 = n539 ^ n424 ^ n228 ;
  assign n1533 = n1532 ^ n521 ^ n473 ;
  assign n1530 = n1148 ^ n363 ^ n190 ;
  assign n1531 = ( n284 & n1444 ) | ( n284 & ~n1530 ) | ( n1444 & ~n1530 ) ;
  assign n1534 = n1533 ^ n1531 ^ n679 ;
  assign n1535 = n1529 & n1534 ;
  assign n1536 = ( ~n1094 & n1526 ) | ( ~n1094 & n1535 ) | ( n1526 & n1535 ) ;
  assign n1537 = ~n154 & n439 ;
  assign n1538 = n1537 ^ n771 ^ n490 ;
  assign n1539 = n585 ^ n563 ^ 1'b0 ;
  assign n1540 = ~n1113 & n1539 ;
  assign n1541 = ( n274 & n1538 ) | ( n274 & n1540 ) | ( n1538 & n1540 ) ;
  assign n1545 = ( x123 & ~n221 ) | ( x123 & n317 ) | ( ~n221 & n317 ) ;
  assign n1542 = n464 ^ x8 ^ 1'b0 ;
  assign n1543 = ~n174 & n1542 ;
  assign n1544 = n1543 ^ n1174 ^ n891 ;
  assign n1546 = n1545 ^ n1544 ^ n859 ;
  assign n1547 = n674 ^ n314 ^ n234 ;
  assign n1548 = n1547 ^ n492 ^ n284 ;
  assign n1549 = ( n572 & n1305 ) | ( n572 & ~n1548 ) | ( n1305 & ~n1548 ) ;
  assign n1550 = ( n698 & ~n1022 ) | ( n698 & n1549 ) | ( ~n1022 & n1549 ) ;
  assign n1551 = ( n1541 & ~n1546 ) | ( n1541 & n1550 ) | ( ~n1546 & n1550 ) ;
  assign n1552 = ( n241 & ~n502 ) | ( n241 & n949 ) | ( ~n502 & n949 ) ;
  assign n1553 = n1552 ^ n732 ^ n574 ;
  assign n1554 = n1017 ^ n878 ^ n465 ;
  assign n1555 = ( n328 & ~n917 ) | ( n328 & n1114 ) | ( ~n917 & n1114 ) ;
  assign n1556 = n1555 ^ n1421 ^ n952 ;
  assign n1557 = ~n356 & n1556 ;
  assign n1558 = n767 | n1557 ;
  assign n1559 = ( n301 & n723 ) | ( n301 & n838 ) | ( n723 & n838 ) ;
  assign n1560 = n165 & n303 ;
  assign n1561 = ~n1559 & n1560 ;
  assign n1562 = n720 & n1561 ;
  assign n1563 = ( n1554 & n1558 ) | ( n1554 & n1562 ) | ( n1558 & n1562 ) ;
  assign n1564 = x95 & n222 ;
  assign n1565 = n1564 ^ n491 ^ 1'b0 ;
  assign n1566 = n287 & n1565 ;
  assign n1567 = n356 & ~n1566 ;
  assign n1568 = n1567 ^ n905 ^ 1'b0 ;
  assign n1569 = x45 & n481 ;
  assign n1580 = n1559 ^ n421 ^ n190 ;
  assign n1581 = ( n200 & n773 ) | ( n200 & ~n1580 ) | ( n773 & ~n1580 ) ;
  assign n1582 = ( ~n290 & n567 ) | ( ~n290 & n1581 ) | ( n567 & n1581 ) ;
  assign n1583 = ( x80 & ~x119 ) | ( x80 & n1135 ) | ( ~x119 & n1135 ) ;
  assign n1584 = ( ~n233 & n1582 ) | ( ~n233 & n1583 ) | ( n1582 & n1583 ) ;
  assign n1575 = n226 ^ n168 ^ x111 ;
  assign n1576 = ( ~n1146 & n1538 ) | ( ~n1146 & n1575 ) | ( n1538 & n1575 ) ;
  assign n1577 = n1576 ^ n463 ^ x106 ;
  assign n1574 = n775 ^ n470 ^ x12 ;
  assign n1578 = n1577 ^ n1574 ^ n386 ;
  assign n1579 = ( n415 & ~n1489 ) | ( n415 & n1578 ) | ( ~n1489 & n1578 ) ;
  assign n1570 = x14 | n409 ;
  assign n1571 = ( ~n205 & n1304 ) | ( ~n205 & n1570 ) | ( n1304 & n1570 ) ;
  assign n1572 = n1571 ^ n662 ^ n176 ;
  assign n1573 = x84 & ~n1572 ;
  assign n1585 = n1584 ^ n1579 ^ n1573 ;
  assign n1586 = ( ~n1491 & n1569 ) | ( ~n1491 & n1585 ) | ( n1569 & n1585 ) ;
  assign n1598 = ( ~n251 & n508 ) | ( ~n251 & n703 ) | ( n508 & n703 ) ;
  assign n1587 = n465 ^ x16 ^ 1'b0 ;
  assign n1588 = ( n637 & n1261 ) | ( n637 & ~n1587 ) | ( n1261 & ~n1587 ) ;
  assign n1589 = ( ~n287 & n319 ) | ( ~n287 & n1588 ) | ( n319 & n1588 ) ;
  assign n1590 = ( n333 & n459 ) | ( n333 & n596 ) | ( n459 & n596 ) ;
  assign n1591 = ( ~n170 & n542 ) | ( ~n170 & n1590 ) | ( n542 & n1590 ) ;
  assign n1592 = n1591 ^ n854 ^ n246 ;
  assign n1593 = ( x2 & n544 ) | ( x2 & n664 ) | ( n544 & n664 ) ;
  assign n1594 = ( ~x70 & n454 ) | ( ~x70 & n1593 ) | ( n454 & n1593 ) ;
  assign n1595 = n1594 ^ n950 ^ n691 ;
  assign n1596 = ( ~n1589 & n1592 ) | ( ~n1589 & n1595 ) | ( n1592 & n1595 ) ;
  assign n1597 = n1596 ^ n1234 ^ n1038 ;
  assign n1599 = n1598 ^ n1597 ^ n1368 ;
  assign n1600 = n460 ^ n357 ^ n355 ;
  assign n1601 = n1367 ^ n444 ^ n253 ;
  assign n1602 = n1343 ^ n157 ^ x75 ;
  assign n1603 = ( n1600 & n1601 ) | ( n1600 & ~n1602 ) | ( n1601 & ~n1602 ) ;
  assign n1604 = n1592 ^ n1375 ^ n375 ;
  assign n1605 = n994 ^ n642 ^ n261 ;
  assign n1606 = n1605 ^ n1517 ^ n154 ;
  assign n1608 = ( n266 & n837 ) | ( n266 & ~n980 ) | ( n837 & ~n980 ) ;
  assign n1609 = n423 & n1608 ;
  assign n1607 = n497 & n621 ;
  assign n1610 = n1609 ^ n1607 ^ 1'b0 ;
  assign n1611 = ( n800 & n1606 ) | ( n800 & ~n1610 ) | ( n1606 & ~n1610 ) ;
  assign n1612 = ( x63 & n814 ) | ( x63 & ~n1346 ) | ( n814 & ~n1346 ) ;
  assign n1613 = n1031 & n1612 ;
  assign n1614 = n1613 ^ n914 ^ 1'b0 ;
  assign n1615 = ( n1604 & n1611 ) | ( n1604 & ~n1614 ) | ( n1611 & ~n1614 ) ;
  assign n1616 = ( n912 & n1603 ) | ( n912 & n1615 ) | ( n1603 & n1615 ) ;
  assign n1617 = n1369 ^ n361 ^ x98 ;
  assign n1618 = n1617 ^ n337 ^ n246 ;
  assign n1619 = ( n300 & ~n589 ) | ( n300 & n903 ) | ( ~n589 & n903 ) ;
  assign n1620 = ( n726 & n909 ) | ( n726 & n1619 ) | ( n909 & n1619 ) ;
  assign n1626 = ( x1 & n310 ) | ( x1 & n498 ) | ( n310 & n498 ) ;
  assign n1621 = ( n309 & n524 ) | ( n309 & ~n1172 ) | ( n524 & ~n1172 ) ;
  assign n1622 = n159 & n1621 ;
  assign n1623 = n1622 ^ n818 ^ 1'b0 ;
  assign n1624 = n1623 ^ n677 ^ n130 ;
  assign n1625 = ( n569 & ~n989 ) | ( n569 & n1624 ) | ( ~n989 & n1624 ) ;
  assign n1627 = n1626 ^ n1625 ^ 1'b0 ;
  assign n1628 = ~n1012 & n1627 ;
  assign n1629 = ( n1618 & n1620 ) | ( n1618 & ~n1628 ) | ( n1620 & ~n1628 ) ;
  assign n1632 = n527 ^ n365 ^ n309 ;
  assign n1633 = ( n196 & ~n633 ) | ( n196 & n1632 ) | ( ~n633 & n1632 ) ;
  assign n1634 = n1633 ^ n541 ^ x75 ;
  assign n1635 = n1634 ^ n713 ^ x74 ;
  assign n1631 = ~n989 & n1042 ;
  assign n1636 = n1635 ^ n1631 ^ 1'b0 ;
  assign n1630 = n1000 ^ n433 ^ x13 ;
  assign n1637 = n1636 ^ n1630 ^ n1287 ;
  assign n1638 = ( n1482 & n1629 ) | ( n1482 & ~n1637 ) | ( n1629 & ~n1637 ) ;
  assign n1639 = ( n833 & ~n881 ) | ( n833 & n910 ) | ( ~n881 & n910 ) ;
  assign n1640 = n1639 ^ n1138 ^ n140 ;
  assign n1641 = n496 | n564 ;
  assign n1642 = n1641 ^ n394 ^ 1'b0 ;
  assign n1643 = ( x87 & n629 ) | ( x87 & n1642 ) | ( n629 & n1642 ) ;
  assign n1644 = n1167 & n1643 ;
  assign n1647 = ( n1173 & ~n1192 ) | ( n1173 & n1367 ) | ( ~n1192 & n1367 ) ;
  assign n1645 = n1171 ^ n444 ^ x105 ;
  assign n1646 = x34 & ~n1645 ;
  assign n1648 = n1647 ^ n1646 ^ 1'b0 ;
  assign n1649 = ~n1515 & n1648 ;
  assign n1650 = x68 & n647 ;
  assign n1651 = n1650 ^ n1426 ^ n732 ;
  assign n1652 = ( n1644 & ~n1649 ) | ( n1644 & n1651 ) | ( ~n1649 & n1651 ) ;
  assign n1654 = x40 & n1463 ;
  assign n1653 = ( x89 & n138 ) | ( x89 & n461 ) | ( n138 & n461 ) ;
  assign n1655 = n1654 ^ n1653 ^ n602 ;
  assign n1656 = x112 & n1408 ;
  assign n1657 = ~n1345 & n1656 ;
  assign n1658 = n1657 ^ n1290 ^ n161 ;
  assign n1660 = n442 ^ n428 ^ n277 ;
  assign n1661 = n1660 ^ n1239 ^ n819 ;
  assign n1662 = n1661 ^ n435 ^ n223 ;
  assign n1659 = n1014 ^ n729 ^ n285 ;
  assign n1663 = n1662 ^ n1659 ^ n706 ;
  assign n1664 = n1545 ^ n1465 ^ n506 ;
  assign n1665 = n1663 | n1664 ;
  assign n1666 = n1270 ^ n1172 ^ x123 ;
  assign n1667 = n773 & ~n1666 ;
  assign n1668 = n1667 ^ n816 ^ n716 ;
  assign n1669 = ~n181 & n1227 ;
  assign n1670 = ( n1425 & ~n1668 ) | ( n1425 & n1669 ) | ( ~n1668 & n1669 ) ;
  assign n1681 = ( x47 & ~n1083 ) | ( x47 & n1260 ) | ( ~n1083 & n1260 ) ;
  assign n1676 = n891 ^ n513 ^ n214 ;
  assign n1677 = ( ~n221 & n1179 ) | ( ~n221 & n1676 ) | ( n1179 & n1676 ) ;
  assign n1678 = n734 & n1677 ;
  assign n1679 = n1678 ^ n478 ^ x113 ;
  assign n1674 = n480 ^ n362 ^ x32 ;
  assign n1675 = n534 | n1674 ;
  assign n1680 = n1679 ^ n1675 ^ 1'b0 ;
  assign n1671 = n620 ^ x102 ^ x15 ;
  assign n1672 = ( n1377 & n1461 ) | ( n1377 & n1610 ) | ( n1461 & n1610 ) ;
  assign n1673 = ( n605 & n1671 ) | ( n605 & n1672 ) | ( n1671 & n1672 ) ;
  assign n1682 = n1681 ^ n1680 ^ n1673 ;
  assign n1683 = x43 & ~n1337 ;
  assign n1684 = ~n1639 & n1683 ;
  assign n1685 = n1662 ^ n952 ^ x125 ;
  assign n1686 = ( n486 & ~n1684 ) | ( n486 & n1685 ) | ( ~n1684 & n1685 ) ;
  assign n1687 = n1061 | n1686 ;
  assign n1689 = n528 ^ n204 ^ x104 ;
  assign n1690 = n1689 ^ n439 ^ n359 ;
  assign n1691 = n1524 ^ n248 ^ 1'b0 ;
  assign n1692 = x74 & n1691 ;
  assign n1693 = ( n242 & ~n1128 ) | ( n242 & n1692 ) | ( ~n1128 & n1692 ) ;
  assign n1694 = n1693 ^ n982 ^ n660 ;
  assign n1695 = ( ~n206 & n1690 ) | ( ~n206 & n1694 ) | ( n1690 & n1694 ) ;
  assign n1688 = n184 & n1087 ;
  assign n1696 = n1695 ^ n1688 ^ 1'b0 ;
  assign n1699 = n439 | n1577 ;
  assign n1700 = n1699 ^ n302 ^ 1'b0 ;
  assign n1697 = n333 ^ n281 ^ x68 ;
  assign n1698 = ( ~n379 & n697 ) | ( ~n379 & n1697 ) | ( n697 & n1697 ) ;
  assign n1701 = n1700 ^ n1698 ^ n349 ;
  assign n1702 = ( ~n1251 & n1682 ) | ( ~n1251 & n1701 ) | ( n1682 & n1701 ) ;
  assign n1703 = ( ~n293 & n1070 ) | ( ~n293 & n1632 ) | ( n1070 & n1632 ) ;
  assign n1704 = n1703 ^ n1303 ^ n223 ;
  assign n1705 = n388 & n646 ;
  assign n1706 = n1463 ^ n769 ^ n142 ;
  assign n1707 = ( n830 & ~n1052 ) | ( n830 & n1706 ) | ( ~n1052 & n1706 ) ;
  assign n1708 = ( ~n357 & n1705 ) | ( ~n357 & n1707 ) | ( n1705 & n1707 ) ;
  assign n1709 = n1403 ^ n760 ^ x97 ;
  assign n1710 = n1709 ^ n920 ^ n574 ;
  assign n1711 = ( n887 & n1318 ) | ( n887 & n1710 ) | ( n1318 & n1710 ) ;
  assign n1712 = n559 & ~n914 ;
  assign n1713 = ( ~n205 & n636 ) | ( ~n205 & n1712 ) | ( n636 & n1712 ) ;
  assign n1714 = n1713 ^ n1298 ^ n686 ;
  assign n1715 = n1714 ^ n1152 ^ n303 ;
  assign n1716 = n1715 ^ n1260 ^ n1147 ;
  assign n1720 = ( ~n157 & n563 ) | ( ~n157 & n861 ) | ( n563 & n861 ) ;
  assign n1721 = ( x29 & x89 ) | ( x29 & n319 ) | ( x89 & n319 ) ;
  assign n1722 = ( n198 & ~n219 ) | ( n198 & n1721 ) | ( ~n219 & n1721 ) ;
  assign n1723 = n1722 ^ n913 ^ 1'b0 ;
  assign n1724 = ( n1140 & n1720 ) | ( n1140 & n1723 ) | ( n1720 & n1723 ) ;
  assign n1717 = ( ~n332 & n516 ) | ( ~n332 & n1036 ) | ( n516 & n1036 ) ;
  assign n1718 = ( n143 & ~n1337 ) | ( n143 & n1538 ) | ( ~n1337 & n1538 ) ;
  assign n1719 = n1717 & n1718 ;
  assign n1725 = n1724 ^ n1719 ^ n1252 ;
  assign n1726 = n1725 ^ n1617 ^ n1285 ;
  assign n1727 = ( n264 & ~n1191 ) | ( n264 & n1238 ) | ( ~n1191 & n1238 ) ;
  assign n1728 = n750 ^ x25 ^ x2 ;
  assign n1729 = ( n477 & n736 ) | ( n477 & ~n1728 ) | ( n736 & ~n1728 ) ;
  assign n1730 = ( n403 & n680 ) | ( n403 & ~n1729 ) | ( n680 & ~n1729 ) ;
  assign n1731 = ( n822 & n1171 ) | ( n822 & n1359 ) | ( n1171 & n1359 ) ;
  assign n1732 = ( n144 & n1706 ) | ( n144 & ~n1731 ) | ( n1706 & ~n1731 ) ;
  assign n1733 = ( n478 & n1730 ) | ( n478 & ~n1732 ) | ( n1730 & ~n1732 ) ;
  assign n1734 = ( n1357 & n1727 ) | ( n1357 & n1733 ) | ( n1727 & n1733 ) ;
  assign n1737 = ( ~n256 & n581 ) | ( ~n256 & n804 ) | ( n581 & n804 ) ;
  assign n1735 = ( ~x85 & n498 ) | ( ~x85 & n506 ) | ( n498 & n506 ) ;
  assign n1736 = n1735 ^ n1068 ^ n361 ;
  assign n1738 = n1737 ^ n1736 ^ n451 ;
  assign n1739 = ( ~x87 & n233 ) | ( ~x87 & n253 ) | ( n233 & n253 ) ;
  assign n1740 = n1739 ^ n1163 ^ 1'b0 ;
  assign n1741 = n1738 & ~n1740 ;
  assign n1742 = ~x92 & x110 ;
  assign n1743 = n1742 ^ n1036 ^ n692 ;
  assign n1744 = n1743 ^ n298 ^ x93 ;
  assign n1745 = n1081 ^ n344 ^ 1'b0 ;
  assign n1746 = n206 & n758 ;
  assign n1747 = n1745 & n1746 ;
  assign n1757 = n387 ^ n212 ^ x127 ;
  assign n1758 = n1757 ^ n1148 ^ n254 ;
  assign n1756 = ~n307 & n633 ;
  assign n1750 = n669 ^ n312 ^ x126 ;
  assign n1751 = ( n294 & ~n559 ) | ( n294 & n1750 ) | ( ~n559 & n1750 ) ;
  assign n1752 = ( x7 & n369 ) | ( x7 & n1594 ) | ( n369 & n1594 ) ;
  assign n1753 = ( n995 & n1751 ) | ( n995 & ~n1752 ) | ( n1751 & ~n1752 ) ;
  assign n1754 = n1753 ^ n1137 ^ n377 ;
  assign n1748 = ( x2 & ~n783 ) | ( x2 & n972 ) | ( ~n783 & n972 ) ;
  assign n1749 = ( n223 & ~n624 ) | ( n223 & n1748 ) | ( ~n624 & n1748 ) ;
  assign n1755 = n1754 ^ n1749 ^ 1'b0 ;
  assign n1759 = n1758 ^ n1756 ^ n1755 ;
  assign n1760 = n1759 ^ n839 ^ 1'b0 ;
  assign n1761 = n1760 ^ n1318 ^ n1009 ;
  assign n1762 = ( x60 & ~n273 ) | ( x60 & n326 ) | ( ~n273 & n326 ) ;
  assign n1763 = n1762 ^ n994 ^ 1'b0 ;
  assign n1764 = n1623 & ~n1763 ;
  assign n1765 = ( n532 & n875 ) | ( n532 & ~n1764 ) | ( n875 & ~n1764 ) ;
  assign n1767 = n853 ^ x59 ^ 1'b0 ;
  assign n1766 = n153 ^ x119 ^ x57 ;
  assign n1768 = n1767 ^ n1766 ^ n1346 ;
  assign n1769 = n1768 ^ n1374 ^ n1034 ;
  assign n1774 = ( ~n845 & n963 ) | ( ~n845 & n1528 ) | ( n963 & n1528 ) ;
  assign n1775 = ( n409 & n1251 ) | ( n409 & n1774 ) | ( n1251 & n1774 ) ;
  assign n1770 = n863 & ~n918 ;
  assign n1771 = ( n148 & n241 ) | ( n148 & n926 ) | ( n241 & n926 ) ;
  assign n1772 = n1248 | n1771 ;
  assign n1773 = n1770 | n1772 ;
  assign n1776 = n1775 ^ n1773 ^ 1'b0 ;
  assign n1777 = ( ~n1765 & n1769 ) | ( ~n1765 & n1776 ) | ( n1769 & n1776 ) ;
  assign n1780 = n368 & ~n381 ;
  assign n1781 = ( n503 & n1102 ) | ( n503 & ~n1780 ) | ( n1102 & ~n1780 ) ;
  assign n1782 = n1781 ^ n1207 ^ n544 ;
  assign n1778 = n506 ^ n394 ^ 1'b0 ;
  assign n1779 = n1778 ^ n1595 ^ n997 ;
  assign n1783 = n1782 ^ n1779 ^ n929 ;
  assign n1791 = x114 & x123 ;
  assign n1792 = n201 ^ x123 ^ x97 ;
  assign n1793 = x67 & ~n1006 ;
  assign n1794 = ( x54 & ~n609 ) | ( x54 & n830 ) | ( ~n609 & n830 ) ;
  assign n1795 = ( n1792 & ~n1793 ) | ( n1792 & n1794 ) | ( ~n1793 & n1794 ) ;
  assign n1796 = n1795 ^ n1345 ^ n1093 ;
  assign n1797 = n1091 ^ n457 ^ 1'b0 ;
  assign n1798 = n1797 ^ x69 ^ 1'b0 ;
  assign n1799 = ( n1791 & n1796 ) | ( n1791 & n1798 ) | ( n1796 & n1798 ) ;
  assign n1790 = ( n387 & n721 ) | ( n387 & ~n1723 ) | ( n721 & ~n1723 ) ;
  assign n1786 = ( x68 & n495 ) | ( x68 & ~n1239 ) | ( n495 & ~n1239 ) ;
  assign n1787 = n1786 ^ n893 ^ n492 ;
  assign n1788 = n1787 ^ n1401 ^ n180 ;
  assign n1784 = ( n176 & ~n210 ) | ( n176 & n876 ) | ( ~n210 & n876 ) ;
  assign n1785 = ( n1277 & n1739 ) | ( n1277 & n1784 ) | ( n1739 & n1784 ) ;
  assign n1789 = n1788 ^ n1785 ^ n1423 ;
  assign n1800 = n1799 ^ n1790 ^ n1789 ;
  assign n1803 = n1576 ^ n1465 ^ x48 ;
  assign n1801 = n597 ^ n433 ^ n175 ;
  assign n1802 = ( n1091 & n1100 ) | ( n1091 & n1801 ) | ( n1100 & n1801 ) ;
  assign n1804 = n1803 ^ n1802 ^ n256 ;
  assign n1805 = ( n369 & n787 ) | ( n369 & n1089 ) | ( n787 & n1089 ) ;
  assign n1806 = ( n854 & ~n1636 ) | ( n854 & n1805 ) | ( ~n1636 & n1805 ) ;
  assign n1807 = ( n1575 & n1804 ) | ( n1575 & n1806 ) | ( n1804 & n1806 ) ;
  assign n1808 = n888 ^ n278 ^ n246 ;
  assign n1809 = ( x97 & ~n676 ) | ( x97 & n1112 ) | ( ~n676 & n1112 ) ;
  assign n1810 = ( n164 & n311 ) | ( n164 & ~n630 ) | ( n311 & ~n630 ) ;
  assign n1811 = ( ~n1808 & n1809 ) | ( ~n1808 & n1810 ) | ( n1809 & n1810 ) ;
  assign n1812 = ( ~n498 & n1147 ) | ( ~n498 & n1811 ) | ( n1147 & n1811 ) ;
  assign n1813 = n1147 ^ n952 ^ n181 ;
  assign n1814 = n1813 ^ n1357 ^ x0 ;
  assign n1815 = ( ~n537 & n1812 ) | ( ~n537 & n1814 ) | ( n1812 & n1814 ) ;
  assign n1825 = n946 ^ x126 ^ x115 ;
  assign n1823 = n374 ^ n271 ^ 1'b0 ;
  assign n1820 = n1617 ^ n160 ^ 1'b0 ;
  assign n1821 = ( ~n369 & n709 ) | ( ~n369 & n1820 ) | ( n709 & n1820 ) ;
  assign n1818 = ( ~n463 & n671 ) | ( ~n463 & n1112 ) | ( n671 & n1112 ) ;
  assign n1817 = ( ~n406 & n839 ) | ( ~n406 & n1632 ) | ( n839 & n1632 ) ;
  assign n1819 = n1818 ^ n1817 ^ 1'b0 ;
  assign n1816 = n1590 ^ n918 ^ 1'b0 ;
  assign n1822 = n1821 ^ n1819 ^ n1816 ;
  assign n1824 = n1823 ^ n1822 ^ x78 ;
  assign n1826 = n1825 ^ n1824 ^ 1'b0 ;
  assign n1827 = n1715 ^ n1263 ^ n244 ;
  assign n1828 = n953 & ~n1827 ;
  assign n1829 = n1828 ^ n605 ^ 1'b0 ;
  assign n1830 = ( n157 & ~n200 ) | ( n157 & n599 ) | ( ~n200 & n599 ) ;
  assign n1831 = n1093 | n1830 ;
  assign n1832 = ( n978 & n1029 ) | ( n978 & ~n1831 ) | ( n1029 & ~n1831 ) ;
  assign n1833 = n131 & n311 ;
  assign n1834 = n586 & ~n1286 ;
  assign n1835 = ( x62 & ~n1833 ) | ( x62 & n1834 ) | ( ~n1833 & n1834 ) ;
  assign n1836 = n1180 ^ n244 ^ x32 ;
  assign n1837 = n1836 ^ n1348 ^ n1146 ;
  assign n1838 = ( ~x2 & n301 ) | ( ~x2 & n913 ) | ( n301 & n913 ) ;
  assign n1839 = ( x56 & ~n197 ) | ( x56 & n1534 ) | ( ~n197 & n1534 ) ;
  assign n1854 = ( n233 & ~n417 ) | ( n233 & n1787 ) | ( ~n417 & n1787 ) ;
  assign n1855 = n1854 ^ n872 ^ x127 ;
  assign n1851 = n1797 ^ n719 ^ 1'b0 ;
  assign n1852 = n818 | n1851 ;
  assign n1853 = n1852 ^ n484 ^ n422 ;
  assign n1847 = n282 ^ n150 ^ x126 ;
  assign n1846 = ( n386 & n1052 ) | ( n386 & ~n1105 ) | ( n1052 & ~n1105 ) ;
  assign n1848 = n1847 ^ n1846 ^ n264 ;
  assign n1845 = n881 ^ x68 ^ 1'b0 ;
  assign n1849 = n1848 ^ n1845 ^ n283 ;
  assign n1840 = n1021 ^ n587 ^ n465 ;
  assign n1841 = n1003 ^ n920 ^ n281 ;
  assign n1842 = n554 ^ n367 ^ n317 ;
  assign n1843 = n1842 ^ n859 ^ x32 ;
  assign n1844 = ( n1840 & n1841 ) | ( n1840 & ~n1843 ) | ( n1841 & ~n1843 ) ;
  assign n1850 = n1849 ^ n1844 ^ n1220 ;
  assign n1856 = n1855 ^ n1853 ^ n1850 ;
  assign n1857 = n1185 & n1505 ;
  assign n1858 = ( n257 & n1856 ) | ( n257 & n1857 ) | ( n1856 & n1857 ) ;
  assign n1859 = ( ~n1838 & n1839 ) | ( ~n1838 & n1858 ) | ( n1839 & n1858 ) ;
  assign n1860 = n932 ^ n789 ^ n258 ;
  assign n1861 = n674 ^ n293 ^ n132 ;
  assign n1863 = ( x125 & n139 ) | ( x125 & ~n147 ) | ( n139 & ~n147 ) ;
  assign n1862 = n719 ^ n295 ^ n251 ;
  assign n1864 = n1863 ^ n1862 ^ 1'b0 ;
  assign n1865 = n255 & n1864 ;
  assign n1866 = n1861 & n1865 ;
  assign n1867 = n1866 ^ n1276 ^ n967 ;
  assign n1871 = ( x75 & ~x103 ) | ( x75 & n247 ) | ( ~x103 & n247 ) ;
  assign n1872 = ( n689 & n1134 ) | ( n689 & n1871 ) | ( n1134 & n1871 ) ;
  assign n1873 = n1345 ^ n1112 ^ 1'b0 ;
  assign n1874 = n1872 & n1873 ;
  assign n1869 = ( n1394 & n1434 ) | ( n1394 & ~n1657 ) | ( n1434 & ~n1657 ) ;
  assign n1868 = n1752 ^ n1293 ^ n949 ;
  assign n1870 = n1869 ^ n1868 ^ n1606 ;
  assign n1875 = n1874 ^ n1870 ^ 1'b0 ;
  assign n1876 = n1867 & n1875 ;
  assign n1877 = ( n352 & n1860 ) | ( n352 & ~n1876 ) | ( n1860 & ~n1876 ) ;
  assign n1878 = n686 | n906 ;
  assign n1879 = ( x41 & n779 ) | ( x41 & n1369 ) | ( n779 & n1369 ) ;
  assign n1880 = ( n417 & n660 ) | ( n417 & n1879 ) | ( n660 & n1879 ) ;
  assign n1881 = n1880 ^ n798 ^ x27 ;
  assign n1882 = ( n607 & ~n1584 ) | ( n607 & n1881 ) | ( ~n1584 & n1881 ) ;
  assign n1883 = n1345 ^ n647 ^ n488 ;
  assign n1884 = ( n1083 & ~n1882 ) | ( n1083 & n1883 ) | ( ~n1882 & n1883 ) ;
  assign n1885 = ( n1877 & ~n1878 ) | ( n1877 & n1884 ) | ( ~n1878 & n1884 ) ;
  assign n1886 = ( x7 & n651 ) | ( x7 & ~n1524 ) | ( n651 & ~n1524 ) ;
  assign n1887 = n1886 ^ n1059 ^ n431 ;
  assign n1888 = ( ~n396 & n1812 ) | ( ~n396 & n1887 ) | ( n1812 & n1887 ) ;
  assign n1889 = n822 ^ n463 ^ n346 ;
  assign n1890 = n1889 ^ n1368 ^ n219 ;
  assign n1892 = n1742 ^ n560 ^ n197 ;
  assign n1891 = n547 ^ x121 ^ x54 ;
  assign n1893 = n1892 ^ n1891 ^ n993 ;
  assign n1894 = ( n345 & n1890 ) | ( n345 & n1893 ) | ( n1890 & n1893 ) ;
  assign n1895 = n912 ^ n371 ^ x4 ;
  assign n1896 = n1895 ^ n745 ^ n448 ;
  assign n1897 = ( n529 & n586 ) | ( n529 & ~n1896 ) | ( n586 & ~n1896 ) ;
  assign n1898 = n1897 ^ n1468 ^ n242 ;
  assign n1899 = ( ~n1218 & n1894 ) | ( ~n1218 & n1898 ) | ( n1894 & n1898 ) ;
  assign n1900 = n583 & ~n912 ;
  assign n1901 = n1403 & n1900 ;
  assign n1902 = n1901 ^ n1097 ^ n246 ;
  assign n1903 = n1552 & n1902 ;
  assign n1904 = ~n1846 & n1903 ;
  assign n1905 = n740 ^ n619 ^ n265 ;
  assign n1906 = ( n343 & n481 ) | ( n343 & n1905 ) | ( n481 & n1905 ) ;
  assign n1907 = n1906 ^ n355 ^ x31 ;
  assign n1908 = x79 & ~n647 ;
  assign n1909 = n1908 ^ n1421 ^ n923 ;
  assign n1910 = ( n214 & n1907 ) | ( n214 & n1909 ) | ( n1907 & n1909 ) ;
  assign n1911 = ( n1411 & n1904 ) | ( n1411 & n1910 ) | ( n1904 & n1910 ) ;
  assign n1912 = n647 ^ n518 ^ x64 ;
  assign n1916 = n524 ^ x99 ^ x18 ;
  assign n1914 = n1363 | n1544 ;
  assign n1915 = n1914 ^ n355 ^ 1'b0 ;
  assign n1917 = n1916 ^ n1915 ^ n1319 ;
  assign n1913 = n1778 ^ n1762 ^ n1203 ;
  assign n1918 = n1917 ^ n1913 ^ n1369 ;
  assign n1922 = n1543 ^ n447 ^ x78 ;
  assign n1920 = n348 ^ n252 ^ 1'b0 ;
  assign n1919 = n1707 ^ n549 ^ n322 ;
  assign n1921 = n1920 ^ n1919 ^ n1175 ;
  assign n1923 = n1922 ^ n1921 ^ n363 ;
  assign n1924 = x92 & ~n1377 ;
  assign n1925 = ~n394 & n1924 ;
  assign n1926 = n1925 ^ n1677 ^ n1128 ;
  assign n1927 = n1403 ^ n1276 ^ n426 ;
  assign n1928 = ~n1926 & n1927 ;
  assign n1929 = ( n1918 & n1923 ) | ( n1918 & n1928 ) | ( n1923 & n1928 ) ;
  assign n1935 = ( n234 & ~n1300 ) | ( n234 & n1752 ) | ( ~n1300 & n1752 ) ;
  assign n1936 = ( ~n492 & n1412 ) | ( ~n492 & n1935 ) | ( n1412 & n1935 ) ;
  assign n1930 = n679 ^ n318 ^ x6 ;
  assign n1931 = ( x111 & n387 ) | ( x111 & n1930 ) | ( n387 & n1930 ) ;
  assign n1932 = n1931 ^ n1460 ^ n369 ;
  assign n1933 = n1932 ^ n373 ^ 1'b0 ;
  assign n1934 = n1933 ^ n1583 ^ x59 ;
  assign n1937 = n1936 ^ n1934 ^ n638 ;
  assign n1938 = n1937 ^ n1815 ^ n838 ;
  assign n1940 = ( n178 & n1368 ) | ( n178 & ~n1465 ) | ( n1368 & ~n1465 ) ;
  assign n1939 = n1434 ^ n894 ^ n810 ;
  assign n1941 = n1940 ^ n1939 ^ x114 ;
  assign n1942 = ( n661 & n1541 ) | ( n661 & n1555 ) | ( n1541 & n1555 ) ;
  assign n1943 = n1942 ^ n1848 ^ n1569 ;
  assign n1944 = n139 & n1932 ;
  assign n1945 = n1944 ^ n1337 ^ 1'b0 ;
  assign n1946 = n1808 ^ n176 ^ 1'b0 ;
  assign n1947 = ( x8 & n322 ) | ( x8 & n339 ) | ( n322 & n339 ) ;
  assign n1948 = n358 | n1947 ;
  assign n1949 = n1946 | n1948 ;
  assign n1950 = n654 & ~n1745 ;
  assign n1951 = ~n1949 & n1950 ;
  assign n1952 = ~n1185 & n1750 ;
  assign n1953 = n1951 & n1952 ;
  assign n1954 = n1866 ^ n351 ^ n186 ;
  assign n1955 = ( n482 & n1764 ) | ( n482 & ~n1954 ) | ( n1764 & ~n1954 ) ;
  assign n1956 = n1955 ^ n743 ^ n292 ;
  assign n1957 = n205 ^ n166 ^ x3 ;
  assign n1958 = n1957 ^ n1480 ^ n248 ;
  assign n1959 = n1958 ^ n292 ^ x3 ;
  assign n1960 = n1959 ^ n1596 ^ n1377 ;
  assign n1961 = ( n1038 & ~n1956 ) | ( n1038 & n1960 ) | ( ~n1956 & n1960 ) ;
  assign n1968 = n827 ^ n710 ^ n428 ;
  assign n1969 = n1968 ^ n885 ^ n709 ;
  assign n1962 = ~n288 & n705 ;
  assign n1963 = ~n646 & n1962 ;
  assign n1964 = n1963 ^ n920 ^ n263 ;
  assign n1965 = n1890 ^ n980 ^ n948 ;
  assign n1966 = n1183 & ~n1965 ;
  assign n1967 = n1964 & n1966 ;
  assign n1970 = n1969 ^ n1967 ^ n580 ;
  assign n1971 = ( n150 & n444 ) | ( n150 & n901 ) | ( n444 & n901 ) ;
  assign n1972 = n1377 ^ n798 ^ n307 ;
  assign n1973 = n789 ^ n603 ^ n587 ;
  assign n1974 = ( n332 & n1252 ) | ( n332 & n1973 ) | ( n1252 & n1973 ) ;
  assign n1975 = n1974 ^ n317 ^ x49 ;
  assign n1976 = ( n1115 & n1972 ) | ( n1115 & ~n1975 ) | ( n1972 & ~n1975 ) ;
  assign n1977 = ( ~n243 & n381 ) | ( ~n243 & n1976 ) | ( n381 & n1976 ) ;
  assign n1982 = n1643 ^ n698 ^ 1'b0 ;
  assign n1983 = ( ~n1276 & n1380 ) | ( ~n1276 & n1982 ) | ( n1380 & n1982 ) ;
  assign n1978 = n1232 ^ n1226 ^ n904 ;
  assign n1979 = n1919 ^ n160 ^ x25 ;
  assign n1980 = ( n1126 & n1883 ) | ( n1126 & n1979 ) | ( n1883 & n1979 ) ;
  assign n1981 = ( n1672 & n1978 ) | ( n1672 & ~n1980 ) | ( n1978 & ~n1980 ) ;
  assign n1984 = n1983 ^ n1981 ^ n1064 ;
  assign n1985 = ( n1971 & n1977 ) | ( n1971 & ~n1984 ) | ( n1977 & ~n1984 ) ;
  assign n1989 = n1359 ^ n248 ^ 1'b0 ;
  assign n1990 = n801 | n1989 ;
  assign n1991 = ( n637 & ~n1227 ) | ( n637 & n1990 ) | ( ~n1227 & n1990 ) ;
  assign n1987 = n495 ^ x26 ^ 1'b0 ;
  assign n1988 = ~n491 & n1987 ;
  assign n1986 = ( x9 & n183 ) | ( x9 & n1806 ) | ( n183 & n1806 ) ;
  assign n1992 = n1991 ^ n1988 ^ n1986 ;
  assign n1993 = ( n218 & n592 ) | ( n218 & n1957 ) | ( n592 & n1957 ) ;
  assign n2000 = ( n608 & n1565 ) | ( n608 & n1731 ) | ( n1565 & n1731 ) ;
  assign n1994 = ( ~n207 & n289 ) | ( ~n207 & n491 ) | ( n289 & n491 ) ;
  assign n1995 = ( x32 & ~n314 ) | ( x32 & n1994 ) | ( ~n314 & n1994 ) ;
  assign n1996 = n1995 ^ n1593 ^ 1'b0 ;
  assign n1997 = n1758 | n1996 ;
  assign n1998 = ( ~x123 & n206 ) | ( ~x123 & n1997 ) | ( n206 & n1997 ) ;
  assign n1999 = ( n510 & n1261 ) | ( n510 & n1998 ) | ( n1261 & n1998 ) ;
  assign n2001 = n2000 ^ n1999 ^ n989 ;
  assign n2002 = n1874 ^ n270 ^ x48 ;
  assign n2003 = ( n1993 & ~n2001 ) | ( n1993 & n2002 ) | ( ~n2001 & n2002 ) ;
  assign n2004 = n640 ^ n314 ^ x93 ;
  assign n2005 = n2004 ^ n1064 ^ n399 ;
  assign n2006 = ~n1697 & n2005 ;
  assign n2007 = n2006 ^ n436 ^ 1'b0 ;
  assign n2008 = ( n502 & ~n560 ) | ( n502 & n1881 ) | ( ~n560 & n1881 ) ;
  assign n2010 = ( ~x78 & n374 ) | ( ~x78 & n1818 ) | ( n374 & n1818 ) ;
  assign n2009 = n1932 ^ n1523 ^ 1'b0 ;
  assign n2011 = n2010 ^ n2009 ^ n1216 ;
  assign n2012 = ( n1990 & ~n2008 ) | ( n1990 & n2011 ) | ( ~n2008 & n2011 ) ;
  assign n2013 = ( n1233 & n1865 ) | ( n1233 & n2012 ) | ( n1865 & n2012 ) ;
  assign n2014 = n2013 ^ n1802 ^ x26 ;
  assign n2025 = n1157 ^ n500 ^ n145 ;
  assign n2015 = ( x44 & x115 ) | ( x44 & n550 ) | ( x115 & n550 ) ;
  assign n2016 = n2015 ^ n1983 ^ n474 ;
  assign n2017 = ( n555 & ~n812 ) | ( n555 & n1046 ) | ( ~n812 & n1046 ) ;
  assign n2018 = n1860 ^ n1163 ^ n713 ;
  assign n2019 = ( n399 & ~n2017 ) | ( n399 & n2018 ) | ( ~n2017 & n2018 ) ;
  assign n2020 = n248 & n853 ;
  assign n2021 = ~n412 & n2020 ;
  assign n2022 = ( n297 & n1571 ) | ( n297 & ~n1908 ) | ( n1571 & ~n1908 ) ;
  assign n2023 = ( n1846 & n2021 ) | ( n1846 & n2022 ) | ( n2021 & n2022 ) ;
  assign n2024 = ( n2016 & n2019 ) | ( n2016 & ~n2023 ) | ( n2019 & ~n2023 ) ;
  assign n2026 = n2025 ^ n2024 ^ 1'b0 ;
  assign n2028 = n743 ^ n522 ^ n406 ;
  assign n2029 = n2028 ^ n876 ^ n539 ;
  assign n2030 = n1313 & ~n2029 ;
  assign n2027 = n1642 ^ n1212 ^ 1'b0 ;
  assign n2031 = n2030 ^ n2027 ^ n906 ;
  assign n2045 = ( ~n144 & n674 ) | ( ~n144 & n901 ) | ( n674 & n901 ) ;
  assign n2041 = n990 ^ n386 ^ n367 ;
  assign n2039 = ( n143 & ~n597 ) | ( n143 & n1271 ) | ( ~n597 & n1271 ) ;
  assign n2040 = ( x94 & ~n1794 ) | ( x94 & n2039 ) | ( ~n1794 & n2039 ) ;
  assign n2038 = ( x57 & ~n986 ) | ( x57 & n1109 ) | ( ~n986 & n1109 ) ;
  assign n2042 = n2041 ^ n2040 ^ n2038 ;
  assign n2034 = ~n164 & n187 ;
  assign n2035 = n2034 ^ n1972 ^ n931 ;
  assign n2036 = n627 & n2035 ;
  assign n2037 = n1346 & n2036 ;
  assign n2043 = n2042 ^ n2037 ^ n833 ;
  assign n2032 = ( n535 & n1002 ) | ( n535 & ~n1609 ) | ( n1002 & ~n1609 ) ;
  assign n2033 = ~n243 & n2032 ;
  assign n2044 = n2043 ^ n2033 ^ 1'b0 ;
  assign n2046 = n2045 ^ n2044 ^ x15 ;
  assign n2047 = ( x114 & n792 ) | ( x114 & ~n1540 ) | ( n792 & ~n1540 ) ;
  assign n2048 = ( n405 & n737 ) | ( n405 & ~n2047 ) | ( n737 & ~n2047 ) ;
  assign n2049 = n178 | n2048 ;
  assign n2050 = n2049 ^ n380 ^ 1'b0 ;
  assign n2051 = n2050 ^ n1310 ^ n438 ;
  assign n2052 = ( x20 & ~n283 ) | ( x20 & n1141 ) | ( ~n283 & n1141 ) ;
  assign n2053 = n2052 ^ n1503 ^ n1205 ;
  assign n2054 = ( n1134 & ~n1690 ) | ( n1134 & n2053 ) | ( ~n1690 & n2053 ) ;
  assign n2055 = x21 & n134 ;
  assign n2056 = n187 ^ n148 ^ x108 ;
  assign n2057 = n2055 & n2056 ;
  assign n2063 = ( n741 & n823 ) | ( n741 & ~n1282 ) | ( n823 & ~n1282 ) ;
  assign n2060 = n232 | n365 ;
  assign n2061 = n2060 ^ n143 ^ 1'b0 ;
  assign n2062 = ~n1021 & n2061 ;
  assign n2058 = ( n339 & n504 ) | ( n339 & ~n1677 ) | ( n504 & ~n1677 ) ;
  assign n2059 = n2058 ^ n1436 ^ n1021 ;
  assign n2064 = n2063 ^ n2062 ^ n2059 ;
  assign n2066 = n1205 ^ n480 ^ x92 ;
  assign n2067 = ( ~n1174 & n1201 ) | ( ~n1174 & n2066 ) | ( n1201 & n2066 ) ;
  assign n2065 = ( ~n631 & n1612 ) | ( ~n631 & n1713 ) | ( n1612 & n1713 ) ;
  assign n2068 = n2067 ^ n2065 ^ x80 ;
  assign n2069 = ( n146 & n812 ) | ( n146 & ~n2017 ) | ( n812 & ~n2017 ) ;
  assign n2070 = n2069 ^ x113 ^ 1'b0 ;
  assign n2071 = n2068 | n2070 ;
  assign n2076 = ( ~n371 & n731 ) | ( ~n371 & n1401 ) | ( n731 & n1401 ) ;
  assign n2075 = n603 ^ x70 ^ x7 ;
  assign n2077 = n2076 ^ n2075 ^ n945 ;
  assign n2073 = n1722 ^ n961 ^ n265 ;
  assign n2072 = ( ~n136 & n193 ) | ( ~n136 & n205 ) | ( n193 & n205 ) ;
  assign n2074 = n2073 ^ n2072 ^ n1444 ;
  assign n2078 = n2077 ^ n2074 ^ 1'b0 ;
  assign n2079 = n1645 ^ n1074 ^ n894 ;
  assign n2080 = ( n157 & n459 ) | ( n157 & n1823 ) | ( n459 & n1823 ) ;
  assign n2081 = ( ~n944 & n2079 ) | ( ~n944 & n2080 ) | ( n2079 & n2080 ) ;
  assign n2082 = n568 & n2081 ;
  assign n2083 = ( n379 & n740 ) | ( n379 & n1181 ) | ( n740 & n1181 ) ;
  assign n2084 = n2083 ^ n341 ^ 1'b0 ;
  assign n2085 = x77 & n2084 ;
  assign n2086 = n2085 ^ n1727 ^ n1134 ;
  assign n2087 = n2086 ^ n567 ^ 1'b0 ;
  assign n2088 = ~n2082 & n2087 ;
  assign n2089 = n2088 ^ n1297 ^ n1238 ;
  assign n2093 = ( n749 & n771 ) | ( n749 & n1969 ) | ( n771 & n1969 ) ;
  assign n2121 = ( ~x30 & n241 ) | ( ~x30 & n2093 ) | ( n241 & n2093 ) ;
  assign n2119 = n1104 ^ n705 ^ x48 ;
  assign n2118 = ( ~x90 & n249 ) | ( ~x90 & n606 ) | ( n249 & n606 ) ;
  assign n2120 = n2119 ^ n2118 ^ n1164 ;
  assign n2122 = n2121 ^ n2120 ^ n986 ;
  assign n2115 = n1879 ^ n1781 ^ n522 ;
  assign n2113 = ~x103 & n1181 ;
  assign n2114 = n2113 ^ n1861 ^ n475 ;
  assign n2116 = n2115 ^ n2114 ^ n1033 ;
  assign n2109 = n1061 ^ n659 ^ n643 ;
  assign n2110 = n1932 ^ n744 ^ n443 ;
  assign n2111 = ( ~n1644 & n2109 ) | ( ~n1644 & n2110 ) | ( n2109 & n2110 ) ;
  assign n2112 = ( n1285 & n1639 ) | ( n1285 & n2111 ) | ( n1639 & n2111 ) ;
  assign n2117 = n2116 ^ n2112 ^ n1532 ;
  assign n2090 = n341 & n578 ;
  assign n2091 = n2090 ^ n1407 ^ n1037 ;
  assign n2092 = ~n203 & n2091 ;
  assign n2095 = ( ~n1588 & n1762 ) | ( ~n1588 & n1802 ) | ( n1762 & n1802 ) ;
  assign n2094 = n2093 ^ n1050 ^ n168 ;
  assign n2096 = n2095 ^ n2094 ^ 1'b0 ;
  assign n2097 = x12 & ~n2096 ;
  assign n2098 = ( ~x49 & n2092 ) | ( ~x49 & n2097 ) | ( n2092 & n2097 ) ;
  assign n2099 = n1088 ^ n214 ^ x56 ;
  assign n2101 = n374 ^ x106 ^ x56 ;
  assign n2100 = n789 ^ n549 ^ n532 ;
  assign n2102 = n2101 ^ n2100 ^ 1'b0 ;
  assign n2103 = n191 & ~n2102 ;
  assign n2104 = ( ~n942 & n1892 ) | ( ~n942 & n2103 ) | ( n1892 & n2103 ) ;
  assign n2105 = n2104 ^ n2103 ^ 1'b0 ;
  assign n2106 = n2105 ^ n340 ^ x23 ;
  assign n2107 = ( n1982 & n2099 ) | ( n1982 & ~n2106 ) | ( n2099 & ~n2106 ) ;
  assign n2108 = ( x36 & n2098 ) | ( x36 & n2107 ) | ( n2098 & n2107 ) ;
  assign n2123 = n2122 ^ n2117 ^ n2108 ;
  assign n2124 = x54 & n457 ;
  assign n2125 = ( ~n251 & n937 ) | ( ~n251 & n2124 ) | ( n937 & n2124 ) ;
  assign n2126 = n464 & n1590 ;
  assign n2127 = n2126 ^ n473 ^ 1'b0 ;
  assign n2128 = n2127 ^ n1494 ^ n1192 ;
  assign n2129 = n215 ^ x29 ^ x22 ;
  assign n2130 = n2129 ^ n1300 ^ 1'b0 ;
  assign n2131 = n1734 & ~n2130 ;
  assign n2147 = ( n321 & n1053 ) | ( n321 & ~n1467 ) | ( n1053 & ~n1467 ) ;
  assign n2133 = ( n768 & n1257 ) | ( n768 & ~n1433 ) | ( n1257 & ~n1433 ) ;
  assign n2137 = ( x89 & n529 ) | ( x89 & n947 ) | ( n529 & n947 ) ;
  assign n2138 = ( n337 & ~n468 ) | ( n337 & n1433 ) | ( ~n468 & n1433 ) ;
  assign n2139 = ( ~x78 & n225 ) | ( ~x78 & n235 ) | ( n225 & n235 ) ;
  assign n2140 = n2139 ^ n1059 ^ n383 ;
  assign n2141 = ( n2137 & n2138 ) | ( n2137 & n2140 ) | ( n2138 & n2140 ) ;
  assign n2142 = n1920 ^ n1752 ^ n1694 ;
  assign n2143 = ( n1052 & ~n2141 ) | ( n1052 & n2142 ) | ( ~n2141 & n2142 ) ;
  assign n2134 = ( ~n664 & n719 ) | ( ~n664 & n1274 ) | ( n719 & n1274 ) ;
  assign n2135 = n2134 ^ n328 ^ x114 ;
  assign n2136 = ( n967 & n1451 ) | ( n967 & n2135 ) | ( n1451 & n2135 ) ;
  assign n2144 = n2143 ^ n2136 ^ n1342 ;
  assign n2145 = ~n2133 & n2144 ;
  assign n2146 = n2145 ^ n249 ^ 1'b0 ;
  assign n2132 = ( n523 & n841 ) | ( n523 & n885 ) | ( n841 & n885 ) ;
  assign n2148 = n2147 ^ n2146 ^ n2132 ;
  assign n2149 = n1925 ^ n1322 ^ n241 ;
  assign n2150 = n2149 ^ n1659 ^ n1076 ;
  assign n2159 = n1765 ^ n1751 ^ n1649 ;
  assign n2157 = n482 ^ n348 ^ n147 ;
  assign n2156 = ( n691 & n1521 ) | ( n691 & ~n1767 ) | ( n1521 & ~n1767 ) ;
  assign n2154 = ( x34 & x44 ) | ( x34 & n890 ) | ( x44 & n890 ) ;
  assign n2152 = n1423 ^ n288 ^ 1'b0 ;
  assign n2151 = n1273 ^ n1028 ^ n824 ;
  assign n2153 = n2152 ^ n2151 ^ n848 ;
  assign n2155 = n2154 ^ n2153 ^ n648 ;
  assign n2158 = n2157 ^ n2156 ^ n2155 ;
  assign n2160 = n2159 ^ n2158 ^ n1894 ;
  assign n2161 = n2160 ^ n228 ^ 1'b0 ;
  assign n2162 = ~n1857 & n2161 ;
  assign n2163 = n1004 | n1353 ;
  assign n2164 = n985 & ~n2163 ;
  assign n2170 = ( ~x2 & n458 ) | ( ~x2 & n687 ) | ( n458 & n687 ) ;
  assign n2168 = x63 & ~n1139 ;
  assign n2169 = ( ~n1181 & n1676 ) | ( ~n1181 & n2168 ) | ( n1676 & n2168 ) ;
  assign n2165 = ( n256 & ~n1369 ) | ( n256 & n1477 ) | ( ~n1369 & n1477 ) ;
  assign n2166 = ( n671 & n1677 ) | ( n671 & ~n2165 ) | ( n1677 & ~n2165 ) ;
  assign n2167 = n2166 ^ n1569 ^ n1034 ;
  assign n2171 = n2170 ^ n2169 ^ n2167 ;
  assign n2172 = n1081 ^ n640 ^ n173 ;
  assign n2173 = n2172 ^ n1957 ^ x114 ;
  assign n2174 = n2173 ^ n1269 ^ n954 ;
  assign n2175 = n1284 ^ n1239 ^ n778 ;
  assign n2176 = ( ~n1730 & n2174 ) | ( ~n1730 & n2175 ) | ( n2174 & n2175 ) ;
  assign n2177 = n2171 | n2176 ;
  assign n2178 = n2101 ^ n1304 ^ n789 ;
  assign n2179 = ( ~n563 & n806 ) | ( ~n563 & n1692 ) | ( n806 & n1692 ) ;
  assign n2180 = n1012 ^ n471 ^ n151 ;
  assign n2181 = n2180 ^ n982 ^ n272 ;
  assign n2182 = n964 & n2181 ;
  assign n2183 = ( n2178 & n2179 ) | ( n2178 & ~n2182 ) | ( n2179 & ~n2182 ) ;
  assign n2184 = ( n1765 & n2177 ) | ( n1765 & ~n2183 ) | ( n2177 & ~n2183 ) ;
  assign n2185 = n1665 ^ n380 ^ 1'b0 ;
  assign n2186 = ( n777 & n2184 ) | ( n777 & n2185 ) | ( n2184 & n2185 ) ;
  assign n2187 = ( n757 & ~n1218 ) | ( n757 & n2186 ) | ( ~n1218 & n2186 ) ;
  assign n2188 = ( x14 & ~n1385 ) | ( x14 & n1753 ) | ( ~n1385 & n1753 ) ;
  assign n2189 = n2188 ^ n428 ^ n409 ;
  assign n2190 = n2189 ^ n1097 ^ 1'b0 ;
  assign n2191 = ~n921 & n2190 ;
  assign n2195 = ( n246 & ~n641 ) | ( n246 & n825 ) | ( ~n641 & n825 ) ;
  assign n2192 = n671 | n833 ;
  assign n2193 = n2192 ^ n429 ^ 1'b0 ;
  assign n2194 = ( n674 & n941 ) | ( n674 & n2193 ) | ( n941 & n2193 ) ;
  assign n2196 = n2195 ^ n2194 ^ n1538 ;
  assign n2197 = n2196 ^ n215 ^ x65 ;
  assign n2198 = n2197 ^ n1840 ^ n360 ;
  assign n2205 = ( n319 & n419 ) | ( n319 & ~n826 ) | ( n419 & ~n826 ) ;
  assign n2203 = n1825 ^ n1083 ^ n244 ;
  assign n2204 = ( ~n536 & n1044 ) | ( ~n536 & n2203 ) | ( n1044 & n2203 ) ;
  assign n2206 = n2205 ^ n2204 ^ n1257 ;
  assign n2207 = n1849 ^ n1791 ^ n1645 ;
  assign n2208 = ( n1269 & n1618 ) | ( n1269 & n1729 ) | ( n1618 & n1729 ) ;
  assign n2209 = n2208 ^ n2129 ^ n1782 ;
  assign n2210 = n692 | n2209 ;
  assign n2211 = n226 | n2210 ;
  assign n2212 = ( n771 & n1033 ) | ( n771 & ~n2211 ) | ( n1033 & ~n2211 ) ;
  assign n2213 = ( ~n2206 & n2207 ) | ( ~n2206 & n2212 ) | ( n2207 & n2212 ) ;
  assign n2199 = n174 | n1244 ;
  assign n2200 = n2199 ^ n260 ^ 1'b0 ;
  assign n2201 = n1786 ^ n891 ^ n311 ;
  assign n2202 = n2200 | n2201 ;
  assign n2214 = n2213 ^ n2202 ^ 1'b0 ;
  assign n2215 = n2214 ^ n1556 ^ n540 ;
  assign n2217 = n373 & n522 ;
  assign n2218 = ( n408 & n443 ) | ( n408 & ~n799 ) | ( n443 & ~n799 ) ;
  assign n2219 = n2218 ^ n729 ^ 1'b0 ;
  assign n2220 = ( n331 & n1737 ) | ( n331 & ~n2219 ) | ( n1737 & ~n2219 ) ;
  assign n2221 = ( n844 & n2217 ) | ( n844 & ~n2220 ) | ( n2217 & ~n2220 ) ;
  assign n2216 = ( n475 & n1064 ) | ( n475 & n2129 ) | ( n1064 & n2129 ) ;
  assign n2222 = n2221 ^ n2216 ^ n1677 ;
  assign n2244 = n133 | n1477 ;
  assign n2245 = n2244 ^ x93 ^ 1'b0 ;
  assign n2246 = n2245 ^ n2218 ^ n1537 ;
  assign n2247 = n1588 ^ n1322 ^ n859 ;
  assign n2248 = ( n328 & n2246 ) | ( n328 & ~n2247 ) | ( n2246 & ~n2247 ) ;
  assign n2249 = n1659 & ~n2248 ;
  assign n2250 = n2249 ^ n946 ^ 1'b0 ;
  assign n2251 = ( n1524 & n2152 ) | ( n1524 & ~n2250 ) | ( n2152 & ~n2250 ) ;
  assign n2252 = n2251 ^ n1637 ^ 1'b0 ;
  assign n2226 = ( n1256 & n1974 ) | ( n1256 & ~n2120 ) | ( n1974 & ~n2120 ) ;
  assign n2238 = n658 & ~n673 ;
  assign n2239 = ( n238 & n387 ) | ( n238 & ~n2238 ) | ( n387 & ~n2238 ) ;
  assign n2240 = n2239 ^ n1982 ^ n1695 ;
  assign n2227 = n2060 ^ n760 ^ n705 ;
  assign n2228 = ( n1000 & ~n1709 ) | ( n1000 & n2227 ) | ( ~n1709 & n2227 ) ;
  assign n2230 = n495 ^ n317 ^ x16 ;
  assign n2231 = n1249 ^ n850 ^ 1'b0 ;
  assign n2232 = n284 & n2231 ;
  assign n2233 = ( n980 & ~n2230 ) | ( n980 & n2232 ) | ( ~n2230 & n2232 ) ;
  assign n2234 = n1840 & ~n2233 ;
  assign n2229 = n1489 ^ n651 ^ n361 ;
  assign n2235 = n2234 ^ n2229 ^ n1872 ;
  assign n2236 = n2235 ^ n1731 ^ n1049 ;
  assign n2237 = ( n1443 & n2228 ) | ( n1443 & n2236 ) | ( n2228 & n2236 ) ;
  assign n2241 = n2240 ^ n2237 ^ n239 ;
  assign n2242 = ~n2226 & n2241 ;
  assign n2243 = ~x67 & n2242 ;
  assign n2223 = ( n311 & n1037 ) | ( n311 & n1146 ) | ( n1037 & n1146 ) ;
  assign n2224 = n1046 ^ n861 ^ x105 ;
  assign n2225 = ( n1538 & n2223 ) | ( n1538 & ~n2224 ) | ( n2223 & ~n2224 ) ;
  assign n2253 = n2252 ^ n2243 ^ n2225 ;
  assign n2254 = n1516 ^ n801 ^ n200 ;
  assign n2255 = n2254 ^ n1267 ^ x100 ;
  assign n2256 = n932 & n2255 ;
  assign n2262 = n1377 ^ n1257 ^ n784 ;
  assign n2263 = n1172 ^ n623 ^ n199 ;
  assign n2264 = ( n214 & n1015 ) | ( n214 & n2263 ) | ( n1015 & n2263 ) ;
  assign n2265 = n2264 ^ n951 ^ n804 ;
  assign n2266 = n958 ^ n889 ^ n650 ;
  assign n2267 = ( n469 & n840 ) | ( n469 & ~n2266 ) | ( n840 & ~n2266 ) ;
  assign n2268 = ~n2265 & n2267 ;
  assign n2269 = ( ~n2220 & n2262 ) | ( ~n2220 & n2268 ) | ( n2262 & n2268 ) ;
  assign n2257 = n1707 ^ n875 ^ x67 ;
  assign n2258 = ~n541 & n2194 ;
  assign n2259 = n2258 ^ n319 ^ 1'b0 ;
  assign n2260 = ( n596 & n2257 ) | ( n596 & ~n2259 ) | ( n2257 & ~n2259 ) ;
  assign n2261 = ~n1108 & n2260 ;
  assign n2270 = n2269 ^ n2261 ^ 1'b0 ;
  assign n2271 = ~n323 & n592 ;
  assign n2272 = n2271 ^ n194 ^ 1'b0 ;
  assign n2273 = n2272 ^ n1288 ^ n871 ;
  assign n2286 = ( x1 & n160 ) | ( x1 & n949 ) | ( n160 & n949 ) ;
  assign n2285 = ( ~x124 & n278 ) | ( ~x124 & n521 ) | ( n278 & n521 ) ;
  assign n2287 = n2286 ^ n2285 ^ n582 ;
  assign n2288 = ( n432 & n914 ) | ( n432 & ~n1537 ) | ( n914 & ~n1537 ) ;
  assign n2289 = n2287 & n2288 ;
  assign n2290 = n1774 & n2289 ;
  assign n2291 = ( n1475 & n1897 ) | ( n1475 & n2290 ) | ( n1897 & n2290 ) ;
  assign n2292 = n2291 ^ n373 ^ 1'b0 ;
  assign n2293 = x108 & ~n2292 ;
  assign n2274 = ~n932 & n1591 ;
  assign n2275 = ( n365 & n797 ) | ( n365 & ~n2274 ) | ( n797 & ~n2274 ) ;
  assign n2276 = ( n547 & n640 ) | ( n547 & ~n2275 ) | ( n640 & ~n2275 ) ;
  assign n2279 = ( n157 & n249 ) | ( n157 & ~n376 ) | ( n249 & ~n376 ) ;
  assign n2277 = ( ~x6 & n341 ) | ( ~x6 & n367 ) | ( n341 & n367 ) ;
  assign n2278 = n2277 ^ n981 ^ n324 ;
  assign n2280 = n2279 ^ n2278 ^ n909 ;
  assign n2281 = ~n816 & n2280 ;
  assign n2282 = n2276 & n2281 ;
  assign n2283 = n2282 ^ n1308 ^ 1'b0 ;
  assign n2284 = ~n2082 & n2283 ;
  assign n2294 = n2293 ^ n2284 ^ 1'b0 ;
  assign n2295 = ( n1226 & n1978 ) | ( n1226 & ~n1980 ) | ( n1978 & ~n1980 ) ;
  assign n2296 = n1403 ^ n932 ^ n779 ;
  assign n2297 = n512 ^ n237 ^ n220 ;
  assign n2298 = n2297 ^ n1752 ^ n340 ;
  assign n2299 = n2298 ^ n1346 ^ 1'b0 ;
  assign n2300 = n2296 & ~n2299 ;
  assign n2301 = n2269 ^ n2245 ^ n1992 ;
  assign n2313 = n608 & ~n936 ;
  assign n2314 = n2313 ^ n1087 ^ 1'b0 ;
  assign n2315 = ( ~n834 & n896 ) | ( ~n834 & n2314 ) | ( n896 & n2314 ) ;
  assign n2316 = n1767 ^ n513 ^ n290 ;
  assign n2317 = ( n2208 & ~n2315 ) | ( n2208 & n2316 ) | ( ~n2315 & n2316 ) ;
  assign n2302 = n1972 ^ n932 ^ 1'b0 ;
  assign n2303 = n281 & n2302 ;
  assign n2304 = n2303 ^ n1483 ^ n352 ;
  assign n2305 = n2304 ^ n1830 ^ n1293 ;
  assign n2307 = n567 | n974 ;
  assign n2308 = n2307 ^ x11 ^ 1'b0 ;
  assign n2309 = n1423 & ~n2308 ;
  assign n2306 = n1124 ^ n789 ^ x105 ;
  assign n2310 = n2309 ^ n2306 ^ n2060 ;
  assign n2311 = n2310 ^ n2209 ^ n530 ;
  assign n2312 = n2305 | n2311 ;
  assign n2318 = n2317 ^ n2312 ^ 1'b0 ;
  assign n2325 = n1171 ^ n210 ^ 1'b0 ;
  assign n2326 = n214 | n2325 ;
  assign n2327 = n2326 ^ n1706 ^ n753 ;
  assign n2320 = ( ~n971 & n1045 ) | ( ~n971 & n1657 ) | ( n1045 & n1657 ) ;
  assign n2321 = ( ~n451 & n805 ) | ( ~n451 & n2320 ) | ( n805 & n2320 ) ;
  assign n2319 = ~n880 & n1407 ;
  assign n2322 = n2321 ^ n2319 ^ 1'b0 ;
  assign n2323 = n2322 ^ n300 ^ 1'b0 ;
  assign n2324 = n905 & n2323 ;
  assign n2328 = n2327 ^ n2324 ^ n139 ;
  assign n2329 = n857 ^ n200 ^ x54 ;
  assign n2330 = n2329 ^ n2184 ^ n1129 ;
  assign n2331 = n2095 | n2133 ;
  assign n2332 = ( n1463 & n2330 ) | ( n1463 & ~n2331 ) | ( n2330 & ~n2331 ) ;
  assign n2333 = ~n169 & n211 ;
  assign n2334 = n1108 & n2333 ;
  assign n2335 = ( n454 & n496 ) | ( n454 & n810 ) | ( n496 & n810 ) ;
  assign n2339 = ( n863 & n924 ) | ( n863 & n1434 ) | ( n924 & n1434 ) ;
  assign n2340 = ( x78 & n2266 ) | ( x78 & n2339 ) | ( n2266 & n2339 ) ;
  assign n2336 = ( x6 & n1113 ) | ( x6 & ~n1645 ) | ( n1113 & ~n1645 ) ;
  assign n2337 = n1771 ^ n732 ^ n722 ;
  assign n2338 = n2336 & ~n2337 ;
  assign n2341 = n2340 ^ n2338 ^ 1'b0 ;
  assign n2342 = n942 ^ n368 ^ x76 ;
  assign n2343 = n2341 & ~n2342 ;
  assign n2344 = ( n1668 & n2335 ) | ( n1668 & n2343 ) | ( n2335 & n2343 ) ;
  assign n2345 = n2344 ^ n1946 ^ n1393 ;
  assign n2346 = n1124 ^ x85 ^ 1'b0 ;
  assign n2347 = n937 | n2346 ;
  assign n2348 = ( ~x16 & n1141 ) | ( ~x16 & n2336 ) | ( n1141 & n2336 ) ;
  assign n2349 = ( n1768 & n2347 ) | ( n1768 & n2348 ) | ( n2347 & n2348 ) ;
  assign n2350 = ( n1046 & n2205 ) | ( n1046 & n2349 ) | ( n2205 & n2349 ) ;
  assign n2351 = n1786 ^ x83 ^ 1'b0 ;
  assign n2352 = n2351 ^ n854 ^ n244 ;
  assign n2353 = n1234 ^ n222 ^ x9 ;
  assign n2354 = n2353 ^ n811 ^ x105 ;
  assign n2355 = ( n1451 & ~n2352 ) | ( n1451 & n2354 ) | ( ~n2352 & n2354 ) ;
  assign n2356 = ( n621 & n709 ) | ( n621 & ~n2355 ) | ( n709 & ~n2355 ) ;
  assign n2357 = ( n1090 & ~n2350 ) | ( n1090 & n2356 ) | ( ~n2350 & n2356 ) ;
  assign n2358 = ( n152 & n183 ) | ( n152 & n253 ) | ( n183 & n253 ) ;
  assign n2359 = ( n287 & n1173 ) | ( n287 & ~n1645 ) | ( n1173 & ~n1645 ) ;
  assign n2360 = n2359 ^ n2093 ^ 1'b0 ;
  assign n2361 = ( n530 & n2358 ) | ( n530 & n2360 ) | ( n2358 & n2360 ) ;
  assign n2362 = n725 & ~n2234 ;
  assign n2363 = n2362 ^ n1207 ^ 1'b0 ;
  assign n2364 = n2363 ^ n1932 ^ n1925 ;
  assign n2371 = ( n243 & n532 ) | ( n243 & ~n944 ) | ( n532 & ~n944 ) ;
  assign n2365 = n792 ^ x65 ^ 1'b0 ;
  assign n2366 = n582 ^ n471 ^ 1'b0 ;
  assign n2367 = n340 | n2366 ;
  assign n2368 = ( n937 & ~n2365 ) | ( n937 & n2367 ) | ( ~n2365 & n2367 ) ;
  assign n2369 = n2368 ^ n1298 ^ 1'b0 ;
  assign n2370 = n2369 ^ n330 ^ 1'b0 ;
  assign n2372 = n2371 ^ n2370 ^ n1445 ;
  assign n2373 = ( n707 & ~n868 ) | ( n707 & n2120 ) | ( ~n868 & n2120 ) ;
  assign n2374 = ( n477 & n1442 ) | ( n477 & ~n2373 ) | ( n1442 & ~n2373 ) ;
  assign n2375 = ( ~n227 & n330 ) | ( ~n227 & n2374 ) | ( n330 & n2374 ) ;
  assign n2376 = n336 & ~n1512 ;
  assign n2377 = ~n1668 & n2376 ;
  assign n2378 = n2377 ^ n2275 ^ n1119 ;
  assign n2379 = ( n542 & ~n1921 ) | ( n542 & n2378 ) | ( ~n1921 & n2378 ) ;
  assign n2380 = n2379 ^ n2113 ^ 1'b0 ;
  assign n2381 = n2063 ^ n1223 ^ n865 ;
  assign n2389 = ~n1172 & n1422 ;
  assign n2390 = ( n1421 & n2091 ) | ( n1421 & n2389 ) | ( n2091 & n2389 ) ;
  assign n2382 = n981 ^ n234 ^ 1'b0 ;
  assign n2383 = n2382 ^ n755 ^ n332 ;
  assign n2384 = x77 & ~n362 ;
  assign n2385 = n2384 ^ n984 ^ 1'b0 ;
  assign n2386 = ( ~x25 & n839 ) | ( ~x25 & n1162 ) | ( n839 & n1162 ) ;
  assign n2387 = ( x127 & n2385 ) | ( x127 & n2386 ) | ( n2385 & n2386 ) ;
  assign n2388 = ( x89 & n2383 ) | ( x89 & ~n2387 ) | ( n2383 & ~n2387 ) ;
  assign n2391 = n2390 ^ n2388 ^ n1452 ;
  assign n2394 = n278 & ~n2382 ;
  assign n2392 = n2347 ^ n1995 ^ n392 ;
  assign n2393 = n2392 ^ n876 ^ n135 ;
  assign n2395 = n2394 ^ n2393 ^ n2172 ;
  assign n2396 = n2314 ^ n1238 ^ n362 ;
  assign n2397 = ( n658 & n1425 ) | ( n658 & n1549 ) | ( n1425 & n1549 ) ;
  assign n2398 = ( n1123 & ~n2396 ) | ( n1123 & n2397 ) | ( ~n2396 & n2397 ) ;
  assign n2399 = ( n2391 & n2395 ) | ( n2391 & n2398 ) | ( n2395 & n2398 ) ;
  assign n2400 = ( n1031 & n2381 ) | ( n1031 & n2399 ) | ( n2381 & n2399 ) ;
  assign n2401 = ( ~n514 & n1736 ) | ( ~n514 & n1816 ) | ( n1736 & n1816 ) ;
  assign n2402 = n2401 ^ n1442 ^ n942 ;
  assign n2403 = n966 ^ n742 ^ n411 ;
  assign n2404 = ~n602 & n1263 ;
  assign n2405 = n1339 & ~n2135 ;
  assign n2406 = ~n688 & n2405 ;
  assign n2407 = n2406 ^ n2121 ^ n1755 ;
  assign n2408 = n1905 ^ n557 ^ n160 ;
  assign n2409 = ( x30 & n416 ) | ( x30 & ~n2408 ) | ( n416 & ~n2408 ) ;
  assign n2410 = n2104 ^ n1940 ^ 1'b0 ;
  assign n2411 = ( n1612 & n2409 ) | ( n1612 & ~n2410 ) | ( n2409 & ~n2410 ) ;
  assign n2412 = ( n2122 & n2407 ) | ( n2122 & ~n2411 ) | ( n2407 & ~n2411 ) ;
  assign n2413 = ( n1482 & n1793 ) | ( n1482 & ~n2298 ) | ( n1793 & ~n2298 ) ;
  assign n2414 = ( n330 & n1035 ) | ( n330 & ~n1593 ) | ( n1035 & ~n1593 ) ;
  assign n2415 = ( n1124 & n1422 ) | ( n1124 & n1581 ) | ( n1422 & n1581 ) ;
  assign n2416 = ( ~n383 & n1942 ) | ( ~n383 & n2415 ) | ( n1942 & n2415 ) ;
  assign n2417 = n1570 ^ n1444 ^ n1152 ;
  assign n2418 = n297 & n2417 ;
  assign n2419 = ( n498 & ~n904 ) | ( n498 & n2418 ) | ( ~n904 & n2418 ) ;
  assign n2420 = ( ~n2414 & n2416 ) | ( ~n2414 & n2419 ) | ( n2416 & n2419 ) ;
  assign n2421 = ~n2413 & n2420 ;
  assign n2422 = ( n783 & ~n878 ) | ( n783 & n2421 ) | ( ~n878 & n2421 ) ;
  assign n2423 = n2298 & ~n2345 ;
  assign n2424 = n2423 ^ n455 ^ 1'b0 ;
  assign n2436 = ( n370 & n474 ) | ( n370 & n606 ) | ( n474 & n606 ) ;
  assign n2437 = n2436 ^ n728 ^ n713 ;
  assign n2433 = n634 ^ n189 ^ x83 ;
  assign n2432 = n1817 ^ n742 ^ x112 ;
  assign n2429 = n1153 ^ x67 ^ 1'b0 ;
  assign n2430 = n421 & n2429 ;
  assign n2431 = n2279 & n2430 ;
  assign n2434 = n2433 ^ n2432 ^ n2431 ;
  assign n2435 = n2434 ^ n963 ^ n524 ;
  assign n2427 = ( x25 & ~n527 ) | ( x25 & n2141 ) | ( ~n527 & n2141 ) ;
  assign n2428 = ( n1276 & n1397 ) | ( n1276 & n2427 ) | ( n1397 & n2427 ) ;
  assign n2438 = n2437 ^ n2435 ^ n2428 ;
  assign n2425 = n1106 ^ n196 ^ 1'b0 ;
  assign n2426 = ( ~n765 & n2007 ) | ( ~n765 & n2425 ) | ( n2007 & n2425 ) ;
  assign n2439 = n2438 ^ n2426 ^ n660 ;
  assign n2441 = n878 ^ n767 ^ n274 ;
  assign n2442 = ( n482 & n517 ) | ( n482 & n1879 ) | ( n517 & n1879 ) ;
  assign n2443 = ( ~n2316 & n2441 ) | ( ~n2316 & n2442 ) | ( n2441 & n2442 ) ;
  assign n2440 = n1994 ^ n1749 ^ n1342 ;
  assign n2444 = n2443 ^ n2440 ^ n1529 ;
  assign n2445 = n573 & n817 ;
  assign n2446 = ~x74 & n2445 ;
  assign n2447 = ( ~n431 & n760 ) | ( ~n431 & n1167 ) | ( n760 & n1167 ) ;
  assign n2448 = ( ~n1173 & n1305 ) | ( ~n1173 & n2351 ) | ( n1305 & n2351 ) ;
  assign n2449 = ( n1024 & n1555 ) | ( n1024 & ~n2221 ) | ( n1555 & ~n2221 ) ;
  assign n2450 = ( n2447 & n2448 ) | ( n2447 & n2449 ) | ( n2448 & n2449 ) ;
  assign n2451 = n2446 & ~n2450 ;
  assign n2452 = ( ~n414 & n577 ) | ( ~n414 & n626 ) | ( n577 & n626 ) ;
  assign n2453 = ~n188 & n771 ;
  assign n2454 = x24 & n716 ;
  assign n2455 = ( n1976 & n2453 ) | ( n1976 & ~n2454 ) | ( n2453 & ~n2454 ) ;
  assign n2456 = ( ~n249 & n1064 ) | ( ~n249 & n2455 ) | ( n1064 & n2455 ) ;
  assign n2457 = ( n967 & ~n2452 ) | ( n967 & n2456 ) | ( ~n2452 & n2456 ) ;
  assign n2458 = ~n1327 & n2457 ;
  assign n2459 = n2458 ^ n2111 ^ n792 ;
  assign n2460 = n370 ^ n356 ^ 1'b0 ;
  assign n2461 = n2460 ^ n2060 ^ n1969 ;
  assign n2462 = n2326 ^ n1554 ^ n315 ;
  assign n2463 = ( x46 & n2274 ) | ( x46 & n2462 ) | ( n2274 & n2462 ) ;
  assign n2464 = n1988 & n2463 ;
  assign n2465 = n2464 ^ n456 ^ 1'b0 ;
  assign n2466 = n2465 ^ n1571 ^ n726 ;
  assign n2467 = n1571 ^ n1303 ^ n757 ;
  assign n2468 = ( n2461 & n2466 ) | ( n2461 & n2467 ) | ( n2466 & n2467 ) ;
  assign n2469 = n1588 & n2468 ;
  assign n2494 = ( n580 & n836 ) | ( n580 & ~n1842 ) | ( n836 & ~n1842 ) ;
  assign n2495 = n2365 | n2494 ;
  assign n2496 = n2267 | n2495 ;
  assign n2492 = n1933 ^ x105 ^ 1'b0 ;
  assign n2493 = ( n1524 & n2095 ) | ( n1524 & ~n2492 ) | ( n2095 & ~n2492 ) ;
  assign n2497 = n2496 ^ n2493 ^ 1'b0 ;
  assign n2498 = n804 & n2497 ;
  assign n2499 = n611 & n2498 ;
  assign n2500 = n2499 ^ n824 ^ 1'b0 ;
  assign n2485 = n2274 ^ n577 ^ n380 ;
  assign n2486 = n2485 ^ n2173 ^ n1283 ;
  assign n2487 = x72 & ~n2314 ;
  assign n2488 = n2487 ^ n465 ^ n280 ;
  assign n2489 = n2488 ^ n1027 ^ n565 ;
  assign n2490 = ( n2303 & n2486 ) | ( n2303 & n2489 ) | ( n2486 & n2489 ) ;
  assign n2483 = ( n139 & n169 ) | ( n139 & n428 ) | ( n169 & n428 ) ;
  assign n2481 = ( ~x65 & n336 ) | ( ~x65 & n1991 ) | ( n336 & n1991 ) ;
  assign n2482 = n946 & n2481 ;
  assign n2484 = n2483 ^ n2482 ^ 1'b0 ;
  assign n2491 = n2490 ^ n2484 ^ 1'b0 ;
  assign n2479 = n1731 ^ n1269 ^ n1124 ;
  assign n2473 = ( n278 & n492 ) | ( n278 & n989 ) | ( n492 & n989 ) ;
  assign n2474 = ( n789 & ~n1061 ) | ( n789 & n2473 ) | ( ~n1061 & n2473 ) ;
  assign n2475 = ( ~n519 & n1908 ) | ( ~n519 & n2474 ) | ( n1908 & n2474 ) ;
  assign n2476 = ( ~n246 & n1895 ) | ( ~n246 & n2475 ) | ( n1895 & n2475 ) ;
  assign n2470 = ( ~n855 & n1369 ) | ( ~n855 & n1901 ) | ( n1369 & n1901 ) ;
  assign n2471 = ( n268 & ~n584 ) | ( n268 & n1042 ) | ( ~n584 & n1042 ) ;
  assign n2472 = ( n494 & n2470 ) | ( n494 & ~n2471 ) | ( n2470 & ~n2471 ) ;
  assign n2477 = n2476 ^ n2472 ^ n1843 ;
  assign n2478 = n638 | n2477 ;
  assign n2480 = n2479 ^ n2478 ^ 1'b0 ;
  assign n2501 = n2500 ^ n2491 ^ n2480 ;
  assign n2502 = ( n941 & n1523 ) | ( n941 & ~n1871 ) | ( n1523 & ~n1871 ) ;
  assign n2503 = n2141 ^ n1906 ^ n1606 ;
  assign n2504 = n2503 ^ n129 ^ x36 ;
  assign n2507 = ( n585 & n1345 ) | ( n585 & n1881 ) | ( n1345 & n1881 ) ;
  assign n2508 = n2507 ^ n1309 ^ n1288 ;
  assign n2505 = ( n200 & n448 ) | ( n200 & n1055 ) | ( n448 & n1055 ) ;
  assign n2506 = n1089 | n2505 ;
  assign n2509 = n2508 ^ n2506 ^ 1'b0 ;
  assign n2510 = n1037 ^ n474 ^ n459 ;
  assign n2511 = n2510 ^ n325 ^ x1 ;
  assign n2512 = n2511 ^ n1198 ^ 1'b0 ;
  assign n2513 = x73 & n2512 ;
  assign n2514 = ( n1161 & ~n1556 ) | ( n1161 & n2513 ) | ( ~n1556 & n2513 ) ;
  assign n2515 = ( ~n1255 & n2278 ) | ( ~n1255 & n2321 ) | ( n2278 & n2321 ) ;
  assign n2516 = n1925 ^ n1133 ^ n131 ;
  assign n2517 = n1646 & n2516 ;
  assign n2518 = n1342 & n2517 ;
  assign n2519 = ( x12 & ~n2515 ) | ( x12 & n2518 ) | ( ~n2515 & n2518 ) ;
  assign n2520 = n2124 & ~n2226 ;
  assign n2521 = ( ~x108 & n2516 ) | ( ~x108 & n2520 ) | ( n2516 & n2520 ) ;
  assign n2522 = n1550 & n2521 ;
  assign n2523 = ( n1619 & n2119 ) | ( n1619 & ~n2522 ) | ( n2119 & ~n2522 ) ;
  assign n2531 = ( n232 & ~n596 ) | ( n232 & n1797 ) | ( ~n596 & n1797 ) ;
  assign n2532 = n2531 ^ n207 ^ n170 ;
  assign n2524 = ( n474 & n524 ) | ( n474 & ~n912 ) | ( n524 & ~n912 ) ;
  assign n2525 = ( n336 & n1794 ) | ( n336 & n2524 ) | ( n1794 & n2524 ) ;
  assign n2526 = n2525 ^ n2141 ^ 1'b0 ;
  assign n2527 = n1963 ^ n660 ^ n256 ;
  assign n2528 = ( ~x14 & n507 ) | ( ~x14 & n2441 ) | ( n507 & n2441 ) ;
  assign n2529 = n2527 | n2528 ;
  assign n2530 = n2526 & ~n2529 ;
  assign n2533 = n2532 ^ n2530 ^ n1330 ;
  assign n2534 = n1634 ^ n1340 ^ n822 ;
  assign n2535 = ( n707 & ~n2108 ) | ( n707 & n2534 ) | ( ~n2108 & n2534 ) ;
  assign n2536 = ( n514 & n872 ) | ( n514 & n1660 ) | ( n872 & n1660 ) ;
  assign n2538 = ~n609 & n1479 ;
  assign n2539 = ( n190 & ~n1584 ) | ( n190 & n2538 ) | ( ~n1584 & n2538 ) ;
  assign n2537 = n1381 ^ n1193 ^ n944 ;
  assign n2540 = n2539 ^ n2537 ^ n1974 ;
  assign n2541 = ( n788 & n1927 ) | ( n788 & n2540 ) | ( n1927 & n2540 ) ;
  assign n2542 = ( n1116 & ~n2536 ) | ( n1116 & n2541 ) | ( ~n2536 & n2541 ) ;
  assign n2543 = ~n1195 & n1793 ;
  assign n2544 = n797 ^ n244 ^ 1'b0 ;
  assign n2545 = n2544 ^ n1157 ^ n603 ;
  assign n2546 = n742 & n1869 ;
  assign n2547 = n2546 ^ n1225 ^ 1'b0 ;
  assign n2548 = n627 & ~n1302 ;
  assign n2549 = n2547 & n2548 ;
  assign n2550 = ( x60 & n674 ) | ( x60 & n1547 ) | ( n674 & n1547 ) ;
  assign n2551 = ( x100 & ~x112 ) | ( x100 & n175 ) | ( ~x112 & n175 ) ;
  assign n2552 = ( x47 & n431 ) | ( x47 & ~n2551 ) | ( n431 & ~n2551 ) ;
  assign n2553 = ( x106 & n1871 ) | ( x106 & ~n2552 ) | ( n1871 & ~n2552 ) ;
  assign n2554 = ( n988 & n2550 ) | ( n988 & n2553 ) | ( n2550 & n2553 ) ;
  assign n2555 = ( ~n1137 & n2549 ) | ( ~n1137 & n2554 ) | ( n2549 & n2554 ) ;
  assign n2564 = n1677 ^ n1515 ^ n304 ;
  assign n2558 = n1855 ^ n482 ^ n381 ;
  assign n2559 = n783 & ~n2558 ;
  assign n2560 = ~n1786 & n2559 ;
  assign n2561 = n859 ^ n478 ^ 1'b0 ;
  assign n2562 = ~n2560 & n2561 ;
  assign n2563 = ( ~n159 & n2280 ) | ( ~n159 & n2562 ) | ( n2280 & n2562 ) ;
  assign n2565 = n2564 ^ n2563 ^ n170 ;
  assign n2556 = n830 & n1845 ;
  assign n2557 = n2556 ^ n2100 ^ n1285 ;
  assign n2566 = n2565 ^ n2557 ^ n978 ;
  assign n2567 = n2539 ^ n1147 ^ x31 ;
  assign n2568 = n155 | n627 ;
  assign n2569 = n2568 ^ n2229 ^ n1550 ;
  assign n2570 = ( n715 & n2567 ) | ( n715 & ~n2569 ) | ( n2567 & ~n2569 ) ;
  assign n2575 = ( ~n228 & n568 ) | ( ~n228 & n913 ) | ( n568 & n913 ) ;
  assign n2574 = ( n242 & n891 ) | ( n242 & n1331 ) | ( n891 & n1331 ) ;
  assign n2572 = ( n855 & n1654 ) | ( n855 & ~n1695 ) | ( n1654 & ~n1695 ) ;
  assign n2571 = ~n1306 & n2316 ;
  assign n2573 = n2572 ^ n2571 ^ 1'b0 ;
  assign n2576 = n2575 ^ n2574 ^ n2573 ;
  assign n2577 = n2576 ^ n1943 ^ x28 ;
  assign n2578 = n1531 & n1872 ;
  assign n2579 = ~n1690 & n2578 ;
  assign n2580 = n1751 ^ n1028 ^ n251 ;
  assign n2581 = ( x59 & ~n1262 ) | ( x59 & n2580 ) | ( ~n1262 & n2580 ) ;
  assign n2582 = ( ~n1038 & n2200 ) | ( ~n1038 & n2581 ) | ( n2200 & n2581 ) ;
  assign n2589 = ( x61 & ~n255 ) | ( x61 & n508 ) | ( ~n255 & n508 ) ;
  assign n2587 = n1645 ^ n759 ^ n540 ;
  assign n2588 = ~n1014 & n2587 ;
  assign n2590 = n2589 ^ n2588 ^ 1'b0 ;
  assign n2583 = ( x63 & ~n549 ) | ( x63 & n792 ) | ( ~n549 & n792 ) ;
  assign n2584 = n1855 ^ n736 ^ 1'b0 ;
  assign n2585 = n2583 & ~n2584 ;
  assign n2586 = n2585 ^ n1290 ^ n752 ;
  assign n2591 = n2590 ^ n2586 ^ n282 ;
  assign n2592 = ( n2327 & n2582 ) | ( n2327 & ~n2591 ) | ( n2582 & ~n2591 ) ;
  assign n2594 = ( x70 & n829 ) | ( x70 & n1184 ) | ( n829 & n1184 ) ;
  assign n2593 = ~n224 & n1618 ;
  assign n2595 = n2594 ^ n2593 ^ 1'b0 ;
  assign n2596 = ( x28 & ~n1273 ) | ( x28 & n2309 ) | ( ~n1273 & n2309 ) ;
  assign n2597 = n2596 ^ n850 ^ n278 ;
  assign n2598 = n2254 ^ n1155 ^ n211 ;
  assign n2599 = ( n637 & n1083 ) | ( n637 & n1587 ) | ( n1083 & n1587 ) ;
  assign n2600 = ( n2220 & ~n2598 ) | ( n2220 & n2599 ) | ( ~n2598 & n2599 ) ;
  assign n2601 = ( n341 & n2597 ) | ( n341 & n2600 ) | ( n2597 & n2600 ) ;
  assign n2602 = ~n2595 & n2601 ;
  assign n2620 = n1594 ^ n559 ^ x89 ;
  assign n2621 = n2238 | n2620 ;
  assign n2622 = n529 | n2621 ;
  assign n2623 = ( ~n189 & n653 ) | ( ~n189 & n2622 ) | ( n653 & n2622 ) ;
  assign n2618 = ( x101 & n692 ) | ( x101 & n937 ) | ( n692 & n937 ) ;
  assign n2619 = ( x6 & n421 ) | ( x6 & n2618 ) | ( n421 & n2618 ) ;
  assign n2624 = n2623 ^ n2619 ^ n2120 ;
  assign n2614 = ( ~x125 & n874 ) | ( ~x125 & n2018 ) | ( n874 & n2018 ) ;
  assign n2615 = n2614 ^ n774 ^ 1'b0 ;
  assign n2610 = ( ~x14 & x25 ) | ( ~x14 & x108 ) | ( x25 & x108 ) ;
  assign n2611 = n829 & n2610 ;
  assign n2612 = n2611 ^ n835 ^ 1'b0 ;
  assign n2607 = n1184 ^ n810 ^ n382 ;
  assign n2605 = ( n161 & n382 ) | ( n161 & n1072 ) | ( n382 & n1072 ) ;
  assign n2603 = ~n381 & n1211 ;
  assign n2604 = n404 & n2603 ;
  assign n2606 = n2605 ^ n2604 ^ n2173 ;
  assign n2608 = n2607 ^ n2606 ^ n2278 ;
  assign n2609 = n2608 ^ n2169 ^ n1822 ;
  assign n2613 = n2612 ^ n2609 ^ n2174 ;
  assign n2616 = n2615 ^ n2613 ^ n373 ;
  assign n2617 = ( n517 & ~n578 ) | ( n517 & n2616 ) | ( ~n578 & n2616 ) ;
  assign n2625 = n2624 ^ n2617 ^ n2234 ;
  assign n2626 = n1755 ^ n1243 ^ n486 ;
  assign n2627 = n1759 ^ n984 ^ n451 ;
  assign n2628 = n646 & n647 ;
  assign n2629 = ~n2308 & n2628 ;
  assign n2630 = ( n560 & n1725 ) | ( n560 & ~n2309 ) | ( n1725 & ~n2309 ) ;
  assign n2631 = n1184 ^ n797 ^ 1'b0 ;
  assign n2632 = n964 | n2631 ;
  assign n2635 = ~n1077 & n1752 ;
  assign n2636 = n2635 ^ n995 ^ 1'b0 ;
  assign n2637 = ( ~n1933 & n1946 ) | ( ~n1933 & n2636 ) | ( n1946 & n2636 ) ;
  assign n2633 = n2618 ^ n644 ^ x12 ;
  assign n2634 = ( n636 & n2447 ) | ( n636 & n2633 ) | ( n2447 & n2633 ) ;
  assign n2638 = n2637 ^ n2634 ^ n1243 ;
  assign n2639 = n999 & ~n2638 ;
  assign n2640 = n2632 & n2639 ;
  assign n2641 = ( ~x25 & n250 ) | ( ~x25 & n1198 ) | ( n250 & n1198 ) ;
  assign n2642 = n2641 ^ n491 ^ n331 ;
  assign n2643 = n879 | n897 ;
  assign n2644 = n2642 & ~n2643 ;
  assign n2645 = ( n267 & n368 ) | ( n267 & ~n1686 ) | ( n368 & ~n1686 ) ;
  assign n2646 = n2645 ^ n1535 ^ n383 ;
  assign n2647 = n1487 ^ x115 ^ 1'b0 ;
  assign n2648 = x111 & n2647 ;
  assign n2649 = ( ~n183 & n537 ) | ( ~n183 & n1244 ) | ( n537 & n1244 ) ;
  assign n2650 = ( n865 & ~n1237 ) | ( n865 & n2649 ) | ( ~n1237 & n2649 ) ;
  assign n2651 = ( n713 & n1302 ) | ( n713 & ~n1856 ) | ( n1302 & ~n1856 ) ;
  assign n2652 = n2651 ^ n2612 ^ n1869 ;
  assign n2656 = n1559 ^ n1147 ^ n140 ;
  assign n2657 = n2656 ^ n2381 ^ n1721 ;
  assign n2653 = ( n160 & n591 ) | ( n160 & ~n1284 ) | ( n591 & ~n1284 ) ;
  assign n2654 = ( ~n1465 & n2194 ) | ( ~n1465 & n2653 ) | ( n2194 & n2653 ) ;
  assign n2655 = n1108 | n2654 ;
  assign n2658 = n2657 ^ n2655 ^ 1'b0 ;
  assign n2659 = ( n563 & n2355 ) | ( n563 & n2658 ) | ( n2355 & n2658 ) ;
  assign n2660 = n826 | n1712 ;
  assign n2661 = n2660 ^ n1556 ^ n982 ;
  assign n2665 = n1384 ^ n438 ^ 1'b0 ;
  assign n2662 = ( ~n305 & n1496 ) | ( ~n305 & n1976 ) | ( n1496 & n1976 ) ;
  assign n2663 = ( n517 & ~n1897 ) | ( n517 & n2662 ) | ( ~n1897 & n2662 ) ;
  assign n2664 = n2663 ^ n1968 ^ n1871 ;
  assign n2666 = n2665 ^ n2664 ^ 1'b0 ;
  assign n2667 = ~n1731 & n2666 ;
  assign n2668 = ~n205 & n1294 ;
  assign n2669 = ( n2661 & n2667 ) | ( n2661 & n2668 ) | ( n2667 & n2668 ) ;
  assign n2670 = ( n2652 & n2659 ) | ( n2652 & ~n2669 ) | ( n2659 & ~n2669 ) ;
  assign n2671 = ( ~n857 & n1337 ) | ( ~n857 & n2670 ) | ( n1337 & n2670 ) ;
  assign n2685 = n137 | n2575 ;
  assign n2686 = n1580 & ~n2685 ;
  assign n2678 = n1731 ^ n1337 ^ n1016 ;
  assign n2679 = n2678 ^ n333 ^ n297 ;
  assign n2680 = ( ~n991 & n1259 ) | ( ~n991 & n2679 ) | ( n1259 & n2679 ) ;
  assign n2681 = n2680 ^ n1143 ^ x15 ;
  assign n2682 = n1821 ^ n1154 ^ n574 ;
  assign n2683 = ( n2443 & ~n2681 ) | ( n2443 & n2682 ) | ( ~n2681 & n2682 ) ;
  assign n2672 = ~n144 & n2245 ;
  assign n2673 = ~x1 & n2672 ;
  assign n2674 = ( n361 & n841 ) | ( n361 & ~n1147 ) | ( n841 & ~n1147 ) ;
  assign n2675 = n679 | n2674 ;
  assign n2676 = n2673 & ~n2675 ;
  assign n2677 = ( ~n360 & n1409 ) | ( ~n360 & n2676 ) | ( n1409 & n2676 ) ;
  assign n2684 = n2683 ^ n2677 ^ n2613 ;
  assign n2687 = n2686 ^ n2684 ^ n1659 ;
  assign n2688 = n732 & ~n2040 ;
  assign n2689 = n2688 ^ n522 ^ 1'b0 ;
  assign n2690 = ( n559 & n1062 ) | ( n559 & ~n2689 ) | ( n1062 & ~n2689 ) ;
  assign n2692 = n2485 ^ n1612 ^ n821 ;
  assign n2691 = ( ~n536 & n2257 ) | ( ~n536 & n2560 ) | ( n2257 & n2560 ) ;
  assign n2693 = n2692 ^ n2691 ^ n1181 ;
  assign n2700 = n1417 ^ n1172 ^ n283 ;
  assign n2694 = n2605 ^ n2058 ^ n1477 ;
  assign n2695 = ( n954 & n1601 ) | ( n954 & ~n1684 ) | ( n1601 & ~n1684 ) ;
  assign n2696 = ( n2017 & ~n2694 ) | ( n2017 & n2695 ) | ( ~n2694 & n2695 ) ;
  assign n2697 = ( n367 & n1162 ) | ( n367 & n2696 ) | ( n1162 & n2696 ) ;
  assign n2698 = n2697 ^ n2021 ^ n1361 ;
  assign n2699 = ( n241 & ~n273 ) | ( n241 & n2698 ) | ( ~n273 & n2698 ) ;
  assign n2701 = n2700 ^ n2699 ^ n2567 ;
  assign n2702 = n1932 & ~n2209 ;
  assign n2703 = n882 & n2702 ;
  assign n2704 = n2703 ^ n2425 ^ n1651 ;
  assign n2705 = ( n453 & n477 ) | ( n453 & n502 ) | ( n477 & n502 ) ;
  assign n2706 = ( n337 & n1282 ) | ( n337 & n1808 ) | ( n1282 & n1808 ) ;
  assign n2707 = n300 & ~n950 ;
  assign n2708 = n2707 ^ n433 ^ 1'b0 ;
  assign n2709 = ( n153 & ~n2706 ) | ( n153 & n2708 ) | ( ~n2706 & n2708 ) ;
  assign n2710 = ( n762 & n1308 ) | ( n762 & n2709 ) | ( n1308 & n2709 ) ;
  assign n2711 = n630 & n2710 ;
  assign n2712 = n2711 ^ n1597 ^ 1'b0 ;
  assign n2713 = ( ~n1783 & n2705 ) | ( ~n1783 & n2712 ) | ( n2705 & n2712 ) ;
  assign n2714 = ( n1300 & n1835 ) | ( n1300 & n2253 ) | ( n1835 & n2253 ) ;
  assign n2725 = x58 & ~n696 ;
  assign n2726 = ~n861 & n2725 ;
  assign n2727 = n2726 ^ n774 ^ 1'b0 ;
  assign n2723 = n1324 ^ n303 ^ x9 ;
  assign n2724 = n2723 ^ n1211 ^ n271 ;
  assign n2718 = n1840 ^ n1269 ^ 1'b0 ;
  assign n2719 = n1907 ^ n1209 ^ n346 ;
  assign n2720 = x24 & ~n2719 ;
  assign n2721 = n2720 ^ n1213 ^ 1'b0 ;
  assign n2722 = ( n1352 & n2718 ) | ( n1352 & ~n2721 ) | ( n2718 & ~n2721 ) ;
  assign n2728 = n2727 ^ n2724 ^ n2722 ;
  assign n2715 = x39 & x76 ;
  assign n2716 = ~n1218 & n2715 ;
  assign n2717 = ( n1592 & n1762 ) | ( n1592 & ~n2716 ) | ( n1762 & ~n2716 ) ;
  assign n2729 = n2728 ^ n2717 ^ n951 ;
  assign n2735 = ( n946 & n1374 ) | ( n946 & n2041 ) | ( n1374 & n2041 ) ;
  assign n2736 = ( n377 & n459 ) | ( n377 & ~n2735 ) | ( n459 & ~n2735 ) ;
  assign n2733 = ( x18 & n1018 ) | ( x18 & n2179 ) | ( n1018 & n2179 ) ;
  assign n2734 = n2733 ^ n1238 ^ n814 ;
  assign n2737 = n2736 ^ n2734 ^ n418 ;
  assign n2730 = n1632 ^ n638 ^ n382 ;
  assign n2731 = n2730 ^ n1844 ^ n1274 ;
  assign n2732 = n2731 ^ n850 ^ x123 ;
  assign n2738 = n2737 ^ n2732 ^ 1'b0 ;
  assign n2739 = ~n2535 & n2738 ;
  assign n2744 = n1692 ^ n424 ^ 1'b0 ;
  assign n2745 = n2744 ^ n745 ^ n738 ;
  assign n2746 = n1537 ^ n427 ^ 1'b0 ;
  assign n2747 = n2745 & ~n2746 ;
  assign n2748 = n2747 ^ n1274 ^ x68 ;
  assign n2749 = ( x109 & n969 ) | ( x109 & ~n2748 ) | ( n969 & ~n2748 ) ;
  assign n2742 = n1363 ^ n368 ^ x101 ;
  assign n2743 = ( n411 & n914 ) | ( n411 & ~n2742 ) | ( n914 & ~n2742 ) ;
  assign n2740 = n1360 ^ n715 ^ n257 ;
  assign n2741 = n2740 ^ x55 ^ 1'b0 ;
  assign n2750 = n2749 ^ n2743 ^ n2741 ;
  assign n2751 = ( n255 & ~n2678 ) | ( n255 & n2750 ) | ( ~n2678 & n2750 ) ;
  assign n2752 = ( n2008 & ~n2091 ) | ( n2008 & n2679 ) | ( ~n2091 & n2679 ) ;
  assign n2753 = ( n305 & n473 ) | ( n305 & n1919 ) | ( n473 & n1919 ) ;
  assign n2754 = ( n200 & n2752 ) | ( n200 & n2753 ) | ( n2752 & n2753 ) ;
  assign n2755 = ( n1444 & n2751 ) | ( n1444 & ~n2754 ) | ( n2751 & ~n2754 ) ;
  assign n2757 = n2453 ^ n191 ^ 1'b0 ;
  assign n2758 = n1887 & n2030 ;
  assign n2759 = n2757 & n2758 ;
  assign n2756 = n2417 ^ n326 ^ 1'b0 ;
  assign n2760 = n2759 ^ n2756 ^ n288 ;
  assign n2761 = n1838 ^ n1676 ^ x14 ;
  assign n2762 = n2761 ^ x77 ^ x8 ;
  assign n2763 = ( n1820 & n2719 ) | ( n1820 & ~n2762 ) | ( n2719 & ~n2762 ) ;
  assign n2764 = n2081 ^ n1102 ^ 1'b0 ;
  assign n2765 = x28 & ~n2764 ;
  assign n2766 = n2765 ^ n937 ^ x49 ;
  assign n2767 = n2066 ^ n1582 ^ 1'b0 ;
  assign n2768 = n1029 & n1531 ;
  assign n2769 = x98 & ~n2768 ;
  assign n2773 = n986 ^ n624 ^ 1'b0 ;
  assign n2770 = ( n291 & n320 ) | ( n291 & n982 ) | ( n320 & n982 ) ;
  assign n2771 = n2770 ^ n532 ^ x20 ;
  assign n2772 = n1391 | n2771 ;
  assign n2774 = n2773 ^ n2772 ^ 1'b0 ;
  assign n2775 = ( n922 & n1614 ) | ( n922 & ~n2774 ) | ( n1614 & ~n2774 ) ;
  assign n2776 = ( n477 & n647 ) | ( n477 & ~n1693 ) | ( n647 & ~n1693 ) ;
  assign n2777 = ( ~n2769 & n2775 ) | ( ~n2769 & n2776 ) | ( n2775 & n2776 ) ;
  assign n2778 = n1626 ^ n1401 ^ n1299 ;
  assign n2779 = ( n873 & n2353 ) | ( n873 & ~n2778 ) | ( n2353 & ~n2778 ) ;
  assign n2780 = n1482 ^ n361 ^ x27 ;
  assign n2781 = n2780 ^ n1403 ^ n1373 ;
  assign n2782 = ( n1695 & n2494 ) | ( n1695 & n2781 ) | ( n2494 & n2781 ) ;
  assign n2783 = n1621 & n2782 ;
  assign n2784 = n2779 & n2783 ;
  assign n2785 = ( ~x124 & n343 ) | ( ~x124 & n1925 ) | ( n343 & n1925 ) ;
  assign n2786 = ( n2018 & n2385 ) | ( n2018 & n2785 ) | ( n2385 & n2785 ) ;
  assign n2787 = ( n2287 & n2661 ) | ( n2287 & n2786 ) | ( n2661 & n2786 ) ;
  assign n2788 = ( n546 & n2784 ) | ( n546 & ~n2787 ) | ( n2784 & ~n2787 ) ;
  assign n2789 = n526 ^ x36 ^ 1'b0 ;
  assign n2790 = ~n1009 & n2789 ;
  assign n2791 = ( n1571 & ~n1849 ) | ( n1571 & n2790 ) | ( ~n1849 & n2790 ) ;
  assign n2792 = n2505 | n2791 ;
  assign n2793 = n2792 ^ n541 ^ 1'b0 ;
  assign n2794 = n2008 ^ n1330 ^ n1261 ;
  assign n2795 = n2597 ^ n1932 ^ n136 ;
  assign n2796 = n2795 ^ n401 ^ n278 ;
  assign n2811 = ( n472 & n783 ) | ( n472 & n1486 ) | ( n783 & n1486 ) ;
  assign n2809 = n1337 | n2726 ;
  assign n2810 = n2809 ^ n1511 ^ 1'b0 ;
  assign n2812 = n2811 ^ n2810 ^ n157 ;
  assign n2806 = n788 ^ n644 ^ n393 ;
  assign n2807 = ( x76 & n969 ) | ( x76 & ~n2806 ) | ( n969 & ~n2806 ) ;
  assign n2808 = ( x64 & n746 ) | ( x64 & ~n2807 ) | ( n746 & ~n2807 ) ;
  assign n2813 = n2812 ^ n2808 ^ n1064 ;
  assign n2814 = n1768 | n2813 ;
  assign n2800 = n1291 ^ n1057 ^ 1'b0 ;
  assign n2801 = ~n2708 & n2800 ;
  assign n2797 = n679 ^ n447 ^ x27 ;
  assign n2798 = ( n1282 & n2221 ) | ( n1282 & n2351 ) | ( n2221 & n2351 ) ;
  assign n2799 = n2797 & n2798 ;
  assign n2802 = n2801 ^ n2799 ^ 1'b0 ;
  assign n2803 = ( ~n274 & n731 ) | ( ~n274 & n949 ) | ( n731 & n949 ) ;
  assign n2804 = ( n147 & n2802 ) | ( n147 & ~n2803 ) | ( n2802 & ~n2803 ) ;
  assign n2805 = ( n762 & n1929 ) | ( n762 & ~n2804 ) | ( n1929 & ~n2804 ) ;
  assign n2815 = n2814 ^ n2805 ^ n2784 ;
  assign n2819 = ( n491 & n1113 ) | ( n491 & ~n2238 ) | ( n1113 & ~n2238 ) ;
  assign n2820 = ( x12 & n244 ) | ( x12 & n2819 ) | ( n244 & n2819 ) ;
  assign n2818 = n305 | n1048 ;
  assign n2821 = n2820 ^ n2818 ^ 1'b0 ;
  assign n2816 = n2663 ^ n1535 ^ n961 ;
  assign n2817 = ~n2538 & n2816 ;
  assign n2822 = n2821 ^ n2817 ^ 1'b0 ;
  assign n2824 = ( ~n191 & n585 ) | ( ~n191 & n1505 ) | ( n585 & n1505 ) ;
  assign n2823 = x79 & ~x114 ;
  assign n2825 = n2824 ^ n2823 ^ n1727 ;
  assign n2826 = ( n1217 & n2633 ) | ( n1217 & ~n2825 ) | ( n2633 & ~n2825 ) ;
  assign n2834 = n628 ^ n168 ^ x16 ;
  assign n2835 = x117 & ~n2834 ;
  assign n2827 = n606 ^ n510 ^ 1'b0 ;
  assign n2828 = n1158 & n2827 ;
  assign n2829 = n874 & n2395 ;
  assign n2830 = ~n2828 & n2829 ;
  assign n2831 = ~n387 & n737 ;
  assign n2832 = n2511 | n2831 ;
  assign n2833 = n2830 & ~n2832 ;
  assign n2836 = n2835 ^ n2833 ^ n1318 ;
  assign n2842 = n1204 ^ n1083 ^ 1'b0 ;
  assign n2843 = n2842 ^ n1709 ^ n595 ;
  assign n2844 = n2843 ^ n1302 ^ n1075 ;
  assign n2837 = n137 & n245 ;
  assign n2838 = ( n1300 & n1994 ) | ( n1300 & n2837 ) | ( n1994 & n2837 ) ;
  assign n2839 = ( n460 & n2263 ) | ( n460 & n2838 ) | ( n2263 & n2838 ) ;
  assign n2840 = n2678 ^ n2657 ^ x83 ;
  assign n2841 = n2839 & ~n2840 ;
  assign n2845 = n2844 ^ n2841 ^ 1'b0 ;
  assign n2852 = n2605 ^ n1047 ^ n137 ;
  assign n2853 = n2852 ^ n1172 ^ n923 ;
  assign n2854 = n2853 ^ n1822 ^ n130 ;
  assign n2850 = ( x116 & ~n1167 ) | ( x116 & n1846 ) | ( ~n1167 & n1846 ) ;
  assign n2847 = n2100 ^ n893 ^ x122 ;
  assign n2848 = n2223 & n2335 ;
  assign n2849 = ( n800 & n2847 ) | ( n800 & ~n2848 ) | ( n2847 & ~n2848 ) ;
  assign n2846 = n1470 ^ n1342 ^ n336 ;
  assign n2851 = n2850 ^ n2849 ^ n2846 ;
  assign n2855 = n2854 ^ n2851 ^ n2732 ;
  assign n2856 = ( ~n747 & n1562 ) | ( ~n747 & n2251 ) | ( n1562 & n2251 ) ;
  assign n2857 = n1718 & ~n1754 ;
  assign n2858 = n2856 & n2857 ;
  assign n2859 = n282 | n1386 ;
  assign n2860 = n2859 ^ n848 ^ 1'b0 ;
  assign n2861 = ( ~x99 & n1321 ) | ( ~x99 & n2860 ) | ( n1321 & n2860 ) ;
  assign n2862 = n2861 ^ n2266 ^ 1'b0 ;
  assign n2863 = n2862 ^ n1764 ^ n1337 ;
  assign n2864 = ( n452 & n705 ) | ( n452 & n880 ) | ( n705 & n880 ) ;
  assign n2865 = ( n628 & n1252 ) | ( n628 & n2864 ) | ( n1252 & n2864 ) ;
  assign n2866 = ( ~n1330 & n2119 ) | ( ~n1330 & n2536 ) | ( n2119 & n2536 ) ;
  assign n2867 = n1172 | n2866 ;
  assign n2868 = n171 | n2867 ;
  assign n2869 = n2000 ^ n1646 ^ n192 ;
  assign n2870 = n2869 ^ n2194 ^ n2160 ;
  assign n2871 = n2868 & n2870 ;
  assign n2872 = n1797 ^ n1178 ^ n436 ;
  assign n2873 = n2872 ^ n987 ^ n212 ;
  assign n2874 = n2227 ^ n400 ^ x91 ;
  assign n2882 = x90 & ~n2257 ;
  assign n2883 = n1703 & ~n2882 ;
  assign n2884 = ~n761 & n2883 ;
  assign n2875 = n1003 ^ n787 ^ n213 ;
  assign n2876 = ( x75 & n219 ) | ( x75 & n616 ) | ( n219 & n616 ) ;
  assign n2877 = ( n1052 & n1147 ) | ( n1052 & n2876 ) | ( n1147 & n2876 ) ;
  assign n2878 = n2877 ^ n1575 ^ n556 ;
  assign n2879 = n2878 ^ n200 ^ n181 ;
  assign n2880 = n1555 ^ n1190 ^ n381 ;
  assign n2881 = ( n2875 & n2879 ) | ( n2875 & ~n2880 ) | ( n2879 & ~n2880 ) ;
  assign n2885 = n2884 ^ n2881 ^ n2489 ;
  assign n2886 = n2885 ^ n1366 ^ 1'b0 ;
  assign n2887 = n2874 | n2886 ;
  assign n2900 = ( ~n490 & n771 ) | ( ~n490 & n1784 ) | ( n771 & n1784 ) ;
  assign n2901 = n2900 ^ n981 ^ n370 ;
  assign n2902 = n2901 ^ n1742 ^ n1569 ;
  assign n2896 = ( x97 & n388 ) | ( x97 & ~n523 ) | ( n388 & ~n523 ) ;
  assign n2897 = n2896 ^ n1137 ^ n662 ;
  assign n2898 = n2897 ^ n2383 ^ 1'b0 ;
  assign n2888 = n791 ^ n432 ^ x112 ;
  assign n2889 = ( x26 & n292 ) | ( x26 & ~n2888 ) | ( n292 & ~n2888 ) ;
  assign n2890 = ( n1580 & ~n1756 ) | ( n1580 & n2510 ) | ( ~n1756 & n2510 ) ;
  assign n2891 = ( ~n220 & n2083 ) | ( ~n220 & n2552 ) | ( n2083 & n2552 ) ;
  assign n2892 = ( n187 & n1533 ) | ( n187 & ~n2891 ) | ( n1533 & ~n2891 ) ;
  assign n2893 = ( n1634 & n2890 ) | ( n1634 & ~n2892 ) | ( n2890 & ~n2892 ) ;
  assign n2894 = n2889 & n2893 ;
  assign n2895 = n2894 ^ n1558 ^ n1269 ;
  assign n2899 = n2898 ^ n2895 ^ n730 ;
  assign n2903 = n2902 ^ n2899 ^ n366 ;
  assign n2904 = ( n2873 & n2887 ) | ( n2873 & n2903 ) | ( n2887 & n2903 ) ;
  assign n2909 = n200 & n2828 ;
  assign n2910 = n2909 ^ n960 ^ 1'b0 ;
  assign n2906 = n291 | n670 ;
  assign n2907 = n2906 ^ n1821 ^ n1715 ;
  assign n2905 = n1653 ^ n238 ^ 1'b0 ;
  assign n2908 = n2907 ^ n2905 ^ n2589 ;
  assign n2911 = n2910 ^ n2908 ^ n821 ;
  assign n2925 = n2441 ^ n2181 ^ n744 ;
  assign n2926 = ~n743 & n2257 ;
  assign n2927 = ~n2925 & n2926 ;
  assign n2923 = ( x104 & n1482 ) | ( x104 & n2180 ) | ( n1482 & n2180 ) ;
  assign n2924 = n2923 ^ n1626 ^ n1178 ;
  assign n2921 = n2172 ^ x114 ^ 1'b0 ;
  assign n2917 = ( n204 & n393 ) | ( n204 & ~n510 ) | ( n393 & ~n510 ) ;
  assign n2918 = ( n632 & n2795 ) | ( n632 & ~n2917 ) | ( n2795 & ~n2917 ) ;
  assign n2919 = ( ~n281 & n639 ) | ( ~n281 & n1664 ) | ( n639 & n1664 ) ;
  assign n2920 = ~n2918 & n2919 ;
  assign n2912 = ( x103 & n273 ) | ( x103 & ~n2745 ) | ( n273 & ~n2745 ) ;
  assign n2913 = ( n1135 & n1246 ) | ( n1135 & ~n2790 ) | ( n1246 & ~n2790 ) ;
  assign n2914 = n2913 ^ n1432 ^ n760 ;
  assign n2915 = ( n2560 & ~n2912 ) | ( n2560 & n2914 ) | ( ~n2912 & n2914 ) ;
  assign n2916 = ( ~n254 & n805 ) | ( ~n254 & n2915 ) | ( n805 & n2915 ) ;
  assign n2922 = n2921 ^ n2920 ^ n2916 ;
  assign n2928 = n2927 ^ n2924 ^ n2922 ;
  assign n2930 = ( n282 & n360 ) | ( n282 & ~n750 ) | ( n360 & ~n750 ) ;
  assign n2931 = n2930 ^ n1752 ^ n637 ;
  assign n2929 = n1759 ^ n1639 ^ x113 ;
  assign n2932 = n2931 ^ n2929 ^ x118 ;
  assign n2933 = ( n2170 & n2592 ) | ( n2170 & n2932 ) | ( n2592 & n2932 ) ;
  assign n2934 = ( n721 & n1324 ) | ( n721 & n1524 ) | ( n1324 & n1524 ) ;
  assign n2935 = ( n499 & n551 ) | ( n499 & ~n2934 ) | ( n551 & ~n2934 ) ;
  assign n2936 = ( ~n513 & n1190 ) | ( ~n513 & n2935 ) | ( n1190 & n2935 ) ;
  assign n2942 = n183 & n1846 ;
  assign n2941 = ( n1080 & ~n2177 ) | ( n1080 & n2581 ) | ( ~n2177 & n2581 ) ;
  assign n2937 = ( n362 & n1788 ) | ( n362 & ~n2094 ) | ( n1788 & ~n2094 ) ;
  assign n2938 = n2937 ^ n2048 ^ n519 ;
  assign n2939 = n1154 & ~n2938 ;
  assign n2940 = n2939 ^ n980 ^ 1'b0 ;
  assign n2943 = n2942 ^ n2941 ^ n2940 ;
  assign n2950 = n1690 ^ n719 ^ 1'b0 ;
  assign n2951 = n245 & ~n2950 ;
  assign n2952 = n2733 ^ n1997 ^ n718 ;
  assign n2953 = ( x126 & ~n2951 ) | ( x126 & n2952 ) | ( ~n2951 & n2952 ) ;
  assign n2944 = ( n617 & n1295 ) | ( n617 & ~n2114 ) | ( n1295 & ~n2114 ) ;
  assign n2945 = n1694 ^ n287 ^ x28 ;
  assign n2946 = n2945 ^ n1791 ^ n1436 ;
  assign n2947 = ( ~n1520 & n1794 ) | ( ~n1520 & n2151 ) | ( n1794 & n2151 ) ;
  assign n2948 = ( n2944 & ~n2946 ) | ( n2944 & n2947 ) | ( ~n2946 & n2947 ) ;
  assign n2949 = ( ~n281 & n2081 ) | ( ~n281 & n2948 ) | ( n2081 & n2948 ) ;
  assign n2954 = n2953 ^ n2949 ^ n705 ;
  assign n2959 = ( n282 & ~n322 ) | ( n282 & n389 ) | ( ~n322 & n389 ) ;
  assign n2958 = n1472 ^ n725 ^ n390 ;
  assign n2960 = n2959 ^ n2958 ^ n2369 ;
  assign n2956 = ( n153 & ~n1964 ) | ( n153 & n1998 ) | ( ~n1964 & n1998 ) ;
  assign n2957 = ( n1205 & ~n2513 ) | ( n1205 & n2956 ) | ( ~n2513 & n2956 ) ;
  assign n2955 = n1616 ^ n657 ^ 1'b0 ;
  assign n2961 = n2960 ^ n2957 ^ n2955 ;
  assign n2962 = ( n722 & n1632 ) | ( n722 & ~n1770 ) | ( n1632 & ~n1770 ) ;
  assign n2963 = n2962 ^ n1306 ^ n601 ;
  assign n2964 = n2963 ^ n1009 ^ n752 ;
  assign n2965 = ( n725 & ~n1425 ) | ( n725 & n2964 ) | ( ~n1425 & n2964 ) ;
  assign n2966 = n1460 ^ n1203 ^ n863 ;
  assign n2967 = ( n1450 & n1630 ) | ( n1450 & n2966 ) | ( n1630 & n2966 ) ;
  assign n2968 = ( n2724 & n2965 ) | ( n2724 & ~n2967 ) | ( n2965 & ~n2967 ) ;
  assign n2969 = n1965 ^ n903 ^ n239 ;
  assign n2971 = n1657 ^ n555 ^ n247 ;
  assign n2972 = n2665 ^ n1632 ^ 1'b0 ;
  assign n2973 = n2971 | n2972 ;
  assign n2970 = n1089 ^ n696 ^ x88 ;
  assign n2974 = n2973 ^ n2970 ^ n2151 ;
  assign n2975 = n499 | n934 ;
  assign n2976 = n937 & n1261 ;
  assign n2977 = ( ~x58 & n394 ) | ( ~x58 & n2976 ) | ( n394 & n2976 ) ;
  assign n2978 = n2977 ^ n2287 ^ n1072 ;
  assign n2979 = n1998 | n2978 ;
  assign n2980 = n2975 & ~n2979 ;
  assign n2981 = n2363 ^ n1968 ^ n469 ;
  assign n2982 = ~n2980 & n2981 ;
  assign n2983 = n2982 ^ n807 ^ 1'b0 ;
  assign n2984 = ~n1664 & n2983 ;
  assign n2985 = ( n2969 & n2974 ) | ( n2969 & ~n2984 ) | ( n2974 & ~n2984 ) ;
  assign n2999 = ( n562 & ~n637 ) | ( n562 & n789 ) | ( ~n637 & n789 ) ;
  assign n2993 = n1146 ^ n938 ^ n261 ;
  assign n2994 = n1730 ^ x6 ^ 1'b0 ;
  assign n2995 = x89 & ~n2994 ;
  assign n2996 = ( n392 & n2993 ) | ( n392 & ~n2995 ) | ( n2993 & ~n2995 ) ;
  assign n2997 = n2996 ^ n1788 ^ n1188 ;
  assign n2998 = n2997 ^ n2219 ^ n376 ;
  assign n3000 = n2999 ^ n2998 ^ n1947 ;
  assign n3001 = n812 | n3000 ;
  assign n3002 = n3001 ^ n2920 ^ 1'b0 ;
  assign n2989 = n960 ^ n834 ^ x48 ;
  assign n2990 = n780 & n2572 ;
  assign n2991 = n2990 ^ n1732 ^ 1'b0 ;
  assign n2992 = ( n1505 & n2989 ) | ( n1505 & ~n2991 ) | ( n2989 & ~n2991 ) ;
  assign n2986 = ( n429 & ~n778 ) | ( n429 & n1087 ) | ( ~n778 & n1087 ) ;
  assign n2987 = n2986 ^ n1490 ^ n1102 ;
  assign n2988 = n2987 ^ n2971 ^ n2171 ;
  assign n3003 = n3002 ^ n2992 ^ n2988 ;
  assign n3004 = ( ~n760 & n848 ) | ( ~n760 & n1819 ) | ( n848 & n1819 ) ;
  assign n3005 = n3004 ^ n2515 ^ 1'b0 ;
  assign n3006 = x34 & n330 ;
  assign n3007 = n3006 ^ x44 ^ 1'b0 ;
  assign n3008 = ( n791 & n2116 ) | ( n791 & ~n3007 ) | ( n2116 & ~n3007 ) ;
  assign n3019 = n2820 ^ n372 ^ n191 ;
  assign n3018 = ( n787 & n1530 ) | ( n787 & n1633 ) | ( n1530 & n1633 ) ;
  assign n3020 = n3019 ^ n3018 ^ n2255 ;
  assign n3009 = n628 | n1548 ;
  assign n3011 = ( n1147 & n1988 ) | ( n1147 & ~n2208 ) | ( n1988 & ~n2208 ) ;
  assign n3012 = n3011 ^ n673 ^ n195 ;
  assign n3010 = ( ~n459 & n1697 ) | ( ~n459 & n2946 ) | ( n1697 & n2946 ) ;
  assign n3013 = n3012 ^ n3010 ^ n1261 ;
  assign n3014 = n3013 ^ n878 ^ 1'b0 ;
  assign n3015 = n3014 ^ n1930 ^ 1'b0 ;
  assign n3016 = n3009 & ~n3015 ;
  assign n3017 = ~n2838 & n3016 ;
  assign n3021 = n3020 ^ n3017 ^ 1'b0 ;
  assign n3028 = ( x11 & ~x65 ) | ( x11 & n342 ) | ( ~x65 & n342 ) ;
  assign n3029 = n1433 ^ n687 ^ n537 ;
  assign n3030 = ( n904 & n3028 ) | ( n904 & n3029 ) | ( n3028 & n3029 ) ;
  assign n3031 = ( ~n475 & n2119 ) | ( ~n475 & n3030 ) | ( n2119 & n3030 ) ;
  assign n3022 = ( n191 & ~n1324 ) | ( n191 & n1580 ) | ( ~n1324 & n1580 ) ;
  assign n3023 = ( n376 & n398 ) | ( n376 & ~n1151 ) | ( n398 & ~n1151 ) ;
  assign n3024 = n953 & ~n2321 ;
  assign n3025 = ~n3023 & n3024 ;
  assign n3026 = ( ~n471 & n3022 ) | ( ~n471 & n3025 ) | ( n3022 & n3025 ) ;
  assign n3027 = ~n1961 & n3026 ;
  assign n3032 = n3031 ^ n3027 ^ 1'b0 ;
  assign n3034 = n1029 ^ n205 ^ n131 ;
  assign n3035 = n3034 ^ n2910 ^ n278 ;
  assign n3033 = ( n258 & n1739 ) | ( n258 & ~n1757 ) | ( n1739 & ~n1757 ) ;
  assign n3036 = n3035 ^ n3033 ^ n195 ;
  assign n3039 = ( n787 & n887 ) | ( n787 & ~n1582 ) | ( n887 & ~n1582 ) ;
  assign n3037 = ( n157 & ~n1103 ) | ( n157 & n2309 ) | ( ~n1103 & n2309 ) ;
  assign n3038 = n777 & n3037 ;
  assign n3040 = n3039 ^ n3038 ^ 1'b0 ;
  assign n3041 = n3040 ^ n2501 ^ n1039 ;
  assign n3042 = ( n1049 & ~n3036 ) | ( n1049 & n3041 ) | ( ~n3036 & n3041 ) ;
  assign n3046 = n791 ^ n584 ^ n578 ;
  assign n3047 = n1581 ^ n456 ^ n261 ;
  assign n3048 = n3047 ^ n739 ^ n608 ;
  assign n3049 = n3048 ^ n1359 ^ n677 ;
  assign n3050 = n3049 ^ n456 ^ 1'b0 ;
  assign n3051 = n3046 | n3050 ;
  assign n3043 = ( n313 & ~n622 ) | ( n313 & n2492 ) | ( ~n622 & n2492 ) ;
  assign n3044 = n3043 ^ n800 ^ n467 ;
  assign n3045 = n2569 & ~n3044 ;
  assign n3052 = n3051 ^ n3045 ^ 1'b0 ;
  assign n3059 = x20 | n838 ;
  assign n3060 = n3059 ^ n2999 ^ n947 ;
  assign n3053 = n400 ^ x16 ^ 1'b0 ;
  assign n3054 = n3053 ^ n3012 ^ n2864 ;
  assign n3055 = ( ~n681 & n1586 ) | ( ~n681 & n3054 ) | ( n1586 & n3054 ) ;
  assign n3056 = n2475 ^ n1264 ^ 1'b0 ;
  assign n3057 = n3056 ^ n2797 ^ n2217 ;
  assign n3058 = ( ~n507 & n3055 ) | ( ~n507 & n3057 ) | ( n3055 & n3057 ) ;
  assign n3061 = n3060 ^ n3058 ^ n3052 ;
  assign n3062 = x62 & n956 ;
  assign n3063 = ~n1261 & n3062 ;
  assign n3064 = n1486 ^ x53 ^ 1'b0 ;
  assign n3065 = ( n2663 & n3063 ) | ( n2663 & ~n3064 ) | ( n3063 & ~n3064 ) ;
  assign n3066 = ( ~x63 & n347 ) | ( ~x63 & n834 ) | ( n347 & n834 ) ;
  assign n3067 = ( n506 & ~n767 ) | ( n506 & n3066 ) | ( ~n767 & n3066 ) ;
  assign n3068 = ( n1786 & n2872 ) | ( n1786 & ~n3067 ) | ( n2872 & ~n3067 ) ;
  assign n3069 = n3068 ^ n409 ^ n320 ;
  assign n3070 = n1161 ^ n242 ^ n146 ;
  assign n3071 = ( n516 & ~n1644 ) | ( n516 & n2652 ) | ( ~n1644 & n2652 ) ;
  assign n3072 = ( n477 & n3070 ) | ( n477 & ~n3071 ) | ( n3070 & ~n3071 ) ;
  assign n3073 = n1758 ^ n785 ^ x56 ;
  assign n3074 = ( n602 & ~n1693 ) | ( n602 & n3073 ) | ( ~n1693 & n3073 ) ;
  assign n3075 = ( ~n1874 & n2473 ) | ( ~n1874 & n2623 ) | ( n2473 & n2623 ) ;
  assign n3076 = n3075 ^ n1596 ^ 1'b0 ;
  assign n3077 = ~n3074 & n3076 ;
  assign n3078 = ( ~n639 & n2913 ) | ( ~n639 & n3077 ) | ( n2913 & n3077 ) ;
  assign n3088 = ( n810 & ~n2140 ) | ( n810 & n2641 ) | ( ~n2140 & n2641 ) ;
  assign n3079 = ( n346 & ~n1270 ) | ( n346 & n2060 ) | ( ~n1270 & n2060 ) ;
  assign n3080 = ( x82 & n232 ) | ( x82 & ~n2369 ) | ( n232 & ~n2369 ) ;
  assign n3081 = n3080 ^ n1494 ^ 1'b0 ;
  assign n3082 = ( n1897 & n2436 ) | ( n1897 & n3081 ) | ( n2436 & n3081 ) ;
  assign n3083 = n3082 ^ n1634 ^ x94 ;
  assign n3084 = n2668 ^ n1081 ^ n472 ;
  assign n3085 = n3084 ^ n1877 ^ 1'b0 ;
  assign n3086 = ( ~n517 & n3083 ) | ( ~n517 & n3085 ) | ( n3083 & n3085 ) ;
  assign n3087 = n3079 | n3086 ;
  assign n3089 = n3088 ^ n3087 ^ 1'b0 ;
  assign n3091 = x84 & ~n494 ;
  assign n3090 = n2664 ^ n2552 ^ n1968 ;
  assign n3092 = n3091 ^ n3090 ^ n1870 ;
  assign n3098 = ( ~n656 & n719 ) | ( ~n656 & n1645 ) | ( n719 & n1645 ) ;
  assign n3093 = ( n258 & ~n464 ) | ( n258 & n878 ) | ( ~n464 & n878 ) ;
  assign n3094 = ( n203 & n1654 ) | ( n203 & ~n2232 ) | ( n1654 & ~n2232 ) ;
  assign n3095 = n3094 ^ n1721 ^ n950 ;
  assign n3096 = ( n1002 & n1207 ) | ( n1002 & n1381 ) | ( n1207 & n1381 ) ;
  assign n3097 = ( n3093 & n3095 ) | ( n3093 & n3096 ) | ( n3095 & n3096 ) ;
  assign n3099 = n3098 ^ n3097 ^ n1647 ;
  assign n3100 = n2673 ^ n1201 ^ n1068 ;
  assign n3101 = ( n416 & n2297 ) | ( n416 & n2806 ) | ( n2297 & n2806 ) ;
  assign n3102 = ( n1198 & n3100 ) | ( n1198 & n3101 ) | ( n3100 & n3101 ) ;
  assign n3103 = ( ~n138 & n362 ) | ( ~n138 & n1577 ) | ( n362 & n1577 ) ;
  assign n3104 = ( ~n1557 & n2139 ) | ( ~n1557 & n3103 ) | ( n2139 & n3103 ) ;
  assign n3107 = n2296 ^ n1043 ^ n480 ;
  assign n3105 = n1642 ^ n137 ^ 1'b0 ;
  assign n3106 = n3105 ^ n1473 ^ n499 ;
  assign n3108 = n3107 ^ n3106 ^ 1'b0 ;
  assign n3109 = ~n3104 & n3108 ;
  assign n3110 = ~n1904 & n3109 ;
  assign n3111 = n3110 ^ n1775 ^ 1'b0 ;
  assign n3114 = n744 ^ n717 ^ n541 ;
  assign n3112 = x109 & n1135 ;
  assign n3113 = n704 | n3112 ;
  assign n3115 = n3114 ^ n3113 ^ n909 ;
  assign n3116 = n3115 ^ n2632 ^ 1'b0 ;
  assign n3117 = ( ~n1788 & n3111 ) | ( ~n1788 & n3116 ) | ( n3111 & n3116 ) ;
  assign n3118 = n2063 ^ n1946 ^ n707 ;
  assign n3119 = n3118 ^ n2004 ^ n256 ;
  assign n3120 = n3119 ^ n996 ^ n683 ;
  assign n3121 = n3120 ^ n2963 ^ 1'b0 ;
  assign n3122 = ( x31 & n930 ) | ( x31 & n1238 ) | ( n930 & n1238 ) ;
  assign n3123 = ( ~n1775 & n3121 ) | ( ~n1775 & n3122 ) | ( n3121 & n3122 ) ;
  assign n3124 = n1832 ^ n1661 ^ n632 ;
  assign n3125 = n3124 ^ n2375 ^ n1750 ;
  assign n3133 = n939 & n1581 ;
  assign n3130 = ~n599 & n608 ;
  assign n3131 = ~x86 & n3130 ;
  assign n3132 = n872 | n3131 ;
  assign n3127 = n1805 ^ x52 ^ 1'b0 ;
  assign n3126 = n1637 ^ n1430 ^ 1'b0 ;
  assign n3128 = n3127 ^ n3126 ^ 1'b0 ;
  assign n3129 = n3128 ^ n2230 ^ n1732 ;
  assign n3134 = n3133 ^ n3132 ^ n3129 ;
  assign n3135 = n2670 ^ n1665 ^ x124 ;
  assign n3144 = n636 ^ n431 ^ x63 ;
  assign n3136 = ( n391 & n612 ) | ( n391 & ~n994 ) | ( n612 & ~n994 ) ;
  assign n3137 = ( x116 & n437 ) | ( x116 & n3136 ) | ( n437 & n3136 ) ;
  assign n3138 = ( ~n492 & n1326 ) | ( ~n492 & n2971 ) | ( n1326 & n2971 ) ;
  assign n3139 = ( n2878 & n3137 ) | ( n2878 & n3138 ) | ( n3137 & n3138 ) ;
  assign n3140 = n1155 ^ n983 ^ 1'b0 ;
  assign n3141 = n1377 | n3140 ;
  assign n3142 = ( ~n704 & n3139 ) | ( ~n704 & n3141 ) | ( n3139 & n3141 ) ;
  assign n3143 = n3142 ^ n2060 ^ n913 ;
  assign n3145 = n3144 ^ n3143 ^ n734 ;
  assign n3146 = n168 & n367 ;
  assign n3147 = ~n295 & n3146 ;
  assign n3148 = ( x102 & n559 ) | ( x102 & ~n1974 ) | ( n559 & ~n1974 ) ;
  assign n3149 = n3148 ^ n1720 ^ n941 ;
  assign n3150 = n3149 ^ n331 ^ n136 ;
  assign n3151 = n2490 & n3150 ;
  assign n3152 = n3147 & n3151 ;
  assign n3163 = n2560 ^ n1407 ^ n257 ;
  assign n3159 = n783 ^ n362 ^ n257 ;
  assign n3160 = n2373 ^ n1240 ^ x74 ;
  assign n3161 = ( x54 & n719 ) | ( x54 & ~n3160 ) | ( n719 & ~n3160 ) ;
  assign n3162 = ( n1192 & n3159 ) | ( n1192 & n3161 ) | ( n3159 & n3161 ) ;
  assign n3158 = n3144 ^ n829 ^ n541 ;
  assign n3164 = n3163 ^ n3162 ^ n3158 ;
  assign n3153 = n1422 ^ n841 ^ x29 ;
  assign n3154 = n3153 ^ n2373 ^ n1710 ;
  assign n3155 = n219 & ~n718 ;
  assign n3156 = ~n2583 & n3155 ;
  assign n3157 = n3154 | n3156 ;
  assign n3165 = n3164 ^ n3157 ^ 1'b0 ;
  assign n3166 = n3165 ^ n1013 ^ n537 ;
  assign n3169 = n414 ^ n320 ^ 1'b0 ;
  assign n3170 = ( x9 & ~n1293 ) | ( x9 & n1619 ) | ( ~n1293 & n1619 ) ;
  assign n3171 = ( ~n1707 & n3169 ) | ( ~n1707 & n3170 ) | ( n3169 & n3170 ) ;
  assign n3172 = ( n175 & n749 ) | ( n175 & n3171 ) | ( n749 & n3171 ) ;
  assign n3167 = n157 & n394 ;
  assign n3168 = ( n1705 & ~n2205 ) | ( n1705 & n3167 ) | ( ~n2205 & n3167 ) ;
  assign n3173 = n3172 ^ n3168 ^ 1'b0 ;
  assign n3174 = ( n2895 & ~n3166 ) | ( n2895 & n3173 ) | ( ~n3166 & n3173 ) ;
  assign n3175 = n221 | n2230 ;
  assign n3176 = ( n238 & n961 ) | ( n238 & ~n968 ) | ( n961 & ~n968 ) ;
  assign n3177 = n2700 ^ x56 ^ 1'b0 ;
  assign n3178 = n227 & ~n3177 ;
  assign n3179 = ( x71 & n3176 ) | ( x71 & n3178 ) | ( n3176 & n3178 ) ;
  assign n3180 = ( n1030 & n2953 ) | ( n1030 & n3179 ) | ( n2953 & n3179 ) ;
  assign n3181 = n1945 ^ n1623 ^ n1400 ;
  assign n3182 = ( n852 & n1204 ) | ( n852 & n2706 ) | ( n1204 & n2706 ) ;
  assign n3183 = n3182 ^ n1294 ^ n871 ;
  assign n3184 = n3183 ^ n1995 ^ n1085 ;
  assign n3186 = ( x23 & n235 ) | ( x23 & n534 ) | ( n235 & n534 ) ;
  assign n3185 = n1879 ^ n1140 ^ 1'b0 ;
  assign n3187 = n3186 ^ n3185 ^ n2730 ;
  assign n3188 = ( ~n1582 & n3184 ) | ( ~n1582 & n3187 ) | ( n3184 & n3187 ) ;
  assign n3189 = n3188 ^ n2184 ^ 1'b0 ;
  assign n3190 = ( n2018 & ~n3181 ) | ( n2018 & n3189 ) | ( ~n3181 & n3189 ) ;
  assign n3191 = n1183 & ~n3190 ;
  assign n3192 = ( ~n3175 & n3180 ) | ( ~n3175 & n3191 ) | ( n3180 & n3191 ) ;
  assign n3193 = n2149 & n3028 ;
  assign n3194 = n3193 ^ n607 ^ 1'b0 ;
  assign n3195 = ( n565 & n751 ) | ( n565 & ~n3194 ) | ( n751 & ~n3194 ) ;
  assign n3196 = ~n3068 & n3195 ;
  assign n3199 = ( n708 & n1692 ) | ( n708 & ~n2082 ) | ( n1692 & ~n2082 ) ;
  assign n3197 = ( n134 & ~n800 ) | ( n134 & n860 ) | ( ~n800 & n860 ) ;
  assign n3198 = n3197 ^ n755 ^ n735 ;
  assign n3200 = n3199 ^ n3198 ^ 1'b0 ;
  assign n3201 = ( n371 & n1281 ) | ( n371 & ~n1477 ) | ( n1281 & ~n1477 ) ;
  assign n3202 = n3201 ^ n1431 ^ 1'b0 ;
  assign n3203 = ( n184 & ~n2747 ) | ( n184 & n3202 ) | ( ~n2747 & n3202 ) ;
  assign n3207 = ( x77 & n214 ) | ( x77 & ~n3186 ) | ( n214 & ~n3186 ) ;
  assign n3205 = n330 ^ n166 ^ 1'b0 ;
  assign n3206 = n1408 & n3205 ;
  assign n3208 = n3207 ^ n3206 ^ n1717 ;
  assign n3204 = n168 ^ n131 ^ x117 ;
  assign n3209 = n3208 ^ n3204 ^ 1'b0 ;
  assign n3210 = n1316 & ~n3209 ;
  assign n3211 = ( n2148 & n2721 ) | ( n2148 & ~n3210 ) | ( n2721 & ~n3210 ) ;
  assign n3212 = n3211 ^ n2336 ^ n1102 ;
  assign n3218 = ( n903 & n1347 ) | ( n903 & ~n2330 ) | ( n1347 & ~n2330 ) ;
  assign n3213 = n2875 ^ n1360 ^ n971 ;
  assign n3214 = n3213 ^ n3179 ^ n1120 ;
  assign n3215 = ( n1686 & n2296 ) | ( n1686 & n3214 ) | ( n2296 & n3214 ) ;
  assign n3216 = ~n1017 & n3215 ;
  assign n3217 = n2094 & n3216 ;
  assign n3219 = n3218 ^ n3217 ^ 1'b0 ;
  assign n3220 = n1531 ^ n725 ^ n595 ;
  assign n3221 = n380 & n3220 ;
  assign n3222 = n1324 & n3221 ;
  assign n3223 = ( n1870 & ~n2580 ) | ( n1870 & n3222 ) | ( ~n2580 & n3222 ) ;
  assign n3224 = n1722 & ~n1770 ;
  assign n3225 = ( n137 & n261 ) | ( n137 & n1963 ) | ( n261 & n1963 ) ;
  assign n3226 = ( n132 & n735 ) | ( n132 & ~n3225 ) | ( n735 & ~n3225 ) ;
  assign n3227 = ( n3223 & ~n3224 ) | ( n3223 & n3226 ) | ( ~n3224 & n3226 ) ;
  assign n3228 = n2516 ^ n1695 ^ n1015 ;
  assign n3229 = ( ~n423 & n767 ) | ( ~n423 & n906 ) | ( n767 & n906 ) ;
  assign n3230 = n560 ^ n341 ^ x67 ;
  assign n3231 = ( n2795 & n3229 ) | ( n2795 & n3230 ) | ( n3229 & n3230 ) ;
  assign n3232 = n2966 ^ n644 ^ n496 ;
  assign n3233 = n3232 ^ n3019 ^ n2110 ;
  assign n3234 = ( n617 & ~n1447 ) | ( n617 & n3233 ) | ( ~n1447 & n3233 ) ;
  assign n3235 = ( n3228 & ~n3231 ) | ( n3228 & n3234 ) | ( ~n3231 & n3234 ) ;
  assign n3236 = ( ~n147 & n161 ) | ( ~n147 & n3235 ) | ( n161 & n3235 ) ;
  assign n3237 = ( n408 & n1511 ) | ( n408 & n3236 ) | ( n1511 & n3236 ) ;
  assign n3238 = n718 ^ n628 ^ x12 ;
  assign n3239 = n3238 ^ n2473 ^ n1724 ;
  assign n3240 = ( ~n1418 & n1802 ) | ( ~n1418 & n3239 ) | ( n1802 & n3239 ) ;
  assign n3241 = n1758 ^ n1310 ^ n223 ;
  assign n3242 = ( ~n1705 & n2434 ) | ( ~n1705 & n3241 ) | ( n2434 & n3241 ) ;
  assign n3243 = ( n1736 & ~n3240 ) | ( n1736 & n3242 ) | ( ~n3240 & n3242 ) ;
  assign n3244 = ~n629 & n1637 ;
  assign n3245 = ( n1302 & n3243 ) | ( n1302 & n3244 ) | ( n3243 & n3244 ) ;
  assign n3246 = n3245 ^ n2659 ^ n956 ;
  assign n3249 = n2710 ^ n1472 ^ n223 ;
  assign n3247 = ( x46 & ~n198 ) | ( x46 & n769 ) | ( ~n198 & n769 ) ;
  assign n3248 = n3247 ^ n2580 ^ n2093 ;
  assign n3250 = n3249 ^ n3248 ^ n1697 ;
  assign n3251 = n3250 ^ n2135 ^ n709 ;
  assign n3254 = ( n430 & n474 ) | ( n430 & ~n549 ) | ( n474 & ~n549 ) ;
  assign n3253 = ( n199 & ~n525 ) | ( n199 & n805 ) | ( ~n525 & n805 ) ;
  assign n3255 = n3254 ^ n3253 ^ n2239 ;
  assign n3256 = ( n195 & n359 ) | ( n195 & ~n3255 ) | ( n359 & ~n3255 ) ;
  assign n3257 = n1376 ^ n800 ^ n460 ;
  assign n3258 = ( ~n242 & n3256 ) | ( ~n242 & n3257 ) | ( n3256 & n3257 ) ;
  assign n3259 = n3258 ^ n2373 ^ n881 ;
  assign n3252 = ( n1461 & n2613 ) | ( n1461 & n3004 ) | ( n2613 & n3004 ) ;
  assign n3260 = n3259 ^ n3252 ^ 1'b0 ;
  assign n3261 = n1973 ^ n568 ^ n474 ;
  assign n3262 = n3261 ^ n936 ^ 1'b0 ;
  assign n3263 = n2315 & ~n3262 ;
  assign n3264 = n1559 ^ n830 ^ n385 ;
  assign n3265 = ( n2243 & n3263 ) | ( n2243 & ~n3264 ) | ( n3263 & ~n3264 ) ;
  assign n3266 = n3265 ^ n1844 ^ n1507 ;
  assign n3268 = ( ~n335 & n799 ) | ( ~n335 & n1819 ) | ( n799 & n1819 ) ;
  assign n3269 = n3268 ^ n393 ^ 1'b0 ;
  assign n3267 = n1370 ^ n1351 ^ n1155 ;
  assign n3270 = n3269 ^ n3267 ^ n1277 ;
  assign n3285 = n137 | n2732 ;
  assign n3271 = n2708 ^ n1273 ^ n977 ;
  assign n3272 = n3271 ^ n2912 ^ n2769 ;
  assign n3273 = n1447 | n3272 ;
  assign n3274 = n3273 ^ n2365 ^ 1'b0 ;
  assign n3279 = ~n468 & n953 ;
  assign n3280 = n2111 & n3279 ;
  assign n3275 = n3093 ^ n2733 ^ n1552 ;
  assign n3276 = n3275 ^ n1161 ^ n1062 ;
  assign n3277 = ( n679 & n2465 ) | ( n679 & n3276 ) | ( n2465 & n3276 ) ;
  assign n3278 = n3277 ^ n506 ^ n250 ;
  assign n3281 = n3280 ^ n3278 ^ n1556 ;
  assign n3282 = ( n706 & n3274 ) | ( n706 & ~n3281 ) | ( n3274 & ~n3281 ) ;
  assign n3283 = n3282 ^ n2813 ^ n2450 ;
  assign n3284 = ( ~n300 & n1509 ) | ( ~n300 & n3283 ) | ( n1509 & n3283 ) ;
  assign n3286 = n3285 ^ n3284 ^ n2440 ;
  assign n3291 = n1369 ^ n1308 ^ n905 ;
  assign n3289 = ( n199 & n298 ) | ( n199 & ~n1124 ) | ( n298 & ~n1124 ) ;
  assign n3287 = n2365 ^ n2320 ^ n1947 ;
  assign n3288 = ( x68 & n2515 ) | ( x68 & n3287 ) | ( n2515 & n3287 ) ;
  assign n3290 = n3289 ^ n3288 ^ n129 ;
  assign n3292 = n3291 ^ n3290 ^ n133 ;
  assign n3293 = n719 ^ n599 ^ x55 ;
  assign n3294 = n3293 ^ n443 ^ 1'b0 ;
  assign n3295 = n1397 | n2040 ;
  assign n3296 = n3295 ^ n1283 ^ 1'b0 ;
  assign n3297 = n3296 ^ n1324 ^ 1'b0 ;
  assign n3298 = ( ~n730 & n1133 ) | ( ~n730 & n1331 ) | ( n1133 & n1331 ) ;
  assign n3299 = n3298 ^ n1619 ^ 1'b0 ;
  assign n3300 = ~n1506 & n3299 ;
  assign n3301 = ~n2377 & n3300 ;
  assign n3302 = ( n414 & ~n3297 ) | ( n414 & n3301 ) | ( ~n3297 & n3301 ) ;
  assign n3303 = ( n1741 & n3294 ) | ( n1741 & ~n3302 ) | ( n3294 & ~n3302 ) ;
  assign n3311 = ( x42 & n747 ) | ( x42 & ~n871 ) | ( n747 & ~n871 ) ;
  assign n3312 = n3311 ^ n841 ^ 1'b0 ;
  assign n3313 = n3312 ^ n787 ^ n193 ;
  assign n3309 = x44 & ~n418 ;
  assign n3310 = ~n207 & n3309 ;
  assign n3314 = n3313 ^ n3310 ^ n1489 ;
  assign n3315 = ( ~n873 & n1118 ) | ( ~n873 & n3314 ) | ( n1118 & n3314 ) ;
  assign n3316 = n3315 ^ n2066 ^ 1'b0 ;
  assign n3304 = ( ~n816 & n1137 ) | ( ~n816 & n2263 ) | ( n1137 & n2263 ) ;
  assign n3305 = n3304 ^ n2452 ^ n727 ;
  assign n3306 = ( n1246 & n1395 ) | ( n1246 & ~n2924 ) | ( n1395 & ~n2924 ) ;
  assign n3307 = n3306 ^ n2149 ^ n1511 ;
  assign n3308 = ( n620 & n3305 ) | ( n620 & n3307 ) | ( n3305 & n3307 ) ;
  assign n3317 = n3316 ^ n3308 ^ 1'b0 ;
  assign n3318 = n1400 ^ n1212 ^ n133 ;
  assign n3319 = ( ~n1091 & n1954 ) | ( ~n1091 & n2723 ) | ( n1954 & n2723 ) ;
  assign n3320 = ( n1609 & ~n3318 ) | ( n1609 & n3319 ) | ( ~n3318 & n3319 ) ;
  assign n3321 = ( x101 & n191 ) | ( x101 & ~n3320 ) | ( n191 & ~n3320 ) ;
  assign n3322 = ~n1426 & n2633 ;
  assign n3323 = ( n134 & n554 ) | ( n134 & ~n685 ) | ( n554 & ~n685 ) ;
  assign n3324 = ( x18 & n539 ) | ( x18 & n2975 ) | ( n539 & n2975 ) ;
  assign n3325 = ( n689 & n3323 ) | ( n689 & ~n3324 ) | ( n3323 & ~n3324 ) ;
  assign n3326 = ~n445 & n3325 ;
  assign n3327 = ~n1647 & n3326 ;
  assign n3328 = n3327 ^ n2727 ^ n2016 ;
  assign n3329 = n2218 ^ n1793 ^ n1376 ;
  assign n3330 = ( ~n213 & n2204 ) | ( ~n213 & n3329 ) | ( n2204 & n3329 ) ;
  assign n3331 = ( n257 & n771 ) | ( n257 & ~n2408 ) | ( n771 & ~n2408 ) ;
  assign n3332 = ( n305 & n1995 ) | ( n305 & n3331 ) | ( n1995 & n3331 ) ;
  assign n3333 = ( n1026 & n3141 ) | ( n1026 & n3332 ) | ( n3141 & n3332 ) ;
  assign n3334 = ( n812 & ~n2962 ) | ( n812 & n3333 ) | ( ~n2962 & n3333 ) ;
  assign n3335 = ( n265 & ~n3330 ) | ( n265 & n3334 ) | ( ~n3330 & n3334 ) ;
  assign n3336 = n3000 ^ n1712 ^ 1'b0 ;
  assign n3337 = n1400 & ~n3336 ;
  assign n3338 = ( n1878 & ~n2793 ) | ( n1878 & n3337 ) | ( ~n2793 & n3337 ) ;
  assign n3339 = n3232 ^ n2913 ^ n1988 ;
  assign n3340 = n1233 & n2600 ;
  assign n3341 = ~n2027 & n3340 ;
  assign n3342 = n3339 & n3341 ;
  assign n3343 = ( n1225 & n3171 ) | ( n1225 & ~n3342 ) | ( n3171 & ~n3342 ) ;
  assign n3344 = ( n3335 & n3338 ) | ( n3335 & n3343 ) | ( n3338 & n3343 ) ;
  assign n3345 = n1016 ^ n543 ^ 1'b0 ;
  assign n3346 = n2842 | n3345 ;
  assign n3347 = ( ~n495 & n1399 ) | ( ~n495 & n3346 ) | ( n1399 & n3346 ) ;
  assign n3362 = n1757 ^ n745 ^ n278 ;
  assign n3360 = n2433 ^ n1012 ^ n333 ;
  assign n3361 = n3360 ^ n1208 ^ n459 ;
  assign n3363 = n3362 ^ n3361 ^ n619 ;
  assign n3355 = n2230 ^ n1797 ^ 1'b0 ;
  assign n3356 = x33 & n3355 ;
  assign n3357 = n1350 ^ n267 ^ 1'b0 ;
  assign n3358 = ( ~n2259 & n3356 ) | ( ~n2259 & n3357 ) | ( n3356 & n3357 ) ;
  assign n3348 = n2589 ^ n471 ^ 1'b0 ;
  assign n3349 = ~n626 & n3348 ;
  assign n3350 = ~n1161 & n3137 ;
  assign n3351 = n980 & n3350 ;
  assign n3352 = ( ~n3066 & n3349 ) | ( ~n3066 & n3351 ) | ( n3349 & n3351 ) ;
  assign n3353 = ( n1888 & n2268 ) | ( n1888 & n3352 ) | ( n2268 & n3352 ) ;
  assign n3354 = ( n1747 & n3156 ) | ( n1747 & n3353 ) | ( n3156 & n3353 ) ;
  assign n3359 = n3358 ^ n3354 ^ n2747 ;
  assign n3364 = n3363 ^ n3359 ^ n1555 ;
  assign n3365 = ( n1385 & n1452 ) | ( n1385 & ~n3054 ) | ( n1452 & ~n3054 ) ;
  assign n3366 = ( x79 & n229 ) | ( x79 & ~n433 ) | ( n229 & ~n433 ) ;
  assign n3367 = n3049 ^ n1983 ^ n1063 ;
  assign n3368 = n3366 & n3367 ;
  assign n3369 = n3368 ^ n1041 ^ 1'b0 ;
  assign n3370 = ( ~n2543 & n3365 ) | ( ~n2543 & n3369 ) | ( n3365 & n3369 ) ;
  assign n3371 = ( n721 & n723 ) | ( n721 & ~n1348 ) | ( n723 & ~n1348 ) ;
  assign n3372 = ( n843 & ~n1590 ) | ( n843 & n3371 ) | ( ~n1590 & n3371 ) ;
  assign n3373 = ( ~n591 & n1069 ) | ( ~n591 & n3372 ) | ( n1069 & n3372 ) ;
  assign n3374 = n1524 ^ n1000 ^ 1'b0 ;
  assign n3375 = n3374 ^ n2671 ^ n2253 ;
  assign n3376 = ( n305 & n3373 ) | ( n305 & n3375 ) | ( n3373 & n3375 ) ;
  assign n3377 = ( n1790 & n1863 ) | ( n1790 & n2393 ) | ( n1863 & n2393 ) ;
  assign n3383 = n3142 ^ n639 ^ n572 ;
  assign n3378 = n1618 ^ n859 ^ n479 ;
  assign n3379 = ( ~x70 & n447 ) | ( ~x70 & n2820 ) | ( n447 & n2820 ) ;
  assign n3380 = n1955 ^ n1840 ^ n1161 ;
  assign n3381 = ( ~x38 & n743 ) | ( ~x38 & n3380 ) | ( n743 & n3380 ) ;
  assign n3382 = ( ~n3378 & n3379 ) | ( ~n3378 & n3381 ) | ( n3379 & n3381 ) ;
  assign n3384 = n3383 ^ n3382 ^ n1677 ;
  assign n3385 = n512 & ~n1090 ;
  assign n3386 = n1403 & n3385 ;
  assign n3387 = ( n446 & ~n1541 ) | ( n446 & n3386 ) | ( ~n1541 & n3386 ) ;
  assign n3391 = ( ~n540 & n1013 ) | ( ~n540 & n1034 ) | ( n1013 & n1034 ) ;
  assign n3388 = n1735 ^ n1383 ^ 1'b0 ;
  assign n3389 = ~n2227 & n3388 ;
  assign n3390 = n3389 ^ n1515 ^ n665 ;
  assign n3392 = n3391 ^ n3390 ^ x24 ;
  assign n3393 = n2228 & n2853 ;
  assign n3394 = n172 & n3393 ;
  assign n3395 = ( n3387 & ~n3392 ) | ( n3387 & n3394 ) | ( ~n3392 & n3394 ) ;
  assign n3404 = ( n461 & n778 ) | ( n461 & ~n1324 ) | ( n778 & ~n1324 ) ;
  assign n3405 = n946 ^ n572 ^ 1'b0 ;
  assign n3406 = n1408 & n3405 ;
  assign n3407 = ( ~n193 & n3404 ) | ( ~n193 & n3406 ) | ( n3404 & n3406 ) ;
  assign n3401 = n3225 ^ n2110 ^ n1014 ;
  assign n3402 = n3401 ^ n373 ^ n169 ;
  assign n3403 = ( x96 & n1114 ) | ( x96 & ~n3402 ) | ( n1114 & ~n3402 ) ;
  assign n3399 = n2144 & n3263 ;
  assign n3400 = ~n1294 & n3399 ;
  assign n3408 = n3407 ^ n3403 ^ n3400 ;
  assign n3409 = n3408 ^ n1736 ^ n1723 ;
  assign n3396 = ( n164 & n677 ) | ( n164 & ~n2385 ) | ( n677 & ~n2385 ) ;
  assign n3397 = n3396 ^ n1443 ^ n972 ;
  assign n3398 = ( n540 & n2804 ) | ( n540 & ~n3397 ) | ( n2804 & ~n3397 ) ;
  assign n3410 = n3409 ^ n3398 ^ n307 ;
  assign n3411 = n3410 ^ n2279 ^ n1026 ;
  assign n3412 = n915 ^ n616 ^ 1'b0 ;
  assign n3413 = ( ~n1457 & n2514 ) | ( ~n1457 & n3412 ) | ( n2514 & n3412 ) ;
  assign n3414 = n2812 ^ n211 ^ 1'b0 ;
  assign n3415 = n3414 ^ n2030 ^ n1549 ;
  assign n3416 = n3415 ^ n3266 ^ n136 ;
  assign n3417 = ( x26 & ~x42 ) | ( x26 & n2651 ) | ( ~x42 & n2651 ) ;
  assign n3418 = n864 | n3417 ;
  assign n3419 = n1975 | n3418 ;
  assign n3420 = n3419 ^ n3390 ^ n2673 ;
  assign n3421 = n2238 ^ n1388 ^ n361 ;
  assign n3422 = ( ~n3131 & n3175 ) | ( ~n3131 & n3421 ) | ( n3175 & n3421 ) ;
  assign n3423 = x29 & ~n2505 ;
  assign n3424 = n3423 ^ n749 ^ 1'b0 ;
  assign n3425 = ( x57 & n1219 ) | ( x57 & ~n3424 ) | ( n1219 & ~n3424 ) ;
  assign n3426 = ( n511 & ~n736 ) | ( n511 & n2714 ) | ( ~n736 & n2714 ) ;
  assign n3428 = ( ~n567 & n571 ) | ( ~n567 & n924 ) | ( n571 & n924 ) ;
  assign n3429 = ( ~n1860 & n2619 ) | ( ~n1860 & n3396 ) | ( n2619 & n3396 ) ;
  assign n3430 = n2223 ^ n788 ^ n771 ;
  assign n3431 = ( n914 & ~n1959 ) | ( n914 & n3430 ) | ( ~n1959 & n3430 ) ;
  assign n3432 = ( ~n3428 & n3429 ) | ( ~n3428 & n3431 ) | ( n3429 & n3431 ) ;
  assign n3427 = n2915 ^ n1651 ^ n150 ;
  assign n3433 = n3432 ^ n3427 ^ n535 ;
  assign n3434 = ~n1589 & n3433 ;
  assign n3435 = n2668 ^ n1819 ^ n1818 ;
  assign n3436 = n3435 ^ n1917 ^ 1'b0 ;
  assign n3437 = n3434 | n3436 ;
  assign n3452 = n838 & ~n868 ;
  assign n3450 = n2034 ^ n662 ^ 1'b0 ;
  assign n3451 = n1081 & ~n3450 ;
  assign n3447 = n3238 ^ n1921 ^ n442 ;
  assign n3448 = ~n2226 & n3447 ;
  assign n3449 = ~n3311 & n3448 ;
  assign n3453 = n3452 ^ n3451 ^ n3449 ;
  assign n3446 = ( ~n1616 & n1665 ) | ( ~n1616 & n1852 ) | ( n1665 & n1852 ) ;
  assign n3438 = n1666 ^ n1534 ^ n240 ;
  assign n3439 = n3438 ^ n2888 ^ n956 ;
  assign n3440 = n1248 ^ n986 ^ 1'b0 ;
  assign n3441 = ( n2240 & ~n3401 ) | ( n2240 & n3440 ) | ( ~n3401 & n3440 ) ;
  assign n3442 = n3441 ^ n2398 ^ 1'b0 ;
  assign n3443 = ( n1563 & ~n3439 ) | ( n1563 & n3442 ) | ( ~n3439 & n3442 ) ;
  assign n3444 = ~n164 & n1153 ;
  assign n3445 = n3443 & n3444 ;
  assign n3454 = n3453 ^ n3446 ^ n3445 ;
  assign n3456 = n1692 ^ n698 ^ n669 ;
  assign n3455 = n2609 ^ n2409 ^ n1286 ;
  assign n3457 = n3456 ^ n3455 ^ n1820 ;
  assign n3458 = ~n809 & n993 ;
  assign n3459 = n3458 ^ n2280 ^ 1'b0 ;
  assign n3460 = n3427 | n3459 ;
  assign n3471 = ( n630 & n1304 ) | ( n630 & n2605 ) | ( n1304 & n2605 ) ;
  assign n3472 = n859 & n3471 ;
  assign n3473 = ~n771 & n3472 ;
  assign n3464 = x114 & ~n764 ;
  assign n3465 = n3464 ^ n635 ^ 1'b0 ;
  assign n3466 = ~n1003 & n3465 ;
  assign n3461 = n1059 ^ n604 ^ n332 ;
  assign n3462 = ( ~n1819 & n1946 ) | ( ~n1819 & n3461 ) | ( n1946 & n3461 ) ;
  assign n3463 = n3462 ^ n3026 ^ n993 ;
  assign n3467 = n3466 ^ n3463 ^ n2813 ;
  assign n3468 = n3467 ^ n3351 ^ n1822 ;
  assign n3469 = ( ~n1457 & n2488 ) | ( ~n1457 & n3468 ) | ( n2488 & n3468 ) ;
  assign n3470 = n3469 ^ n2962 ^ n696 ;
  assign n3474 = n3473 ^ n3470 ^ n768 ;
  assign n3484 = n1771 ^ n1108 ^ n718 ;
  assign n3477 = n1106 ^ n274 ^ 1'b0 ;
  assign n3478 = ~n2392 & n3477 ;
  assign n3475 = n357 & ~n3357 ;
  assign n3476 = ~n281 & n3475 ;
  assign n3479 = n3478 ^ n3476 ^ n3051 ;
  assign n3480 = ( n164 & ~n174 ) | ( n164 & n360 ) | ( ~n174 & n360 ) ;
  assign n3481 = n3480 ^ n1485 ^ n1021 ;
  assign n3482 = n3481 ^ n2776 ^ n1401 ;
  assign n3483 = ( n1116 & n3479 ) | ( n1116 & ~n3482 ) | ( n3479 & ~n3482 ) ;
  assign n3485 = n3484 ^ n3483 ^ n887 ;
  assign n3486 = n2689 ^ n583 ^ 1'b0 ;
  assign n3487 = ~n3229 & n3486 ;
  assign n3488 = ( x99 & n3471 ) | ( x99 & ~n3487 ) | ( n3471 & ~n3487 ) ;
  assign n3489 = n2475 ^ n1731 ^ n1121 ;
  assign n3490 = ( n1557 & n3421 ) | ( n1557 & n3489 ) | ( n3421 & n3489 ) ;
  assign n3493 = n2151 ^ n1080 ^ n333 ;
  assign n3491 = ( n334 & ~n363 ) | ( n334 & n3401 ) | ( ~n363 & n3401 ) ;
  assign n3492 = ~n1437 & n3491 ;
  assign n3494 = n3493 ^ n3492 ^ 1'b0 ;
  assign n3495 = ~n2157 & n2435 ;
  assign n3496 = n1544 & n3495 ;
  assign n3497 = n1998 ^ n1171 ^ x117 ;
  assign n3498 = n1425 & ~n3497 ;
  assign n3500 = n1920 & ~n2433 ;
  assign n3499 = ( n2229 & n3106 ) | ( n2229 & n3178 ) | ( n3106 & n3178 ) ;
  assign n3501 = n3500 ^ n3499 ^ n2234 ;
  assign n3502 = ( ~n3387 & n3498 ) | ( ~n3387 & n3501 ) | ( n3498 & n3501 ) ;
  assign n3503 = ( ~n1850 & n3496 ) | ( ~n1850 & n3502 ) | ( n3496 & n3502 ) ;
  assign n3504 = n2279 ^ n1446 ^ n1253 ;
  assign n3505 = n3504 ^ n664 ^ x122 ;
  assign n3506 = ( n336 & ~n673 ) | ( n336 & n3505 ) | ( ~n673 & n3505 ) ;
  assign n3507 = n3503 & ~n3506 ;
  assign n3508 = n1031 ^ n931 ^ 1'b0 ;
  assign n3509 = n1008 | n3508 ;
  assign n3510 = ( n845 & n1549 ) | ( n845 & n3509 ) | ( n1549 & n3509 ) ;
  assign n3512 = x47 & ~n2913 ;
  assign n3513 = ~n263 & n3512 ;
  assign n3511 = n289 & ~n3440 ;
  assign n3514 = n3513 ^ n3511 ^ 1'b0 ;
  assign n3515 = ( n1386 & ~n3510 ) | ( n1386 & n3514 ) | ( ~n3510 & n3514 ) ;
  assign n3517 = ( n699 & n790 ) | ( n699 & n2230 ) | ( n790 & n2230 ) ;
  assign n3516 = n1793 ^ n1358 ^ 1'b0 ;
  assign n3518 = n3517 ^ n3516 ^ n2335 ;
  assign n3527 = ( n2029 & n2466 ) | ( n2029 & n3358 ) | ( n2466 & n3358 ) ;
  assign n3521 = n2975 ^ n2352 ^ n264 ;
  assign n3522 = n3521 ^ x97 ^ x11 ;
  assign n3523 = n3522 ^ n1341 ^ n868 ;
  assign n3519 = ( x20 & n189 ) | ( x20 & n1473 ) | ( n189 & n1473 ) ;
  assign n3520 = n3519 ^ n1242 ^ 1'b0 ;
  assign n3524 = n3523 ^ n3520 ^ n2964 ;
  assign n3525 = ( ~n427 & n2425 ) | ( ~n427 & n3524 ) | ( n2425 & n3524 ) ;
  assign n3526 = n3525 ^ n2920 ^ n898 ;
  assign n3528 = n3527 ^ n3526 ^ n2141 ;
  assign n3529 = ( n1558 & n3518 ) | ( n1558 & ~n3528 ) | ( n3518 & ~n3528 ) ;
  assign n3530 = n1990 ^ n1530 ^ n383 ;
  assign n3534 = n254 & n3230 ;
  assign n3535 = n3534 ^ n2454 ^ 1'b0 ;
  assign n3536 = n3535 ^ n1520 ^ n738 ;
  assign n3537 = ( ~n2019 & n2022 ) | ( ~n2019 & n3536 ) | ( n2022 & n3536 ) ;
  assign n3531 = ( n676 & ~n1209 ) | ( n676 & n2101 ) | ( ~n1209 & n2101 ) ;
  assign n3532 = ( n2171 & n2958 ) | ( n2171 & ~n3531 ) | ( n2958 & ~n3531 ) ;
  assign n3533 = n3532 ^ n2205 ^ n1232 ;
  assign n3538 = n3537 ^ n3533 ^ n1211 ;
  assign n3539 = ( n1393 & n1799 ) | ( n1393 & ~n3538 ) | ( n1799 & ~n3538 ) ;
  assign n3540 = n3539 ^ n2680 ^ 1'b0 ;
  assign n3541 = ~n3530 & n3540 ;
  assign n3544 = ( n1977 & n2390 ) | ( n1977 & ~n2866 ) | ( n2390 & ~n2866 ) ;
  assign n3542 = n196 & n1707 ;
  assign n3543 = n3542 ^ n2342 ^ 1'b0 ;
  assign n3545 = n3544 ^ n3543 ^ n2410 ;
  assign n3550 = n3372 ^ n2995 ^ n2591 ;
  assign n3549 = n2695 ^ n1886 ^ n722 ;
  assign n3546 = n1786 ^ n1069 ^ 1'b0 ;
  assign n3547 = n1681 & n3546 ;
  assign n3548 = n3547 ^ n1125 ^ n1122 ;
  assign n3551 = n3550 ^ n3549 ^ n3548 ;
  assign n3552 = n3551 ^ n2320 ^ n2024 ;
  assign n3557 = ( ~x125 & n160 ) | ( ~x125 & n380 ) | ( n160 & n380 ) ;
  assign n3558 = n3557 ^ x63 ^ x0 ;
  assign n3556 = n2568 ^ n2151 ^ n1226 ;
  assign n3555 = ( n178 & ~n1848 ) | ( n178 & n3012 ) | ( ~n1848 & n3012 ) ;
  assign n3559 = n3558 ^ n3556 ^ n3555 ;
  assign n3554 = n455 ^ x103 ^ 1'b0 ;
  assign n3553 = ( n949 & n2347 ) | ( n949 & ~n2770 ) | ( n2347 & ~n2770 ) ;
  assign n3560 = n3559 ^ n3554 ^ n3553 ;
  assign n3562 = ( n856 & ~n1813 ) | ( n856 & n2837 ) | ( ~n1813 & n2837 ) ;
  assign n3561 = ( ~n438 & n1620 ) | ( ~n438 & n2998 ) | ( n1620 & n2998 ) ;
  assign n3563 = n3562 ^ n3561 ^ n1742 ;
  assign n3565 = ( ~n468 & n1771 ) | ( ~n468 & n2238 ) | ( n1771 & n2238 ) ;
  assign n3566 = n3565 ^ n1511 ^ n1140 ;
  assign n3564 = n1927 ^ n1912 ^ n1290 ;
  assign n3567 = n3566 ^ n3564 ^ n1917 ;
  assign n3585 = n2178 ^ n777 ^ 1'b0 ;
  assign n3586 = n594 & ~n3585 ;
  assign n3582 = n3500 ^ n1612 ^ n1282 ;
  assign n3579 = ~n2140 & n2995 ;
  assign n3580 = n3579 ^ n1350 ^ 1'b0 ;
  assign n3577 = ( x62 & ~n205 ) | ( x62 & n1407 ) | ( ~n205 & n1407 ) ;
  assign n3578 = ( ~n661 & n2446 ) | ( ~n661 & n3577 ) | ( n2446 & n3577 ) ;
  assign n3581 = n3580 ^ n3578 ^ n1440 ;
  assign n3576 = ( n639 & n2878 ) | ( n639 & ~n3022 ) | ( n2878 & ~n3022 ) ;
  assign n3583 = n3582 ^ n3581 ^ n3576 ;
  assign n3584 = n3583 ^ n2393 ^ n409 ;
  assign n3568 = n3034 ^ n1727 ^ n276 ;
  assign n3569 = n2610 ^ n1662 ^ 1'b0 ;
  assign n3570 = n628 & n3569 ;
  assign n3571 = ( ~n1311 & n1612 ) | ( ~n1311 & n2774 ) | ( n1612 & n2774 ) ;
  assign n3572 = ( n761 & ~n3570 ) | ( n761 & n3571 ) | ( ~n3570 & n3571 ) ;
  assign n3573 = ( x90 & n1991 ) | ( x90 & ~n2149 ) | ( n1991 & ~n2149 ) ;
  assign n3574 = ( n3568 & ~n3572 ) | ( n3568 & n3573 ) | ( ~n3572 & n3573 ) ;
  assign n3575 = n3574 ^ n2735 ^ n627 ;
  assign n3587 = n3586 ^ n3584 ^ n3575 ;
  assign n3588 = ( n1257 & n2662 ) | ( n1257 & n3568 ) | ( n2662 & n3568 ) ;
  assign n3589 = n1650 | n3588 ;
  assign n3590 = n3589 ^ n1823 ^ n978 ;
  assign n3591 = n3590 ^ n3369 ^ n2691 ;
  assign n3594 = n951 ^ n605 ^ 1'b0 ;
  assign n3595 = n2735 ^ n270 ^ 1'b0 ;
  assign n3596 = ~n921 & n3595 ;
  assign n3597 = ( n1898 & n2613 ) | ( n1898 & n3596 ) | ( n2613 & n3596 ) ;
  assign n3602 = n2993 ^ n1845 ^ x46 ;
  assign n3599 = ( n348 & ~n1098 ) | ( n348 & n2742 ) | ( ~n1098 & n2742 ) ;
  assign n3598 = ( x63 & x65 ) | ( x63 & ~n855 ) | ( x65 & ~n855 ) ;
  assign n3600 = n3599 ^ n3598 ^ n3578 ;
  assign n3601 = ( n933 & n2338 ) | ( n933 & n3600 ) | ( n2338 & n3600 ) ;
  assign n3603 = n3602 ^ n3601 ^ n2091 ;
  assign n3604 = ( ~n3118 & n3597 ) | ( ~n3118 & n3603 ) | ( n3597 & n3603 ) ;
  assign n3605 = ( ~n1309 & n3594 ) | ( ~n1309 & n3604 ) | ( n3594 & n3604 ) ;
  assign n3592 = ~n458 & n3178 ;
  assign n3593 = n3592 ^ n3028 ^ 1'b0 ;
  assign n3606 = n3605 ^ n3593 ^ n147 ;
  assign n3608 = x20 & n1081 ;
  assign n3609 = n3250 & n3608 ;
  assign n3607 = ~n1731 & n3077 ;
  assign n3610 = n3609 ^ n3607 ^ 1'b0 ;
  assign n3611 = ( ~n524 & n994 ) | ( ~n524 & n1929 ) | ( n994 & n1929 ) ;
  assign n3612 = n1876 & ~n3611 ;
  assign n3613 = n2287 ^ n1173 ^ 1'b0 ;
  assign n3614 = n3613 ^ n2100 ^ n1517 ;
  assign n3621 = ( n530 & ~n817 ) | ( n530 & n1762 ) | ( ~n817 & n1762 ) ;
  assign n3615 = n3028 ^ n367 ^ 1'b0 ;
  assign n3616 = ( n1535 & n2155 ) | ( n1535 & n3615 ) | ( n2155 & n3615 ) ;
  assign n3617 = n1557 ^ n903 ^ n737 ;
  assign n3618 = ( n684 & n1975 ) | ( n684 & n2876 ) | ( n1975 & n2876 ) ;
  assign n3619 = ( n332 & n2337 ) | ( n332 & ~n3618 ) | ( n2337 & ~n3618 ) ;
  assign n3620 = ( ~n3616 & n3617 ) | ( ~n3616 & n3619 ) | ( n3617 & n3619 ) ;
  assign n3622 = n3621 ^ n3620 ^ n676 ;
  assign n3623 = n3622 ^ n3531 ^ n2144 ;
  assign n3624 = ( n674 & n1486 ) | ( n674 & n1862 ) | ( n1486 & n1862 ) ;
  assign n3625 = n3624 ^ n2839 ^ n1021 ;
  assign n3626 = ( n3614 & n3623 ) | ( n3614 & ~n3625 ) | ( n3623 & ~n3625 ) ;
  assign n3631 = ( n850 & ~n2541 ) | ( n850 & n3288 ) | ( ~n2541 & n3288 ) ;
  assign n3629 = ( n253 & n289 ) | ( n253 & n1581 ) | ( n289 & n1581 ) ;
  assign n3627 = n1316 ^ n867 ^ 1'b0 ;
  assign n3628 = n3627 ^ n2716 ^ n1889 ;
  assign n3630 = n3629 ^ n3628 ^ n1610 ;
  assign n3632 = n3631 ^ n3630 ^ 1'b0 ;
  assign n3633 = n1395 & n2257 ;
  assign n3634 = ( n1352 & n2664 ) | ( n1352 & n3633 ) | ( n2664 & n3633 ) ;
  assign n3635 = ( n628 & ~n822 ) | ( n628 & n2297 ) | ( ~n822 & n2297 ) ;
  assign n3636 = n3311 ^ n1846 ^ n1644 ;
  assign n3637 = ( ~n1926 & n2890 ) | ( ~n1926 & n3636 ) | ( n2890 & n3636 ) ;
  assign n3638 = n1099 ^ n864 ^ n301 ;
  assign n3639 = n3638 ^ n1543 ^ n967 ;
  assign n3640 = n3639 ^ n1780 ^ n426 ;
  assign n3641 = ( n3635 & n3637 ) | ( n3635 & n3640 ) | ( n3637 & n3640 ) ;
  assign n3642 = n3641 ^ n2011 ^ x81 ;
  assign n3643 = n3642 ^ n801 ^ 1'b0 ;
  assign n3664 = n1081 ^ n765 ^ 1'b0 ;
  assign n3665 = ~n221 & n3664 ;
  assign n3661 = n1044 ^ n451 ^ n365 ;
  assign n3662 = n2513 & n3661 ;
  assign n3663 = ( ~n150 & n923 ) | ( ~n150 & n3662 ) | ( n923 & n3662 ) ;
  assign n3656 = ( ~x75 & n651 ) | ( ~x75 & n1081 ) | ( n651 & n1081 ) ;
  assign n3654 = n2680 ^ n2320 ^ n1476 ;
  assign n3651 = ( n850 & ~n1559 ) | ( n850 & n2139 ) | ( ~n1559 & n2139 ) ;
  assign n3649 = x104 & n494 ;
  assign n3650 = n3649 ^ n3220 ^ 1'b0 ;
  assign n3652 = n3651 ^ n3650 ^ n986 ;
  assign n3653 = n3652 ^ n3568 ^ n3138 ;
  assign n3648 = ( ~n649 & n1582 ) | ( ~n649 & n2615 ) | ( n1582 & n2615 ) ;
  assign n3655 = n3654 ^ n3653 ^ n3648 ;
  assign n3644 = ( ~n287 & n834 ) | ( ~n287 & n2901 ) | ( n834 & n2901 ) ;
  assign n3645 = ( x36 & x90 ) | ( x36 & ~n1538 ) | ( x90 & ~n1538 ) ;
  assign n3646 = n2915 & n3645 ;
  assign n3647 = ( n1077 & n3644 ) | ( n1077 & n3646 ) | ( n3644 & n3646 ) ;
  assign n3657 = n3656 ^ n3655 ^ n3647 ;
  assign n3658 = ( n530 & ~n2612 ) | ( n530 & n3657 ) | ( ~n2612 & n3657 ) ;
  assign n3659 = n3658 ^ n3533 ^ 1'b0 ;
  assign n3660 = ~n852 & n3659 ;
  assign n3666 = n3665 ^ n3663 ^ n3660 ;
  assign n3669 = n326 & ~n913 ;
  assign n3667 = n2607 ^ n334 ^ x31 ;
  assign n3668 = n3667 ^ n2645 ^ n703 ;
  assign n3670 = n3669 ^ n3668 ^ n2301 ;
  assign n3671 = n3670 ^ n2452 ^ n1970 ;
  assign n3672 = n939 ^ n646 ^ n310 ;
  assign n3673 = ( n289 & n678 ) | ( n289 & n3672 ) | ( n678 & n3672 ) ;
  assign n3674 = n3673 ^ n2975 ^ n678 ;
  assign n3675 = n3674 ^ n2306 ^ n1454 ;
  assign n3676 = n3207 ^ n2838 ^ n286 ;
  assign n3677 = ( ~n358 & n2579 ) | ( ~n358 & n3676 ) | ( n2579 & n3676 ) ;
  assign n3678 = n3677 ^ n2513 ^ n1960 ;
  assign n3685 = n3366 ^ n1538 ^ n719 ;
  assign n3679 = n2558 ^ n1889 ^ n1874 ;
  assign n3680 = ( n2141 & n3280 ) | ( n2141 & n3679 ) | ( n3280 & n3679 ) ;
  assign n3681 = ( n847 & n1201 ) | ( n847 & n2015 ) | ( n1201 & n2015 ) ;
  assign n3682 = ( n1644 & n1881 ) | ( n1644 & n3681 ) | ( n1881 & n3681 ) ;
  assign n3683 = ( n1397 & n2083 ) | ( n1397 & n3682 ) | ( n2083 & n3682 ) ;
  assign n3684 = ( n3238 & n3680 ) | ( n3238 & n3683 ) | ( n3680 & n3683 ) ;
  assign n3686 = n3685 ^ n3684 ^ n1039 ;
  assign n3687 = n3529 ^ n3430 ^ n679 ;
  assign n3688 = ( n890 & n1178 ) | ( n890 & ~n2806 ) | ( n1178 & ~n2806 ) ;
  assign n3689 = n3688 ^ n3390 ^ n188 ;
  assign n3690 = n3689 ^ n1197 ^ 1'b0 ;
  assign n3691 = ( ~n184 & n582 ) | ( ~n184 & n847 ) | ( n582 & n847 ) ;
  assign n3692 = n3691 ^ n2808 ^ 1'b0 ;
  assign n3693 = n3692 ^ x68 ^ 1'b0 ;
  assign n3694 = ( x5 & n1513 ) | ( x5 & n3693 ) | ( n1513 & n3693 ) ;
  assign n3695 = n2727 ^ n2055 ^ x5 ;
  assign n3696 = ~n2097 & n3695 ;
  assign n3697 = n697 ^ n690 ^ n133 ;
  assign n3698 = ( n2264 & n3547 ) | ( n2264 & n3697 ) | ( n3547 & n3697 ) ;
  assign n3699 = n2884 & n3698 ;
  assign n3700 = n305 | n1566 ;
  assign n3701 = n1841 & ~n3700 ;
  assign n3702 = n3701 ^ n241 ^ n202 ;
  assign n3703 = n3702 ^ n436 ^ x97 ;
  assign n3704 = ( n1036 & ~n1762 ) | ( n1036 & n3703 ) | ( ~n1762 & n3703 ) ;
  assign n3705 = ( ~n1158 & n1961 ) | ( ~n1158 & n3704 ) | ( n1961 & n3704 ) ;
  assign n3710 = n2572 ^ n726 ^ n234 ;
  assign n3707 = n961 ^ n697 ^ n284 ;
  assign n3708 = ( ~n1991 & n3327 ) | ( ~n1991 & n3707 ) | ( n3327 & n3707 ) ;
  assign n3709 = n3708 ^ n1716 ^ n1522 ;
  assign n3706 = n1479 ^ n678 ^ n554 ;
  assign n3711 = n3710 ^ n3709 ^ n3706 ;
  assign n3712 = n2294 | n3711 ;
  assign n3719 = ( ~n1845 & n2353 ) | ( ~n1845 & n3661 ) | ( n2353 & n3661 ) ;
  assign n3720 = n2093 ^ n1467 ^ n191 ;
  assign n3721 = n3720 ^ n2604 ^ x6 ;
  assign n3722 = ( n1049 & ~n3103 ) | ( n1049 & n3721 ) | ( ~n3103 & n3721 ) ;
  assign n3723 = ( n497 & n2338 ) | ( n497 & ~n3722 ) | ( n2338 & ~n3722 ) ;
  assign n3724 = n1706 ^ n890 ^ n769 ;
  assign n3725 = ~n1698 & n3724 ;
  assign n3726 = n3725 ^ n947 ^ n844 ;
  assign n3727 = ( ~n3719 & n3723 ) | ( ~n3719 & n3726 ) | ( n3723 & n3726 ) ;
  assign n3715 = n1797 ^ n1650 ^ n694 ;
  assign n3716 = n3715 ^ n1787 ^ n454 ;
  assign n3714 = n3229 ^ n1625 ^ n1069 ;
  assign n3717 = n3716 ^ n3714 ^ 1'b0 ;
  assign n3713 = ( ~n666 & n1205 ) | ( ~n666 & n2320 ) | ( n1205 & n2320 ) ;
  assign n3718 = n3717 ^ n3713 ^ 1'b0 ;
  assign n3728 = n3727 ^ n3718 ^ n3121 ;
  assign n3730 = n717 ^ n261 ^ 1'b0 ;
  assign n3731 = n1947 | n3730 ;
  assign n3732 = n467 & n512 ;
  assign n3733 = n3731 & n3732 ;
  assign n3734 = ( ~x115 & n1237 ) | ( ~x115 & n3733 ) | ( n1237 & n3733 ) ;
  assign n3729 = n1922 ^ n1779 ^ n1046 ;
  assign n3735 = n3734 ^ n3729 ^ n965 ;
  assign n3736 = n1559 ^ n734 ^ 1'b0 ;
  assign n3737 = n3736 ^ n2712 ^ n1017 ;
  assign n3738 = ( ~n213 & n2057 ) | ( ~n213 & n3639 ) | ( n2057 & n3639 ) ;
  assign n3739 = n3738 ^ n3614 ^ n1934 ;
  assign n3740 = n2479 ^ n2456 ^ n1718 ;
  assign n3741 = n3740 ^ n2698 ^ n2186 ;
  assign n3742 = ( ~n268 & n656 ) | ( ~n268 & n1813 ) | ( n656 & n1813 ) ;
  assign n3743 = n3742 ^ n2775 ^ n2264 ;
  assign n3744 = ( ~n1258 & n3051 ) | ( ~n1258 & n3743 ) | ( n3051 & n3743 ) ;
  assign n3745 = ( n990 & n3741 ) | ( n990 & n3744 ) | ( n3741 & n3744 ) ;
  assign n3746 = ( ~n1183 & n1201 ) | ( ~n1183 & n2022 ) | ( n1201 & n2022 ) ;
  assign n3748 = ( n383 & n460 ) | ( n383 & ~n3360 ) | ( n460 & ~n3360 ) ;
  assign n3749 = n3748 ^ n929 ^ n744 ;
  assign n3750 = n3749 ^ n1226 ^ n379 ;
  assign n3751 = ( ~x84 & n1479 ) | ( ~x84 & n3750 ) | ( n1479 & n3750 ) ;
  assign n3747 = n3111 ^ n1945 ^ n313 ;
  assign n3752 = n3751 ^ n3747 ^ n3276 ;
  assign n3753 = n3752 ^ n524 ^ 1'b0 ;
  assign n3754 = ( n2442 & n3746 ) | ( n2442 & ~n3753 ) | ( n3746 & ~n3753 ) ;
  assign n3755 = ( ~n216 & n534 ) | ( ~n216 & n3093 ) | ( n534 & n3093 ) ;
  assign n3756 = n3755 ^ n2665 ^ 1'b0 ;
  assign n3762 = ( n498 & n896 ) | ( n498 & n1491 ) | ( n896 & n1491 ) ;
  assign n3761 = ( n1386 & n2492 ) | ( n1386 & ~n3688 ) | ( n2492 & ~n3688 ) ;
  assign n3763 = n3762 ^ n3761 ^ n328 ;
  assign n3757 = n3570 ^ n1147 ^ n700 ;
  assign n3758 = ( n1558 & n1993 ) | ( n1558 & n3331 ) | ( n1993 & n3331 ) ;
  assign n3759 = ( n738 & n848 ) | ( n738 & ~n3758 ) | ( n848 & ~n3758 ) ;
  assign n3760 = ( n2881 & n3757 ) | ( n2881 & n3759 ) | ( n3757 & n3759 ) ;
  assign n3764 = n3763 ^ n3760 ^ 1'b0 ;
  assign n3765 = n2478 & n3764 ;
  assign n3766 = n3765 ^ x59 ^ 1'b0 ;
  assign n3767 = n3756 & ~n3766 ;
  assign n3768 = ( n814 & ~n1444 ) | ( n814 & n1997 ) | ( ~n1444 & n1997 ) ;
  assign n3769 = n174 | n404 ;
  assign n3770 = n3769 ^ n1280 ^ 1'b0 ;
  assign n3771 = n240 & ~n3770 ;
  assign n3772 = n1768 ^ n1630 ^ n1212 ;
  assign n3773 = ( ~n1364 & n1528 ) | ( ~n1364 & n2322 ) | ( n1528 & n2322 ) ;
  assign n3774 = ( ~n3771 & n3772 ) | ( ~n3771 & n3773 ) | ( n3772 & n3773 ) ;
  assign n3775 = ~n3768 & n3774 ;
  assign n3776 = n2768 ^ n1309 ^ n549 ;
  assign n3777 = n3776 ^ n3535 ^ n323 ;
  assign n3778 = n3777 ^ n3316 ^ x102 ;
  assign n3779 = n2080 ^ n1411 ^ n748 ;
  assign n3780 = ( n459 & n2260 ) | ( n459 & n3779 ) | ( n2260 & n3779 ) ;
  assign n3782 = ( ~n343 & n455 ) | ( ~n343 & n1664 ) | ( n455 & n1664 ) ;
  assign n3783 = n3782 ^ n1818 ^ n619 ;
  assign n3784 = n3783 ^ n2067 ^ n447 ;
  assign n3781 = n3760 ^ n1867 ^ n1238 ;
  assign n3785 = n3784 ^ n3781 ^ 1'b0 ;
  assign n3786 = n2123 | n3785 ;
  assign n3792 = n1754 ^ n1589 ^ n160 ;
  assign n3788 = n2780 ^ n1124 ^ n983 ;
  assign n3789 = n3788 ^ n3521 ^ n525 ;
  assign n3790 = ~n1172 & n1889 ;
  assign n3791 = ~n3789 & n3790 ;
  assign n3787 = n3580 ^ n2316 ^ n2007 ;
  assign n3793 = n3792 ^ n3791 ^ n3787 ;
  assign n3796 = n1110 | n1547 ;
  assign n3794 = ( x71 & n731 ) | ( x71 & ~n1511 ) | ( n731 & ~n1511 ) ;
  assign n3795 = n3794 ^ n1774 ^ n1113 ;
  assign n3797 = n3796 ^ n3795 ^ n1692 ;
  assign n3798 = n3797 ^ n2942 ^ n1716 ;
  assign n3799 = n2814 ^ n1122 ^ 1'b0 ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3801 = ( n2929 & ~n3793 ) | ( n2929 & n3800 ) | ( ~n3793 & n3800 ) ;
  assign n3802 = ( ~x3 & n1543 ) | ( ~x3 & n2976 ) | ( n1543 & n2976 ) ;
  assign n3810 = n910 | n2133 ;
  assign n3808 = ( n647 & n736 ) | ( n647 & ~n934 ) | ( n736 & ~n934 ) ;
  assign n3805 = n347 & ~n1574 ;
  assign n3806 = ~n603 & n3805 ;
  assign n3807 = n3806 ^ n3688 ^ 1'b0 ;
  assign n3803 = n957 ^ n657 ^ n604 ;
  assign n3804 = n3803 ^ n3638 ^ n2708 ;
  assign n3809 = n3808 ^ n3807 ^ n3804 ;
  assign n3811 = n3810 ^ n3809 ^ n1351 ;
  assign n3812 = n3802 & ~n3811 ;
  assign n3813 = ~n2744 & n3812 ;
  assign n3817 = ( n679 & n884 ) | ( n679 & n2524 ) | ( n884 & n2524 ) ;
  assign n3814 = n3187 ^ n2730 ^ n2395 ;
  assign n3815 = ( n391 & n1449 ) | ( n391 & n3814 ) | ( n1449 & n3814 ) ;
  assign n3816 = n3736 | n3815 ;
  assign n3818 = n3817 ^ n3816 ^ n2998 ;
  assign n3821 = ( ~n588 & n2091 ) | ( ~n588 & n2180 ) | ( n2091 & n2180 ) ;
  assign n3822 = ( x67 & n181 ) | ( x67 & n3821 ) | ( n181 & n3821 ) ;
  assign n3819 = n1671 ^ n910 ^ n369 ;
  assign n3820 = n3819 ^ n3602 ^ x113 ;
  assign n3823 = n3822 ^ n3820 ^ n2359 ;
  assign n3824 = n3514 ^ n1690 ^ 1'b0 ;
  assign n3825 = n3824 ^ n2837 ^ 1'b0 ;
  assign n3834 = n2619 ^ n1714 ^ n1454 ;
  assign n3835 = ( n1601 & n2733 ) | ( n1601 & ~n3834 ) | ( n2733 & ~n3834 ) ;
  assign n3836 = n3835 ^ n2712 ^ n1719 ;
  assign n3826 = ( n1306 & ~n1670 ) | ( n1306 & n2582 ) | ( ~n1670 & n2582 ) ;
  assign n3827 = ( n588 & n1246 ) | ( n588 & ~n3826 ) | ( n1246 & ~n3826 ) ;
  assign n3828 = n3827 ^ n2392 ^ n1175 ;
  assign n3829 = n3689 | n3828 ;
  assign n3830 = n1657 ^ n1064 ^ x43 ;
  assign n3831 = n3830 ^ n2167 ^ n775 ;
  assign n3832 = x29 & ~n225 ;
  assign n3833 = ( ~n3829 & n3831 ) | ( ~n3829 & n3832 ) | ( n3831 & n3832 ) ;
  assign n3837 = n3836 ^ n3833 ^ n707 ;
  assign n3845 = n2120 ^ n1867 ^ x120 ;
  assign n3846 = ( n1167 & ~n3119 ) | ( n1167 & n3845 ) | ( ~n3119 & n3845 ) ;
  assign n3847 = ~n1335 & n1526 ;
  assign n3848 = n3846 & ~n3847 ;
  assign n3849 = n2658 & n3848 ;
  assign n3842 = n276 ^ x114 ^ 1'b0 ;
  assign n3843 = n699 | n3842 ;
  assign n3841 = ( n847 & n918 ) | ( n847 & n2303 ) | ( n918 & n2303 ) ;
  assign n3839 = ( n780 & n1164 ) | ( n780 & n1905 ) | ( n1164 & n1905 ) ;
  assign n3840 = ( ~n439 & n3792 ) | ( ~n439 & n3839 ) | ( n3792 & n3839 ) ;
  assign n3844 = n3843 ^ n3841 ^ n3840 ;
  assign n3838 = ( n221 & n429 ) | ( n221 & ~n2256 ) | ( n429 & ~n2256 ) ;
  assign n3850 = n3849 ^ n3844 ^ n3838 ;
  assign n3851 = n3850 ^ n2730 ^ 1'b0 ;
  assign n3852 = n417 ^ n396 ^ 1'b0 ;
  assign n3853 = n246 & ~n3852 ;
  assign n3854 = ( n1845 & n2012 ) | ( n1845 & n3853 ) | ( n2012 & n3853 ) ;
  assign n3855 = n1777 ^ n1686 ^ n1523 ;
  assign n3856 = n479 & n1263 ;
  assign n3857 = ~x51 & n3856 ;
  assign n3858 = n2288 ^ n541 ^ 1'b0 ;
  assign n3859 = n3857 | n3858 ;
  assign n3860 = n2139 ^ n486 ^ x68 ;
  assign n3861 = n3860 ^ n1491 ^ n1139 ;
  assign n3862 = ~n3859 & n3861 ;
  assign n3863 = n1527 & n2308 ;
  assign n3864 = ~n2134 & n3863 ;
  assign n3865 = n2217 ^ n1825 ^ n1465 ;
  assign n3866 = ( n648 & n3864 ) | ( n648 & ~n3865 ) | ( n3864 & ~n3865 ) ;
  assign n3867 = ( ~n1306 & n1384 ) | ( ~n1306 & n2963 ) | ( n1384 & n2963 ) ;
  assign n3868 = n1787 ^ n383 ^ x66 ;
  assign n3869 = ( ~n1141 & n3758 ) | ( ~n1141 & n3868 ) | ( n3758 & n3868 ) ;
  assign n3870 = ( n1820 & n3867 ) | ( n1820 & n3869 ) | ( n3867 & n3869 ) ;
  assign n3871 = ( ~n344 & n1664 ) | ( ~n344 & n3870 ) | ( n1664 & n3870 ) ;
  assign n3872 = ( n396 & n3866 ) | ( n396 & ~n3871 ) | ( n3866 & ~n3871 ) ;
  assign n3873 = n3872 ^ n2983 ^ x8 ;
  assign n3874 = n2580 ^ n2262 ^ n1174 ;
  assign n3875 = n2141 ^ n686 ^ n473 ;
  assign n3876 = n1556 | n3278 ;
  assign n3877 = ~n3875 & n3876 ;
  assign n3878 = n904 ^ n698 ^ n130 ;
  assign n3879 = ( n3874 & n3877 ) | ( n3874 & n3878 ) | ( n3877 & n3878 ) ;
  assign n3882 = n2507 ^ n2322 ^ n1495 ;
  assign n3880 = ~n756 & n1729 ;
  assign n3881 = n3880 ^ n1929 ^ 1'b0 ;
  assign n3883 = n3882 ^ n3881 ^ n3182 ;
  assign n3884 = n3030 ^ n321 ^ 1'b0 ;
  assign n3885 = n3884 ^ n1224 ^ n1131 ;
  assign n3886 = ( n2424 & ~n3173 ) | ( n2424 & n3885 ) | ( ~n3173 & n3885 ) ;
  assign n3887 = n2308 ^ n1021 ^ n676 ;
  assign n3888 = n3887 ^ n3748 ^ n2397 ;
  assign n3889 = n3888 ^ n3191 ^ n274 ;
  assign n3890 = ( ~n579 & n932 ) | ( ~n579 & n3051 ) | ( n932 & n3051 ) ;
  assign n3891 = ~n1013 & n1603 ;
  assign n3892 = n3891 ^ n2429 ^ x13 ;
  assign n3893 = n3892 ^ n1386 ^ n507 ;
  assign n3894 = ( n2989 & n3770 ) | ( n2989 & ~n3893 ) | ( n3770 & ~n3893 ) ;
  assign n3895 = n2383 ^ n2121 ^ n834 ;
  assign n3896 = x50 & n240 ;
  assign n3897 = ~n1654 & n3896 ;
  assign n3898 = ( ~n508 & n812 ) | ( ~n508 & n3897 ) | ( n812 & n3897 ) ;
  assign n3899 = ( ~n974 & n3895 ) | ( ~n974 & n3898 ) | ( n3895 & n3898 ) ;
  assign n3900 = ~n1941 & n3899 ;
  assign n3901 = n3900 ^ n873 ^ 1'b0 ;
  assign n3902 = ( n3890 & n3894 ) | ( n3890 & ~n3901 ) | ( n3894 & ~n3901 ) ;
  assign n3931 = n3120 ^ n2564 ^ x99 ;
  assign n3930 = n2279 ^ n1739 ^ n1342 ;
  assign n3922 = ( n175 & n1801 ) | ( n175 & n2609 ) | ( n1801 & n2609 ) ;
  assign n3923 = n3922 ^ n482 ^ 1'b0 ;
  assign n3925 = ( ~n449 & n647 ) | ( ~n449 & n1577 ) | ( n647 & n1577 ) ;
  assign n3924 = n3520 ^ n3318 ^ n2399 ;
  assign n3926 = n3925 ^ n3924 ^ n238 ;
  assign n3927 = n3923 & n3926 ;
  assign n3928 = n3927 ^ n2248 ^ 1'b0 ;
  assign n3903 = n1116 ^ x93 ^ 1'b0 ;
  assign n3904 = n258 & ~n3903 ;
  assign n3913 = ~n2133 & n2452 ;
  assign n3914 = n1309 & n3913 ;
  assign n3915 = n132 | n3762 ;
  assign n3916 = n3914 & ~n3915 ;
  assign n3917 = n3916 ^ n3056 ^ n1297 ;
  assign n3918 = ~n502 & n3917 ;
  assign n3919 = n3918 ^ n3810 ^ 1'b0 ;
  assign n3905 = ( ~n990 & n1848 ) | ( ~n990 & n2709 ) | ( n1848 & n2709 ) ;
  assign n3906 = n183 | n620 ;
  assign n3907 = n3906 ^ n996 ^ 1'b0 ;
  assign n3908 = ( n752 & ~n2194 ) | ( n752 & n3907 ) | ( ~n2194 & n3907 ) ;
  assign n3909 = ~n348 & n3908 ;
  assign n3910 = n2955 & ~n3909 ;
  assign n3911 = ~n3905 & n3910 ;
  assign n3912 = ( n3071 & n3250 ) | ( n3071 & n3911 ) | ( n3250 & n3911 ) ;
  assign n3920 = n3919 ^ n3912 ^ n2981 ;
  assign n3921 = n3904 & ~n3920 ;
  assign n3929 = n3928 ^ n3921 ^ 1'b0 ;
  assign n3932 = n3931 ^ n3930 ^ n3929 ;
  assign n3933 = n1540 ^ n950 ^ n578 ;
  assign n3934 = n1643 ^ n1479 ^ x42 ;
  assign n3935 = ( n1619 & n3933 ) | ( n1619 & n3934 ) | ( n3933 & n3934 ) ;
  assign n3936 = ~n2106 & n3935 ;
  assign n3937 = n3936 ^ n1543 ^ 1'b0 ;
  assign n3942 = n3465 ^ n2479 ^ n967 ;
  assign n3943 = n3942 ^ n1849 ^ n507 ;
  assign n3944 = n2183 ^ n1993 ^ n1264 ;
  assign n3945 = ( n875 & ~n1098 ) | ( n875 & n3944 ) | ( ~n1098 & n3944 ) ;
  assign n3946 = ( n240 & ~n3943 ) | ( n240 & n3945 ) | ( ~n3943 & n3945 ) ;
  assign n3938 = n1818 ^ n555 ^ 1'b0 ;
  assign n3939 = n3938 ^ n2804 ^ n1161 ;
  assign n3940 = ( n2174 & n2975 ) | ( n2174 & ~n3939 ) | ( n2975 & ~n3939 ) ;
  assign n3941 = n3940 ^ n757 ^ 1'b0 ;
  assign n3947 = n3946 ^ n3941 ^ n2625 ;
  assign n3953 = n1968 ^ n1163 ^ n1146 ;
  assign n3954 = ( n1508 & n2238 ) | ( n1508 & n3953 ) | ( n2238 & n3953 ) ;
  assign n3955 = n3954 ^ n1442 ^ 1'b0 ;
  assign n3956 = n1295 & ~n3955 ;
  assign n3951 = n857 ^ n562 ^ n332 ;
  assign n3952 = n2193 | n3951 ;
  assign n3948 = n1949 ^ n737 ^ 1'b0 ;
  assign n3949 = ( n2358 & n2745 ) | ( n2358 & ~n3948 ) | ( n2745 & ~n3948 ) ;
  assign n3950 = n3949 ^ n2203 ^ x21 ;
  assign n3957 = n3956 ^ n3952 ^ n3950 ;
  assign n3958 = n3957 ^ n456 ^ 1'b0 ;
  assign n3959 = ( n1062 & n2487 ) | ( n1062 & ~n3131 ) | ( n2487 & ~n3131 ) ;
  assign n3960 = n271 | n1480 ;
  assign n3961 = n3960 ^ n393 ^ 1'b0 ;
  assign n3962 = ( x107 & n3618 ) | ( x107 & ~n3961 ) | ( n3618 & ~n3961 ) ;
  assign n3963 = ( n1364 & n3959 ) | ( n1364 & n3962 ) | ( n3959 & n3962 ) ;
  assign n3971 = ( ~n426 & n745 ) | ( ~n426 & n1176 ) | ( n745 & n1176 ) ;
  assign n3964 = n1830 ^ n1252 ^ n857 ;
  assign n3965 = ( x51 & ~n1147 ) | ( x51 & n3022 ) | ( ~n1147 & n3022 ) ;
  assign n3966 = n2847 ^ n821 ^ n469 ;
  assign n3967 = n3965 & ~n3966 ;
  assign n3968 = n2220 & n3967 ;
  assign n3969 = ( n845 & ~n3964 ) | ( n845 & n3968 ) | ( ~n3964 & n3968 ) ;
  assign n3970 = n3969 ^ n1424 ^ n528 ;
  assign n3972 = n3971 ^ n3970 ^ n754 ;
  assign n3973 = ( n361 & n1322 ) | ( n361 & ~n1405 ) | ( n1322 & ~n1405 ) ;
  assign n3974 = ~n774 & n1140 ;
  assign n3975 = n3974 ^ n2180 ^ 1'b0 ;
  assign n3976 = ( n984 & n1823 ) | ( n984 & ~n3975 ) | ( n1823 & ~n3975 ) ;
  assign n3977 = ( n414 & n747 ) | ( n414 & n3976 ) | ( n747 & n3976 ) ;
  assign n3978 = n3977 ^ n954 ^ 1'b0 ;
  assign n3979 = n2010 ^ n745 ^ n554 ;
  assign n3980 = ( n3548 & n3978 ) | ( n3548 & ~n3979 ) | ( n3978 & ~n3979 ) ;
  assign n3987 = n1727 ^ n882 ^ 1'b0 ;
  assign n3982 = ( n1446 & ~n1480 ) | ( n1446 & n1605 ) | ( ~n1480 & n1605 ) ;
  assign n3983 = n3982 ^ n3748 ^ n290 ;
  assign n3984 = ( ~n349 & n1674 ) | ( ~n349 & n3983 ) | ( n1674 & n3983 ) ;
  assign n3981 = x115 & ~n1995 ;
  assign n3985 = n3984 ^ n3981 ^ 1'b0 ;
  assign n3986 = n3985 ^ n915 ^ n716 ;
  assign n3988 = n3987 ^ n3986 ^ n2773 ;
  assign n3989 = n1706 ^ n1593 ^ 1'b0 ;
  assign n3990 = ( x105 & ~n597 ) | ( x105 & n3989 ) | ( ~n597 & n3989 ) ;
  assign n3991 = n3360 & ~n3990 ;
  assign n3992 = n496 & n3991 ;
  assign n3993 = n3992 ^ n2959 ^ n801 ;
  assign n3994 = n1246 ^ n1083 ^ 1'b0 ;
  assign n3995 = n3938 ^ n1710 ^ n200 ;
  assign n3996 = ( n985 & n2298 ) | ( n985 & ~n3995 ) | ( n2298 & ~n3995 ) ;
  assign n3997 = ( ~n556 & n1264 ) | ( ~n556 & n3996 ) | ( n1264 & n3996 ) ;
  assign n3998 = ( n907 & n3441 ) | ( n907 & n3997 ) | ( n3441 & n3997 ) ;
  assign n4000 = n131 & n646 ;
  assign n4001 = n4000 ^ n799 ^ 1'b0 ;
  assign n4002 = ( n714 & n1707 ) | ( n714 & n4001 ) | ( n1707 & n4001 ) ;
  assign n4003 = n4002 ^ n1135 ^ n524 ;
  assign n3999 = ( n1126 & n2475 ) | ( n1126 & ~n3673 ) | ( n2475 & ~n3673 ) ;
  assign n4004 = n4003 ^ n3999 ^ n3521 ;
  assign n4005 = ( ~n1440 & n3187 ) | ( ~n1440 & n4004 ) | ( n3187 & n4004 ) ;
  assign n4006 = ( n3994 & n3998 ) | ( n3994 & n4005 ) | ( n3998 & n4005 ) ;
  assign n4007 = ( n1138 & ~n3993 ) | ( n1138 & n4006 ) | ( ~n3993 & n4006 ) ;
  assign n4011 = ( n300 & n2094 ) | ( n300 & ~n2298 ) | ( n2094 & ~n2298 ) ;
  assign n4009 = ( n267 & ~n1065 ) | ( n267 & n2326 ) | ( ~n1065 & n2326 ) ;
  assign n4010 = n4009 ^ n1445 ^ n841 ;
  assign n4008 = n1953 ^ n1618 ^ n809 ;
  assign n4012 = n4011 ^ n4010 ^ n4008 ;
  assign n4013 = ( ~n945 & n1351 ) | ( ~n945 & n2500 ) | ( n1351 & n2500 ) ;
  assign n4014 = ( n674 & ~n1012 ) | ( n674 & n3362 ) | ( ~n1012 & n3362 ) ;
  assign n4015 = n4014 ^ n832 ^ x12 ;
  assign n4016 = ( n641 & n2563 ) | ( n641 & n2730 ) | ( n2563 & n2730 ) ;
  assign n4017 = ( n514 & ~n2035 ) | ( n514 & n4016 ) | ( ~n2035 & n4016 ) ;
  assign n4018 = ( n1035 & n4015 ) | ( n1035 & ~n4017 ) | ( n4015 & ~n4017 ) ;
  assign n4019 = ( ~n3830 & n4013 ) | ( ~n3830 & n4018 ) | ( n4013 & n4018 ) ;
  assign n4022 = ( n383 & ~n2347 ) | ( n383 & n2473 ) | ( ~n2347 & n2473 ) ;
  assign n4021 = ( ~n623 & n1437 ) | ( ~n623 & n1876 ) | ( n1437 & n1876 ) ;
  assign n4020 = n1529 ^ n1074 ^ 1'b0 ;
  assign n4023 = n4022 ^ n4021 ^ n4020 ;
  assign n4024 = ( n332 & n3750 ) | ( n332 & n4023 ) | ( n3750 & n4023 ) ;
  assign n4025 = ( n597 & ~n1346 ) | ( n597 & n1723 ) | ( ~n1346 & n1723 ) ;
  assign n4026 = n424 & n4025 ;
  assign n4027 = ~n4024 & n4026 ;
  assign n4028 = n3484 ^ n2039 ^ n651 ;
  assign n4029 = n3674 ^ n2831 ^ n1119 ;
  assign n4030 = ( ~n819 & n1456 ) | ( ~n819 & n3596 ) | ( n1456 & n3596 ) ;
  assign n4031 = ~n3520 & n4030 ;
  assign n4032 = ~n2363 & n4031 ;
  assign n4033 = n4032 ^ n1850 ^ 1'b0 ;
  assign n4034 = ~n4029 & n4033 ;
  assign n4035 = ( n1436 & n4028 ) | ( n1436 & ~n4034 ) | ( n4028 & ~n4034 ) ;
  assign n4036 = ( n510 & ~n723 ) | ( n510 & n758 ) | ( ~n723 & n758 ) ;
  assign n4039 = n4036 ^ n3386 ^ n1443 ;
  assign n4038 = n2882 ^ n1491 ^ n332 ;
  assign n4037 = ( ~n1437 & n2864 ) | ( ~n1437 & n4036 ) | ( n2864 & n4036 ) ;
  assign n4040 = n4039 ^ n4038 ^ n4037 ;
  assign n4044 = n1395 ^ n825 ^ n737 ;
  assign n4045 = n718 & n4044 ;
  assign n4041 = ( ~n2046 & n3832 ) | ( ~n2046 & n3839 ) | ( n3832 & n3839 ) ;
  assign n4042 = n3282 ^ n2600 ^ 1'b0 ;
  assign n4043 = ( n2610 & ~n4041 ) | ( n2610 & n4042 ) | ( ~n4041 & n4042 ) ;
  assign n4046 = n4045 ^ n4043 ^ n1487 ;
  assign n4066 = n991 & n3178 ;
  assign n4051 = n2178 ^ n465 ^ n200 ;
  assign n4052 = n1105 ^ n1100 ^ n555 ;
  assign n4053 = ( n1106 & n4051 ) | ( n1106 & ~n4052 ) | ( n4051 & ~n4052 ) ;
  assign n4047 = ( ~n606 & n2286 ) | ( ~n606 & n4022 ) | ( n2286 & n4022 ) ;
  assign n4048 = n2279 ^ n1208 ^ 1'b0 ;
  assign n4049 = ( n1252 & n4047 ) | ( n1252 & n4048 ) | ( n4047 & n4048 ) ;
  assign n4050 = ( ~n733 & n1554 ) | ( ~n733 & n4049 ) | ( n1554 & n4049 ) ;
  assign n4054 = n4053 ^ n4050 ^ x103 ;
  assign n4055 = ( ~x21 & n1861 ) | ( ~x21 & n4054 ) | ( n1861 & n4054 ) ;
  assign n4056 = ( n387 & n2204 ) | ( n387 & n4055 ) | ( n2204 & n4055 ) ;
  assign n4057 = n2880 ^ n2322 ^ 1'b0 ;
  assign n4058 = n4057 ^ n3673 ^ n3048 ;
  assign n4059 = n4058 ^ n3289 ^ n974 ;
  assign n4060 = ( ~n271 & n2136 ) | ( ~n271 & n4059 ) | ( n2136 & n4059 ) ;
  assign n4061 = ( n649 & ~n1387 ) | ( n649 & n2010 ) | ( ~n1387 & n2010 ) ;
  assign n4062 = n4061 ^ n3476 ^ n2975 ;
  assign n4063 = n4062 ^ n2583 ^ n658 ;
  assign n4064 = n4063 ^ n2694 ^ n1089 ;
  assign n4065 = ( n4056 & n4060 ) | ( n4056 & ~n4064 ) | ( n4060 & ~n4064 ) ;
  assign n4067 = n4066 ^ n4065 ^ n1589 ;
  assign n4068 = ( ~n1477 & n2274 ) | ( ~n1477 & n3275 ) | ( n2274 & n3275 ) ;
  assign n4069 = n4068 ^ n1323 ^ n232 ;
  assign n4070 = n1904 ^ n880 ^ 1'b0 ;
  assign n4071 = ~n452 & n4070 ;
  assign n4072 = ( ~n3623 & n4069 ) | ( ~n3623 & n4071 ) | ( n4069 & n4071 ) ;
  assign n4073 = ( n442 & n1845 ) | ( n442 & ~n4072 ) | ( n1845 & ~n4072 ) ;
  assign n4082 = ( n2315 & ~n2775 ) | ( n2315 & n3271 ) | ( ~n2775 & n3271 ) ;
  assign n4080 = n3105 ^ n2479 ^ 1'b0 ;
  assign n4081 = n1160 | n4080 ;
  assign n4083 = n4082 ^ n4081 ^ 1'b0 ;
  assign n4074 = n3164 ^ n2786 ^ n1494 ;
  assign n4075 = n1036 & n3255 ;
  assign n4076 = n1806 ^ n1313 ^ n999 ;
  assign n4077 = n4076 ^ n1784 ^ n1036 ;
  assign n4078 = n4077 ^ n2011 ^ 1'b0 ;
  assign n4079 = ( ~n4074 & n4075 ) | ( ~n4074 & n4078 ) | ( n4075 & n4078 ) ;
  assign n4084 = n4083 ^ n4079 ^ n2907 ;
  assign n4085 = n2618 ^ n1775 ^ n1756 ;
  assign n4086 = n1380 ^ n1273 ^ n596 ;
  assign n4087 = ( x55 & ~n1541 ) | ( x55 & n4086 ) | ( ~n1541 & n4086 ) ;
  assign n4088 = ( ~n2509 & n4085 ) | ( ~n2509 & n4087 ) | ( n4085 & n4087 ) ;
  assign n4089 = n3957 ^ n2895 ^ n1976 ;
  assign n4090 = n2682 ^ n1901 ^ n450 ;
  assign n4091 = ( n282 & n411 ) | ( n282 & n814 ) | ( n411 & n814 ) ;
  assign n4092 = n3661 & ~n4091 ;
  assign n4093 = n4092 ^ n3965 ^ 1'b0 ;
  assign n4094 = n4093 ^ n750 ^ n500 ;
  assign n4095 = n296 | n4094 ;
  assign n4099 = ( n535 & n999 ) | ( n535 & n3827 ) | ( n999 & n3827 ) ;
  assign n4096 = ( ~n222 & n3049 ) | ( ~n222 & n3519 ) | ( n3049 & n3519 ) ;
  assign n4097 = ( ~n1295 & n2413 ) | ( ~n1295 & n4096 ) | ( n2413 & n4096 ) ;
  assign n4098 = ( n711 & n826 ) | ( n711 & n4097 ) | ( n826 & n4097 ) ;
  assign n4100 = n4099 ^ n4098 ^ 1'b0 ;
  assign n4101 = n4100 ^ n3633 ^ n3494 ;
  assign n4103 = n2060 ^ n726 ^ 1'b0 ;
  assign n4104 = n1324 | n4103 ;
  assign n4105 = ( n627 & ~n858 ) | ( n627 & n4104 ) | ( ~n858 & n4104 ) ;
  assign n4102 = n3139 ^ n1366 ^ n721 ;
  assign n4106 = n4105 ^ n4102 ^ n537 ;
  assign n4123 = n3255 ^ n2177 ^ n1088 ;
  assign n4120 = ( ~n717 & n1191 ) | ( ~n717 & n3070 ) | ( n1191 & n3070 ) ;
  assign n4121 = n4120 ^ n3392 ^ n646 ;
  assign n4118 = n2513 ^ n408 ^ 1'b0 ;
  assign n4119 = ~n2220 & n4118 ;
  assign n4122 = n4121 ^ n4119 ^ 1'b0 ;
  assign n4114 = n1215 & ~n1460 ;
  assign n4115 = n4114 ^ n3777 ^ 1'b0 ;
  assign n4116 = n4115 ^ n2083 ^ n474 ;
  assign n4109 = n1606 ^ n676 ^ 1'b0 ;
  assign n4110 = n884 & n4109 ;
  assign n4111 = n4110 ^ x0 ^ 1'b0 ;
  assign n4112 = n3547 & n4111 ;
  assign n4113 = ( n2144 & n2706 ) | ( n2144 & ~n4112 ) | ( n2706 & ~n4112 ) ;
  assign n4107 = ( n1808 & n2876 ) | ( n1808 & ~n3447 ) | ( n2876 & ~n3447 ) ;
  assign n4108 = ( n1380 & n3808 ) | ( n1380 & n4107 ) | ( n3808 & n4107 ) ;
  assign n4117 = n4116 ^ n4113 ^ n4108 ;
  assign n4124 = n4123 ^ n4122 ^ n4117 ;
  assign n4130 = n432 ^ n321 ^ n313 ;
  assign n4128 = n2098 ^ n1050 ^ n796 ;
  assign n4129 = ( n2511 & ~n3751 ) | ( n2511 & n4128 ) | ( ~n3751 & n4128 ) ;
  assign n4126 = n3845 ^ n3428 ^ n3136 ;
  assign n4125 = ~n997 & n2017 ;
  assign n4127 = n4126 ^ n4125 ^ 1'b0 ;
  assign n4131 = n4130 ^ n4129 ^ n4127 ;
  assign n4132 = n4131 ^ n354 ^ x26 ;
  assign n4133 = n2525 & ~n3792 ;
  assign n4134 = ( n3839 & n4132 ) | ( n3839 & ~n4133 ) | ( n4132 & ~n4133 ) ;
  assign n4135 = ~n1100 & n4134 ;
  assign n4136 = ~n2948 & n3550 ;
  assign n4145 = n2612 ^ n1735 ^ n1677 ;
  assign n4144 = n1057 ^ n824 ^ n791 ;
  assign n4141 = ( n218 & n980 ) | ( n218 & ~n1848 ) | ( n980 & ~n1848 ) ;
  assign n4142 = n4141 ^ n3139 ^ n1588 ;
  assign n4139 = ( n1436 & ~n2226 ) | ( n1436 & n3048 ) | ( ~n2226 & n3048 ) ;
  assign n4140 = n4139 ^ n1179 ^ n325 ;
  assign n4137 = n3046 ^ n717 ^ x42 ;
  assign n4138 = n4137 ^ n1466 ^ n686 ;
  assign n4143 = n4142 ^ n4140 ^ n4138 ;
  assign n4146 = n4145 ^ n4144 ^ n4143 ;
  assign n4147 = n3597 & ~n4146 ;
  assign n4148 = n4136 & n4147 ;
  assign n4149 = ( ~n2035 & n2306 ) | ( ~n2035 & n3491 ) | ( n2306 & n3491 ) ;
  assign n4153 = n2572 ^ n1610 ^ x123 ;
  assign n4150 = ( ~n1693 & n2082 ) | ( ~n1693 & n3938 ) | ( n2082 & n3938 ) ;
  assign n4151 = ~n1380 & n4150 ;
  assign n4152 = n4151 ^ n4074 ^ n799 ;
  assign n4154 = n4153 ^ n4152 ^ x81 ;
  assign n4155 = ( n1442 & n4149 ) | ( n1442 & ~n4154 ) | ( n4149 & ~n4154 ) ;
  assign n4156 = ( n181 & n421 ) | ( n181 & n1052 ) | ( n421 & n1052 ) ;
  assign n4157 = ( n1063 & n1120 ) | ( n1063 & n2951 ) | ( n1120 & n2951 ) ;
  assign n4158 = n4156 & n4157 ;
  assign n4159 = ( n1452 & n4155 ) | ( n1452 & ~n4158 ) | ( n4155 & ~n4158 ) ;
  assign n4160 = ( ~n471 & n549 ) | ( ~n471 & n1328 ) | ( n549 & n1328 ) ;
  assign n4161 = n940 ^ n676 ^ n524 ;
  assign n4162 = ( x57 & n621 ) | ( x57 & n2243 ) | ( n621 & n2243 ) ;
  assign n4163 = ( n4160 & n4161 ) | ( n4160 & n4162 ) | ( n4161 & n4162 ) ;
  assign n4164 = n2465 ^ n1647 ^ 1'b0 ;
  assign n4165 = n256 & n4164 ;
  assign n4166 = ( n594 & ~n3840 ) | ( n594 & n4165 ) | ( ~n3840 & n4165 ) ;
  assign n4169 = n1933 ^ n351 ^ 1'b0 ;
  assign n4170 = n1442 & n4169 ;
  assign n4167 = ( ~n506 & n1470 ) | ( ~n506 & n3390 ) | ( n1470 & n3390 ) ;
  assign n4168 = n4167 ^ n3481 ^ n1034 ;
  assign n4171 = n4170 ^ n4168 ^ n988 ;
  assign n4178 = ( n296 & ~n1029 ) | ( n296 & n1304 ) | ( ~n1029 & n1304 ) ;
  assign n4179 = n1991 & n4178 ;
  assign n4180 = n4179 ^ n438 ^ 1'b0 ;
  assign n4173 = ( ~x41 & n1570 ) | ( ~x41 & n2487 ) | ( n1570 & n2487 ) ;
  assign n4174 = ( ~x51 & n1855 ) | ( ~x51 & n4173 ) | ( n1855 & n4173 ) ;
  assign n4175 = n4174 ^ n3887 ^ n3163 ;
  assign n4176 = n4175 ^ n3204 ^ n665 ;
  assign n4172 = n3807 ^ n3602 ^ n535 ;
  assign n4177 = n4176 ^ n4172 ^ 1'b0 ;
  assign n4181 = n4180 ^ n4177 ^ n2373 ;
  assign n4182 = ( n4166 & ~n4171 ) | ( n4166 & n4181 ) | ( ~n4171 & n4181 ) ;
  assign n4192 = n3361 ^ n2045 ^ x20 ;
  assign n4190 = ( n324 & n671 ) | ( n324 & ~n2101 ) | ( n671 & ~n2101 ) ;
  assign n4191 = ( n173 & ~n1941 ) | ( n173 & n4190 ) | ( ~n1941 & n4190 ) ;
  assign n4186 = ( ~n206 & n377 ) | ( ~n206 & n1571 ) | ( n377 & n1571 ) ;
  assign n4187 = ( n1258 & n2066 ) | ( n1258 & ~n4186 ) | ( n2066 & ~n4186 ) ;
  assign n4184 = ( n731 & n2360 ) | ( n731 & n2623 ) | ( n2360 & n2623 ) ;
  assign n4185 = n2721 & n4184 ;
  assign n4188 = n4187 ^ n4185 ^ 1'b0 ;
  assign n4183 = ( x34 & ~n942 ) | ( x34 & n3199 ) | ( ~n942 & n3199 ) ;
  assign n4189 = n4188 ^ n4183 ^ n3827 ;
  assign n4193 = n4192 ^ n4191 ^ n4189 ;
  assign n4199 = n3500 ^ n1442 ^ n410 ;
  assign n4196 = n2075 & ~n2703 ;
  assign n4194 = n1546 ^ n1056 ^ 1'b0 ;
  assign n4195 = ( n726 & ~n1920 ) | ( n726 & n4194 ) | ( ~n1920 & n4194 ) ;
  assign n4197 = n4196 ^ n4195 ^ n661 ;
  assign n4198 = n4197 ^ n2624 ^ n1960 ;
  assign n4200 = n4199 ^ n4198 ^ n1198 ;
  assign n4215 = n1748 ^ n864 ^ 1'b0 ;
  assign n4216 = ~n1477 & n4215 ;
  assign n4201 = ~x43 & n2564 ;
  assign n4202 = n692 | n1473 ;
  assign n4203 = n3783 & ~n4202 ;
  assign n4204 = n482 | n3137 ;
  assign n4207 = ( n374 & n1976 ) | ( n374 & ~n3366 ) | ( n1976 & ~n3366 ) ;
  assign n4205 = n2463 ^ n334 ^ 1'b0 ;
  assign n4206 = n4205 ^ n1537 ^ n1137 ;
  assign n4208 = n4207 ^ n4206 ^ 1'b0 ;
  assign n4209 = ~n527 & n4208 ;
  assign n4210 = ( n3661 & n4204 ) | ( n3661 & ~n4209 ) | ( n4204 & ~n4209 ) ;
  assign n4211 = ( n3847 & ~n4203 ) | ( n3847 & n4210 ) | ( ~n4203 & n4210 ) ;
  assign n4212 = ( n2214 & ~n4201 ) | ( n2214 & n4211 ) | ( ~n4201 & n4211 ) ;
  assign n4213 = ( n1808 & n2766 ) | ( n1808 & ~n4212 ) | ( n2766 & ~n4212 ) ;
  assign n4214 = ~n3392 & n4213 ;
  assign n4217 = n4216 ^ n4214 ^ 1'b0 ;
  assign n4218 = n4217 ^ n2015 ^ 1'b0 ;
  assign n4219 = n1230 ^ n854 ^ n765 ;
  assign n4220 = ( ~n1085 & n1710 ) | ( ~n1085 & n4219 ) | ( n1710 & n4219 ) ;
  assign n4221 = n3201 ^ n1257 ^ n877 ;
  assign n4222 = ( n3141 & ~n4220 ) | ( n3141 & n4221 ) | ( ~n4220 & n4221 ) ;
  assign n4223 = n1387 | n4222 ;
  assign n4224 = n1163 | n1352 ;
  assign n4225 = n4224 ^ n2930 ^ 1'b0 ;
  assign n4226 = n3594 ^ n996 ^ 1'b0 ;
  assign n4227 = n4226 ^ n2481 ^ 1'b0 ;
  assign n4228 = n2617 | n4227 ;
  assign n4229 = ( n1682 & n3516 ) | ( n1682 & n4228 ) | ( n3516 & n4228 ) ;
  assign n4230 = ( n1010 & ~n4225 ) | ( n1010 & n4229 ) | ( ~n4225 & n4229 ) ;
  assign n4231 = n655 | n1684 ;
  assign n4232 = n4231 ^ n3861 ^ n2469 ;
  assign n4233 = ( n377 & n511 ) | ( n377 & ~n1249 ) | ( n511 & ~n1249 ) ;
  assign n4234 = ( n1991 & n3386 ) | ( n1991 & ~n4233 ) | ( n3386 & ~n4233 ) ;
  assign n4235 = ( n1400 & n3150 ) | ( n1400 & ~n4234 ) | ( n3150 & ~n4234 ) ;
  assign n4236 = n4235 ^ n2960 ^ n910 ;
  assign n4237 = n4236 ^ n2918 ^ n1732 ;
  assign n4238 = n4237 ^ n734 ^ n256 ;
  assign n4239 = ~n4232 & n4238 ;
  assign n4240 = ~n4230 & n4239 ;
  assign n4241 = ( n304 & ~n2436 ) | ( n304 & n3144 ) | ( ~n2436 & n3144 ) ;
  assign n4242 = n1391 ^ n214 ^ 1'b0 ;
  assign n4243 = n4242 ^ n235 ^ x64 ;
  assign n4244 = ( n2987 & n4241 ) | ( n2987 & n4243 ) | ( n4241 & n4243 ) ;
  assign n4245 = n4244 ^ n4178 ^ n3172 ;
  assign n4246 = n3028 ^ n860 ^ n350 ;
  assign n4247 = n2599 & ~n4246 ;
  assign n4248 = n2203 ^ n1787 ^ n1349 ;
  assign n4249 = n1973 ^ n958 ^ n753 ;
  assign n4250 = ( n359 & n482 ) | ( n359 & ~n1437 ) | ( n482 & ~n1437 ) ;
  assign n4251 = ( ~n4094 & n4249 ) | ( ~n4094 & n4250 ) | ( n4249 & n4250 ) ;
  assign n4252 = ( n2762 & n4248 ) | ( n2762 & n4251 ) | ( n4248 & n4251 ) ;
  assign n4253 = ( n1729 & ~n3779 ) | ( n1729 & n4252 ) | ( ~n3779 & n4252 ) ;
  assign n4254 = ( n2080 & n4247 ) | ( n2080 & ~n4253 ) | ( n4247 & ~n4253 ) ;
  assign n4255 = ( n2392 & n3271 ) | ( n2392 & n4130 ) | ( n3271 & n4130 ) ;
  assign n4256 = n2605 ^ n2486 ^ n2385 ;
  assign n4257 = n4256 ^ n3762 ^ n1129 ;
  assign n4258 = ( n174 & n3247 ) | ( n174 & n3300 ) | ( n3247 & n3300 ) ;
  assign n4259 = n4258 ^ n1321 ^ x111 ;
  assign n4260 = ~n4257 & n4259 ;
  assign n4261 = n4150 & n4260 ;
  assign n4265 = n4057 ^ n977 ^ 1'b0 ;
  assign n4266 = ( n1928 & n2443 ) | ( n1928 & n3537 ) | ( n2443 & n3537 ) ;
  assign n4267 = ( n1943 & n4265 ) | ( n1943 & n4266 ) | ( n4265 & n4266 ) ;
  assign n4262 = ( ~n214 & n657 ) | ( ~n214 & n914 ) | ( n657 & n914 ) ;
  assign n4263 = ( ~n1044 & n2427 ) | ( ~n1044 & n3168 ) | ( n2427 & n3168 ) ;
  assign n4264 = ~n4262 & n4263 ;
  assign n4268 = n4267 ^ n4264 ^ n1088 ;
  assign n4276 = ~n1888 & n1921 ;
  assign n4277 = n3655 & n4276 ;
  assign n4274 = ( ~n544 & n1041 ) | ( ~n544 & n1890 ) | ( n1041 & n1890 ) ;
  assign n4275 = ( n3239 & n3520 ) | ( n3239 & n4274 ) | ( n3520 & n4274 ) ;
  assign n4269 = n466 ^ n387 ^ x48 ;
  assign n4270 = n4269 ^ n1516 ^ 1'b0 ;
  assign n4271 = ( n1619 & ~n2948 ) | ( n1619 & n4270 ) | ( ~n2948 & n4270 ) ;
  assign n4272 = n3280 | n4271 ;
  assign n4273 = n4272 ^ n178 ^ 1'b0 ;
  assign n4278 = n4277 ^ n4275 ^ n4273 ;
  assign n4279 = ( ~n623 & n3387 ) | ( ~n623 & n4278 ) | ( n3387 & n4278 ) ;
  assign n4280 = n4279 ^ n4081 ^ x25 ;
  assign n4283 = n2806 ^ n661 ^ x47 ;
  assign n4284 = n3791 ^ n1123 ^ 1'b0 ;
  assign n4285 = ~n4283 & n4284 ;
  assign n4281 = n2575 ^ n749 ^ 1'b0 ;
  assign n4282 = n4281 ^ n3225 ^ n189 ;
  assign n4286 = n4285 ^ n4282 ^ n1104 ;
  assign n4289 = n1278 ^ n679 ^ n186 ;
  assign n4288 = n2733 ^ n1226 ^ n845 ;
  assign n4290 = n4289 ^ n4288 ^ n1185 ;
  assign n4291 = ( n638 & n1652 ) | ( n638 & ~n4290 ) | ( n1652 & ~n4290 ) ;
  assign n4287 = n4199 ^ n1844 ^ n948 ;
  assign n4292 = n4291 ^ n4287 ^ n1689 ;
  assign n4293 = n2787 ^ n1725 ^ n150 ;
  assign n4294 = n4293 ^ n3556 ^ n1759 ;
  assign n4295 = n4294 ^ n4117 ^ n1644 ;
  assign n4296 = ( ~n863 & n2607 ) | ( ~n863 & n2960 ) | ( n2607 & n2960 ) ;
  assign n4297 = ( n2224 & n2541 ) | ( n2224 & n3136 ) | ( n2541 & n3136 ) ;
  assign n4298 = n4297 ^ n2476 ^ n877 ;
  assign n4299 = ( ~n3806 & n4296 ) | ( ~n3806 & n4298 ) | ( n4296 & n4298 ) ;
  assign n4300 = ~n2151 & n4299 ;
  assign n4301 = n4300 ^ n1059 ^ 1'b0 ;
  assign n4302 = ( ~n610 & n1109 ) | ( ~n610 & n1801 ) | ( n1109 & n1801 ) ;
  assign n4303 = ( n1473 & n1540 ) | ( n1473 & n4302 ) | ( n1540 & n4302 ) ;
  assign n4312 = n2622 ^ x53 ^ 1'b0 ;
  assign n4313 = ~n1503 & n4312 ;
  assign n4308 = n2580 ^ n2397 ^ 1'b0 ;
  assign n4309 = n2980 | n4308 ;
  assign n4310 = n4309 ^ n3187 ^ n1386 ;
  assign n4311 = n4310 ^ n470 ^ n174 ;
  assign n4306 = ( n356 & ~n2710 ) | ( n356 & n3075 ) | ( ~n2710 & n3075 ) ;
  assign n4304 = n1597 ^ n1002 ^ x44 ;
  assign n4305 = ~n3582 & n4304 ;
  assign n4307 = n4306 ^ n4305 ^ 1'b0 ;
  assign n4314 = n4313 ^ n4311 ^ n4307 ;
  assign n4315 = n4303 & n4314 ;
  assign n4316 = n3401 ^ n2293 ^ 1'b0 ;
  assign n4317 = n1213 | n4316 ;
  assign n4318 = ( ~n3071 & n3870 ) | ( ~n3071 & n4317 ) | ( n3870 & n4317 ) ;
  assign n4329 = n1271 ^ n478 ^ x18 ;
  assign n4330 = n545 & ~n4329 ;
  assign n4331 = n4330 ^ n2627 ^ 1'b0 ;
  assign n4326 = ( ~n958 & n1182 ) | ( ~n958 & n2314 ) | ( n1182 & n2314 ) ;
  assign n4327 = n3919 ^ n1783 ^ n382 ;
  assign n4328 = ( ~n2776 & n4326 ) | ( ~n2776 & n4327 ) | ( n4326 & n4327 ) ;
  assign n4319 = ( ~n1822 & n2813 ) | ( ~n1822 & n4145 ) | ( n2813 & n4145 ) ;
  assign n4320 = n235 & n4319 ;
  assign n4321 = n4320 ^ n4020 ^ 1'b0 ;
  assign n4322 = ( x63 & ~n324 ) | ( x63 & n2806 ) | ( ~n324 & n2806 ) ;
  assign n4323 = ( n443 & n4321 ) | ( n443 & n4322 ) | ( n4321 & n4322 ) ;
  assign n4324 = n4323 ^ n751 ^ 1'b0 ;
  assign n4325 = n1761 & n4324 ;
  assign n4332 = n4331 ^ n4328 ^ n4325 ;
  assign n4333 = n3965 ^ n3125 ^ n2608 ;
  assign n4337 = ~n2143 & n3100 ;
  assign n4338 = n634 & n4337 ;
  assign n4339 = n4338 ^ n3159 ^ n1562 ;
  assign n4335 = ( n419 & n426 ) | ( n419 & n1863 ) | ( n426 & n1863 ) ;
  assign n4336 = n4335 ^ n2708 ^ n1488 ;
  assign n4334 = n4278 ^ n2382 ^ n1466 ;
  assign n4340 = n4339 ^ n4336 ^ n4334 ;
  assign n4353 = n643 | n2726 ;
  assign n4354 = n4353 ^ n3287 ^ 1'b0 ;
  assign n4355 = ( ~n2329 & n3401 ) | ( ~n2329 & n4354 ) | ( n3401 & n4354 ) ;
  assign n4356 = ( n602 & ~n2810 ) | ( n602 & n4355 ) | ( ~n2810 & n4355 ) ;
  assign n4349 = n2958 ^ n2247 ^ n2208 ;
  assign n4347 = ( x10 & ~n175 ) | ( x10 & n2080 ) | ( ~n175 & n2080 ) ;
  assign n4348 = ( n1608 & n3310 ) | ( n1608 & ~n4347 ) | ( n3310 & ~n4347 ) ;
  assign n4350 = n4349 ^ n4348 ^ n785 ;
  assign n4341 = n1154 & ~n3313 ;
  assign n4342 = n1012 & n4341 ;
  assign n4343 = ( ~n1479 & n1642 ) | ( ~n1479 & n2009 ) | ( n1642 & n2009 ) ;
  assign n4344 = n4343 ^ n3876 ^ n3479 ;
  assign n4345 = ~n4342 & n4344 ;
  assign n4346 = n4345 ^ n1362 ^ 1'b0 ;
  assign n4351 = n4350 ^ n4346 ^ n1091 ;
  assign n4352 = ( ~n235 & n3740 ) | ( ~n235 & n4351 ) | ( n3740 & n4351 ) ;
  assign n4357 = n4356 ^ n4352 ^ n1044 ;
  assign n4358 = n4357 ^ n4034 ^ n621 ;
  assign n4369 = n2112 ^ n879 ^ x2 ;
  assign n4370 = n4369 ^ n1772 ^ n573 ;
  assign n4368 = ( n334 & ~n1316 ) | ( n334 & n2703 ) | ( ~n1316 & n2703 ) ;
  assign n4371 = n4370 ^ n4368 ^ n2235 ;
  assign n4362 = n1114 | n2081 ;
  assign n4363 = ~n995 & n4362 ;
  assign n4364 = n3281 & n4363 ;
  assign n4365 = n4364 ^ n2531 ^ 1'b0 ;
  assign n4359 = ( n650 & n2086 ) | ( n650 & n3934 ) | ( n2086 & n3934 ) ;
  assign n4360 = n4359 ^ n3570 ^ 1'b0 ;
  assign n4361 = n4360 ^ n3977 ^ n852 ;
  assign n4366 = n4365 ^ n4361 ^ 1'b0 ;
  assign n4367 = n3280 | n4366 ;
  assign n4372 = n4371 ^ n4367 ^ n2176 ;
  assign n4373 = n641 & n1587 ;
  assign n4374 = n4373 ^ n2966 ^ 1'b0 ;
  assign n4375 = n4374 ^ n2123 ^ n198 ;
  assign n4376 = n2674 ^ n1609 ^ 1'b0 ;
  assign n4377 = ( n175 & n1628 ) | ( n175 & ~n4376 ) | ( n1628 & ~n4376 ) ;
  assign n4378 = ( n2415 & ~n2894 ) | ( n2415 & n4377 ) | ( ~n2894 & n4377 ) ;
  assign n4379 = n623 ^ n445 ^ x57 ;
  assign n4387 = ( n2590 & ~n2993 ) | ( n2590 & n4137 ) | ( ~n2993 & n4137 ) ;
  assign n4380 = ( n985 & n2266 ) | ( n985 & ~n2383 ) | ( n2266 & ~n2383 ) ;
  assign n4381 = n1931 ^ n517 ^ 1'b0 ;
  assign n4382 = n4381 ^ n1410 ^ n674 ;
  assign n4383 = ( ~x3 & n3462 ) | ( ~x3 & n4382 ) | ( n3462 & n4382 ) ;
  assign n4384 = ~n4380 & n4383 ;
  assign n4385 = ( n534 & n3656 ) | ( n534 & ~n4384 ) | ( n3656 & ~n4384 ) ;
  assign n4386 = ( n1486 & n2876 ) | ( n1486 & ~n4385 ) | ( n2876 & ~n4385 ) ;
  assign n4388 = n4387 ^ n4386 ^ n1576 ;
  assign n4389 = n4388 ^ n3699 ^ 1'b0 ;
  assign n4390 = ~n4379 & n4389 ;
  assign n4407 = n3581 ^ n2035 ^ 1'b0 ;
  assign n4408 = n2834 | n4407 ;
  assign n4409 = n4408 ^ n1880 ^ x34 ;
  assign n4410 = n261 | n4409 ;
  assign n4411 = n4410 ^ n385 ^ 1'b0 ;
  assign n4397 = n1894 ^ n1749 ^ n1154 ;
  assign n4394 = n1931 ^ n575 ^ n435 ;
  assign n4395 = n4394 ^ n1667 ^ n774 ;
  assign n4396 = n4395 ^ n745 ^ x2 ;
  assign n4391 = n966 ^ n871 ^ n463 ;
  assign n4392 = n2256 ^ n2120 ^ n900 ;
  assign n4393 = ( n1354 & ~n4391 ) | ( n1354 & n4392 ) | ( ~n4391 & n4392 ) ;
  assign n4398 = n4397 ^ n4396 ^ n4393 ;
  assign n4399 = ( n1302 & ~n3043 ) | ( n1302 & n4091 ) | ( ~n3043 & n4091 ) ;
  assign n4400 = ( n646 & ~n1407 ) | ( n646 & n4050 ) | ( ~n1407 & n4050 ) ;
  assign n4401 = ( n1940 & ~n4399 ) | ( n1940 & n4400 ) | ( ~n4399 & n4400 ) ;
  assign n4402 = ( ~n521 & n606 ) | ( ~n521 & n875 ) | ( n606 & n875 ) ;
  assign n4403 = n3758 ^ n3396 ^ n2860 ;
  assign n4404 = ( n2677 & n4402 ) | ( n2677 & ~n4403 ) | ( n4402 & ~n4403 ) ;
  assign n4405 = ~n4401 & n4404 ;
  assign n4406 = ~n4398 & n4405 ;
  assign n4412 = n4411 ^ n4406 ^ n1366 ;
  assign n4416 = n2466 ^ n390 ^ 1'b0 ;
  assign n4413 = ( n480 & ~n818 ) | ( n480 & n1452 ) | ( ~n818 & n1452 ) ;
  assign n4414 = ( n2741 & n4399 ) | ( n2741 & ~n4413 ) | ( n4399 & ~n4413 ) ;
  assign n4415 = ( n1287 & n4107 ) | ( n1287 & n4414 ) | ( n4107 & n4414 ) ;
  assign n4417 = n4416 ^ n4415 ^ n254 ;
  assign n4418 = n2811 ^ n2079 ^ n1429 ;
  assign n4419 = ( n1711 & n4401 ) | ( n1711 & n4418 ) | ( n4401 & n4418 ) ;
  assign n4420 = ( n428 & n575 ) | ( n428 & n2287 ) | ( n575 & n2287 ) ;
  assign n4421 = n697 & n1414 ;
  assign n4422 = ~n4420 & n4421 ;
  assign n4423 = ( n1796 & n1901 ) | ( n1796 & n4422 ) | ( n1901 & n4422 ) ;
  assign n4424 = n4423 ^ n2251 ^ n504 ;
  assign n4425 = ( ~n3138 & n4419 ) | ( ~n3138 & n4424 ) | ( n4419 & n4424 ) ;
  assign n4426 = ( ~n2478 & n2496 ) | ( ~n2478 & n4344 ) | ( n2496 & n4344 ) ;
  assign n4427 = n4426 ^ n3642 ^ 1'b0 ;
  assign n4429 = ( ~n339 & n1534 ) | ( ~n339 & n2442 ) | ( n1534 & n2442 ) ;
  assign n4430 = ( n584 & ~n2601 ) | ( n584 & n4429 ) | ( ~n2601 & n4429 ) ;
  assign n4428 = n895 | n903 ;
  assign n4431 = n4430 ^ n4428 ^ 1'b0 ;
  assign n4432 = n4431 ^ n1625 ^ n1316 ;
  assign n4440 = n3352 ^ n2449 ^ x23 ;
  assign n4433 = n1931 ^ n692 ^ n405 ;
  assign n4434 = n4433 ^ n2905 ^ n1689 ;
  assign n4435 = ( n884 & n1818 ) | ( n884 & ~n2515 ) | ( n1818 & ~n2515 ) ;
  assign n4436 = n519 | n788 ;
  assign n4437 = n4436 ^ n3429 ^ n1359 ;
  assign n4438 = n4435 & n4437 ;
  assign n4439 = n4434 & ~n4438 ;
  assign n4441 = n4440 ^ n4439 ^ n2810 ;
  assign n4442 = ( n411 & n981 ) | ( n411 & n1133 ) | ( n981 & n1133 ) ;
  assign n4443 = n986 ^ n465 ^ n325 ;
  assign n4444 = n4443 ^ n2907 ^ n1181 ;
  assign n4445 = ( ~n319 & n3218 ) | ( ~n319 & n4444 ) | ( n3218 & n4444 ) ;
  assign n4446 = ( n474 & n514 ) | ( n474 & ~n2761 ) | ( n514 & ~n2761 ) ;
  assign n4447 = ( n1566 & n4002 ) | ( n1566 & n4053 ) | ( n4002 & n4053 ) ;
  assign n4448 = ( n4068 & ~n4446 ) | ( n4068 & n4447 ) | ( ~n4446 & n4447 ) ;
  assign n4449 = ( n1569 & n4445 ) | ( n1569 & ~n4448 ) | ( n4445 & ~n4448 ) ;
  assign n4450 = ( ~n2414 & n4139 ) | ( ~n2414 & n4449 ) | ( n4139 & n4449 ) ;
  assign n4451 = ( ~n578 & n843 ) | ( ~n578 & n890 ) | ( n843 & n890 ) ;
  assign n4452 = ( n1349 & n2262 ) | ( n1349 & ~n4451 ) | ( n2262 & ~n4451 ) ;
  assign n4453 = n917 & n4452 ;
  assign n4454 = n4453 ^ n2398 ^ 1'b0 ;
  assign n4455 = n2203 ^ n160 ^ 1'b0 ;
  assign n4456 = n4455 ^ n4298 ^ n487 ;
  assign n4457 = ( n1401 & ~n4454 ) | ( n1401 & n4456 ) | ( ~n4454 & n4456 ) ;
  assign n4458 = n4457 ^ n2806 ^ n1000 ;
  assign n4463 = n3550 ^ n1342 ^ n1210 ;
  assign n4459 = ( n954 & n1410 ) | ( n954 & ~n1706 ) | ( n1410 & ~n1706 ) ;
  assign n4460 = n2310 ^ n1634 ^ 1'b0 ;
  assign n4461 = ( n2534 & n2591 ) | ( n2534 & n4460 ) | ( n2591 & n4460 ) ;
  assign n4462 = n4459 & n4461 ;
  assign n4464 = n4463 ^ n4462 ^ 1'b0 ;
  assign n4465 = n4285 ^ n479 ^ 1'b0 ;
  assign n4466 = ( ~n1774 & n4464 ) | ( ~n1774 & n4465 ) | ( n4464 & n4465 ) ;
  assign n4467 = ( ~n1847 & n2668 ) | ( ~n1847 & n4466 ) | ( n2668 & n4466 ) ;
  assign n4475 = n2729 ^ n1892 ^ n832 ;
  assign n4472 = n2605 ^ n861 ^ n212 ;
  assign n4473 = ( ~n2013 & n2918 ) | ( ~n2013 & n4472 ) | ( n2918 & n4472 ) ;
  assign n4474 = ( ~n626 & n968 ) | ( ~n626 & n4473 ) | ( n968 & n4473 ) ;
  assign n4469 = ( n999 & n1528 ) | ( n999 & ~n2195 ) | ( n1528 & ~n2195 ) ;
  assign n4470 = n4469 ^ n3639 ^ n1367 ;
  assign n4468 = ( ~n1300 & n1716 ) | ( ~n1300 & n4258 ) | ( n1716 & n4258 ) ;
  assign n4471 = n4470 ^ n4468 ^ n4343 ;
  assign n4476 = n4475 ^ n4474 ^ n4471 ;
  assign n4477 = n4155 ^ n2590 ^ n2508 ;
  assign n4478 = n1274 ^ n1043 ^ 1'b0 ;
  assign n4479 = n4478 ^ n3618 ^ n2514 ;
  assign n4480 = ( ~n1503 & n2473 ) | ( ~n1503 & n4479 ) | ( n2473 & n4479 ) ;
  assign n4481 = ( n2254 & ~n4477 ) | ( n2254 & n4480 ) | ( ~n4477 & n4480 ) ;
  assign n4482 = n3362 ^ n973 ^ 1'b0 ;
  assign n4483 = ( n1267 & n1279 ) | ( n1267 & n4482 ) | ( n1279 & n4482 ) ;
  assign n4484 = n4483 ^ n1953 ^ 1'b0 ;
  assign n4493 = n3827 ^ n2332 ^ n2275 ;
  assign n4494 = ( n1456 & ~n4444 ) | ( n1456 & n4493 ) | ( ~n4444 & n4493 ) ;
  assign n4487 = n1661 ^ n1039 ^ n900 ;
  assign n4488 = n4487 ^ n2032 ^ x89 ;
  assign n4485 = ( n689 & ~n1690 ) | ( n689 & n1813 ) | ( ~n1690 & n1813 ) ;
  assign n4486 = n4485 ^ n2298 ^ x86 ;
  assign n4489 = n4488 ^ n4486 ^ 1'b0 ;
  assign n4490 = n2652 & n4489 ;
  assign n4491 = n4490 ^ n2804 ^ n2365 ;
  assign n4492 = ( n2274 & ~n3105 ) | ( n2274 & n4491 ) | ( ~n3105 & n4491 ) ;
  assign n4495 = n4494 ^ n4492 ^ n2209 ;
  assign n4496 = n474 & n2046 ;
  assign n4497 = n1906 & n1939 ;
  assign n4498 = n4497 ^ n3519 ^ n1172 ;
  assign n4499 = n4180 ^ n3310 ^ n386 ;
  assign n4500 = n4499 ^ n3056 ^ n2136 ;
  assign n4501 = n4498 & ~n4500 ;
  assign n4502 = n4496 & ~n4501 ;
  assign n4503 = n4502 ^ n3923 ^ 1'b0 ;
  assign n4504 = n3721 ^ n3633 ^ n1681 ;
  assign n4505 = ( ~n1753 & n1757 ) | ( ~n1753 & n4504 ) | ( n1757 & n4504 ) ;
  assign n4506 = n4505 ^ n1596 ^ n1443 ;
  assign n4507 = n3094 ^ n3071 ^ 1'b0 ;
  assign n4508 = n4480 & ~n4507 ;
  assign n4509 = n2659 & ~n3902 ;
  assign n4510 = n4509 ^ n865 ^ 1'b0 ;
  assign n4513 = n1014 ^ n795 ^ n694 ;
  assign n4514 = ( n1327 & ~n2595 ) | ( n1327 & n4513 ) | ( ~n2595 & n4513 ) ;
  assign n4511 = ( n251 & ~n1686 ) | ( n251 & n2029 ) | ( ~n1686 & n2029 ) ;
  assign n4512 = n4511 ^ n3349 ^ n354 ;
  assign n4515 = n4514 ^ n4512 ^ n2060 ;
  assign n4516 = n3905 & n4515 ;
  assign n4521 = n3476 ^ n1886 ^ n1523 ;
  assign n4518 = ( n588 & ~n1148 ) | ( n588 & n1990 ) | ( ~n1148 & n1990 ) ;
  assign n4519 = ( n215 & n659 ) | ( n215 & n4518 ) | ( n659 & n4518 ) ;
  assign n4517 = ( x72 & n819 ) | ( x72 & ~n1301 ) | ( n819 & ~n1301 ) ;
  assign n4520 = n4519 ^ n4517 ^ n4066 ;
  assign n4522 = n4521 ^ n4520 ^ n2058 ;
  assign n4523 = ~n2037 & n4522 ;
  assign n4524 = n4516 & n4523 ;
  assign n4525 = ~n1602 & n4154 ;
  assign n4526 = n4525 ^ n3234 ^ n3100 ;
  assign n4528 = ( n1124 & n1543 ) | ( n1124 & n3580 ) | ( n1543 & n3580 ) ;
  assign n4527 = n2810 | n3044 ;
  assign n4529 = n4528 ^ n4527 ^ n3907 ;
  assign n4532 = ( n287 & ~n1274 ) | ( n287 & n1644 ) | ( ~n1274 & n1644 ) ;
  assign n4533 = n4532 ^ n1684 ^ 1'b0 ;
  assign n4534 = n4533 ^ n4120 ^ 1'b0 ;
  assign n4535 = n664 | n4534 ;
  assign n4530 = ( n740 & n800 ) | ( n740 & n3645 ) | ( n800 & n3645 ) ;
  assign n4531 = ~n2978 & n4530 ;
  assign n4536 = n4535 ^ n4531 ^ 1'b0 ;
  assign n4537 = n807 ^ n504 ^ n420 ;
  assign n4538 = ~n1770 & n4537 ;
  assign n4539 = n181 & n4538 ;
  assign n4541 = ( n1035 & n1386 ) | ( n1035 & ~n2267 ) | ( n1386 & ~n2267 ) ;
  assign n4540 = n3867 ^ n2520 ^ n965 ;
  assign n4542 = n4541 ^ n4540 ^ 1'b0 ;
  assign n4543 = ~n4539 & n4542 ;
  assign n4544 = n4543 ^ n4265 ^ n132 ;
  assign n4545 = ( n159 & n4536 ) | ( n159 & ~n4544 ) | ( n4536 & ~n4544 ) ;
  assign n4546 = x20 & ~n1522 ;
  assign n4547 = ( ~n783 & n1193 ) | ( ~n783 & n4546 ) | ( n1193 & n4546 ) ;
  assign n4548 = n2156 ^ n566 ^ 1'b0 ;
  assign n4549 = n1264 & ~n4548 ;
  assign n4550 = ( ~n1087 & n1357 ) | ( ~n1087 & n1399 ) | ( n1357 & n1399 ) ;
  assign n4551 = n1497 ^ n1345 ^ 1'b0 ;
  assign n4552 = ( ~n1126 & n3892 ) | ( ~n1126 & n4551 ) | ( n3892 & n4551 ) ;
  assign n4553 = ( n1806 & ~n4550 ) | ( n1806 & n4552 ) | ( ~n4550 & n4552 ) ;
  assign n4554 = ( n3724 & n4549 ) | ( n3724 & n4553 ) | ( n4549 & n4553 ) ;
  assign n4557 = ( n207 & ~n1686 ) | ( n207 & n2030 ) | ( ~n1686 & n2030 ) ;
  assign n4555 = n714 ^ n300 ^ n181 ;
  assign n4556 = ( n1459 & n1805 ) | ( n1459 & ~n4555 ) | ( n1805 & ~n4555 ) ;
  assign n4558 = n4557 ^ n4556 ^ n1633 ;
  assign n4559 = n2265 ^ n1942 ^ n387 ;
  assign n4560 = n559 & ~n4487 ;
  assign n4561 = ~n4559 & n4560 ;
  assign n4562 = ( n2040 & n4558 ) | ( n2040 & ~n4561 ) | ( n4558 & ~n4561 ) ;
  assign n4563 = n2008 ^ n1444 ^ n639 ;
  assign n4564 = n3661 & ~n4563 ;
  assign n4565 = n4562 & n4564 ;
  assign n4568 = n257 & ~n1302 ;
  assign n4569 = n4568 ^ n202 ^ 1'b0 ;
  assign n4570 = n4569 ^ n4410 ^ n2273 ;
  assign n4566 = ( n707 & ~n989 ) | ( n707 & n2186 ) | ( ~n989 & n2186 ) ;
  assign n4567 = ( n3369 & n3431 ) | ( n3369 & n4566 ) | ( n3431 & n4566 ) ;
  assign n4571 = n4570 ^ n4567 ^ 1'b0 ;
  assign n4572 = n4571 ^ n1143 ^ 1'b0 ;
  assign n4573 = n4556 ^ n4093 ^ n758 ;
  assign n4574 = ( n264 & ~n4262 ) | ( n264 & n4451 ) | ( ~n4262 & n4451 ) ;
  assign n4575 = ( ~n1549 & n1612 ) | ( ~n1549 & n3414 ) | ( n1612 & n3414 ) ;
  assign n4576 = ( n1395 & n1822 ) | ( n1395 & ~n2614 ) | ( n1822 & ~n2614 ) ;
  assign n4577 = n4576 ^ n1762 ^ n440 ;
  assign n4578 = ( ~n2854 & n3214 ) | ( ~n2854 & n4577 ) | ( n3214 & n4577 ) ;
  assign n4579 = ~n4575 & n4578 ;
  assign n4580 = n4574 & n4579 ;
  assign n4581 = ( x53 & n913 ) | ( x53 & ~n3325 ) | ( n913 & ~n3325 ) ;
  assign n4582 = n3167 ^ n985 ^ n186 ;
  assign n4583 = ( ~n237 & n3166 ) | ( ~n237 & n4582 ) | ( n3166 & n4582 ) ;
  assign n4584 = ~n4077 & n4583 ;
  assign n4585 = n4581 & n4584 ;
  assign n4586 = n3312 ^ n1695 ^ n577 ;
  assign n4587 = n4586 ^ n2527 ^ n312 ;
  assign n4588 = n4587 ^ n839 ^ 1'b0 ;
  assign n4589 = n4044 ^ n2761 ^ n2414 ;
  assign n4590 = n4589 ^ n2912 ^ n705 ;
  assign n4591 = n1854 ^ n1507 ^ 1'b0 ;
  assign n4592 = ~n4590 & n4591 ;
  assign n4593 = ~n877 & n4592 ;
  assign n4594 = n4593 ^ n2700 ^ n1283 ;
  assign n4595 = n758 & ~n1663 ;
  assign n4596 = ( x108 & n725 ) | ( x108 & n2209 ) | ( n725 & n2209 ) ;
  assign n4597 = ( ~n3066 & n3791 ) | ( ~n3066 & n4596 ) | ( n3791 & n4596 ) ;
  assign n4598 = ( n198 & n1747 ) | ( n198 & n4597 ) | ( n1747 & n4597 ) ;
  assign n4599 = ( n4594 & ~n4595 ) | ( n4594 & n4598 ) | ( ~n4595 & n4598 ) ;
  assign n4600 = ( n3504 & n4588 ) | ( n3504 & n4599 ) | ( n4588 & n4599 ) ;
  assign n4601 = ( n707 & n1211 ) | ( n707 & n4205 ) | ( n1211 & n4205 ) ;
  assign n4614 = ( n478 & n1303 ) | ( n478 & n3939 ) | ( n1303 & n3939 ) ;
  assign n4611 = n1377 ^ n986 ^ n621 ;
  assign n4610 = ( ~n2054 & n2195 ) | ( ~n2054 & n2619 ) | ( n2195 & n2619 ) ;
  assign n4612 = n4611 ^ n4610 ^ n2522 ;
  assign n4613 = x88 & ~n4612 ;
  assign n4606 = n930 | n2528 ;
  assign n4607 = n4606 ^ n3669 ^ 1'b0 ;
  assign n4605 = ( n1411 & n1635 ) | ( n1411 & n1867 ) | ( n1635 & n1867 ) ;
  assign n4602 = n4586 ^ n1009 ^ n826 ;
  assign n4603 = n2558 ^ n2251 ^ 1'b0 ;
  assign n4604 = n4602 & ~n4603 ;
  assign n4608 = n4607 ^ n4605 ^ n4604 ;
  assign n4609 = ( n1202 & ~n1680 ) | ( n1202 & n4608 ) | ( ~n1680 & n4608 ) ;
  assign n4615 = n4614 ^ n4613 ^ n4609 ;
  assign n4628 = ( n465 & ~n985 ) | ( n465 & n1017 ) | ( ~n985 & n1017 ) ;
  assign n4629 = x89 & ~n4628 ;
  assign n4630 = ~n3762 & n4629 ;
  assign n4631 = n4630 ^ n4302 ^ n1639 ;
  assign n4626 = n2110 ^ n1041 ^ n879 ;
  assign n4624 = n4016 ^ n2727 ^ n607 ;
  assign n4623 = ( ~x104 & n2076 ) | ( ~x104 & n2703 ) | ( n2076 & n2703 ) ;
  assign n4625 = n4624 ^ n4623 ^ n2769 ;
  assign n4617 = n2382 ^ n1849 ^ n655 ;
  assign n4616 = n131 & ~n405 ;
  assign n4618 = n4617 ^ n4616 ^ 1'b0 ;
  assign n4619 = n4618 ^ n1123 ^ n265 ;
  assign n4620 = n3094 ^ n1907 ^ n1700 ;
  assign n4621 = n4620 ^ n4619 ^ n734 ;
  assign n4622 = ( ~n2677 & n4619 ) | ( ~n2677 & n4621 ) | ( n4619 & n4621 ) ;
  assign n4627 = n4626 ^ n4625 ^ n4622 ;
  assign n4632 = n4631 ^ n4627 ^ n602 ;
  assign n4637 = n3427 ^ n2804 ^ n1774 ;
  assign n4638 = n2456 ^ n2117 ^ n595 ;
  assign n4639 = ~x99 & n4638 ;
  assign n4640 = n4639 ^ n2434 ^ n651 ;
  assign n4641 = n4637 & ~n4640 ;
  assign n4635 = ( n1174 & n2047 ) | ( n1174 & ~n2115 ) | ( n2047 & ~n2115 ) ;
  assign n4633 = x123 & ~n737 ;
  assign n4634 = ( n448 & n1825 ) | ( n448 & n4633 ) | ( n1825 & n4633 ) ;
  assign n4636 = n4635 ^ n4634 ^ n4500 ;
  assign n4642 = n4641 ^ n4636 ^ n3481 ;
  assign n4643 = n1890 & ~n1982 ;
  assign n4644 = ( n422 & ~n1474 ) | ( n422 & n2279 ) | ( ~n1474 & n2279 ) ;
  assign n4645 = ( x18 & n1362 ) | ( x18 & n3403 ) | ( n1362 & n3403 ) ;
  assign n4646 = ( n1315 & n4644 ) | ( n1315 & ~n4645 ) | ( n4644 & ~n4645 ) ;
  assign n4647 = n4646 ^ n3493 ^ n2023 ;
  assign n4648 = ( n4294 & ~n4643 ) | ( n4294 & n4647 ) | ( ~n4643 & n4647 ) ;
  assign n4649 = ( ~n1544 & n2116 ) | ( ~n1544 & n2408 ) | ( n2116 & n2408 ) ;
  assign n4650 = n4649 ^ n1967 ^ n1929 ;
  assign n4651 = ( ~n1304 & n1963 ) | ( ~n1304 & n3928 ) | ( n1963 & n3928 ) ;
  assign n4652 = ( n1269 & ~n4650 ) | ( n1269 & n4651 ) | ( ~n4650 & n4651 ) ;
  assign n4674 = n2604 ^ n2239 ^ n1654 ;
  assign n4666 = n1077 ^ n997 ^ n623 ;
  assign n4659 = n256 & ~n3504 ;
  assign n4660 = n966 & n4659 ;
  assign n4661 = n4660 ^ n2212 ^ n474 ;
  assign n4662 = n4661 ^ n2872 ^ 1'b0 ;
  assign n4663 = n224 | n4662 ;
  assign n4664 = n897 | n4663 ;
  assign n4665 = n4664 ^ n1230 ^ 1'b0 ;
  assign n4667 = n4666 ^ n4665 ^ n1028 ;
  assign n4668 = ( n1512 & n1594 ) | ( n1512 & n3163 ) | ( n1594 & n3163 ) ;
  assign n4669 = n4668 ^ n2881 ^ n307 ;
  assign n4670 = ( ~n2912 & n3749 ) | ( ~n2912 & n4669 ) | ( n3749 & n4669 ) ;
  assign n4671 = n3866 | n4670 ;
  assign n4672 = n1588 | n4671 ;
  assign n4673 = ( x49 & n4667 ) | ( x49 & ~n4672 ) | ( n4667 & ~n4672 ) ;
  assign n4657 = n1205 ^ n197 ^ x115 ;
  assign n4655 = ( n1653 & ~n1930 ) | ( n1653 & n2052 ) | ( ~n1930 & n2052 ) ;
  assign n4656 = n4655 ^ n1986 ^ n147 ;
  assign n4653 = n1182 & ~n2121 ;
  assign n4654 = n3638 & n4653 ;
  assign n4658 = n4657 ^ n4656 ^ n4654 ;
  assign n4675 = n4674 ^ n4673 ^ n4658 ;
  assign n4676 = n2447 ^ n291 ^ x70 ;
  assign n4677 = n4676 ^ n2391 ^ n1237 ;
  assign n4678 = ( ~n2368 & n3439 ) | ( ~n2368 & n3636 ) | ( n3439 & n3636 ) ;
  assign n4679 = ( n1985 & ~n4127 ) | ( n1985 & n4678 ) | ( ~n4127 & n4678 ) ;
  assign n4680 = ( n2474 & ~n4183 ) | ( n2474 & n4679 ) | ( ~n4183 & n4679 ) ;
  assign n4681 = n4680 ^ n2935 ^ 1'b0 ;
  assign n4682 = n2181 ^ n1174 ^ n914 ;
  assign n4683 = n4682 ^ n4196 ^ n4178 ;
  assign n4684 = ( n958 & n1278 ) | ( n958 & ~n4683 ) | ( n1278 & ~n4683 ) ;
  assign n4685 = n2925 ^ n2735 ^ 1'b0 ;
  assign n4686 = ( n1417 & n4682 ) | ( n1417 & n4685 ) | ( n4682 & n4685 ) ;
  assign n4687 = ( n781 & n963 ) | ( n781 & ~n4686 ) | ( n963 & ~n4686 ) ;
  assign n4688 = ( ~n474 & n4684 ) | ( ~n474 & n4687 ) | ( n4684 & n4687 ) ;
  assign n4689 = n3517 & n3703 ;
  assign n4690 = ~n3080 & n4689 ;
  assign n4691 = n3319 ^ x70 ^ 1'b0 ;
  assign n4692 = n1651 & n4691 ;
  assign n4693 = ( n3243 & n4690 ) | ( n3243 & n4692 ) | ( n4690 & n4692 ) ;
  assign n4694 = ( ~n1951 & n4688 ) | ( ~n1951 & n4693 ) | ( n4688 & n4693 ) ;
  assign n4695 = ( n1753 & n2211 ) | ( n1753 & n2723 ) | ( n2211 & n2723 ) ;
  assign n4696 = ( x102 & n442 ) | ( x102 & ~n3372 ) | ( n442 & ~n3372 ) ;
  assign n4697 = n3287 ^ n1784 ^ 1'b0 ;
  assign n4698 = ( n2135 & n4696 ) | ( n2135 & n4697 ) | ( n4696 & n4697 ) ;
  assign n4699 = n4249 | n4698 ;
  assign n4700 = n4695 | n4699 ;
  assign n4709 = n2377 ^ n812 ^ 1'b0 ;
  assign n4701 = n635 & n1339 ;
  assign n4702 = n4701 ^ n2236 ^ n270 ;
  assign n4703 = n4702 ^ n2198 ^ 1'b0 ;
  assign n4704 = n2853 ^ n352 ^ 1'b0 ;
  assign n4705 = n609 & ~n2873 ;
  assign n4706 = n4705 ^ n4180 ^ 1'b0 ;
  assign n4707 = ( n1210 & n3188 ) | ( n1210 & ~n4706 ) | ( n3188 & ~n4706 ) ;
  assign n4708 = ( n4703 & n4704 ) | ( n4703 & n4707 ) | ( n4704 & n4707 ) ;
  assign n4710 = n4709 ^ n4708 ^ n3175 ;
  assign n4711 = n1476 ^ n1393 ^ n130 ;
  assign n4712 = n689 & ~n4711 ;
  assign n4713 = n623 | n3133 ;
  assign n4714 = ( n1895 & n2181 ) | ( n1895 & ~n4713 ) | ( n2181 & ~n4713 ) ;
  assign n4715 = ( n1223 & n3726 ) | ( n1223 & n4714 ) | ( n3726 & n4714 ) ;
  assign n4724 = ( ~n1705 & n2503 ) | ( ~n1705 & n3784 ) | ( n2503 & n3784 ) ;
  assign n4725 = ( n2553 & n4409 ) | ( n2553 & n4724 ) | ( n4409 & n4724 ) ;
  assign n4721 = ( n313 & n1211 ) | ( n313 & ~n2839 ) | ( n1211 & ~n2839 ) ;
  assign n4722 = ( n646 & n1173 ) | ( n646 & n4721 ) | ( n1173 & n4721 ) ;
  assign n4723 = n2013 & n4722 ;
  assign n4717 = n4001 ^ n3026 ^ n2834 ;
  assign n4716 = n379 | n2370 ;
  assign n4718 = n4717 ^ n4716 ^ 1'b0 ;
  assign n4719 = n4718 ^ n719 ^ 1'b0 ;
  assign n4720 = ~n2695 & n4719 ;
  assign n4726 = n4725 ^ n4723 ^ n4720 ;
  assign n4727 = n1345 & n1619 ;
  assign n4728 = n4727 ^ n1585 ^ n196 ;
  assign n4729 = n1667 | n3939 ;
  assign n4730 = n4728 & ~n4729 ;
  assign n4731 = ( n4093 & ~n4520 ) | ( n4093 & n4730 ) | ( ~n4520 & n4730 ) ;
  assign n4732 = ( ~n1912 & n4145 ) | ( ~n1912 & n4515 ) | ( n4145 & n4515 ) ;
  assign n4733 = ( x30 & ~n804 ) | ( x30 & n2052 ) | ( ~n804 & n2052 ) ;
  assign n4734 = n4478 ^ n3744 ^ 1'b0 ;
  assign n4735 = n1230 | n4734 ;
  assign n4736 = ( n3452 & n4733 ) | ( n3452 & n4735 ) | ( n4733 & n4735 ) ;
  assign n4737 = n3824 ^ n1352 ^ n319 ;
  assign n4751 = n2581 ^ n1990 ^ n978 ;
  assign n4748 = n2383 ^ n385 ^ 1'b0 ;
  assign n4749 = n2000 & ~n4748 ;
  assign n4750 = n4749 ^ n2862 ^ 1'b0 ;
  assign n4745 = n4394 ^ n1968 ^ n1804 ;
  assign n4746 = n4745 ^ n3819 ^ 1'b0 ;
  assign n4738 = ( ~n197 & n523 ) | ( ~n197 & n1140 ) | ( n523 & n1140 ) ;
  assign n4739 = n1593 ^ n929 ^ 1'b0 ;
  assign n4740 = n4739 ^ n2553 ^ 1'b0 ;
  assign n4741 = n2539 & n4740 ;
  assign n4742 = ( n3351 & ~n4738 ) | ( n3351 & n4741 ) | ( ~n4738 & n4741 ) ;
  assign n4743 = n2122 & n4742 ;
  assign n4744 = n4743 ^ n1732 ^ 1'b0 ;
  assign n4747 = n4746 ^ n4744 ^ n292 ;
  assign n4752 = n4751 ^ n4750 ^ n4747 ;
  assign n4756 = n304 & n455 ;
  assign n4753 = n751 & n784 ;
  assign n4754 = ~n1208 & n4753 ;
  assign n4755 = n4754 ^ n2878 ^ n1788 ;
  assign n4757 = n4756 ^ n4755 ^ n1943 ;
  assign n4758 = ( n3175 & ~n4701 ) | ( n3175 & n4757 ) | ( ~n4701 & n4757 ) ;
  assign n4761 = n2410 ^ n2337 ^ n2139 ;
  assign n4759 = ( ~n290 & n742 ) | ( ~n290 & n2889 ) | ( n742 & n2889 ) ;
  assign n4760 = ( ~n521 & n2703 ) | ( ~n521 & n4759 ) | ( n2703 & n4759 ) ;
  assign n4762 = n4761 ^ n4760 ^ n487 ;
  assign n4763 = n4762 ^ n1399 ^ 1'b0 ;
  assign n4764 = n2409 ^ n2093 ^ n523 ;
  assign n4765 = n4764 ^ n3839 ^ n3069 ;
  assign n4770 = n2207 ^ n1048 ^ n984 ;
  assign n4769 = n3112 ^ n2286 ^ n151 ;
  assign n4771 = n4770 ^ n4769 ^ n840 ;
  assign n4766 = n1571 ^ n950 ^ x63 ;
  assign n4767 = ( x112 & n2023 ) | ( x112 & n4766 ) | ( n2023 & n4766 ) ;
  assign n4768 = ( n1444 & n3378 ) | ( n1444 & n4767 ) | ( n3378 & n4767 ) ;
  assign n4772 = n4771 ^ n4768 ^ n3562 ;
  assign n4773 = n2334 ^ n1645 ^ n223 ;
  assign n4775 = ( n183 & n204 ) | ( n183 & n691 ) | ( n204 & n691 ) ;
  assign n4774 = ( ~n273 & n1997 ) | ( ~n273 & n2149 ) | ( n1997 & n2149 ) ;
  assign n4776 = n4775 ^ n4774 ^ n1795 ;
  assign n4777 = n4490 ^ n3049 ^ 1'b0 ;
  assign n4778 = n4776 & n4777 ;
  assign n4779 = ( n1692 & n2217 ) | ( n1692 & ~n4141 ) | ( n2217 & ~n4141 ) ;
  assign n4780 = n1238 ^ n994 ^ 1'b0 ;
  assign n4781 = ( n2273 & n4779 ) | ( n2273 & n4780 ) | ( n4779 & n4780 ) ;
  assign n4783 = ~n1326 & n1963 ;
  assign n4782 = n1983 ^ n1545 ^ n1242 ;
  assign n4784 = n4783 ^ n4782 ^ 1'b0 ;
  assign n4785 = ~n4781 & n4784 ;
  assign n4786 = ( ~n4365 & n4778 ) | ( ~n4365 & n4785 ) | ( n4778 & n4785 ) ;
  assign n4787 = n2466 ^ n1530 ^ 1'b0 ;
  assign n4788 = n4787 ^ n4384 ^ n1584 ;
  assign n4789 = n2649 ^ n1098 ^ 1'b0 ;
  assign n4790 = n3843 ^ n2272 ^ n1685 ;
  assign n4791 = ( ~n4561 & n4789 ) | ( ~n4561 & n4790 ) | ( n4789 & n4790 ) ;
  assign n4792 = n1993 ^ n1233 ^ 1'b0 ;
  assign n4793 = n1756 ^ n985 ^ 1'b0 ;
  assign n4794 = ( x23 & ~n1797 ) | ( x23 & n4302 ) | ( ~n1797 & n4302 ) ;
  assign n4796 = ( n936 & ~n1768 ) | ( n936 & n2597 ) | ( ~n1768 & n2597 ) ;
  assign n4795 = ( ~n1347 & n1599 ) | ( ~n1347 & n2275 ) | ( n1599 & n2275 ) ;
  assign n4797 = n4796 ^ n4795 ^ n1479 ;
  assign n4798 = n2077 ^ n1634 ^ n452 ;
  assign n4799 = ( n737 & ~n767 ) | ( n737 & n4798 ) | ( ~n767 & n4798 ) ;
  assign n4800 = ( ~n4794 & n4797 ) | ( ~n4794 & n4799 ) | ( n4797 & n4799 ) ;
  assign n4801 = ( ~n474 & n1265 ) | ( ~n474 & n1333 ) | ( n1265 & n1333 ) ;
  assign n4802 = n4801 ^ n1381 ^ n1036 ;
  assign n4803 = n4802 ^ x25 ^ 1'b0 ;
  assign n4804 = ~n2248 & n4803 ;
  assign n4805 = ( n4793 & n4800 ) | ( n4793 & n4804 ) | ( n4800 & n4804 ) ;
  assign n4806 = ( n2129 & ~n3392 ) | ( n2129 & n3502 ) | ( ~n3392 & n3502 ) ;
  assign n4815 = n4319 ^ n799 ^ 1'b0 ;
  assign n4816 = ~n387 & n4815 ;
  assign n4811 = ( ~x105 & n233 ) | ( ~x105 & n1549 ) | ( n233 & n1549 ) ;
  assign n4812 = n4811 ^ n2118 ^ n720 ;
  assign n4813 = n4676 & n4812 ;
  assign n4814 = n4813 ^ n4269 ^ 1'b0 ;
  assign n4807 = n1140 ^ n207 ^ 1'b0 ;
  assign n4808 = n4807 ^ n4160 ^ n1635 ;
  assign n4809 = ( n1477 & ~n1609 ) | ( n1477 & n2776 ) | ( ~n1609 & n2776 ) ;
  assign n4810 = ( ~n2924 & n4808 ) | ( ~n2924 & n4809 ) | ( n4808 & n4809 ) ;
  assign n4817 = n4816 ^ n4814 ^ n4810 ;
  assign n4818 = ( n390 & n2440 ) | ( n390 & n4817 ) | ( n2440 & n4817 ) ;
  assign n4819 = n3878 & ~n4818 ;
  assign n4825 = n4569 ^ n4518 ^ n1213 ;
  assign n4821 = x97 & ~n1964 ;
  assign n4822 = n4821 ^ n1263 ^ 1'b0 ;
  assign n4823 = ~n1506 & n3510 ;
  assign n4824 = n4822 & n4823 ;
  assign n4820 = ( n454 & n1658 ) | ( n454 & n3088 ) | ( n1658 & n3088 ) ;
  assign n4826 = n4825 ^ n4824 ^ n4820 ;
  assign n4827 = n3369 ^ n2474 ^ n2044 ;
  assign n4828 = n4827 ^ n1603 ^ n203 ;
  assign n4829 = n260 ^ n203 ^ 1'b0 ;
  assign n4830 = n4829 ^ n3777 ^ n2113 ;
  assign n4831 = n2957 ^ n442 ^ 1'b0 ;
  assign n4832 = n4830 | n4831 ;
  assign n4848 = n4110 ^ n1561 ^ x89 ;
  assign n4837 = n2265 ^ n921 ^ 1'b0 ;
  assign n4838 = n1659 & n4837 ;
  assign n4839 = ( ~n2931 & n4569 ) | ( ~n2931 & n4838 ) | ( n4569 & n4838 ) ;
  assign n4841 = ( n187 & ~n893 ) | ( n187 & n1056 ) | ( ~n893 & n1056 ) ;
  assign n4842 = n4841 ^ n876 ^ n200 ;
  assign n4840 = n4219 ^ n2475 ^ n2106 ;
  assign n4843 = n4842 ^ n4840 ^ n462 ;
  assign n4844 = n4843 ^ n1520 ^ n233 ;
  assign n4845 = n4844 ^ n3277 ^ 1'b0 ;
  assign n4846 = n4839 & n4845 ;
  assign n4834 = ( n257 & ~n2065 ) | ( n257 & n3079 ) | ( ~n2065 & n3079 ) ;
  assign n4835 = ( n214 & n854 ) | ( n214 & ~n4834 ) | ( n854 & ~n4834 ) ;
  assign n4833 = n4607 ^ n2283 ^ n2144 ;
  assign n4836 = n4835 ^ n4833 ^ n2645 ;
  assign n4847 = n4846 ^ n4836 ^ n2427 ;
  assign n4849 = n4848 ^ n4847 ^ n1615 ;
  assign n4850 = ( x20 & ~n242 ) | ( x20 & n2977 ) | ( ~n242 & n2977 ) ;
  assign n4851 = n4850 ^ n993 ^ n816 ;
  assign n4852 = ( n3747 & n3782 ) | ( n3747 & ~n4851 ) | ( n3782 & ~n4851 ) ;
  assign n4853 = n3945 ^ n1980 ^ n651 ;
  assign n4854 = ( n3956 & n4852 ) | ( n3956 & n4853 ) | ( n4852 & n4853 ) ;
  assign n4856 = ( n297 & n2656 ) | ( n297 & ~n4129 ) | ( n2656 & ~n4129 ) ;
  assign n4855 = ( ~n246 & n344 ) | ( ~n246 & n3925 ) | ( n344 & n3925 ) ;
  assign n4857 = n4856 ^ n4855 ^ n1587 ;
  assign n4860 = n3366 ^ n2473 ^ n1629 ;
  assign n4861 = n4860 ^ n4704 ^ n1085 ;
  assign n4858 = ( ~n1583 & n2326 ) | ( ~n1583 & n3048 ) | ( n2326 & n3048 ) ;
  assign n4859 = ( n2719 & ~n3866 ) | ( n2719 & n4858 ) | ( ~n3866 & n4858 ) ;
  assign n4862 = n4861 ^ n4859 ^ n1569 ;
  assign n4867 = n1706 ^ n449 ^ 1'b0 ;
  assign n4868 = ( n423 & ~n1629 ) | ( n423 & n4867 ) | ( ~n1629 & n4867 ) ;
  assign n4865 = ( n1491 & n2306 ) | ( n1491 & ~n4289 ) | ( n2306 & ~n4289 ) ;
  assign n4866 = n4865 ^ n1008 ^ n173 ;
  assign n4869 = n4868 ^ n4866 ^ 1'b0 ;
  assign n4863 = n3509 ^ n574 ^ n184 ;
  assign n4864 = n4863 ^ n2171 ^ n2000 ;
  assign n4870 = n4869 ^ n4864 ^ n4816 ;
  assign n4871 = ( n151 & n603 ) | ( n151 & n4288 ) | ( n603 & n4288 ) ;
  assign n4872 = n3948 ^ n3372 ^ 1'b0 ;
  assign n4873 = ~n1238 & n2810 ;
  assign n4874 = n1391 & n4873 ;
  assign n4875 = ( n135 & n2230 ) | ( n135 & n4874 ) | ( n2230 & n4874 ) ;
  assign n4876 = ( n500 & n639 ) | ( n500 & n2286 ) | ( n639 & n2286 ) ;
  assign n4877 = n4876 ^ n4416 ^ n2218 ;
  assign n4878 = ( n391 & ~n1578 ) | ( n391 & n4877 ) | ( ~n1578 & n4877 ) ;
  assign n4879 = ( ~n4872 & n4875 ) | ( ~n4872 & n4878 ) | ( n4875 & n4878 ) ;
  assign n4880 = ( n3516 & ~n4871 ) | ( n3516 & n4879 ) | ( ~n4871 & n4879 ) ;
  assign n4881 = ( n953 & n1831 ) | ( n953 & n4880 ) | ( n1831 & n4880 ) ;
  assign n4891 = n3238 ^ n1715 ^ n280 ;
  assign n4892 = ( n2367 & ~n2677 ) | ( n2367 & n4891 ) | ( ~n2677 & n4891 ) ;
  assign n4888 = n1140 ^ n288 ^ x122 ;
  assign n4882 = n2483 ^ n2304 ^ n704 ;
  assign n4883 = ( n762 & ~n1022 ) | ( n762 & n1363 ) | ( ~n1022 & n1363 ) ;
  assign n4884 = n2442 ^ n380 ^ n290 ;
  assign n4885 = n1588 & n4884 ;
  assign n4886 = ~x86 & n4885 ;
  assign n4887 = ( ~n4882 & n4883 ) | ( ~n4882 & n4886 ) | ( n4883 & n4886 ) ;
  assign n4889 = n4888 ^ n4887 ^ 1'b0 ;
  assign n4890 = n829 & n4889 ;
  assign n4893 = n4892 ^ n4890 ^ n2233 ;
  assign n4894 = n1629 & n3731 ;
  assign n4895 = n4894 ^ n668 ^ n644 ;
  assign n4896 = ( ~n1442 & n2993 ) | ( ~n1442 & n4895 ) | ( n2993 & n4895 ) ;
  assign n4897 = ( x47 & ~n881 ) | ( x47 & n1201 ) | ( ~n881 & n1201 ) ;
  assign n4898 = n4897 ^ n2700 ^ n2490 ;
  assign n4899 = n4898 ^ n845 ^ 1'b0 ;
  assign n4900 = n4899 ^ n668 ^ 1'b0 ;
  assign n4901 = ~n1245 & n4900 ;
  assign n4902 = ( n2573 & n4896 ) | ( n2573 & n4901 ) | ( n4896 & n4901 ) ;
  assign n4903 = n2706 ^ n915 ^ 1'b0 ;
  assign n4904 = ~n2748 & n4903 ;
  assign n4905 = ( n406 & n2342 ) | ( n406 & n4904 ) | ( n2342 & n4904 ) ;
  assign n4906 = ( x28 & ~n732 ) | ( x28 & n1993 ) | ( ~n732 & n1993 ) ;
  assign n4907 = n3748 ^ n905 ^ x120 ;
  assign n4908 = ( ~n1015 & n1173 ) | ( ~n1015 & n4907 ) | ( n1173 & n4907 ) ;
  assign n4909 = n2369 ^ n744 ^ 1'b0 ;
  assign n4910 = n4908 & ~n4909 ;
  assign n4911 = n4906 & n4910 ;
  assign n4912 = ~n1104 & n4911 ;
  assign n4913 = ( n1247 & ~n4905 ) | ( n1247 & n4912 ) | ( ~n4905 & n4912 ) ;
  assign n4915 = n1993 & n2610 ;
  assign n4916 = ~n1647 & n4915 ;
  assign n4914 = ( ~n2193 & n4220 ) | ( ~n2193 & n4839 ) | ( n4220 & n4839 ) ;
  assign n4917 = n4916 ^ n4914 ^ 1'b0 ;
  assign n4918 = ~n4913 & n4917 ;
  assign n4925 = n2172 ^ n1068 ^ n934 ;
  assign n4923 = n3442 ^ n2523 ^ 1'b0 ;
  assign n4924 = n1057 | n4923 ;
  assign n4919 = ~n1405 & n2075 ;
  assign n4920 = ( n1262 & n2117 ) | ( n1262 & ~n3112 ) | ( n2117 & ~n3112 ) ;
  assign n4921 = n4920 ^ n3669 ^ 1'b0 ;
  assign n4922 = n4919 | n4921 ;
  assign n4926 = n4925 ^ n4924 ^ n4922 ;
  assign n4927 = n1517 ^ n711 ^ 1'b0 ;
  assign n4928 = n4287 | n4927 ;
  assign n4934 = n4306 ^ n909 ^ 1'b0 ;
  assign n4929 = ~n3272 & n3721 ;
  assign n4930 = n4303 ^ n1353 ^ n165 ;
  assign n4931 = n4930 ^ n3689 ^ n3513 ;
  assign n4932 = ( n3865 & n4929 ) | ( n3865 & n4931 ) | ( n4929 & n4931 ) ;
  assign n4933 = n4932 ^ n3328 ^ n1112 ;
  assign n4935 = n4934 ^ n4933 ^ n2569 ;
  assign n4939 = n2678 ^ n1249 ^ n1121 ;
  assign n4940 = ( n1743 & n1781 ) | ( n1743 & n4939 ) | ( n1781 & n4939 ) ;
  assign n4936 = ( n685 & n1802 ) | ( n685 & n2819 ) | ( n1802 & n2819 ) ;
  assign n4937 = ( n1762 & n1781 ) | ( n1762 & ~n4936 ) | ( n1781 & ~n4936 ) ;
  assign n4938 = n3518 & ~n4937 ;
  assign n4941 = n4940 ^ n4938 ^ 1'b0 ;
  assign n4945 = ~n1558 & n2429 ;
  assign n4943 = n2348 ^ n1405 ^ n500 ;
  assign n4942 = n2178 ^ n1253 ^ 1'b0 ;
  assign n4944 = n4943 ^ n4942 ^ n1103 ;
  assign n4946 = n4945 ^ n4944 ^ n2401 ;
  assign n4969 = ~n4381 & n4738 ;
  assign n4970 = ( n1173 & ~n4099 ) | ( n1173 & n4969 ) | ( ~n4099 & n4969 ) ;
  assign n4958 = ( ~n843 & n1572 ) | ( ~n843 & n2040 ) | ( n1572 & n2040 ) ;
  assign n4961 = n438 & n990 ;
  assign n4962 = n4961 ^ n1600 ^ n896 ;
  assign n4959 = n4422 ^ n3182 ^ n2116 ;
  assign n4960 = ( n1490 & n2542 ) | ( n1490 & ~n4959 ) | ( n2542 & ~n4959 ) ;
  assign n4963 = n4962 ^ n4960 ^ 1'b0 ;
  assign n4964 = ( ~n2679 & n4958 ) | ( ~n2679 & n4963 ) | ( n4958 & n4963 ) ;
  assign n4947 = ( n726 & ~n1343 ) | ( n726 & n2365 ) | ( ~n1343 & n2365 ) ;
  assign n4948 = n4947 ^ n2429 ^ n2035 ;
  assign n4954 = ( n470 & n1397 ) | ( n470 & n1422 ) | ( n1397 & n1422 ) ;
  assign n4949 = ( n379 & ~n399 ) | ( n379 & n1110 ) | ( ~n399 & n1110 ) ;
  assign n4950 = x71 & n467 ;
  assign n4951 = n4950 ^ n272 ^ 1'b0 ;
  assign n4952 = n4951 ^ n4718 ^ 1'b0 ;
  assign n4953 = ~n4949 & n4952 ;
  assign n4955 = n4954 ^ n4953 ^ n4195 ;
  assign n4956 = ( n1301 & n2385 ) | ( n1301 & ~n4955 ) | ( n2385 & ~n4955 ) ;
  assign n4957 = n4948 & ~n4956 ;
  assign n4965 = n4964 ^ n4957 ^ 1'b0 ;
  assign n4966 = n3975 ^ n1955 ^ n342 ;
  assign n4967 = n4966 ^ n2471 ^ n2358 ;
  assign n4968 = n4965 & n4967 ;
  assign n4971 = n4970 ^ n4968 ^ 1'b0 ;
  assign n4972 = n1240 ^ n656 ^ n164 ;
  assign n4973 = ( n3274 & ~n3449 ) | ( n3274 & n4972 ) | ( ~n3449 & n4972 ) ;
  assign n4974 = n1205 & n2334 ;
  assign n4975 = ( n307 & ~n2191 ) | ( n307 & n4974 ) | ( ~n2191 & n4974 ) ;
  assign n4976 = n4975 ^ n2048 ^ 1'b0 ;
  assign n4977 = ( n750 & n1433 ) | ( n750 & n3289 ) | ( n1433 & n3289 ) ;
  assign n4979 = n2581 ^ n2013 ^ n252 ;
  assign n4978 = n4660 ^ n3184 ^ n2728 ;
  assign n4980 = n4979 ^ n4978 ^ n2139 ;
  assign n4981 = ~n4977 & n4980 ;
  assign n4982 = ( n872 & ~n3247 ) | ( n872 & n4091 ) | ( ~n3247 & n4091 ) ;
  assign n4983 = n343 ^ x108 ^ x42 ;
  assign n4984 = ( n2150 & ~n3677 ) | ( n2150 & n4983 ) | ( ~n3677 & n4983 ) ;
  assign n4985 = n4984 ^ n1806 ^ 1'b0 ;
  assign n4986 = n3413 ^ n359 ^ 1'b0 ;
  assign n4987 = ~n4368 & n4986 ;
  assign n4988 = n4071 & n4987 ;
  assign n4989 = n4988 ^ n1615 ^ 1'b0 ;
  assign n4990 = n4725 ^ n1544 ^ n536 ;
  assign n4991 = n4990 ^ n3680 ^ n640 ;
  assign n4996 = n3810 ^ n449 ^ n256 ;
  assign n4997 = ( n739 & n1442 ) | ( n739 & n4996 ) | ( n1442 & n4996 ) ;
  assign n4995 = ( n938 & n4339 ) | ( n938 & ~n4539 ) | ( n4339 & ~n4539 ) ;
  assign n4992 = n1201 ^ n1083 ^ x16 ;
  assign n4993 = n4992 ^ n1316 ^ n665 ;
  assign n4994 = n4993 ^ n4482 ^ n2277 ;
  assign n4998 = n4997 ^ n4995 ^ n4994 ;
  assign n4999 = ( ~n716 & n1215 ) | ( ~n716 & n4998 ) | ( n1215 & n4998 ) ;
  assign n5000 = ( n977 & ~n3055 ) | ( n977 & n3803 ) | ( ~n3055 & n3803 ) ;
  assign n5001 = n3571 ^ n2670 ^ 1'b0 ;
  assign n5002 = n4278 & n5001 ;
  assign n5003 = n700 ^ n439 ^ x110 ;
  assign n5004 = n5003 ^ n1551 ^ n778 ;
  assign n5005 = ( ~n2336 & n4830 ) | ( ~n2336 & n5004 ) | ( n4830 & n5004 ) ;
  assign n5007 = ( n187 & n1178 ) | ( n187 & n2705 ) | ( n1178 & n2705 ) ;
  assign n5008 = ( n2216 & ~n2562 ) | ( n2216 & n5007 ) | ( ~n2562 & n5007 ) ;
  assign n5009 = ( n3312 & ~n4183 ) | ( n3312 & n5008 ) | ( ~n4183 & n5008 ) ;
  assign n5006 = ( x80 & ~n2288 ) | ( x80 & n3396 ) | ( ~n2288 & n3396 ) ;
  assign n5010 = n5009 ^ n5006 ^ x81 ;
  assign n5011 = n1371 ^ n1140 ^ n355 ;
  assign n5012 = ( n1923 & n4262 ) | ( n1923 & n5011 ) | ( n4262 & n5011 ) ;
  assign n5013 = ( ~n5005 & n5010 ) | ( ~n5005 & n5012 ) | ( n5010 & n5012 ) ;
  assign n5024 = n2574 ^ n1176 ^ x109 ;
  assign n5020 = n1990 ^ n1601 ^ 1'b0 ;
  assign n5021 = ( n1865 & ~n2587 ) | ( n1865 & n5020 ) | ( ~n2587 & n5020 ) ;
  assign n5022 = ( n1267 & n2064 ) | ( n1267 & n5021 ) | ( n2064 & n5021 ) ;
  assign n5023 = ( n1441 & n4920 ) | ( n1441 & n5022 ) | ( n4920 & n5022 ) ;
  assign n5014 = ( n930 & n1842 ) | ( n930 & n2278 ) | ( n1842 & n2278 ) ;
  assign n5015 = n1968 ^ x119 ^ x15 ;
  assign n5016 = n5015 ^ n3000 ^ n1788 ;
  assign n5017 = ( n1320 & n2267 ) | ( n1320 & n5016 ) | ( n2267 & n5016 ) ;
  assign n5018 = n229 & ~n1949 ;
  assign n5019 = ( n5014 & n5017 ) | ( n5014 & ~n5018 ) | ( n5017 & ~n5018 ) ;
  assign n5025 = n5024 ^ n5023 ^ n5019 ;
  assign n5026 = ( n458 & n1895 ) | ( n458 & n4904 ) | ( n1895 & n4904 ) ;
  assign n5027 = n3803 ^ n782 ^ n421 ;
  assign n5028 = n4551 ^ n203 ^ 1'b0 ;
  assign n5029 = n5027 | n5028 ;
  assign n5030 = n5026 | n5029 ;
  assign n5031 = n5030 ^ n1333 ^ 1'b0 ;
  assign n5032 = ( n154 & n311 ) | ( n154 & n1395 ) | ( n311 & n1395 ) ;
  assign n5033 = ( ~n163 & n629 ) | ( ~n163 & n2183 ) | ( n629 & n2183 ) ;
  assign n5034 = n5033 ^ n2960 ^ n942 ;
  assign n5035 = ~n5032 & n5034 ;
  assign n5048 = n720 & n2877 ;
  assign n5049 = n431 & n5048 ;
  assign n5045 = n1594 & n2976 ;
  assign n5046 = n5045 ^ n1049 ^ 1'b0 ;
  assign n5047 = n5046 ^ n2115 ^ n967 ;
  assign n5041 = n1027 ^ n787 ^ n286 ;
  assign n5040 = ( n1146 & ~n1161 ) | ( n1146 & n1333 ) | ( ~n1161 & n1333 ) ;
  assign n5042 = n5041 ^ n5040 ^ n803 ;
  assign n5039 = n4259 ^ n2981 ^ 1'b0 ;
  assign n5036 = ( n384 & ~n768 ) | ( n384 & n4380 ) | ( ~n768 & n4380 ) ;
  assign n5037 = ( n394 & n4386 ) | ( n394 & ~n5036 ) | ( n4386 & ~n5036 ) ;
  assign n5038 = ( n584 & n1342 ) | ( n584 & ~n5037 ) | ( n1342 & ~n5037 ) ;
  assign n5043 = n5042 ^ n5039 ^ n5038 ;
  assign n5044 = n5043 ^ n3494 ^ n207 ;
  assign n5050 = n5049 ^ n5047 ^ n5044 ;
  assign n5051 = n3621 ^ n3187 ^ n351 ;
  assign n5052 = ( n450 & n1151 ) | ( n450 & ~n4234 ) | ( n1151 & ~n4234 ) ;
  assign n5053 = n3113 & n5052 ;
  assign n5054 = ( n2690 & ~n3561 ) | ( n2690 & n5053 ) | ( ~n3561 & n5053 ) ;
  assign n5055 = ( n3059 & ~n5051 ) | ( n3059 & n5054 ) | ( ~n5051 & n5054 ) ;
  assign n5056 = ( n3447 & ~n5050 ) | ( n3447 & n5055 ) | ( ~n5050 & n5055 ) ;
  assign n5057 = n1215 & n5056 ;
  assign n5058 = ~n1110 & n2344 ;
  assign n5062 = n1182 ^ n350 ^ n267 ;
  assign n5063 = n5062 ^ n2973 ^ n1433 ;
  assign n5064 = ( ~n1024 & n3352 ) | ( ~n1024 & n5063 ) | ( n3352 & n5063 ) ;
  assign n5059 = n3114 ^ n1810 ^ n1068 ;
  assign n5060 = n5059 ^ n233 ^ 1'b0 ;
  assign n5061 = ( n2462 & n3471 ) | ( n2462 & ~n5060 ) | ( n3471 & ~n5060 ) ;
  assign n5065 = n5064 ^ n5061 ^ n2343 ;
  assign n5066 = ( n543 & n5058 ) | ( n543 & n5065 ) | ( n5058 & n5065 ) ;
  assign n5067 = ~n4438 & n4724 ;
  assign n5068 = n5067 ^ n4244 ^ n2189 ;
  assign n5069 = n1041 ^ x58 ^ x33 ;
  assign n5070 = n3310 ^ n163 ^ 1'b0 ;
  assign n5071 = ~n1940 & n5070 ;
  assign n5072 = n5071 ^ n1350 ^ 1'b0 ;
  assign n5073 = ( ~n2069 & n5069 ) | ( ~n2069 & n5072 ) | ( n5069 & n5072 ) ;
  assign n5074 = n4329 ^ n1897 ^ n1545 ;
  assign n5084 = ( n607 & n1088 ) | ( n607 & n2460 ) | ( n1088 & n2460 ) ;
  assign n5081 = ( n1384 & ~n2114 ) | ( n1384 & n2286 ) | ( ~n2114 & n2286 ) ;
  assign n5082 = ~n2069 & n5081 ;
  assign n5083 = n5082 ^ n4118 ^ 1'b0 ;
  assign n5079 = n1494 ^ n1446 ^ n1060 ;
  assign n5075 = n504 & n1400 ;
  assign n5076 = ~n889 & n5075 ;
  assign n5077 = n5076 ^ n349 ^ n250 ;
  assign n5078 = n5077 ^ n3136 ^ n2028 ;
  assign n5080 = n5079 ^ n5078 ^ 1'b0 ;
  assign n5085 = n5084 ^ n5083 ^ n5080 ;
  assign n5086 = ~n4372 & n5085 ;
  assign n5087 = ~n5074 & n5086 ;
  assign n5088 = n984 ^ x50 ^ 1'b0 ;
  assign n5089 = ( ~n333 & n1595 ) | ( ~n333 & n5088 ) | ( n1595 & n5088 ) ;
  assign n5090 = n3527 ^ n756 ^ n522 ;
  assign n5095 = n2787 ^ n2038 ^ n848 ;
  assign n5091 = n2723 ^ n580 ^ n535 ;
  assign n5092 = n5091 ^ n3525 ^ n3035 ;
  assign n5093 = n5092 ^ n1969 ^ n1139 ;
  assign n5094 = n2844 | n5093 ;
  assign n5096 = n5095 ^ n5094 ^ 1'b0 ;
  assign n5097 = n5090 | n5096 ;
  assign n5100 = ~n2314 & n2718 ;
  assign n5101 = n5100 ^ n3644 ^ 1'b0 ;
  assign n5102 = n5101 ^ n4709 ^ n3481 ;
  assign n5098 = n1706 ^ n867 ^ n803 ;
  assign n5099 = n5098 ^ n3551 ^ 1'b0 ;
  assign n5103 = n5102 ^ n5099 ^ n1729 ;
  assign n5104 = n5103 ^ n943 ^ n473 ;
  assign n5105 = n1109 ^ n494 ^ n487 ;
  assign n5106 = n5105 ^ n3860 ^ n2855 ;
  assign n5107 = ( n2136 & n3951 ) | ( n2136 & n5106 ) | ( n3951 & n5106 ) ;
  assign n5108 = n4545 ^ n2617 ^ n1309 ;
  assign n5109 = ( x48 & n4882 ) | ( x48 & ~n4993 ) | ( n4882 & ~n4993 ) ;
  assign n5110 = ( n1274 & n2903 ) | ( n1274 & n4558 ) | ( n2903 & n4558 ) ;
  assign n5111 = n2228 ^ n875 ^ n130 ;
  assign n5112 = ( ~n341 & n942 ) | ( ~n341 & n5111 ) | ( n942 & n5111 ) ;
  assign n5113 = n5112 ^ n1858 ^ n657 ;
  assign n5114 = ( n761 & n1247 ) | ( n761 & ~n1400 ) | ( n1247 & ~n1400 ) ;
  assign n5115 = ( ~n1995 & n4309 ) | ( ~n1995 & n5114 ) | ( n4309 & n5114 ) ;
  assign n5116 = ( x8 & n2038 ) | ( x8 & n5115 ) | ( n2038 & n5115 ) ;
  assign n5117 = ( ~n5110 & n5113 ) | ( ~n5110 & n5116 ) | ( n5113 & n5116 ) ;
  assign n5118 = n4665 ^ n1239 ^ 1'b0 ;
  assign n5119 = ( ~n750 & n1575 ) | ( ~n750 & n2397 ) | ( n1575 & n2397 ) ;
  assign n5120 = n5119 ^ n4440 ^ n3729 ;
  assign n5121 = n5120 ^ n4338 ^ n1660 ;
  assign n5122 = n3707 ^ n2287 ^ n268 ;
  assign n5123 = n5121 | n5122 ;
  assign n5130 = n1871 ^ n1433 ^ n819 ;
  assign n5131 = n5130 ^ n2233 ^ n1006 ;
  assign n5132 = n3452 ^ n1086 ^ n172 ;
  assign n5133 = ( n237 & n5131 ) | ( n237 & n5132 ) | ( n5131 & n5132 ) ;
  assign n5134 = ( ~n4844 & n5092 ) | ( ~n4844 & n5133 ) | ( n5092 & n5133 ) ;
  assign n5129 = ( ~n1264 & n1516 ) | ( ~n1264 & n4703 ) | ( n1516 & n4703 ) ;
  assign n5135 = n5134 ^ n5129 ^ n4887 ;
  assign n5124 = ( n1036 & ~n1713 ) | ( n1036 & n2683 ) | ( ~n1713 & n2683 ) ;
  assign n5125 = n2173 ^ n1520 ^ x62 ;
  assign n5126 = ( ~n2079 & n4591 ) | ( ~n2079 & n5125 ) | ( n4591 & n5125 ) ;
  assign n5127 = ( n1330 & n5124 ) | ( n1330 & ~n5126 ) | ( n5124 & ~n5126 ) ;
  assign n5128 = n917 | n5127 ;
  assign n5136 = n5135 ^ n5128 ^ x64 ;
  assign n5137 = n3935 ^ n2027 ^ n1775 ;
  assign n5138 = ( n1643 & ~n2477 ) | ( n1643 & n5137 ) | ( ~n2477 & n5137 ) ;
  assign n5139 = ~n493 & n1997 ;
  assign n5140 = ( ~n4115 & n4505 ) | ( ~n4115 & n5139 ) | ( n4505 & n5139 ) ;
  assign n5141 = ( ~n250 & n5138 ) | ( ~n250 & n5140 ) | ( n5138 & n5140 ) ;
  assign n5145 = n1284 & n2550 ;
  assign n5142 = n2099 ^ n330 ^ 1'b0 ;
  assign n5143 = n5142 ^ n3661 ^ n242 ;
  assign n5144 = n5143 ^ n2640 ^ n2277 ;
  assign n5146 = n5145 ^ n5144 ^ n3412 ;
  assign n5147 = n3953 ^ n2487 ^ n1858 ;
  assign n5148 = ( n1840 & n1857 ) | ( n1840 & ~n5147 ) | ( n1857 & ~n5147 ) ;
  assign n5149 = ( n1169 & n1975 ) | ( n1169 & ~n2779 ) | ( n1975 & ~n2779 ) ;
  assign n5150 = n5149 ^ n1371 ^ n166 ;
  assign n5151 = n633 ^ n296 ^ n280 ;
  assign n5152 = ~n3282 & n5151 ;
  assign n5153 = ~n1949 & n5152 ;
  assign n5154 = n3826 ^ n232 ^ 1'b0 ;
  assign n5155 = ( n5150 & ~n5153 ) | ( n5150 & n5154 ) | ( ~n5153 & n5154 ) ;
  assign n5156 = n1227 & ~n3351 ;
  assign n5157 = ( n2316 & n4440 ) | ( n2316 & n5156 ) | ( n4440 & n5156 ) ;
  assign n5158 = n5157 ^ n848 ^ n405 ;
  assign n5159 = ( ~n375 & n417 ) | ( ~n375 & n4566 ) | ( n417 & n4566 ) ;
  assign n5160 = n5159 ^ n2805 ^ n742 ;
  assign n5161 = n5160 ^ n4082 ^ n3239 ;
  assign n5162 = n5161 ^ n2787 ^ 1'b0 ;
  assign n5163 = n3312 ^ n1407 ^ 1'b0 ;
  assign n5164 = ~n5162 & n5163 ;
  assign n5165 = ( ~n5155 & n5158 ) | ( ~n5155 & n5164 ) | ( n5158 & n5164 ) ;
  assign n5167 = n731 ^ n504 ^ n200 ;
  assign n5168 = n5167 ^ n689 ^ x64 ;
  assign n5166 = n1108 ^ n1008 ^ n346 ;
  assign n5169 = n5168 ^ n5166 ^ n1351 ;
  assign n5170 = n347 & ~n5169 ;
  assign n5171 = n5170 ^ n3614 ^ 1'b0 ;
  assign n5172 = ( n1372 & ~n4795 ) | ( n1372 & n5171 ) | ( ~n4795 & n5171 ) ;
  assign n5173 = ( ~n1804 & n3895 ) | ( ~n1804 & n5172 ) | ( n3895 & n5172 ) ;
  assign n5174 = ( n2542 & ~n2594 ) | ( n2542 & n5173 ) | ( ~n2594 & n5173 ) ;
  assign n5175 = n3453 ^ n2592 ^ n765 ;
  assign n5176 = n5175 ^ n610 ^ 1'b0 ;
  assign n5177 = n5174 & ~n5176 ;
  assign n5178 = n3975 ^ n2705 ^ n1982 ;
  assign n5180 = ( n412 & ~n1393 ) | ( n412 & n4241 ) | ( ~n1393 & n4241 ) ;
  assign n5181 = ~n3860 & n5180 ;
  assign n5182 = n5181 ^ n1784 ^ 1'b0 ;
  assign n5179 = x21 & ~n857 ;
  assign n5183 = n5182 ^ n5179 ^ 1'b0 ;
  assign n5184 = n5178 & n5183 ;
  assign n5185 = ~n5177 & n5184 ;
  assign n5186 = n1997 | n4545 ;
  assign n5187 = n5186 ^ n1586 ^ n442 ;
  assign n5188 = n5187 ^ n2983 ^ 1'b0 ;
  assign n5189 = ( n169 & n924 ) | ( n169 & ~n1077 ) | ( n924 & ~n1077 ) ;
  assign n5190 = n5189 ^ n880 ^ n178 ;
  assign n5191 = n4028 ^ n1211 ^ 1'b0 ;
  assign n5192 = ( n1672 & n5190 ) | ( n1672 & ~n5191 ) | ( n5190 & ~n5191 ) ;
  assign n5193 = ~n168 & n1594 ;
  assign n5194 = n4587 ^ n1555 ^ n1384 ;
  assign n5195 = n5194 ^ n1023 ^ n522 ;
  assign n5197 = n832 ^ x91 ^ 1'b0 ;
  assign n5196 = x42 | n3096 ;
  assign n5198 = n5197 ^ n5196 ^ n960 ;
  assign n5199 = n5195 | n5198 ;
  assign n5203 = n628 & ~n4750 ;
  assign n5204 = n5203 ^ n744 ^ 1'b0 ;
  assign n5200 = n1992 ^ n859 ^ x124 ;
  assign n5201 = ( ~n2712 & n4511 ) | ( ~n2712 & n5200 ) | ( n4511 & n5200 ) ;
  assign n5202 = n5201 ^ n4613 ^ n1055 ;
  assign n5205 = n5204 ^ n5202 ^ 1'b0 ;
  assign n5206 = n4010 ^ n3888 ^ n173 ;
  assign n5207 = n3648 ^ n2433 ^ 1'b0 ;
  assign n5208 = n5207 ^ n953 ^ 1'b0 ;
  assign n5209 = ( ~n142 & n960 ) | ( ~n142 & n1410 ) | ( n960 & n1410 ) ;
  assign n5210 = n1770 ^ n822 ^ n627 ;
  assign n5211 = ( n583 & n995 ) | ( n583 & ~n4044 ) | ( n995 & ~n4044 ) ;
  assign n5212 = n2398 ^ n254 ^ 1'b0 ;
  assign n5213 = n4281 & ~n5212 ;
  assign n5214 = ( ~n5210 & n5211 ) | ( ~n5210 & n5213 ) | ( n5211 & n5213 ) ;
  assign n5215 = ( n917 & ~n5209 ) | ( n917 & n5214 ) | ( ~n5209 & n5214 ) ;
  assign n5216 = ( n163 & ~n5208 ) | ( n163 & n5215 ) | ( ~n5208 & n5215 ) ;
  assign n5217 = n5216 ^ n1752 ^ 1'b0 ;
  assign n5218 = ( ~n3669 & n5206 ) | ( ~n3669 & n5217 ) | ( n5206 & n5217 ) ;
  assign n5225 = ( ~x109 & x121 ) | ( ~x109 & n2466 ) | ( x121 & n2466 ) ;
  assign n5224 = n3443 ^ n2791 ^ n354 ;
  assign n5226 = n5225 ^ n5224 ^ 1'b0 ;
  assign n5227 = ~n1895 & n5226 ;
  assign n5220 = ( n161 & ~n1262 ) | ( n161 & n2569 ) | ( ~n1262 & n2569 ) ;
  assign n5221 = n5220 ^ n1741 ^ 1'b0 ;
  assign n5222 = n152 & n5221 ;
  assign n5223 = n5222 ^ n2963 ^ n2786 ;
  assign n5228 = n5227 ^ n5223 ^ n3116 ;
  assign n5219 = n3815 ^ n2144 ^ n1715 ;
  assign n5229 = n5228 ^ n5219 ^ n1526 ;
  assign n5230 = n2239 ^ n1249 ^ n383 ;
  assign n5231 = n5206 ^ n428 ^ n386 ;
  assign n5232 = ( n1895 & n5230 ) | ( n1895 & n5231 ) | ( n5230 & n5231 ) ;
  assign n5233 = ( x109 & n817 ) | ( x109 & ~n4262 ) | ( n817 & ~n4262 ) ;
  assign n5234 = n5233 ^ n3445 ^ n272 ;
  assign n5235 = n2729 ^ n2164 ^ 1'b0 ;
  assign n5236 = n2017 ^ n1749 ^ 1'b0 ;
  assign n5237 = ( ~n1580 & n3066 ) | ( ~n1580 & n5236 ) | ( n3066 & n5236 ) ;
  assign n5238 = n655 & ~n1403 ;
  assign n5239 = n5238 ^ x17 ^ 1'b0 ;
  assign n5240 = ( n3710 & n4797 ) | ( n3710 & ~n5239 ) | ( n4797 & ~n5239 ) ;
  assign n5241 = ( n340 & n1789 ) | ( n340 & ~n5240 ) | ( n1789 & ~n5240 ) ;
  assign n5242 = n5241 ^ n3712 ^ n433 ;
  assign n5243 = ~n5237 & n5242 ;
  assign n5244 = ~n5235 & n5243 ;
  assign n5245 = n4085 ^ n3895 ^ n3520 ;
  assign n5246 = ( n3637 & ~n4004 ) | ( n3637 & n5245 ) | ( ~n4004 & n5245 ) ;
  assign n5251 = ( n3281 & ~n4850 ) | ( n3281 & n4908 ) | ( ~n4850 & n4908 ) ;
  assign n5252 = ( n1065 & n2570 ) | ( n1065 & ~n5251 ) | ( n2570 & ~n5251 ) ;
  assign n5247 = ~n322 & n3175 ;
  assign n5248 = n5247 ^ n797 ^ 1'b0 ;
  assign n5249 = ( n4044 & n5088 ) | ( n4044 & n5248 ) | ( n5088 & n5248 ) ;
  assign n5250 = n5249 ^ n5092 ^ n1735 ;
  assign n5253 = n5252 ^ n5250 ^ n4174 ;
  assign n5256 = n4711 ^ n1708 ^ n433 ;
  assign n5257 = n5256 ^ n2489 ^ n2368 ;
  assign n5254 = n4001 ^ n1844 ^ n163 ;
  assign n5255 = ~n954 & n5254 ;
  assign n5258 = n5257 ^ n5255 ^ 1'b0 ;
  assign n5259 = n5258 ^ n3626 ^ n3040 ;
  assign n5260 = n5259 ^ n997 ^ n289 ;
  assign n5261 = n2961 ^ n2213 ^ n1379 ;
  assign n5262 = n2683 ^ n694 ^ n224 ;
  assign n5263 = n5262 ^ n1241 ^ n810 ;
  assign n5264 = n5263 ^ n737 ^ 1'b0 ;
  assign n5265 = ~n5261 & n5264 ;
  assign n5266 = n2103 ^ n910 ^ n634 ;
  assign n5267 = n5266 ^ n2993 ^ n2600 ;
  assign n5268 = ( ~n1033 & n1850 ) | ( ~n1033 & n4639 ) | ( n1850 & n4639 ) ;
  assign n5269 = n1791 ^ n271 ^ 1'b0 ;
  assign n5270 = n1466 ^ n1281 ^ 1'b0 ;
  assign n5271 = ( n2322 & n3421 ) | ( n2322 & ~n5270 ) | ( n3421 & ~n5270 ) ;
  assign n5272 = n5271 ^ n4338 ^ n1345 ;
  assign n5273 = ( n1672 & n5269 ) | ( n1672 & ~n5272 ) | ( n5269 & ~n5272 ) ;
  assign n5274 = n4231 ^ n2371 ^ n1660 ;
  assign n5275 = ( ~n3742 & n5273 ) | ( ~n3742 & n5274 ) | ( n5273 & n5274 ) ;
  assign n5276 = ( n352 & n2220 ) | ( n352 & ~n3253 ) | ( n2220 & ~n3253 ) ;
  assign n5277 = n5276 ^ n678 ^ 1'b0 ;
  assign n5278 = n1170 & ~n2597 ;
  assign n5279 = n5278 ^ n410 ^ 1'b0 ;
  assign n5280 = n5277 & ~n5279 ;
  assign n5281 = n4704 ^ n3136 ^ n1374 ;
  assign n5282 = n5281 ^ n2582 ^ n2381 ;
  assign n5283 = n5282 ^ n4304 ^ n292 ;
  assign n5284 = n3404 ^ n2816 ^ 1'b0 ;
  assign n5285 = n5284 ^ n4283 ^ n3070 ;
  assign n5286 = n5285 ^ n3874 ^ n897 ;
  assign n5287 = ( n1374 & ~n3782 ) | ( n1374 & n4834 ) | ( ~n3782 & n4834 ) ;
  assign n5288 = ( n3035 & n3719 ) | ( n3035 & n5287 ) | ( n3719 & n5287 ) ;
  assign n5289 = n5288 ^ n3838 ^ n222 ;
  assign n5290 = n4802 ^ n2294 ^ 1'b0 ;
  assign n5291 = n5290 ^ n4396 ^ n1589 ;
  assign n5292 = ( n211 & n343 ) | ( n211 & ~n641 ) | ( n343 & ~n641 ) ;
  assign n5301 = ( n232 & n2124 ) | ( n232 & n3049 ) | ( n2124 & n3049 ) ;
  assign n5293 = n4154 ^ n2463 ^ x109 ;
  assign n5294 = n5293 ^ n5016 ^ n333 ;
  assign n5295 = n5294 ^ n2478 ^ n1543 ;
  assign n5296 = n2492 ^ n1185 ^ n495 ;
  assign n5297 = n2525 & n5296 ;
  assign n5298 = n5297 ^ n2947 ^ 1'b0 ;
  assign n5299 = ( n4830 & n5295 ) | ( n4830 & ~n5298 ) | ( n5295 & ~n5298 ) ;
  assign n5300 = ( n3942 & ~n3968 ) | ( n3942 & n5299 ) | ( ~n3968 & n5299 ) ;
  assign n5302 = n5301 ^ n5300 ^ n3539 ;
  assign n5303 = ( ~n187 & n419 ) | ( ~n187 & n1197 ) | ( n419 & n1197 ) ;
  assign n5304 = n5303 ^ n2365 ^ n871 ;
  assign n5307 = ( n1478 & n4061 ) | ( n1478 & ~n4794 ) | ( n4061 & ~n4794 ) ;
  assign n5308 = n5307 ^ n4977 ^ n4297 ;
  assign n5305 = ( n633 & n2580 ) | ( n633 & ~n3276 ) | ( n2580 & ~n3276 ) ;
  assign n5306 = ( n3133 & n4947 ) | ( n3133 & ~n5305 ) | ( n4947 & ~n5305 ) ;
  assign n5309 = n5308 ^ n5306 ^ n3825 ;
  assign n5310 = ( ~n2632 & n5304 ) | ( ~n2632 & n5309 ) | ( n5304 & n5309 ) ;
  assign n5317 = n3208 ^ n2927 ^ 1'b0 ;
  assign n5318 = n493 | n5317 ;
  assign n5316 = n4051 ^ n2633 ^ n1705 ;
  assign n5319 = n5318 ^ n5316 ^ n1971 ;
  assign n5320 = n5319 ^ n5215 ^ 1'b0 ;
  assign n5311 = ~n237 & n1702 ;
  assign n5312 = n2037 & n5311 ;
  assign n5313 = n5312 ^ n3114 ^ n2007 ;
  assign n5314 = n5313 ^ n4742 ^ n4588 ;
  assign n5315 = n2010 | n5314 ;
  assign n5321 = n5320 ^ n5315 ^ n438 ;
  assign n5322 = n825 & n2582 ;
  assign n5323 = ( ~n366 & n3740 ) | ( ~n366 & n4877 ) | ( n3740 & n4877 ) ;
  assign n5324 = n2227 | n5323 ;
  assign n5325 = n2953 & ~n5324 ;
  assign n5326 = ( n3888 & n4051 ) | ( n3888 & ~n5325 ) | ( n4051 & ~n5325 ) ;
  assign n5327 = n1106 ^ n756 ^ n728 ;
  assign n5328 = ( n1497 & n1772 ) | ( n1497 & ~n3746 ) | ( n1772 & ~n3746 ) ;
  assign n5329 = n5327 & n5328 ;
  assign n5330 = n5329 ^ n3239 ^ 1'b0 ;
  assign n5331 = n5330 ^ n1035 ^ n927 ;
  assign n5332 = ( n3914 & n5326 ) | ( n3914 & n5331 ) | ( n5326 & n5331 ) ;
  assign n5333 = ( n2549 & n5322 ) | ( n2549 & n5332 ) | ( n5322 & n5332 ) ;
  assign n5334 = ( ~n2851 & n3487 ) | ( ~n2851 & n5333 ) | ( n3487 & n5333 ) ;
  assign n5335 = n2981 ^ n939 ^ 1'b0 ;
  assign n5336 = ( n204 & n903 ) | ( n204 & ~n5335 ) | ( n903 & ~n5335 ) ;
  assign n5337 = n1143 | n4661 ;
  assign n5338 = ( n1576 & ~n2322 ) | ( n1576 & n5337 ) | ( ~n2322 & n5337 ) ;
  assign n5339 = n3133 ^ n2119 ^ n659 ;
  assign n5340 = n5339 ^ n3643 ^ 1'b0 ;
  assign n5341 = n3724 ^ n2486 ^ n567 ;
  assign n5342 = ~n3335 & n4618 ;
  assign n5343 = ~n5341 & n5342 ;
  assign n5344 = n5343 ^ n4354 ^ n3875 ;
  assign n5345 = ( n5338 & n5340 ) | ( n5338 & n5344 ) | ( n5340 & n5344 ) ;
  assign n5347 = n5088 ^ n1228 ^ 1'b0 ;
  assign n5348 = n1978 & ~n5347 ;
  assign n5349 = ( n472 & ~n4936 ) | ( n472 & n5348 ) | ( ~n4936 & n5348 ) ;
  assign n5346 = ( n393 & n795 ) | ( n393 & n4270 ) | ( n795 & n4270 ) ;
  assign n5350 = n5349 ^ n5346 ^ n431 ;
  assign n5359 = ( ~x95 & n922 ) | ( ~x95 & n1589 ) | ( n922 & n1589 ) ;
  assign n5351 = n4947 ^ n2695 ^ n1505 ;
  assign n5352 = n1753 | n3953 ;
  assign n5353 = n5352 ^ n439 ^ 1'b0 ;
  assign n5354 = n992 & ~n5353 ;
  assign n5355 = n5354 ^ n2490 ^ 1'b0 ;
  assign n5356 = n5355 ^ n1896 ^ 1'b0 ;
  assign n5357 = n5351 | n5356 ;
  assign n5358 = n4141 & n5357 ;
  assign n5360 = n5359 ^ n5358 ^ 1'b0 ;
  assign n5361 = ( x88 & ~n2104 ) | ( x88 & n4071 ) | ( ~n2104 & n4071 ) ;
  assign n5365 = n2810 ^ n364 ^ 1'b0 ;
  assign n5366 = n2770 & ~n5365 ;
  assign n5367 = n5366 ^ n3294 ^ 1'b0 ;
  assign n5368 = n5367 ^ n1263 ^ n204 ;
  assign n5362 = ( x0 & n176 ) | ( x0 & n1571 ) | ( n176 & n1571 ) ;
  assign n5363 = ( x2 & n2394 ) | ( x2 & n5362 ) | ( n2394 & n5362 ) ;
  assign n5364 = n5363 ^ n821 ^ n305 ;
  assign n5369 = n5368 ^ n5364 ^ n4167 ;
  assign n5370 = n3367 & ~n5369 ;
  assign n5371 = n5157 ^ n3633 ^ 1'b0 ;
  assign n5372 = ~n3162 & n5371 ;
  assign n5373 = n4115 & ~n5372 ;
  assign n5374 = ( ~n5020 & n5370 ) | ( ~n5020 & n5373 ) | ( n5370 & n5373 ) ;
  assign n5375 = ( ~n3898 & n4257 ) | ( ~n3898 & n4701 ) | ( n4257 & n4701 ) ;
  assign n5376 = n2912 ^ n2306 ^ n1497 ;
  assign n5377 = n5376 ^ n2359 ^ n1335 ;
  assign n5378 = n5377 ^ n4834 ^ n1988 ;
  assign n5379 = n5301 ^ n4303 ^ n1650 ;
  assign n5380 = ( n690 & n1004 ) | ( n690 & n1273 ) | ( n1004 & n1273 ) ;
  assign n5381 = n5380 ^ n2026 ^ n1246 ;
  assign n5382 = ( n1888 & n3762 ) | ( n1888 & n5381 ) | ( n3762 & n5381 ) ;
  assign n5383 = ( n5378 & n5379 ) | ( n5378 & n5382 ) | ( n5379 & n5382 ) ;
  assign n5384 = ( n833 & n4062 ) | ( n833 & n5383 ) | ( n4062 & n5383 ) ;
  assign n5388 = x42 & x47 ;
  assign n5389 = n361 & n5388 ;
  assign n5385 = ( n478 & ~n823 ) | ( n478 & n1423 ) | ( ~n823 & n1423 ) ;
  assign n5386 = ( ~n1982 & n3459 ) | ( ~n1982 & n4904 ) | ( n3459 & n4904 ) ;
  assign n5387 = ( n2510 & ~n5385 ) | ( n2510 & n5386 ) | ( ~n5385 & n5386 ) ;
  assign n5390 = n5389 ^ n5387 ^ n641 ;
  assign n5391 = ( n5375 & n5384 ) | ( n5375 & ~n5390 ) | ( n5384 & ~n5390 ) ;
  assign n5392 = n5391 ^ n4299 ^ n2610 ;
  assign n5393 = ( n540 & n1022 ) | ( n540 & n2113 ) | ( n1022 & n2113 ) ;
  assign n5394 = n4963 ^ n4809 ^ n3493 ;
  assign n5395 = ( ~n211 & n900 ) | ( ~n211 & n1086 ) | ( n900 & n1086 ) ;
  assign n5396 = ( ~n1933 & n2996 ) | ( ~n1933 & n5395 ) | ( n2996 & n5395 ) ;
  assign n5397 = n3159 & ~n5396 ;
  assign n5398 = n4907 ^ n2489 ^ n574 ;
  assign n5399 = n5398 ^ n405 ^ 1'b0 ;
  assign n5400 = ~n5014 & n5399 ;
  assign n5401 = n4799 ^ x84 ^ 1'b0 ;
  assign n5402 = n1712 & ~n5401 ;
  assign n5408 = n3995 ^ n3836 ^ x108 ;
  assign n5405 = ~n568 & n4910 ;
  assign n5406 = n5405 ^ n809 ^ x113 ;
  assign n5403 = ( x112 & ~n349 ) | ( x112 & n669 ) | ( ~n349 & n669 ) ;
  assign n5404 = n1715 & n5403 ;
  assign n5407 = n5406 ^ n5404 ^ 1'b0 ;
  assign n5409 = n5408 ^ n5407 ^ n2678 ;
  assign n5410 = ( n136 & n764 ) | ( n136 & n1463 ) | ( n764 & n1463 ) ;
  assign n5411 = n2278 ^ n1657 ^ n629 ;
  assign n5412 = ( n284 & n1280 ) | ( n284 & ~n5411 ) | ( n1280 & ~n5411 ) ;
  assign n5413 = n5410 & ~n5412 ;
  assign n5414 = ~n5409 & n5413 ;
  assign n5415 = n5402 & ~n5414 ;
  assign n5417 = ( x109 & n365 ) | ( x109 & n757 ) | ( n365 & n757 ) ;
  assign n5416 = n637 ^ x44 ^ 1'b0 ;
  assign n5418 = n5417 ^ n5416 ^ n4383 ;
  assign n5419 = n5418 ^ n2722 ^ n257 ;
  assign n5420 = n5419 ^ n3494 ^ n1803 ;
  assign n5421 = n5420 ^ n3994 ^ 1'b0 ;
  assign n5430 = n3002 ^ n339 ^ 1'b0 ;
  assign n5431 = n5430 ^ n4517 ^ n716 ;
  assign n5433 = n3073 ^ n2360 ^ n1738 ;
  assign n5434 = n5433 ^ n1618 ^ n721 ;
  assign n5432 = ( n3289 & n3562 ) | ( n3289 & ~n3616 ) | ( n3562 & ~n3616 ) ;
  assign n5435 = n5434 ^ n5432 ^ 1'b0 ;
  assign n5436 = n5431 | n5435 ;
  assign n5437 = n5436 ^ n5419 ^ n1556 ;
  assign n5422 = n1463 & n1866 ;
  assign n5423 = ~n457 & n5422 ;
  assign n5424 = ( n393 & ~n2097 ) | ( n393 & n3102 ) | ( ~n2097 & n3102 ) ;
  assign n5425 = n157 & ~n3819 ;
  assign n5426 = ( n1116 & n4256 ) | ( n1116 & n5425 ) | ( n4256 & n5425 ) ;
  assign n5427 = n5426 ^ n2476 ^ n435 ;
  assign n5428 = ( ~n3230 & n4673 ) | ( ~n3230 & n5427 ) | ( n4673 & n5427 ) ;
  assign n5429 = ( n5423 & n5424 ) | ( n5423 & ~n5428 ) | ( n5424 & ~n5428 ) ;
  assign n5438 = n5437 ^ n5429 ^ 1'b0 ;
  assign n5439 = ( ~n487 & n1308 ) | ( ~n487 & n2391 ) | ( n1308 & n2391 ) ;
  assign n5440 = n755 & ~n914 ;
  assign n5441 = n5440 ^ n3520 ^ 1'b0 ;
  assign n5442 = ( n4497 & ~n5439 ) | ( n4497 & n5441 ) | ( ~n5439 & n5441 ) ;
  assign n5443 = n5442 ^ n5385 ^ n1470 ;
  assign n5444 = n3478 ^ n2064 ^ 1'b0 ;
  assign n5445 = ( n4073 & ~n5443 ) | ( n4073 & n5444 ) | ( ~n5443 & n5444 ) ;
  assign n5446 = n3179 ^ n2930 ^ n1808 ;
  assign n5453 = n984 ^ n921 ^ 1'b0 ;
  assign n5454 = n4519 & ~n5453 ;
  assign n5456 = ( n879 & ~n1241 ) | ( n879 & n4633 ) | ( ~n1241 & n4633 ) ;
  assign n5455 = n2288 & ~n3835 ;
  assign n5457 = n5456 ^ n5455 ^ 1'b0 ;
  assign n5458 = n5457 ^ n732 ^ n145 ;
  assign n5459 = n5458 ^ n2970 ^ n1369 ;
  assign n5460 = ( n2515 & n5454 ) | ( n2515 & ~n5459 ) | ( n5454 & ~n5459 ) ;
  assign n5447 = x67 & ~n4620 ;
  assign n5448 = n3500 ^ n2286 ^ n130 ;
  assign n5449 = n5448 ^ n4015 ^ n330 ;
  assign n5450 = ( n2402 & n3429 ) | ( n2402 & n5449 ) | ( n3429 & n5449 ) ;
  assign n5451 = n4983 | n5450 ;
  assign n5452 = n5447 & ~n5451 ;
  assign n5461 = n5460 ^ n5452 ^ n190 ;
  assign n5463 = ( ~n405 & n2115 ) | ( ~n405 & n2604 ) | ( n2115 & n2604 ) ;
  assign n5462 = n3510 ^ n3179 ^ n252 ;
  assign n5464 = n5463 ^ n5462 ^ n5195 ;
  assign n5465 = n5464 ^ n2853 ^ n2052 ;
  assign n5466 = n807 ^ n586 ^ n446 ;
  assign n5467 = ( n525 & ~n1003 ) | ( n525 & n3342 ) | ( ~n1003 & n3342 ) ;
  assign n5468 = ~n5466 & n5467 ;
  assign n5470 = n982 & ~n4676 ;
  assign n5469 = n4068 ^ n1563 ^ x7 ;
  assign n5471 = n5470 ^ n5469 ^ n773 ;
  assign n5472 = ( ~n1155 & n2645 ) | ( ~n1155 & n4949 ) | ( n2645 & n4949 ) ;
  assign n5473 = n5472 ^ n5361 ^ 1'b0 ;
  assign n5474 = n3057 & ~n5473 ;
  assign n5475 = n5088 ^ n1823 ^ n146 ;
  assign n5476 = n5475 ^ n5231 ^ n2923 ;
  assign n5477 = ( n1342 & ~n2486 ) | ( n1342 & n5476 ) | ( ~n2486 & n5476 ) ;
  assign n5478 = n3394 ^ n2454 ^ n1069 ;
  assign n5489 = n1726 ^ n328 ^ 1'b0 ;
  assign n5490 = n5489 ^ n1744 ^ 1'b0 ;
  assign n5491 = ( ~n2108 & n5040 ) | ( ~n2108 & n5490 ) | ( n5040 & n5490 ) ;
  assign n5483 = n2032 ^ n271 ^ x76 ;
  assign n5484 = ( ~n1261 & n1710 ) | ( ~n1261 & n1819 ) | ( n1710 & n1819 ) ;
  assign n5485 = n2877 ^ n556 ^ n170 ;
  assign n5486 = ( n5483 & n5484 ) | ( n5483 & ~n5485 ) | ( n5484 & ~n5485 ) ;
  assign n5480 = ( x126 & n1304 ) | ( x126 & n2556 ) | ( n1304 & n2556 ) ;
  assign n5481 = n1605 ^ n901 ^ 1'b0 ;
  assign n5482 = n5480 & ~n5481 ;
  assign n5479 = n3220 ^ n2041 ^ n491 ;
  assign n5487 = n5486 ^ n5482 ^ n5479 ;
  assign n5488 = n5487 ^ n4418 ^ n2262 ;
  assign n5492 = n5491 ^ n5488 ^ n588 ;
  assign n5493 = ( n1507 & n3172 ) | ( n1507 & ~n5492 ) | ( n3172 & ~n5492 ) ;
  assign n5496 = ( ~n428 & n549 ) | ( ~n428 & n1515 ) | ( n549 & n1515 ) ;
  assign n5494 = n3404 ^ n1181 ^ 1'b0 ;
  assign n5495 = n5494 ^ n1524 ^ n578 ;
  assign n5497 = n5496 ^ n5495 ^ n604 ;
  assign n5498 = n3758 | n5497 ;
  assign n5499 = n4315 ^ n3692 ^ n1182 ;
  assign n5500 = ( n679 & ~n3936 ) | ( n679 & n5499 ) | ( ~n3936 & n5499 ) ;
  assign n5501 = ( n360 & n2498 ) | ( n360 & ~n3256 ) | ( n2498 & ~n3256 ) ;
  assign n5502 = n4485 ^ n250 ^ 1'b0 ;
  assign n5503 = ( ~n268 & n2831 ) | ( ~n268 & n4770 ) | ( n2831 & n4770 ) ;
  assign n5504 = n4811 ^ n4555 ^ n3761 ;
  assign n5505 = ( n2721 & n3944 ) | ( n2721 & ~n5504 ) | ( n3944 & ~n5504 ) ;
  assign n5506 = n5503 & n5505 ;
  assign n5507 = n5506 ^ n1614 ^ 1'b0 ;
  assign n5508 = n5507 ^ n4800 ^ n887 ;
  assign n5509 = ~n1768 & n5508 ;
  assign n5510 = n5502 & n5509 ;
  assign n5511 = n1791 ^ n1353 ^ 1'b0 ;
  assign n5512 = n3670 | n5511 ;
  assign n5513 = ( n692 & n1780 ) | ( n692 & ~n5512 ) | ( n1780 & ~n5512 ) ;
  assign n5514 = n2958 ^ n2716 ^ n1697 ;
  assign n5515 = ( n2989 & n3037 ) | ( n2989 & n5514 ) | ( n3037 & n5514 ) ;
  assign n5516 = ( ~n1788 & n3374 ) | ( ~n1788 & n5515 ) | ( n3374 & n5515 ) ;
  assign n5517 = n3942 ^ n1052 ^ 1'b0 ;
  assign n5518 = n5517 ^ n1650 ^ 1'b0 ;
  assign n5519 = n1225 & ~n5518 ;
  assign n5520 = n5519 ^ n500 ^ 1'b0 ;
  assign n5521 = n5516 & n5520 ;
  assign n5522 = n3562 ^ n2791 ^ n1486 ;
  assign n5523 = n3843 | n5522 ;
  assign n5524 = n249 & ~n5523 ;
  assign n5525 = n5524 ^ n4930 ^ n3792 ;
  assign n5526 = ( n621 & ~n3185 ) | ( n621 & n5525 ) | ( ~n3185 & n5525 ) ;
  assign n5527 = ( n2110 & n5521 ) | ( n2110 & n5526 ) | ( n5521 & n5526 ) ;
  assign n5528 = n4016 ^ n3734 ^ 1'b0 ;
  assign n5529 = ~n1079 & n1717 ;
  assign n5530 = ~n1175 & n5529 ;
  assign n5531 = ( x58 & n811 ) | ( x58 & n2309 ) | ( n811 & n2309 ) ;
  assign n5532 = ( ~n1845 & n4674 ) | ( ~n1845 & n5531 ) | ( n4674 & n5531 ) ;
  assign n5533 = ( n825 & n5530 ) | ( n825 & n5532 ) | ( n5530 & n5532 ) ;
  assign n5534 = ( n264 & n3028 ) | ( n264 & n5533 ) | ( n3028 & n5533 ) ;
  assign n5539 = n2276 ^ n2147 ^ n139 ;
  assign n5535 = ( n669 & n772 ) | ( n669 & n1421 ) | ( n772 & n1421 ) ;
  assign n5536 = n5535 ^ n3956 ^ n947 ;
  assign n5537 = n5536 ^ n1830 ^ n506 ;
  assign n5538 = n3199 | n5537 ;
  assign n5540 = n5539 ^ n5538 ^ n1618 ;
  assign n5541 = n5540 ^ n5123 ^ n4264 ;
  assign n5559 = n3589 ^ n1083 ^ 1'b0 ;
  assign n5560 = ~n694 & n5559 ;
  assign n5550 = n1999 ^ n398 ^ n290 ;
  assign n5547 = ( n934 & ~n1491 ) | ( n934 & n2326 ) | ( ~n1491 & n2326 ) ;
  assign n5548 = n1147 & ~n5547 ;
  assign n5549 = ( n1000 & ~n1559 ) | ( n1000 & n5548 ) | ( ~n1559 & n5548 ) ;
  assign n5545 = n1612 ^ n1331 ^ n566 ;
  assign n5542 = ( n180 & n2264 ) | ( n180 & ~n3046 ) | ( n2264 & ~n3046 ) ;
  assign n5543 = n3275 ^ n1353 ^ 1'b0 ;
  assign n5544 = ( ~n2563 & n5542 ) | ( ~n2563 & n5543 ) | ( n5542 & n5543 ) ;
  assign n5546 = n5545 ^ n5544 ^ n4259 ;
  assign n5551 = n5550 ^ n5549 ^ n5546 ;
  assign n5553 = n2106 ^ n1537 ^ n603 ;
  assign n5554 = ( ~n781 & n985 ) | ( ~n781 & n5553 ) | ( n985 & n5553 ) ;
  assign n5552 = ( ~n2360 & n3439 ) | ( ~n2360 & n3615 ) | ( n3439 & n3615 ) ;
  assign n5555 = n5554 ^ n5552 ^ n1298 ;
  assign n5556 = n3998 ^ n3369 ^ n3311 ;
  assign n5557 = n5556 ^ n3726 ^ n759 ;
  assign n5558 = ( n5551 & ~n5555 ) | ( n5551 & n5557 ) | ( ~n5555 & n5557 ) ;
  assign n5561 = n5560 ^ n5558 ^ n4052 ;
  assign n5562 = ( n744 & n1597 ) | ( n744 & n3120 ) | ( n1597 & n3120 ) ;
  assign n5563 = n880 | n2367 ;
  assign n5564 = n2304 & ~n5563 ;
  assign n5565 = ( n2159 & ~n5562 ) | ( n2159 & n5564 ) | ( ~n5562 & n5564 ) ;
  assign n5569 = n2726 ^ n2019 ^ n1438 ;
  assign n5568 = n2308 ^ x108 ^ 1'b0 ;
  assign n5570 = n5569 ^ n5568 ^ n4023 ;
  assign n5566 = ( n1800 & n2385 ) | ( n1800 & n2457 ) | ( n2385 & n2457 ) ;
  assign n5567 = n5566 ^ n2541 ^ n557 ;
  assign n5571 = n5570 ^ n5567 ^ 1'b0 ;
  assign n5572 = n4447 ^ n2619 ^ n735 ;
  assign n5573 = n205 & n5230 ;
  assign n5574 = n5572 & n5573 ;
  assign n5575 = n4798 ^ n2406 ^ x95 ;
  assign n5576 = n5575 ^ n2182 ^ n571 ;
  assign n5577 = ( x41 & n4242 ) | ( x41 & ~n5576 ) | ( n4242 & ~n5576 ) ;
  assign n5578 = ( n714 & ~n985 ) | ( n714 & n3131 ) | ( ~n985 & n3131 ) ;
  assign n5579 = ( n971 & n3801 ) | ( n971 & ~n5578 ) | ( n3801 & ~n5578 ) ;
  assign n5580 = n5579 ^ n610 ^ n313 ;
  assign n5581 = n5486 ^ n2925 ^ n2197 ;
  assign n5582 = n277 & ~n5581 ;
  assign n5583 = n2421 & n5582 ;
  assign n5584 = n1282 ^ n951 ^ n826 ;
  assign n5585 = ~n3104 & n5584 ;
  assign n5586 = ~n822 & n5585 ;
  assign n5587 = ( n3120 & n5583 ) | ( n3120 & n5586 ) | ( n5583 & n5586 ) ;
  assign n5588 = ( ~x100 & n1366 ) | ( ~x100 & n2209 ) | ( n1366 & n2209 ) ;
  assign n5589 = n5167 ^ n1043 ^ x86 ;
  assign n5590 = ( n5543 & ~n5588 ) | ( n5543 & n5589 ) | ( ~n5588 & n5589 ) ;
  assign n5591 = ( ~n165 & n1083 ) | ( ~n165 & n3404 ) | ( n1083 & n3404 ) ;
  assign n5592 = n4751 ^ n679 ^ 1'b0 ;
  assign n5593 = n5591 | n5592 ;
  assign n5594 = n5590 | n5593 ;
  assign n5595 = ( n5580 & ~n5587 ) | ( n5580 & n5594 ) | ( ~n5587 & n5594 ) ;
  assign n5596 = n877 & n3747 ;
  assign n5597 = ~n4083 & n5596 ;
  assign n5598 = n482 ^ n403 ^ 1'b0 ;
  assign n5599 = ~n4790 & n5598 ;
  assign n5600 = ( n2453 & n3178 ) | ( n2453 & ~n5599 ) | ( n3178 & ~n5599 ) ;
  assign n5601 = ( n1836 & n5597 ) | ( n1836 & n5600 ) | ( n5597 & n5600 ) ;
  assign n5602 = ( n966 & n2879 ) | ( n966 & ~n3943 ) | ( n2879 & ~n3943 ) ;
  assign n5603 = n5602 ^ n5474 ^ n405 ;
  assign n5606 = ( ~x84 & n1487 ) | ( ~x84 & n5530 ) | ( n1487 & n5530 ) ;
  assign n5607 = ( n1353 & n2582 ) | ( n1353 & ~n5606 ) | ( n2582 & ~n5606 ) ;
  assign n5608 = n5607 ^ n1070 ^ n606 ;
  assign n5605 = n4014 ^ n3647 ^ n2038 ;
  assign n5604 = n2010 ^ n989 ^ 1'b0 ;
  assign n5609 = n5608 ^ n5605 ^ n5604 ;
  assign n5610 = n5077 ^ n1689 ^ n1594 ;
  assign n5611 = n5610 ^ n4409 ^ n2490 ;
  assign n5612 = n344 & ~n5611 ;
  assign n5613 = n1330 ^ n885 ^ 1'b0 ;
  assign n5614 = ( n811 & ~n2562 ) | ( n811 & n5613 ) | ( ~n2562 & n5613 ) ;
  assign n5615 = n4014 ^ n1305 ^ n1254 ;
  assign n5616 = ( n188 & ~n5614 ) | ( n188 & n5615 ) | ( ~n5614 & n5615 ) ;
  assign n5617 = n3643 ^ n3409 ^ n3223 ;
  assign n5618 = ( n857 & n2389 ) | ( n857 & ~n3982 ) | ( n2389 & ~n3982 ) ;
  assign n5619 = ( n2898 & ~n3035 ) | ( n2898 & n5618 ) | ( ~n3035 & n5618 ) ;
  assign n5620 = n5619 ^ n5223 ^ n858 ;
  assign n5621 = ( n2964 & n5617 ) | ( n2964 & n5620 ) | ( n5617 & n5620 ) ;
  assign n5622 = ( ~n1174 & n2211 ) | ( ~n1174 & n2466 ) | ( n2211 & n2466 ) ;
  assign n5623 = n5622 ^ n529 ^ n304 ;
  assign n5624 = ( n800 & ~n4818 ) | ( n800 & n5623 ) | ( ~n4818 & n5623 ) ;
  assign n5625 = n4897 ^ n4517 ^ n3677 ;
  assign n5626 = ( n3808 & ~n3897 ) | ( n3808 & n5625 ) | ( ~n3897 & n5625 ) ;
  assign n5627 = n5626 ^ n780 ^ 1'b0 ;
  assign n5628 = n1758 ^ n645 ^ x48 ;
  assign n5629 = n5628 ^ n1297 ^ x109 ;
  assign n5630 = ( n2040 & ~n4289 ) | ( n2040 & n5629 ) | ( ~n4289 & n5629 ) ;
  assign n5631 = n1563 ^ n470 ^ 1'b0 ;
  assign n5632 = n5630 | n5631 ;
  assign n5633 = n5632 ^ n5239 ^ n4418 ;
  assign n5634 = n4796 ^ n2963 ^ n399 ;
  assign n5635 = ( n477 & ~n3390 ) | ( n477 & n5634 ) | ( ~n3390 & n5634 ) ;
  assign n5639 = n879 | n1139 ;
  assign n5637 = ( n1986 & n2105 ) | ( n1986 & ~n2774 ) | ( n2105 & ~n2774 ) ;
  assign n5636 = ( n1328 & ~n3982 ) | ( n1328 & n4248 ) | ( ~n3982 & n4248 ) ;
  assign n5638 = n5637 ^ n5636 ^ n2079 ;
  assign n5640 = n5639 ^ n5638 ^ n628 ;
  assign n5641 = ( n5114 & ~n5635 ) | ( n5114 & n5640 ) | ( ~n5635 & n5640 ) ;
  assign n5645 = n861 ^ n574 ^ x66 ;
  assign n5646 = n5645 ^ n2027 ^ n1791 ;
  assign n5644 = ( n1297 & n2595 ) | ( n1297 & ~n4692 ) | ( n2595 & ~n4692 ) ;
  assign n5642 = n3265 ^ x61 ^ 1'b0 ;
  assign n5643 = ( n3788 & ~n3820 ) | ( n3788 & n5642 ) | ( ~n3820 & n5642 ) ;
  assign n5647 = n5646 ^ n5644 ^ n5643 ;
  assign n5648 = n5647 ^ n5369 ^ n475 ;
  assign n5654 = n2314 ^ n1586 ^ n1259 ;
  assign n5649 = n3992 ^ n3392 ^ x21 ;
  assign n5650 = n3325 ^ n171 ^ 1'b0 ;
  assign n5651 = ~n1997 & n5650 ;
  assign n5652 = ~n5649 & n5651 ;
  assign n5653 = n2073 & n5652 ;
  assign n5655 = n5654 ^ n5653 ^ 1'b0 ;
  assign n5660 = n2419 ^ n599 ^ n209 ;
  assign n5659 = ( n512 & ~n2025 ) | ( n512 & n3776 ) | ( ~n2025 & n3776 ) ;
  assign n5656 = n4834 ^ n2297 ^ n1203 ;
  assign n5657 = n5656 ^ n2252 ^ n2134 ;
  assign n5658 = n5657 ^ n3964 ^ n3167 ;
  assign n5661 = n5660 ^ n5659 ^ n5658 ;
  assign n5662 = n5661 ^ n3290 ^ x11 ;
  assign n5663 = n3141 | n5662 ;
  assign n5664 = n5655 & ~n5663 ;
  assign n5665 = ( ~n3652 & n5648 ) | ( ~n3652 & n5664 ) | ( n5648 & n5664 ) ;
  assign n5666 = n3523 ^ n1990 ^ n1782 ;
  assign n5667 = n4951 ^ n3114 ^ n2159 ;
  assign n5668 = ( ~n2449 & n5666 ) | ( ~n2449 & n5667 ) | ( n5666 & n5667 ) ;
  assign n5684 = n5349 ^ n1574 ^ n197 ;
  assign n5678 = n881 & n4751 ;
  assign n5679 = n5678 ^ n1759 ^ n1657 ;
  assign n5680 = ( ~n1692 & n2246 ) | ( ~n1692 & n5466 ) | ( n2246 & n5466 ) ;
  assign n5681 = n5680 ^ n2641 ^ 1'b0 ;
  assign n5682 = ~n5679 & n5681 ;
  assign n5683 = n5682 ^ n2009 ^ n1278 ;
  assign n5685 = n5684 ^ n5683 ^ n5619 ;
  assign n5674 = ( n734 & n1269 ) | ( n734 & n4961 ) | ( n1269 & n4961 ) ;
  assign n5675 = ( n883 & n1131 ) | ( n883 & ~n5674 ) | ( n1131 & ~n5674 ) ;
  assign n5670 = ( n244 & ~n1112 ) | ( n244 & n1802 ) | ( ~n1112 & n1802 ) ;
  assign n5671 = n5670 ^ n601 ^ n469 ;
  assign n5669 = n4446 ^ n2139 ^ 1'b0 ;
  assign n5672 = n5671 ^ n5669 ^ n2295 ;
  assign n5673 = n5672 ^ n4834 ^ n863 ;
  assign n5676 = n5675 ^ n5673 ^ 1'b0 ;
  assign n5677 = ~n3449 & n5676 ;
  assign n5686 = n5685 ^ n5677 ^ n4769 ;
  assign n5687 = n5642 & ~n5686 ;
  assign n5688 = ~n5668 & n5687 ;
  assign n5695 = ( ~n2686 & n3127 ) | ( ~n2686 & n4843 ) | ( n3127 & n4843 ) ;
  assign n5696 = n5695 ^ n3274 ^ n1339 ;
  assign n5693 = n1515 ^ n1510 ^ n153 ;
  assign n5694 = n5693 ^ n2983 ^ n1044 ;
  assign n5697 = n5696 ^ n5694 ^ n719 ;
  assign n5689 = n3556 & ~n5578 ;
  assign n5690 = n5689 ^ n4236 ^ 1'b0 ;
  assign n5691 = ( n2424 & ~n4240 ) | ( n2424 & n5690 ) | ( ~n4240 & n5690 ) ;
  assign n5692 = n5691 ^ n2826 ^ n365 ;
  assign n5698 = n5697 ^ n5692 ^ n1751 ;
  assign n5701 = ( n438 & ~n1106 ) | ( n438 & n2034 ) | ( ~n1106 & n2034 ) ;
  assign n5702 = ( n1612 & n5124 ) | ( n1612 & ~n5701 ) | ( n5124 & ~n5701 ) ;
  assign n5703 = ( n558 & ~n2010 ) | ( n558 & n5702 ) | ( ~n2010 & n5702 ) ;
  assign n5699 = n649 ^ x6 ^ 1'b0 ;
  assign n5700 = n5699 ^ n4802 ^ n2624 ;
  assign n5704 = n5703 ^ n5700 ^ n1013 ;
  assign n5705 = n3738 ^ n749 ^ 1'b0 ;
  assign n5706 = ( ~n3543 & n3802 ) | ( ~n3543 & n5051 ) | ( n3802 & n5051 ) ;
  assign n5707 = n5482 ^ n4905 ^ 1'b0 ;
  assign n5708 = ~n5706 & n5707 ;
  assign n5709 = n5708 ^ n3386 ^ n977 ;
  assign n5710 = n5705 & n5709 ;
  assign n5711 = ~n5704 & n5710 ;
  assign n5712 = n1065 & ~n2217 ;
  assign n5713 = n5712 ^ n1076 ^ 1'b0 ;
  assign n5714 = n5713 ^ n3694 ^ 1'b0 ;
  assign n5715 = n2727 & n5714 ;
  assign n5716 = ( n361 & n2797 ) | ( n361 & n4074 ) | ( n2797 & n4074 ) ;
  assign n5717 = ( n848 & n2139 ) | ( n848 & n4775 ) | ( n2139 & n4775 ) ;
  assign n5721 = ( x50 & ~n167 ) | ( x50 & n2166 ) | ( ~n167 & n2166 ) ;
  assign n5722 = n5721 ^ n1543 ^ n939 ;
  assign n5723 = n5722 ^ n1862 ^ x127 ;
  assign n5718 = n2770 ^ n595 ^ n229 ;
  assign n5719 = ( x16 & n215 ) | ( x16 & ~n5084 ) | ( n215 & ~n5084 ) ;
  assign n5720 = ( n1506 & ~n5718 ) | ( n1506 & n5719 ) | ( ~n5718 & n5719 ) ;
  assign n5724 = n5723 ^ n5720 ^ n452 ;
  assign n5725 = n588 & n1729 ;
  assign n5726 = x13 & ~n5725 ;
  assign n5727 = ~n5724 & n5726 ;
  assign n5728 = ( n3830 & ~n5717 ) | ( n3830 & n5727 ) | ( ~n5717 & n5727 ) ;
  assign n5729 = ( n5116 & ~n5716 ) | ( n5116 & n5728 ) | ( ~n5716 & n5728 ) ;
  assign n5730 = n1277 | n5194 ;
  assign n5731 = n4149 | n5730 ;
  assign n5732 = n5731 ^ n1448 ^ n867 ;
  assign n5733 = n5095 ^ n3836 ^ n2456 ;
  assign n5734 = ( n1557 & ~n4645 ) | ( n1557 & n5733 ) | ( ~n4645 & n5733 ) ;
  assign n5739 = ( n1331 & ~n2875 ) | ( n1331 & n3118 ) | ( ~n2875 & n3118 ) ;
  assign n5740 = ( n676 & n3276 ) | ( n676 & n5739 ) | ( n3276 & n5739 ) ;
  assign n5741 = n5740 ^ n3172 ^ n502 ;
  assign n5737 = ( n335 & ~n2719 ) | ( n335 & n3278 ) | ( ~n2719 & n3278 ) ;
  assign n5738 = n5737 ^ n2335 ^ n314 ;
  assign n5735 = ( n1282 & n2741 ) | ( n1282 & n3555 ) | ( n2741 & n3555 ) ;
  assign n5736 = n5735 ^ n4838 ^ n2937 ;
  assign n5742 = n5741 ^ n5738 ^ n5736 ;
  assign n5743 = ( n322 & ~n1546 ) | ( n322 & n4313 ) | ( ~n1546 & n4313 ) ;
  assign n5744 = n5743 ^ n5379 ^ n4221 ;
  assign n5745 = n1762 ^ n1209 ^ n1065 ;
  assign n5746 = n4091 ^ n973 ^ n896 ;
  assign n5747 = n5745 & n5746 ;
  assign n5748 = n5747 ^ n4041 ^ n1750 ;
  assign n5749 = n5430 ^ n4211 ^ n3028 ;
  assign n5750 = ( ~n3150 & n5748 ) | ( ~n3150 & n5749 ) | ( n5748 & n5749 ) ;
  assign n5751 = n2757 & ~n5750 ;
  assign n5752 = n5744 & n5751 ;
  assign n5753 = ( ~n5734 & n5742 ) | ( ~n5734 & n5752 ) | ( n5742 & n5752 ) ;
  assign n5754 = ( n274 & n2889 ) | ( n274 & ~n3094 ) | ( n2889 & ~n3094 ) ;
  assign n5755 = ( n2915 & n3289 ) | ( n2915 & ~n5754 ) | ( n3289 & ~n5754 ) ;
  assign n5756 = n5755 ^ n5626 ^ n1794 ;
  assign n5757 = n3572 ^ n2132 ^ n760 ;
  assign n5758 = n5757 ^ n5418 ^ n3165 ;
  assign n5759 = n5133 & ~n5758 ;
  assign n5760 = n5756 & n5759 ;
  assign n5768 = ( n206 & n2069 ) | ( n206 & ~n2291 ) | ( n2069 & ~n2291 ) ;
  assign n5763 = n3905 ^ n1224 ^ n164 ;
  assign n5764 = n2999 | n5763 ;
  assign n5765 = n136 | n5764 ;
  assign n5761 = ( ~n309 & n1245 ) | ( ~n309 & n1461 ) | ( n1245 & n1461 ) ;
  assign n5762 = n5761 ^ n4463 ^ n344 ;
  assign n5766 = n5765 ^ n5762 ^ n3085 ;
  assign n5767 = ( ~n2401 & n4067 ) | ( ~n2401 & n5766 ) | ( n4067 & n5766 ) ;
  assign n5769 = n5768 ^ n5767 ^ n3316 ;
  assign n5770 = n1587 ^ n1429 ^ n250 ;
  assign n5774 = n2218 ^ n1808 ^ n614 ;
  assign n5775 = ( n989 & ~n1605 ) | ( n989 & n5774 ) | ( ~n1605 & n5774 ) ;
  assign n5776 = ( n496 & n2388 ) | ( n496 & ~n5775 ) | ( n2388 & ~n5775 ) ;
  assign n5771 = ( ~n2391 & n4733 ) | ( ~n2391 & n4794 ) | ( n4733 & n4794 ) ;
  assign n5772 = n5771 ^ n3022 ^ 1'b0 ;
  assign n5773 = n3410 | n5772 ;
  assign n5777 = n5776 ^ n5773 ^ n3230 ;
  assign n5778 = ( n3188 & n5770 ) | ( n3188 & ~n5777 ) | ( n5770 & ~n5777 ) ;
  assign n5782 = n4233 ^ n4056 ^ n1559 ;
  assign n5779 = n3159 ^ n1689 ^ n779 ;
  assign n5780 = n5779 ^ n192 ^ 1'b0 ;
  assign n5781 = ( n194 & ~n2024 ) | ( n194 & n5780 ) | ( ~n2024 & n5780 ) ;
  assign n5783 = n5782 ^ n5781 ^ n3037 ;
  assign n5784 = ( ~n1226 & n1295 ) | ( ~n1226 & n3930 ) | ( n1295 & n3930 ) ;
  assign n5785 = ( ~n3319 & n4761 ) | ( ~n3319 & n5784 ) | ( n4761 & n5784 ) ;
  assign n5786 = n5785 ^ n1695 ^ n246 ;
  assign n5787 = ( x79 & ~n879 ) | ( x79 & n2673 ) | ( ~n879 & n2673 ) ;
  assign n5788 = ( n1727 & ~n5786 ) | ( n1727 & n5787 ) | ( ~n5786 & n5787 ) ;
  assign n5794 = n890 ^ n382 ^ n209 ;
  assign n5793 = n1301 ^ n974 ^ x6 ;
  assign n5795 = n5794 ^ n5793 ^ n1870 ;
  assign n5789 = n170 & ~n2060 ;
  assign n5790 = ~n2257 & n5789 ;
  assign n5791 = n3562 ^ n2874 ^ n276 ;
  assign n5792 = ( n2391 & ~n5790 ) | ( n2391 & n5791 ) | ( ~n5790 & n5791 ) ;
  assign n5796 = n5795 ^ n5792 ^ n4607 ;
  assign n5797 = n5078 ^ n1141 ^ n398 ;
  assign n5798 = n5363 ^ n2155 ^ n780 ;
  assign n5811 = n4232 ^ n2129 ^ n1951 ;
  assign n5810 = n4282 ^ n4186 ^ n1868 ;
  assign n5799 = n3010 ^ n880 ^ 1'b0 ;
  assign n5800 = n1965 ^ n624 ^ n278 ;
  assign n5801 = n1035 ^ n433 ^ 1'b0 ;
  assign n5802 = n5800 & n5801 ;
  assign n5803 = ( ~n2737 & n4878 ) | ( ~n2737 & n5802 ) | ( n4878 & n5802 ) ;
  assign n5804 = ( n506 & ~n3707 ) | ( n506 & n4519 ) | ( ~n3707 & n4519 ) ;
  assign n5805 = ( n2245 & n3691 ) | ( n2245 & ~n5804 ) | ( n3691 & ~n5804 ) ;
  assign n5806 = ( n1482 & n1970 ) | ( n1482 & n5755 ) | ( n1970 & n5755 ) ;
  assign n5807 = n5806 ^ n1754 ^ n1575 ;
  assign n5808 = ( n2227 & ~n5805 ) | ( n2227 & n5807 ) | ( ~n5805 & n5807 ) ;
  assign n5809 = ( n5799 & n5803 ) | ( n5799 & n5808 ) | ( n5803 & n5808 ) ;
  assign n5812 = n5811 ^ n5810 ^ n5809 ;
  assign n5813 = ~n1472 & n5041 ;
  assign n5814 = n5813 ^ n403 ^ 1'b0 ;
  assign n5815 = ( n611 & n2037 ) | ( n611 & ~n5814 ) | ( n2037 & ~n5814 ) ;
  assign n5820 = n2484 & ~n4249 ;
  assign n5819 = ( ~n1771 & n2353 ) | ( ~n1771 & n3567 ) | ( n2353 & n3567 ) ;
  assign n5816 = ( n1047 & n1302 ) | ( n1047 & ~n2600 ) | ( n1302 & ~n2600 ) ;
  assign n5817 = ( n263 & ~n2678 ) | ( n263 & n5816 ) | ( ~n2678 & n5816 ) ;
  assign n5818 = ( n4865 & ~n5288 ) | ( n4865 & n5817 ) | ( ~n5288 & n5817 ) ;
  assign n5821 = n5820 ^ n5819 ^ n5818 ;
  assign n5828 = n3983 ^ n3171 ^ n1430 ;
  assign n5825 = ( n507 & n1532 ) | ( n507 & n1931 ) | ( n1532 & n1931 ) ;
  assign n5829 = n5828 ^ n5825 ^ 1'b0 ;
  assign n5830 = n5829 ^ n3566 ^ n701 ;
  assign n5822 = ( n972 & n1565 ) | ( n972 & ~n2740 ) | ( n1565 & ~n2740 ) ;
  assign n5823 = ( ~n392 & n5411 ) | ( ~n392 & n5822 ) | ( n5411 & n5822 ) ;
  assign n5824 = n206 & n283 ;
  assign n5826 = n5825 ^ n5824 ^ 1'b0 ;
  assign n5827 = ( n225 & n5823 ) | ( n225 & ~n5826 ) | ( n5823 & ~n5826 ) ;
  assign n5831 = n5830 ^ n5827 ^ n688 ;
  assign n5832 = ( n767 & n2407 ) | ( n767 & n5831 ) | ( n2407 & n5831 ) ;
  assign n5833 = n3294 ^ n2165 ^ n1809 ;
  assign n5846 = n783 & n1427 ;
  assign n5847 = n5846 ^ n3953 ^ n3055 ;
  assign n5842 = n2958 ^ n1461 ^ 1'b0 ;
  assign n5843 = n1847 & ~n5842 ;
  assign n5841 = x20 & ~n3060 ;
  assign n5844 = n5843 ^ n5841 ^ n2309 ;
  assign n5845 = n5844 ^ n5807 ^ n1599 ;
  assign n5834 = n1931 ^ n773 ^ n729 ;
  assign n5835 = n5834 ^ n4452 ^ n232 ;
  assign n5836 = n3112 ^ n1694 ^ n812 ;
  assign n5837 = n5836 ^ n1089 ^ n387 ;
  assign n5838 = n5837 ^ n4875 ^ n1809 ;
  assign n5839 = n2094 | n5838 ;
  assign n5840 = n5835 | n5839 ;
  assign n5848 = n5847 ^ n5845 ^ n5840 ;
  assign n5849 = n2255 ^ n1162 ^ n1080 ;
  assign n5850 = ( n1739 & n3723 ) | ( n1739 & n3808 ) | ( n3723 & n3808 ) ;
  assign n5851 = n246 & n719 ;
  assign n5852 = ( n5849 & n5850 ) | ( n5849 & n5851 ) | ( n5850 & n5851 ) ;
  assign n5853 = ( n569 & ~n729 ) | ( n569 & n2388 ) | ( ~n729 & n2388 ) ;
  assign n5854 = ~n1771 & n5853 ;
  assign n5855 = n5852 & n5854 ;
  assign n5856 = n971 & n4843 ;
  assign n5857 = n5856 ^ n1180 ^ 1'b0 ;
  assign n5858 = ( n3079 & n4257 ) | ( n3079 & ~n5857 ) | ( n4257 & ~n5857 ) ;
  assign n5859 = ~n4765 & n5858 ;
  assign n5860 = n800 & n1036 ;
  assign n5861 = n5860 ^ n3537 ^ n1767 ;
  assign n5862 = n5861 ^ n4632 ^ n455 ;
  assign n5863 = ( ~n1500 & n3969 ) | ( ~n1500 & n5862 ) | ( n3969 & n5862 ) ;
  assign n5864 = ( n1534 & n3864 ) | ( n1534 & ~n4835 ) | ( n3864 & ~n4835 ) ;
  assign n5867 = n5555 ^ n2956 ^ n1848 ;
  assign n5865 = ( n2174 & ~n3056 ) | ( n2174 & n3697 ) | ( ~n3056 & n3697 ) ;
  assign n5866 = n5865 ^ n4951 ^ n1545 ;
  assign n5868 = n5867 ^ n5866 ^ n2144 ;
  assign n5869 = n3533 ^ n733 ^ n596 ;
  assign n5870 = ( n1890 & n2153 ) | ( n1890 & n3796 ) | ( n2153 & n3796 ) ;
  assign n5871 = ( ~n591 & n5869 ) | ( ~n591 & n5870 ) | ( n5869 & n5870 ) ;
  assign n5872 = n3687 ^ n2052 ^ n714 ;
  assign n5873 = n1657 ^ n1287 ^ 1'b0 ;
  assign n5874 = x68 & ~n5873 ;
  assign n5875 = ( n2617 & ~n3751 ) | ( n2617 & n4075 ) | ( ~n3751 & n4075 ) ;
  assign n5876 = n5875 ^ n5672 ^ n2585 ;
  assign n5877 = n1284 ^ n1028 ^ n669 ;
  assign n5878 = n5877 ^ n5288 ^ n431 ;
  assign n5886 = n4004 ^ n3408 ^ n154 ;
  assign n5887 = ~n3681 & n5886 ;
  assign n5879 = n1283 ^ n731 ^ x40 ;
  assign n5880 = ( n733 & ~n3748 ) | ( n733 & n5879 ) | ( ~n3748 & n5879 ) ;
  assign n5881 = n5880 ^ n1681 ^ 1'b0 ;
  assign n5882 = n5881 ^ n5835 ^ n5049 ;
  assign n5883 = ( n4009 & ~n5248 ) | ( n4009 & n5882 ) | ( ~n5248 & n5882 ) ;
  assign n5884 = ( ~n1803 & n5380 ) | ( ~n1803 & n5883 ) | ( n5380 & n5883 ) ;
  assign n5885 = ~n3500 & n5884 ;
  assign n5888 = n5887 ^ n5885 ^ n4682 ;
  assign n5889 = ( ~n1608 & n5878 ) | ( ~n1608 & n5888 ) | ( n5878 & n5888 ) ;
  assign n5895 = n5137 ^ n1915 ^ n1544 ;
  assign n5892 = n5542 ^ n3679 ^ n1351 ;
  assign n5893 = ( n351 & ~n5883 ) | ( n351 & n5892 ) | ( ~n5883 & n5892 ) ;
  assign n5894 = ( n2540 & n4850 ) | ( n2540 & n5893 ) | ( n4850 & n5893 ) ;
  assign n5896 = n5895 ^ n5894 ^ 1'b0 ;
  assign n5890 = n3798 ^ n360 ^ 1'b0 ;
  assign n5891 = ( ~n681 & n4380 ) | ( ~n681 & n5890 ) | ( n4380 & n5890 ) ;
  assign n5897 = n5896 ^ n5891 ^ n1386 ;
  assign n5898 = ( n1698 & n1848 ) | ( n1698 & n3656 ) | ( n1848 & n3656 ) ;
  assign n5899 = n5898 ^ n2396 ^ 1'b0 ;
  assign n5924 = n2885 ^ n2507 ^ n2389 ;
  assign n5922 = n1909 ^ n1423 ^ n1175 ;
  assign n5914 = n1097 ^ n628 ^ n319 ;
  assign n5911 = n2034 ^ n1932 ^ x19 ;
  assign n5912 = ( n545 & n1468 ) | ( n545 & n1820 ) | ( n1468 & n1820 ) ;
  assign n5913 = ( ~n3183 & n5911 ) | ( ~n3183 & n5912 ) | ( n5911 & n5912 ) ;
  assign n5915 = n5914 ^ n5913 ^ 1'b0 ;
  assign n5916 = n559 & ~n5915 ;
  assign n5918 = n2314 ^ n1098 ^ n968 ;
  assign n5917 = n3011 ^ n238 ^ n201 ;
  assign n5919 = n5918 ^ n5917 ^ n499 ;
  assign n5920 = ( n3581 & ~n5916 ) | ( n3581 & n5919 ) | ( ~n5916 & n5919 ) ;
  assign n5900 = ( n165 & n2785 ) | ( n165 & n3187 ) | ( n2785 & n3187 ) ;
  assign n5901 = ( ~n850 & n1125 ) | ( ~n850 & n5362 ) | ( n1125 & n5362 ) ;
  assign n5902 = ( n764 & n2807 ) | ( n764 & n5901 ) | ( n2807 & n5901 ) ;
  assign n5903 = n3894 ^ n1224 ^ n1170 ;
  assign n5904 = n2484 & n5903 ;
  assign n5905 = ( n5900 & n5902 ) | ( n5900 & n5904 ) | ( n5902 & n5904 ) ;
  assign n5906 = ( n1901 & n3582 ) | ( n1901 & n3631 ) | ( n3582 & n3631 ) ;
  assign n5907 = n2486 & ~n5906 ;
  assign n5908 = ~n5770 & n5907 ;
  assign n5909 = n5908 ^ n4056 ^ 1'b0 ;
  assign n5910 = n5905 & ~n5909 ;
  assign n5921 = n5920 ^ n5910 ^ n1594 ;
  assign n5923 = n5922 ^ n5921 ^ n3778 ;
  assign n5925 = n5924 ^ n5923 ^ 1'b0 ;
  assign n5926 = ~n4211 & n5925 ;
  assign n5927 = ( n1909 & n5899 ) | ( n1909 & ~n5926 ) | ( n5899 & ~n5926 ) ;
  assign n5928 = ( n1233 & ~n2700 ) | ( n1233 & n3530 ) | ( ~n2700 & n3530 ) ;
  assign n5929 = n1642 ^ n1000 ^ 1'b0 ;
  assign n5930 = n1671 & n5929 ;
  assign n5931 = n2938 ^ n2937 ^ n1501 ;
  assign n5932 = ( n2427 & ~n5930 ) | ( n2427 & n5931 ) | ( ~n5930 & n5931 ) ;
  assign n5933 = ( n689 & n5785 ) | ( n689 & n5932 ) | ( n5785 & n5932 ) ;
  assign n5934 = n4288 ^ n4186 ^ n680 ;
  assign n5935 = n5934 ^ n3020 ^ 1'b0 ;
  assign n5936 = n2878 ^ n1306 ^ n1128 ;
  assign n5937 = ( n1185 & n4770 ) | ( n1185 & n5936 ) | ( n4770 & n5936 ) ;
  assign n5938 = ( n5933 & n5935 ) | ( n5933 & ~n5937 ) | ( n5935 & ~n5937 ) ;
  assign n5939 = n2217 ^ n983 ^ 1'b0 ;
  assign n5940 = ( n169 & n495 ) | ( n169 & ~n5939 ) | ( n495 & ~n5939 ) ;
  assign n5941 = n5940 ^ n3254 ^ 1'b0 ;
  assign n5942 = n2179 ^ n563 ^ n241 ;
  assign n5943 = n242 & n5942 ;
  assign n5944 = ~n5941 & n5943 ;
  assign n5945 = n4141 ^ n1140 ^ n228 ;
  assign n5949 = x11 | n3213 ;
  assign n5950 = ( x83 & ~n212 ) | ( x83 & n5949 ) | ( ~n212 & n5949 ) ;
  assign n5951 = ( n1018 & ~n4385 ) | ( n1018 & n5950 ) | ( ~n4385 & n5950 ) ;
  assign n5946 = ( n2544 & n4197 ) | ( n2544 & ~n4754 ) | ( n4197 & ~n4754 ) ;
  assign n5947 = ( n980 & n3702 ) | ( n980 & ~n5946 ) | ( n3702 & ~n5946 ) ;
  assign n5948 = n5947 ^ n3908 ^ 1'b0 ;
  assign n5952 = n5951 ^ n5948 ^ 1'b0 ;
  assign n5953 = n5895 & ~n5952 ;
  assign n5954 = n5953 ^ n4634 ^ n2212 ;
  assign n5955 = ( n326 & n5945 ) | ( n326 & ~n5954 ) | ( n5945 & ~n5954 ) ;
  assign n5956 = n5454 ^ n1975 ^ n1690 ;
  assign n5962 = n2326 ^ n1090 ^ x13 ;
  assign n5957 = ( ~n260 & n370 ) | ( ~n260 & n383 ) | ( n370 & n383 ) ;
  assign n5958 = ( n759 & n1239 ) | ( n759 & ~n5957 ) | ( n1239 & ~n5957 ) ;
  assign n5959 = ( n190 & n1502 ) | ( n190 & ~n2853 ) | ( n1502 & ~n2853 ) ;
  assign n5960 = ( n1930 & n5958 ) | ( n1930 & ~n5959 ) | ( n5958 & ~n5959 ) ;
  assign n5961 = ( n762 & n5486 ) | ( n762 & n5960 ) | ( n5486 & n5960 ) ;
  assign n5963 = n5962 ^ n5961 ^ n2732 ;
  assign n5965 = n3759 ^ n1995 ^ n1712 ;
  assign n5966 = ( n2169 & ~n5826 ) | ( n2169 & n5965 ) | ( ~n5826 & n5965 ) ;
  assign n5964 = ~n4862 & n4875 ;
  assign n5967 = n5966 ^ n5964 ^ 1'b0 ;
  assign n5972 = n4399 ^ n4022 ^ 1'b0 ;
  assign n5968 = ~n493 & n740 ;
  assign n5969 = n354 & n5968 ;
  assign n5970 = ( n1854 & n2587 ) | ( n1854 & n5969 ) | ( n2587 & n5969 ) ;
  assign n5971 = ~n261 & n5970 ;
  assign n5973 = n5972 ^ n5971 ^ n2286 ;
  assign n5974 = n1649 ^ n214 ^ x27 ;
  assign n5975 = ( n2613 & ~n4391 ) | ( n2613 & n5974 ) | ( ~n4391 & n5974 ) ;
  assign n5976 = n5326 ^ n1289 ^ n474 ;
  assign n5977 = n1531 ^ n1467 ^ n215 ;
  assign n5978 = ( n924 & n5976 ) | ( n924 & ~n5977 ) | ( n5976 & ~n5977 ) ;
  assign n5979 = ( ~n1708 & n2782 ) | ( ~n1708 & n4388 ) | ( n2782 & n4388 ) ;
  assign n5980 = ( n180 & n655 ) | ( n180 & ~n2777 ) | ( n655 & ~n2777 ) ;
  assign n5981 = n5980 ^ n1881 ^ n733 ;
  assign n5983 = n4846 ^ n4249 ^ n2309 ;
  assign n5982 = ( n966 & ~n1660 ) | ( n966 & n4819 ) | ( ~n1660 & n4819 ) ;
  assign n5984 = n5983 ^ n5982 ^ n5628 ;
  assign n5985 = ( n2015 & n2779 ) | ( n2015 & ~n3162 ) | ( n2779 & ~n3162 ) ;
  assign n5986 = n5985 ^ n3622 ^ 1'b0 ;
  assign n5987 = n5986 ^ n3697 ^ n3532 ;
  assign n5990 = n5403 ^ n1366 ^ n705 ;
  assign n5991 = ( ~n1932 & n2023 ) | ( ~n1932 & n5990 ) | ( n2023 & n5990 ) ;
  assign n5988 = ~n800 & n2607 ;
  assign n5989 = n5988 ^ n1978 ^ 1'b0 ;
  assign n5992 = n5991 ^ n5989 ^ n2168 ;
  assign n5993 = n5992 ^ n2967 ^ n199 ;
  assign n5994 = ( n1838 & ~n5607 ) | ( n1838 & n5993 ) | ( ~n5607 & n5993 ) ;
  assign n5995 = n3712 & ~n5588 ;
  assign n5996 = n5994 & n5995 ;
  assign n6008 = ( ~n305 & n414 ) | ( ~n305 & n981 ) | ( n414 & n981 ) ;
  assign n5997 = ( n848 & ~n967 ) | ( n848 & n3547 ) | ( ~n967 & n3547 ) ;
  assign n5998 = n3601 ^ n2000 ^ n887 ;
  assign n5999 = n5997 & ~n5998 ;
  assign n6000 = n4229 ^ n145 ^ 1'b0 ;
  assign n6001 = ~n5999 & n6000 ;
  assign n6002 = ( n814 & n1026 ) | ( n814 & ~n2807 ) | ( n1026 & ~n2807 ) ;
  assign n6003 = n5370 ^ n874 ^ 1'b0 ;
  assign n6004 = ~n1380 & n6003 ;
  assign n6005 = ( n2671 & n6002 ) | ( n2671 & ~n6004 ) | ( n6002 & ~n6004 ) ;
  assign n6006 = n6005 ^ n3786 ^ 1'b0 ;
  assign n6007 = ( n1533 & n6001 ) | ( n1533 & ~n6006 ) | ( n6001 & ~n6006 ) ;
  assign n6009 = n6008 ^ n6007 ^ n4665 ;
  assign n6011 = ( n1262 & ~n3582 ) | ( n1262 & n4775 ) | ( ~n3582 & n4775 ) ;
  assign n6012 = n2897 ^ n1738 ^ n989 ;
  assign n6013 = n4944 & n6012 ;
  assign n6014 = ~n6011 & n6013 ;
  assign n6010 = n5154 ^ n2617 ^ n604 ;
  assign n6015 = n6014 ^ n6010 ^ n1427 ;
  assign n6016 = n3158 ^ n206 ^ 1'b0 ;
  assign n6017 = ( n2390 & n4100 ) | ( n2390 & n6016 ) | ( n4100 & n6016 ) ;
  assign n6020 = n5411 ^ n2193 ^ 1'b0 ;
  assign n6018 = n3456 | n5746 ;
  assign n6019 = n6018 ^ n780 ^ 1'b0 ;
  assign n6021 = n6020 ^ n6019 ^ n1863 ;
  assign n6022 = ~n2676 & n6021 ;
  assign n6023 = n5444 ^ n2615 ^ n1254 ;
  assign n6024 = ( n1895 & ~n6022 ) | ( n1895 & n6023 ) | ( ~n6022 & n6023 ) ;
  assign n6027 = n2550 ^ n2473 ^ n977 ;
  assign n6028 = ( n167 & n1329 ) | ( n167 & n6027 ) | ( n1329 & n6027 ) ;
  assign n6029 = ( n1172 & ~n3828 ) | ( n1172 & n6028 ) | ( ~n3828 & n6028 ) ;
  assign n6025 = n2331 & n5568 ;
  assign n6026 = n6025 ^ n1554 ^ 1'b0 ;
  assign n6030 = n6029 ^ n6026 ^ n2868 ;
  assign n6031 = n850 ^ n351 ^ 1'b0 ;
  assign n6032 = n6031 ^ n5405 ^ n676 ;
  assign n6033 = n6032 ^ n1685 ^ n1270 ;
  assign n6034 = n1525 ^ n357 ^ n328 ;
  assign n6035 = n2437 ^ n2387 ^ n1816 ;
  assign n6036 = ( ~n2378 & n6034 ) | ( ~n2378 & n6035 ) | ( n6034 & n6035 ) ;
  assign n6037 = n4781 ^ n4495 ^ n2138 ;
  assign n6038 = ( n1818 & n6036 ) | ( n1818 & ~n6037 ) | ( n6036 & ~n6037 ) ;
  assign n6041 = ( n307 & n704 ) | ( n307 & ~n3535 ) | ( n704 & ~n3535 ) ;
  assign n6042 = ( n596 & n1322 ) | ( n596 & n6041 ) | ( n1322 & n6041 ) ;
  assign n6039 = n2948 ^ n1843 ^ n1426 ;
  assign n6040 = n6039 ^ n3022 ^ n2241 ;
  assign n6043 = n6042 ^ n6040 ^ n566 ;
  assign n6044 = n1587 ^ n918 ^ 1'b0 ;
  assign n6045 = n6044 ^ n4039 ^ n1337 ;
  assign n6048 = ( n825 & ~n1558 ) | ( n825 & n1574 ) | ( ~n1558 & n1574 ) ;
  assign n6049 = ( ~n725 & n1511 ) | ( ~n725 & n4396 ) | ( n1511 & n4396 ) ;
  assign n6050 = ( n5671 & n6048 ) | ( n5671 & n6049 ) | ( n6048 & n6049 ) ;
  assign n6046 = n3907 | n4745 ;
  assign n6047 = n6046 ^ n495 ^ 1'b0 ;
  assign n6051 = n6050 ^ n6047 ^ n582 ;
  assign n6052 = n6051 ^ n1747 ^ 1'b0 ;
  assign n6053 = ~n6045 & n6052 ;
  assign n6055 = ( n1023 & n1311 ) | ( n1023 & n1466 ) | ( n1311 & n1466 ) ;
  assign n6056 = ( n1425 & ~n1480 ) | ( n1425 & n6055 ) | ( ~n1480 & n6055 ) ;
  assign n6057 = n6056 ^ n1752 ^ x10 ;
  assign n6054 = n3293 ^ n876 ^ 1'b0 ;
  assign n6058 = n6057 ^ n6054 ^ 1'b0 ;
  assign n6059 = ~n1004 & n6058 ;
  assign n6060 = n6059 ^ n2848 ^ n569 ;
  assign n6061 = n6060 ^ n4475 ^ n2881 ;
  assign n6062 = n6061 ^ n2344 ^ n2164 ;
  assign n6067 = n685 & n3547 ;
  assign n6068 = n5791 & n6067 ;
  assign n6069 = n6068 ^ n4771 ^ 1'b0 ;
  assign n6070 = ( ~n291 & n5700 ) | ( ~n291 & n6069 ) | ( n5700 & n6069 ) ;
  assign n6063 = n1636 & n2156 ;
  assign n6064 = n6063 ^ n462 ^ 1'b0 ;
  assign n6065 = n6064 ^ n2218 ^ n1713 ;
  assign n6066 = n6065 ^ n2526 ^ n1521 ;
  assign n6071 = n6070 ^ n6066 ^ n2649 ;
  assign n6072 = n5098 ^ n4501 ^ n2374 ;
  assign n6073 = n6072 ^ n3763 ^ n1477 ;
  assign n6074 = n6073 ^ n879 ^ 1'b0 ;
  assign n6075 = n5682 ^ n4793 ^ 1'b0 ;
  assign n6077 = ( n906 & n1892 ) | ( n906 & ~n3707 ) | ( n1892 & ~n3707 ) ;
  assign n6076 = ( x46 & n1252 ) | ( x46 & n2160 ) | ( n1252 & n2160 ) ;
  assign n6078 = n6077 ^ n6076 ^ x30 ;
  assign n6079 = ( n3362 & n5189 ) | ( n3362 & ~n6078 ) | ( n5189 & ~n6078 ) ;
  assign n6080 = n2607 & n6079 ;
  assign n6081 = n6080 ^ n1167 ^ 1'b0 ;
  assign n6082 = n6075 | n6081 ;
  assign n6083 = n5070 ^ n2075 ^ 1'b0 ;
  assign n6084 = n2471 & ~n6083 ;
  assign n6085 = n6084 ^ n4594 ^ 1'b0 ;
  assign n6086 = n2721 ^ n1541 ^ n774 ;
  assign n6087 = ( ~n2471 & n2992 ) | ( ~n2471 & n6086 ) | ( n2992 & n6086 ) ;
  assign n6088 = n1630 ^ n638 ^ n602 ;
  assign n6089 = n5836 ^ n1628 ^ n634 ;
  assign n6090 = ( n697 & n1616 ) | ( n697 & n1723 ) | ( n1616 & n1723 ) ;
  assign n6091 = ( n5827 & ~n6089 ) | ( n5827 & n6090 ) | ( ~n6089 & n6090 ) ;
  assign n6093 = ( ~n2194 & n2566 ) | ( ~n2194 & n3654 ) | ( n2566 & n3654 ) ;
  assign n6094 = n6093 ^ n5835 ^ n2761 ;
  assign n6092 = n4014 ^ n2390 ^ n133 ;
  assign n6095 = n6094 ^ n6092 ^ n238 ;
  assign n6096 = ( n6088 & n6091 ) | ( n6088 & n6095 ) | ( n6091 & n6095 ) ;
  assign n6097 = n6096 ^ n3164 ^ n2186 ;
  assign n6098 = n2471 ^ n1275 ^ n647 ;
  assign n6099 = n6098 ^ n6094 ^ n3124 ;
  assign n6100 = ( ~n1580 & n6002 ) | ( ~n1580 & n6099 ) | ( n6002 & n6099 ) ;
  assign n6101 = n5808 ^ n3807 ^ 1'b0 ;
  assign n6102 = ~n6100 & n6101 ;
  assign n6109 = n493 | n1562 ;
  assign n6106 = n5774 ^ n3049 ^ 1'b0 ;
  assign n6104 = n3520 ^ n2286 ^ n678 ;
  assign n6105 = ( x113 & n2570 ) | ( x113 & n6104 ) | ( n2570 & n6104 ) ;
  assign n6107 = n6106 ^ n6105 ^ n2569 ;
  assign n6108 = n6107 ^ n1909 ^ n1345 ;
  assign n6103 = n5562 ^ n1857 ^ 1'b0 ;
  assign n6110 = n6109 ^ n6108 ^ n6103 ;
  assign n6111 = n4420 ^ n2932 ^ n956 ;
  assign n6112 = ( n993 & n3401 ) | ( n993 & ~n6111 ) | ( n3401 & ~n6111 ) ;
  assign n6121 = n4302 ^ n1798 ^ 1'b0 ;
  assign n6122 = n6121 ^ n4228 ^ n2676 ;
  assign n6114 = n3740 ^ n1120 ^ n341 ;
  assign n6115 = ( n1940 & ~n4907 ) | ( n1940 & n6114 ) | ( ~n4907 & n6114 ) ;
  assign n6116 = n6115 ^ n5083 ^ x71 ;
  assign n6117 = n3291 & n6116 ;
  assign n6118 = n2157 & n6117 ;
  assign n6113 = n530 & n2280 ;
  assign n6119 = n6118 ^ n6113 ^ 1'b0 ;
  assign n6120 = ( n1841 & ~n4199 ) | ( n1841 & n6119 ) | ( ~n4199 & n6119 ) ;
  assign n6123 = n6122 ^ n6120 ^ n1533 ;
  assign n6124 = ( n3237 & ~n6112 ) | ( n3237 & n6123 ) | ( ~n6112 & n6123 ) ;
  assign n6125 = ( ~n317 & n514 ) | ( ~n317 & n5723 ) | ( n514 & n5723 ) ;
  assign n6126 = ( n2426 & ~n2505 ) | ( n2426 & n2987 ) | ( ~n2505 & n2987 ) ;
  assign n6127 = ( n1074 & n2005 ) | ( n1074 & ~n3287 ) | ( n2005 & ~n3287 ) ;
  assign n6128 = n6127 ^ n3167 ^ 1'b0 ;
  assign n6129 = n6126 | n6128 ;
  assign n6130 = ( n1901 & n4041 ) | ( n1901 & n6129 ) | ( n4041 & n6129 ) ;
  assign n6131 = n4706 ^ n3882 ^ 1'b0 ;
  assign n6132 = ~n6130 & n6131 ;
  assign n6133 = ( n2875 & ~n6125 ) | ( n2875 & n6132 ) | ( ~n6125 & n6132 ) ;
  assign n6134 = n6133 ^ n4087 ^ n3571 ;
  assign n6139 = n2970 ^ n1981 ^ n440 ;
  assign n6135 = ( x33 & ~n1095 ) | ( x33 & n2034 ) | ( ~n1095 & n2034 ) ;
  assign n6136 = ( ~n565 & n758 ) | ( ~n565 & n6135 ) | ( n758 & n6135 ) ;
  assign n6137 = ( n3339 & n5836 ) | ( n3339 & n6136 ) | ( n5836 & n6136 ) ;
  assign n6138 = n6137 ^ n5042 ^ n1714 ;
  assign n6140 = n6139 ^ n6138 ^ 1'b0 ;
  assign n6141 = n5287 ^ n859 ^ 1'b0 ;
  assign n6142 = n4003 & n6141 ;
  assign n6143 = n933 | n6142 ;
  assign n6144 = n6143 ^ n3204 ^ n905 ;
  assign n6145 = n2451 ^ n1981 ^ 1'b0 ;
  assign n6146 = n6145 ^ n5119 ^ n1682 ;
  assign n6147 = n6146 ^ n2932 ^ 1'b0 ;
  assign n6148 = n3673 & ~n6147 ;
  assign n6149 = ( n164 & n910 ) | ( n164 & n913 ) | ( n910 & n913 ) ;
  assign n6150 = n6149 ^ n2086 ^ n1057 ;
  assign n6151 = ( x101 & n1816 ) | ( x101 & ~n4572 ) | ( n1816 & ~n4572 ) ;
  assign n6157 = n1803 ^ x33 ^ 1'b0 ;
  assign n6158 = n2938 ^ n2653 ^ n2147 ;
  assign n6159 = ( ~n616 & n6157 ) | ( ~n616 & n6158 ) | ( n6157 & n6158 ) ;
  assign n6153 = n3644 ^ n2141 ^ n551 ;
  assign n6152 = ( ~x22 & n1167 ) | ( ~x22 & n1650 ) | ( n1167 & n1650 ) ;
  assign n6154 = n6153 ^ n6152 ^ 1'b0 ;
  assign n6155 = n6154 ^ n2055 ^ x32 ;
  assign n6156 = n1041 & ~n6155 ;
  assign n6160 = n6159 ^ n6156 ^ 1'b0 ;
  assign n6161 = n3374 ^ n491 ^ 1'b0 ;
  assign n6162 = n3869 & ~n6161 ;
  assign n6163 = n691 ^ n601 ^ x37 ;
  assign n6164 = n6163 ^ n3827 ^ n1406 ;
  assign n6165 = ( ~n131 & n6162 ) | ( ~n131 & n6164 ) | ( n6162 & n6164 ) ;
  assign n6166 = ( n1809 & n6160 ) | ( n1809 & n6165 ) | ( n6160 & n6165 ) ;
  assign n6167 = ( ~n1928 & n4231 ) | ( ~n1928 & n6166 ) | ( n4231 & n6166 ) ;
  assign n6168 = ( x12 & n1434 ) | ( x12 & n5355 ) | ( n1434 & n5355 ) ;
  assign n6169 = n6168 ^ n5432 ^ n4750 ;
  assign n6170 = ( n383 & n1065 ) | ( n383 & ~n5304 ) | ( n1065 & ~n5304 ) ;
  assign n6171 = n2556 ^ x50 ^ 1'b0 ;
  assign n6172 = ( n6169 & ~n6170 ) | ( n6169 & n6171 ) | ( ~n6170 & n6171 ) ;
  assign n6173 = n4360 | n6172 ;
  assign n6174 = ( n5269 & n6012 ) | ( n5269 & ~n6173 ) | ( n6012 & ~n6173 ) ;
  assign n6175 = n6174 ^ n5664 ^ n5136 ;
  assign n6184 = n706 ^ x32 ^ 1'b0 ;
  assign n6185 = ( n2736 & n4013 ) | ( n2736 & ~n6184 ) | ( n4013 & ~n6184 ) ;
  assign n6183 = n2035 ^ n1043 ^ n822 ;
  assign n6181 = n2925 ^ n1637 ^ n1561 ;
  assign n6179 = n5098 ^ n2112 ^ n1239 ;
  assign n6180 = ( n354 & n5348 ) | ( n354 & ~n6179 ) | ( n5348 & ~n6179 ) ;
  assign n6177 = ( ~n352 & n658 ) | ( ~n352 & n1030 ) | ( n658 & n1030 ) ;
  assign n6176 = ~n4113 & n4635 ;
  assign n6178 = n6177 ^ n6176 ^ n603 ;
  assign n6182 = n6181 ^ n6180 ^ n6178 ;
  assign n6186 = n6185 ^ n6183 ^ n6182 ;
  assign n6188 = ( ~n811 & n2172 ) | ( ~n811 & n2442 ) | ( n2172 & n2442 ) ;
  assign n6189 = ( n1417 & ~n4558 ) | ( n1417 & n6188 ) | ( ~n4558 & n6188 ) ;
  assign n6187 = n647 & n5459 ;
  assign n6190 = n6189 ^ n6187 ^ 1'b0 ;
  assign n6191 = n1728 | n1818 ;
  assign n6192 = n3378 ^ n2816 ^ n1614 ;
  assign n6193 = ( n3094 & n4801 ) | ( n3094 & n6192 ) | ( n4801 & n6192 ) ;
  assign n6194 = n6193 ^ n5969 ^ n5083 ;
  assign n6195 = n6194 ^ n4251 ^ n2114 ;
  assign n6196 = ( n5118 & ~n6014 ) | ( n5118 & n6032 ) | ( ~n6014 & n6032 ) ;
  assign n6197 = n495 & ~n3716 ;
  assign n6201 = n3090 ^ n992 ^ x122 ;
  assign n6198 = n198 & ~n5739 ;
  assign n6199 = n6198 ^ n5180 ^ 1'b0 ;
  assign n6200 = n6199 ^ n5784 ^ n2851 ;
  assign n6202 = n6201 ^ n6200 ^ n4283 ;
  assign n6203 = ( n3778 & n6197 ) | ( n3778 & ~n6202 ) | ( n6197 & ~n6202 ) ;
  assign n6205 = ( ~n227 & n2479 ) | ( ~n227 & n2853 ) | ( n2479 & n2853 ) ;
  assign n6206 = ( n1822 & n2204 ) | ( n1822 & ~n6205 ) | ( n2204 & ~n6205 ) ;
  assign n6204 = ( n4895 & n5186 ) | ( n4895 & n5983 ) | ( n5186 & n5983 ) ;
  assign n6207 = n6206 ^ n6204 ^ n5503 ;
  assign n6208 = n4492 ^ n2842 ^ n1806 ;
  assign n6209 = ( n300 & ~n3548 ) | ( n300 & n6208 ) | ( ~n3548 & n6208 ) ;
  assign n6210 = n3141 ^ n1490 ^ n1067 ;
  assign n6211 = ( ~n332 & n4231 ) | ( ~n332 & n6210 ) | ( n4231 & n6210 ) ;
  assign n6212 = n6211 ^ n4045 ^ 1'b0 ;
  assign n6213 = n6212 ^ n3808 ^ n2352 ;
  assign n6216 = n1863 & n2999 ;
  assign n6217 = ( n1252 & n4156 ) | ( n1252 & ~n6216 ) | ( n4156 & ~n6216 ) ;
  assign n6218 = n3524 ^ n642 ^ 1'b0 ;
  assign n6219 = n6217 | n6218 ;
  assign n6220 = ( ~n1563 & n3033 ) | ( ~n1563 & n6219 ) | ( n3033 & n6219 ) ;
  assign n6221 = ( n1447 & n3354 ) | ( n1447 & n6220 ) | ( n3354 & n6220 ) ;
  assign n6214 = ( n699 & ~n1120 ) | ( n699 & n4110 ) | ( ~n1120 & n4110 ) ;
  assign n6215 = ( n920 & n3215 ) | ( n920 & ~n6214 ) | ( n3215 & ~n6214 ) ;
  assign n6222 = n6221 ^ n6215 ^ n4138 ;
  assign n6223 = ( n3499 & ~n4105 ) | ( n3499 & n6222 ) | ( ~n4105 & n6222 ) ;
  assign n6224 = ( n780 & n6213 ) | ( n780 & ~n6223 ) | ( n6213 & ~n6223 ) ;
  assign n6225 = ( n4562 & n6209 ) | ( n4562 & n6224 ) | ( n6209 & n6224 ) ;
  assign n6239 = ~n1430 & n2373 ;
  assign n6230 = n4203 ^ n3971 ^ n1676 ;
  assign n6231 = n5463 ^ n734 ^ 1'b0 ;
  assign n6232 = n1105 | n3144 ;
  assign n6233 = n836 | n6232 ;
  assign n6234 = ( ~n529 & n2993 ) | ( ~n529 & n6233 ) | ( n2993 & n6233 ) ;
  assign n6235 = ( n1529 & n2109 ) | ( n1529 & n6234 ) | ( n2109 & n6234 ) ;
  assign n6236 = ( n6230 & ~n6231 ) | ( n6230 & n6235 ) | ( ~n6231 & n6235 ) ;
  assign n6226 = n274 | n4617 ;
  assign n6227 = n220 | n6226 ;
  assign n6228 = ( n761 & n1795 ) | ( n761 & ~n5110 ) | ( n1795 & ~n5110 ) ;
  assign n6229 = ( ~n3953 & n6227 ) | ( ~n3953 & n6228 ) | ( n6227 & n6228 ) ;
  assign n6237 = n6236 ^ n6229 ^ n640 ;
  assign n6238 = ( ~n4192 & n5517 ) | ( ~n4192 & n6237 ) | ( n5517 & n6237 ) ;
  assign n6240 = n6239 ^ n6238 ^ n1915 ;
  assign n6241 = n5755 ^ n4641 ^ n1643 ;
  assign n6243 = ( n1195 & n2045 ) | ( n1195 & n4044 ) | ( n2045 & n4044 ) ;
  assign n6242 = ( n991 & ~n1719 ) | ( n991 & n3584 ) | ( ~n1719 & n3584 ) ;
  assign n6244 = n6243 ^ n6242 ^ n793 ;
  assign n6245 = n4437 ^ n2322 ^ n753 ;
  assign n6246 = ( n6241 & ~n6244 ) | ( n6241 & n6245 ) | ( ~n6244 & n6245 ) ;
  assign n6249 = n2452 ^ n1397 ^ n1034 ;
  assign n6250 = n2443 ^ x9 ^ 1'b0 ;
  assign n6251 = n6249 & ~n6250 ;
  assign n6247 = n5746 ^ n4549 ^ x70 ;
  assign n6248 = n4385 & n6247 ;
  assign n6252 = n6251 ^ n6248 ^ 1'b0 ;
  assign n6253 = ~n1457 & n6252 ;
  assign n6254 = ~n2686 & n2744 ;
  assign n6255 = n6254 ^ n1098 ^ 1'b0 ;
  assign n6256 = ~n758 & n1670 ;
  assign n6257 = n4173 ^ n3466 ^ n1672 ;
  assign n6258 = n6257 ^ n4808 ^ n4086 ;
  assign n6259 = ( n188 & ~n6256 ) | ( n188 & n6258 ) | ( ~n6256 & n6258 ) ;
  assign n6260 = ( n1108 & ~n6255 ) | ( n1108 & n6259 ) | ( ~n6255 & n6259 ) ;
  assign n6261 = n6260 ^ n543 ^ 1'b0 ;
  assign n6262 = ~n6253 & n6261 ;
  assign n6263 = ~n498 & n2164 ;
  assign n6264 = n2391 & ~n6263 ;
  assign n6265 = n6264 ^ n4769 ^ 1'b0 ;
  assign n6266 = ( n3120 & n5682 ) | ( n3120 & n6265 ) | ( n5682 & n6265 ) ;
  assign n6279 = n3454 | n4163 ;
  assign n6267 = ( x102 & n3150 ) | ( x102 & ~n4577 ) | ( n3150 & ~n4577 ) ;
  assign n6268 = n6267 ^ n4651 ^ n2784 ;
  assign n6269 = n6268 ^ n2203 ^ 1'b0 ;
  assign n6271 = ( n1452 & ~n1965 ) | ( n1452 & n6251 ) | ( ~n1965 & n6251 ) ;
  assign n6272 = ( n1355 & n4871 ) | ( n1355 & ~n6271 ) | ( n4871 & ~n6271 ) ;
  assign n6273 = n4434 | n6272 ;
  assign n6270 = n4207 ^ n1430 ^ n1421 ;
  assign n6274 = n6273 ^ n6270 ^ n5750 ;
  assign n6275 = n2149 & n3961 ;
  assign n6276 = n3840 ^ n1578 ^ x95 ;
  assign n6277 = ( n2608 & n6275 ) | ( n2608 & ~n6276 ) | ( n6275 & ~n6276 ) ;
  assign n6278 = ( n6269 & ~n6274 ) | ( n6269 & n6277 ) | ( ~n6274 & n6277 ) ;
  assign n6280 = n6279 ^ n6278 ^ n1446 ;
  assign n6281 = ~n2123 & n6280 ;
  assign n6282 = n2239 ^ n1342 ^ 1'b0 ;
  assign n6283 = ( ~x31 & n863 ) | ( ~x31 & n2897 ) | ( n863 & n2897 ) ;
  assign n6284 = ( ~n1908 & n6282 ) | ( ~n1908 & n6283 ) | ( n6282 & n6283 ) ;
  assign n6285 = ( ~x90 & n3372 ) | ( ~x90 & n6284 ) | ( n3372 & n6284 ) ;
  assign n6286 = ( n408 & n3236 ) | ( n408 & ~n6285 ) | ( n3236 & ~n6285 ) ;
  assign n6287 = ( ~n174 & n439 ) | ( ~n174 & n5076 ) | ( n439 & n5076 ) ;
  assign n6288 = ( n3517 & n4451 ) | ( n3517 & ~n6287 ) | ( n4451 & ~n6287 ) ;
  assign n6289 = n6288 ^ n3414 ^ n3406 ;
  assign n6290 = ( n881 & ~n4727 ) | ( n881 & n5197 ) | ( ~n4727 & n5197 ) ;
  assign n6291 = n6290 ^ n6078 ^ 1'b0 ;
  assign n6292 = n6289 & n6291 ;
  assign n6293 = n3660 & n6292 ;
  assign n6294 = n6293 ^ n3371 ^ 1'b0 ;
  assign n6295 = n6286 & ~n6294 ;
  assign n6318 = n5007 ^ n3962 ^ n848 ;
  assign n6313 = n1369 & n2260 ;
  assign n6314 = n3547 ^ n2073 ^ n227 ;
  assign n6315 = n6314 ^ n1999 ^ n1461 ;
  assign n6316 = ( ~n6044 & n6313 ) | ( ~n6044 & n6315 ) | ( n6313 & n6315 ) ;
  assign n6317 = ( n1907 & n5865 ) | ( n1907 & n6316 ) | ( n5865 & n6316 ) ;
  assign n6310 = ( n1012 & n1323 ) | ( n1012 & ~n5645 ) | ( n1323 & ~n5645 ) ;
  assign n6311 = ( n3275 & ~n5318 ) | ( n3275 & n6310 ) | ( ~n5318 & n6310 ) ;
  assign n6309 = n5046 ^ n4875 ^ x104 ;
  assign n6306 = n692 | n1881 ;
  assign n6307 = n2166 | n6306 ;
  assign n6298 = ~n700 & n1422 ;
  assign n6299 = n1782 & n6298 ;
  assign n6300 = n6299 ^ n3197 ^ n1482 ;
  assign n6301 = n1737 ^ n1580 ^ n1479 ;
  assign n6302 = n6301 ^ n457 ^ x19 ;
  assign n6303 = n3581 ^ n1642 ^ 1'b0 ;
  assign n6304 = n6302 & ~n6303 ;
  assign n6305 = ( n2763 & n6300 ) | ( n2763 & n6304 ) | ( n6300 & n6304 ) ;
  assign n6296 = ( n1852 & n5120 ) | ( n1852 & n5912 ) | ( n5120 & n5912 ) ;
  assign n6297 = n6296 ^ n3723 ^ n1906 ;
  assign n6308 = n6307 ^ n6305 ^ n6297 ;
  assign n6312 = n6311 ^ n6309 ^ n6308 ;
  assign n6319 = n6318 ^ n6317 ^ n6312 ;
  assign n6320 = n3841 ^ n604 ^ n295 ;
  assign n6321 = ~n4688 & n6320 ;
  assign n6326 = n5167 ^ n637 ^ n189 ;
  assign n6322 = ( ~n1334 & n2575 ) | ( ~n1334 & n3550 ) | ( n2575 & n3550 ) ;
  assign n6323 = ( n1224 & ~n1358 ) | ( n1224 & n6322 ) | ( ~n1358 & n6322 ) ;
  assign n6324 = n6323 ^ n4411 ^ n707 ;
  assign n6325 = n6324 ^ n3735 ^ n1162 ;
  assign n6327 = n6326 ^ n6325 ^ n4234 ;
  assign n6328 = ( n539 & n853 ) | ( n539 & ~n3386 ) | ( n853 & ~n3386 ) ;
  assign n6329 = ~n5553 & n6328 ;
  assign n6330 = n1348 | n2705 ;
  assign n6331 = n6330 ^ n4343 ^ n2544 ;
  assign n6332 = ( n4155 & n4769 ) | ( n4155 & n6331 ) | ( n4769 & n6331 ) ;
  assign n6333 = n6332 ^ n2662 ^ 1'b0 ;
  assign n6334 = ( n222 & n6329 ) | ( n222 & n6333 ) | ( n6329 & n6333 ) ;
  assign n6338 = ( ~n1181 & n1435 ) | ( ~n1181 & n2195 ) | ( n1435 & n2195 ) ;
  assign n6339 = ( n3113 & n6255 ) | ( n3113 & n6338 ) | ( n6255 & n6338 ) ;
  assign n6335 = ( n463 & ~n2697 ) | ( n463 & n4868 ) | ( ~n2697 & n4868 ) ;
  assign n6336 = n6335 ^ n4695 ^ n4113 ;
  assign n6337 = n3758 & ~n6336 ;
  assign n6340 = n6339 ^ n6337 ^ 1'b0 ;
  assign n6341 = n2447 & n4953 ;
  assign n6342 = n6341 ^ n2039 ^ 1'b0 ;
  assign n6343 = n6342 ^ n3532 ^ n1584 ;
  assign n6344 = ( n2835 & ~n6302 ) | ( n2835 & n6343 ) | ( ~n6302 & n6343 ) ;
  assign n6345 = ( n1334 & ~n6340 ) | ( n1334 & n6344 ) | ( ~n6340 & n6344 ) ;
  assign n6346 = n6311 ^ n5102 ^ n4958 ;
  assign n6347 = n6346 ^ n1269 ^ n668 ;
  assign n6348 = ( n1447 & n4649 ) | ( n1447 & n6347 ) | ( n4649 & n6347 ) ;
  assign n6349 = n6348 ^ n2278 ^ n1503 ;
  assign n6350 = n342 & ~n617 ;
  assign n6351 = n6350 ^ n785 ^ 1'b0 ;
  assign n6352 = ~n1157 & n6351 ;
  assign n6353 = n6352 ^ n6110 ^ n4201 ;
  assign n6354 = n6002 ^ n2142 ^ 1'b0 ;
  assign n6355 = n6354 ^ n3936 ^ 1'b0 ;
  assign n6356 = n4586 ^ n3782 ^ n270 ;
  assign n6357 = n4556 ^ n3925 ^ x89 ;
  assign n6358 = ( n2050 & n4187 ) | ( n2050 & n6357 ) | ( n4187 & n6357 ) ;
  assign n6359 = n6087 ^ n4289 ^ 1'b0 ;
  assign n6360 = n6358 & ~n6359 ;
  assign n6361 = ( ~n1371 & n3235 ) | ( ~n1371 & n4025 ) | ( n3235 & n4025 ) ;
  assign n6362 = ( n1039 & n1709 ) | ( n1039 & ~n6361 ) | ( n1709 & ~n6361 ) ;
  assign n6363 = ( ~n1461 & n6229 ) | ( ~n1461 & n6362 ) | ( n6229 & n6362 ) ;
  assign n6364 = ( x20 & n753 ) | ( x20 & n3835 ) | ( n753 & n3835 ) ;
  assign n6365 = ( n2797 & n3479 ) | ( n2797 & ~n6227 ) | ( n3479 & ~n6227 ) ;
  assign n6366 = n6365 ^ n2286 ^ 1'b0 ;
  assign n6367 = ( ~n4469 & n6364 ) | ( ~n4469 & n6366 ) | ( n6364 & n6366 ) ;
  assign n6368 = n6367 ^ n5211 ^ n1939 ;
  assign n6370 = ( n1080 & n3600 ) | ( n1080 & n5088 ) | ( n3600 & n5088 ) ;
  assign n6371 = n4929 | n6370 ;
  assign n6372 = n2038 & ~n6371 ;
  assign n6369 = ( x25 & ~n1049 ) | ( x25 & n1400 ) | ( ~n1049 & n1400 ) ;
  assign n6373 = n6372 ^ n6369 ^ n1491 ;
  assign n6374 = ~n305 & n2646 ;
  assign n6375 = ~n6373 & n6374 ;
  assign n6376 = n6375 ^ n901 ^ 1'b0 ;
  assign n6377 = n3931 ^ n1209 ^ 1'b0 ;
  assign n6378 = ~n2406 & n6377 ;
  assign n6379 = n6378 ^ n2197 ^ n255 ;
  assign n6380 = n5675 ^ n4184 ^ x102 ;
  assign n6381 = n206 & ~n1929 ;
  assign n6382 = n4674 & n6381 ;
  assign n6383 = ( n1796 & n4002 ) | ( n1796 & n6008 ) | ( n4002 & n6008 ) ;
  assign n6384 = n6383 ^ n6029 ^ n2073 ;
  assign n6385 = n6384 ^ n5551 ^ n3794 ;
  assign n6386 = ( ~n1371 & n2241 ) | ( ~n1371 & n5258 ) | ( n2241 & n5258 ) ;
  assign n6387 = n5785 ^ n5684 ^ n2542 ;
  assign n6388 = ( n2110 & n6386 ) | ( n2110 & ~n6387 ) | ( n6386 & ~n6387 ) ;
  assign n6389 = ( n4334 & n5088 ) | ( n4334 & n6388 ) | ( n5088 & n6388 ) ;
  assign n6390 = ~n137 & n745 ;
  assign n6391 = n2047 ^ n1429 ^ n614 ;
  assign n6392 = ( n2288 & n4888 ) | ( n2288 & ~n6391 ) | ( n4888 & ~n6391 ) ;
  assign n6393 = n3740 ^ n3544 ^ n2067 ;
  assign n6394 = ( n3264 & n4233 ) | ( n3264 & ~n6393 ) | ( n4233 & ~n6393 ) ;
  assign n6395 = ( x7 & ~n1617 ) | ( x7 & n6394 ) | ( ~n1617 & n6394 ) ;
  assign n6396 = ( ~n5785 & n6392 ) | ( ~n5785 & n6395 ) | ( n6392 & n6395 ) ;
  assign n6397 = ( n3768 & n6390 ) | ( n3768 & n6396 ) | ( n6390 & n6396 ) ;
  assign n6405 = n2427 ^ n2218 ^ n317 ;
  assign n6406 = ( n1490 & n2152 ) | ( n1490 & ~n6405 ) | ( n2152 & ~n6405 ) ;
  assign n6407 = ( n3356 & n6119 ) | ( n3356 & n6406 ) | ( n6119 & n6406 ) ;
  assign n6403 = n5514 ^ n2436 ^ n962 ;
  assign n6404 = ( n919 & n5090 ) | ( n919 & n6403 ) | ( n5090 & n6403 ) ;
  assign n6398 = ( x99 & n160 ) | ( x99 & n910 ) | ( n160 & n910 ) ;
  assign n6399 = n3600 ^ n3114 ^ 1'b0 ;
  assign n6400 = n3710 ^ n3269 ^ x107 ;
  assign n6401 = ( n6398 & n6399 ) | ( n6398 & n6400 ) | ( n6399 & n6400 ) ;
  assign n6402 = n6401 ^ n4153 ^ n1707 ;
  assign n6408 = n6407 ^ n6404 ^ n6402 ;
  assign n6411 = ( n232 & n1377 ) | ( n232 & n1861 ) | ( n1377 & n1861 ) ;
  assign n6412 = ( n834 & n4394 ) | ( n834 & n5007 ) | ( n4394 & n5007 ) ;
  assign n6413 = ( n1345 & n6411 ) | ( n1345 & ~n6412 ) | ( n6411 & ~n6412 ) ;
  assign n6409 = ( ~n2833 & n3035 ) | ( ~n2833 & n3359 ) | ( n3035 & n3359 ) ;
  assign n6410 = ( n2201 & n3305 ) | ( n2201 & ~n6409 ) | ( n3305 & ~n6409 ) ;
  assign n6414 = n6413 ^ n6410 ^ n3127 ;
  assign n6415 = ( ~n1399 & n2991 ) | ( ~n1399 & n3839 ) | ( n2991 & n3839 ) ;
  assign n6416 = ( n2684 & ~n5015 ) | ( n2684 & n6415 ) | ( ~n5015 & n6415 ) ;
  assign n6417 = n6352 ^ n3724 ^ n1602 ;
  assign n6418 = n6417 ^ n4751 ^ 1'b0 ;
  assign n6419 = n6416 & n6418 ;
  assign n6420 = n4344 ^ n3698 ^ n1754 ;
  assign n6425 = n6415 ^ n2188 ^ x15 ;
  assign n6426 = ( n254 & n4136 ) | ( n254 & ~n6425 ) | ( n4136 & ~n6425 ) ;
  assign n6423 = n4684 ^ n4231 ^ n1404 ;
  assign n6421 = ( ~n2429 & n3154 ) | ( ~n2429 & n3366 ) | ( n3154 & n3366 ) ;
  assign n6422 = n6421 ^ n3256 ^ n1609 ;
  assign n6424 = n6423 ^ n6422 ^ n4955 ;
  assign n6427 = n6426 ^ n6424 ^ n2278 ;
  assign n6428 = n4433 & ~n5838 ;
  assign n6429 = n6428 ^ n6233 ^ n4201 ;
  assign n6430 = n6429 ^ n5006 ^ n904 ;
  assign n6431 = n6430 ^ n1494 ^ n1361 ;
  assign n6432 = n4717 | n6431 ;
  assign n6433 = ( n6420 & ~n6427 ) | ( n6420 & n6432 ) | ( ~n6427 & n6432 ) ;
  assign n6442 = ( n523 & n545 ) | ( n523 & n822 ) | ( n545 & n822 ) ;
  assign n6443 = ( n673 & n1274 ) | ( n673 & ~n6442 ) | ( n1274 & ~n6442 ) ;
  assign n6444 = n6443 ^ n4013 ^ n2179 ;
  assign n6434 = n4709 ^ n2493 ^ n1799 ;
  assign n6435 = n6434 ^ n3046 ^ n298 ;
  assign n6436 = n3792 ^ n2660 ^ n926 ;
  assign n6437 = ( x69 & ~n1075 ) | ( x69 & n1674 ) | ( ~n1075 & n1674 ) ;
  assign n6438 = ~n3064 & n6437 ;
  assign n6439 = n6438 ^ x111 ^ 1'b0 ;
  assign n6440 = ( ~n5201 & n6436 ) | ( ~n5201 & n6439 ) | ( n6436 & n6439 ) ;
  assign n6441 = ~n6435 & n6440 ;
  assign n6445 = n6444 ^ n6441 ^ 1'b0 ;
  assign n6449 = ( n133 & ~n2581 ) | ( n133 & n3082 ) | ( ~n2581 & n3082 ) ;
  assign n6450 = ( n6057 & n6184 ) | ( n6057 & ~n6449 ) | ( n6184 & ~n6449 ) ;
  assign n6446 = n5774 ^ n4201 ^ n761 ;
  assign n6447 = ( ~n856 & n3562 ) | ( ~n856 & n6446 ) | ( n3562 & n6446 ) ;
  assign n6448 = n6447 ^ n4068 ^ n4049 ;
  assign n6451 = n6450 ^ n6448 ^ n2462 ;
  assign n6452 = ( n152 & n362 ) | ( n152 & ~n1994 ) | ( n362 & ~n1994 ) ;
  assign n6453 = n6452 ^ n2697 ^ n2120 ;
  assign n6454 = n6453 ^ n3653 ^ n2460 ;
  assign n6455 = n793 & ~n1002 ;
  assign n6456 = n2030 & ~n6455 ;
  assign n6457 = ~n5245 & n6456 ;
  assign n6458 = n2283 ^ n643 ^ 1'b0 ;
  assign n6459 = n1661 ^ n1573 ^ n617 ;
  assign n6460 = ( ~n1336 & n3665 ) | ( ~n1336 & n6459 ) | ( n3665 & n6459 ) ;
  assign n6461 = ( n1574 & n6458 ) | ( n1574 & ~n6460 ) | ( n6458 & ~n6460 ) ;
  assign n6462 = ( ~n456 & n6457 ) | ( ~n456 & n6461 ) | ( n6457 & n6461 ) ;
  assign n6463 = n6454 & ~n6462 ;
  assign n6464 = ~n4251 & n6463 ;
  assign n6469 = ~n1928 & n2985 ;
  assign n6470 = n6469 ^ n6118 ^ n2769 ;
  assign n6465 = n2892 ^ n555 ^ 1'b0 ;
  assign n6466 = n4663 ^ n2331 ^ n2326 ;
  assign n6467 = ( ~n1463 & n3238 ) | ( ~n1463 & n6466 ) | ( n3238 & n6466 ) ;
  assign n6468 = ( n2034 & n6465 ) | ( n2034 & n6467 ) | ( n6465 & n6467 ) ;
  assign n6471 = n6470 ^ n6468 ^ n4965 ;
  assign n6472 = ( n2349 & ~n6129 ) | ( n2349 & n6471 ) | ( ~n6129 & n6471 ) ;
  assign n6479 = ( n374 & ~n1137 ) | ( n374 & n2575 ) | ( ~n1137 & n2575 ) ;
  assign n6480 = n6479 ^ n2340 ^ n2183 ;
  assign n6473 = ( x90 & ~n153 ) | ( x90 & n4128 ) | ( ~n153 & n4128 ) ;
  assign n6474 = n1623 & ~n1909 ;
  assign n6475 = n6474 ^ n1454 ^ 1'b0 ;
  assign n6476 = ( ~n1726 & n1804 ) | ( ~n1726 & n3670 ) | ( n1804 & n3670 ) ;
  assign n6477 = ( n760 & n6475 ) | ( n760 & ~n6476 ) | ( n6475 & ~n6476 ) ;
  assign n6478 = n6473 | n6477 ;
  assign n6481 = n6480 ^ n6478 ^ 1'b0 ;
  assign n6482 = n1489 ^ n1157 ^ n637 ;
  assign n6483 = ( n498 & n1371 ) | ( n498 & ~n2153 ) | ( n1371 & ~n2153 ) ;
  assign n6484 = ( n5416 & ~n6482 ) | ( n5416 & n6483 ) | ( ~n6482 & n6483 ) ;
  assign n6485 = n6484 ^ n4066 ^ n2649 ;
  assign n6496 = n2733 ^ n2665 ^ n2166 ;
  assign n6492 = n5695 ^ n2511 ^ n882 ;
  assign n6493 = n4058 & n6492 ;
  assign n6489 = ( x76 & n559 ) | ( x76 & ~n639 ) | ( n559 & ~n639 ) ;
  assign n6490 = ( ~n734 & n992 ) | ( ~n734 & n6489 ) | ( n992 & n6489 ) ;
  assign n6491 = n6490 ^ n1241 ^ 1'b0 ;
  assign n6494 = n6493 ^ n6491 ^ n3783 ;
  assign n6495 = n4219 & ~n6494 ;
  assign n6497 = n6496 ^ n6495 ^ 1'b0 ;
  assign n6486 = n2971 ^ n2457 ^ n2322 ;
  assign n6487 = ( ~n1331 & n2180 ) | ( ~n1331 & n4456 ) | ( n2180 & n4456 ) ;
  assign n6488 = ( n3404 & n6486 ) | ( n3404 & n6487 ) | ( n6486 & n6487 ) ;
  assign n6498 = n6497 ^ n6488 ^ 1'b0 ;
  assign n6499 = ~n6485 & n6498 ;
  assign n6500 = ( n2598 & n6344 ) | ( n2598 & n6499 ) | ( n6344 & n6499 ) ;
  assign n6506 = n1703 & ~n2176 ;
  assign n6502 = n4793 ^ n1623 ^ n1264 ;
  assign n6503 = n1121 & n1625 ;
  assign n6504 = n6502 & n6503 ;
  assign n6505 = n6504 ^ n930 ^ n257 ;
  assign n6501 = n4122 ^ x7 ^ 1'b0 ;
  assign n6507 = n6506 ^ n6505 ^ n6501 ;
  assign n6508 = n3056 & n4802 ;
  assign n6509 = ~n1524 & n6508 ;
  assign n6510 = x124 & n1849 ;
  assign n6511 = n6510 ^ x112 ^ 1'b0 ;
  assign n6512 = ( n3281 & ~n6509 ) | ( n3281 & n6511 ) | ( ~n6509 & n6511 ) ;
  assign n6513 = n6289 ^ n4274 ^ n2147 ;
  assign n6514 = ( n4265 & n6512 ) | ( n4265 & n6513 ) | ( n6512 & n6513 ) ;
  assign n6515 = ( n1427 & n6460 ) | ( n1427 & ~n6514 ) | ( n6460 & ~n6514 ) ;
  assign n6516 = ( n2661 & n5139 ) | ( n2661 & ~n6515 ) | ( n5139 & ~n6515 ) ;
  assign n6517 = n4518 ^ n2063 ^ n440 ;
  assign n6518 = n1327 | n6517 ;
  assign n6519 = n6518 ^ n5997 ^ 1'b0 ;
  assign n6520 = ( n2488 & n5187 ) | ( n2488 & n6519 ) | ( n5187 & n6519 ) ;
  assign n6521 = ( x11 & n1152 ) | ( x11 & ~n3239 ) | ( n1152 & ~n3239 ) ;
  assign n6522 = n6521 ^ n5186 ^ 1'b0 ;
  assign n6529 = n640 | n3272 ;
  assign n6530 = n414 & ~n6529 ;
  assign n6531 = n2296 ^ n2283 ^ 1'b0 ;
  assign n6532 = ~n1235 & n1474 ;
  assign n6533 = ( n6530 & n6531 ) | ( n6530 & n6532 ) | ( n6531 & n6532 ) ;
  assign n6534 = n6533 ^ n2821 ^ n2705 ;
  assign n6527 = ( n3254 & ~n3760 ) | ( n3254 & n5607 ) | ( ~n3760 & n5607 ) ;
  assign n6528 = n6527 ^ n3338 ^ n2343 ;
  assign n6523 = ( n1623 & ~n4532 ) | ( n1623 & n6370 ) | ( ~n4532 & n6370 ) ;
  assign n6524 = ( ~n2727 & n3339 ) | ( ~n2727 & n6523 ) | ( n3339 & n6523 ) ;
  assign n6525 = n6450 ^ n4886 ^ n3061 ;
  assign n6526 = ( n3613 & n6524 ) | ( n3613 & n6525 ) | ( n6524 & n6525 ) ;
  assign n6535 = n6534 ^ n6528 ^ n6526 ;
  assign n6547 = n2389 ^ n2025 ^ n245 ;
  assign n6544 = ( n440 & ~n909 ) | ( n440 & n1496 ) | ( ~n909 & n1496 ) ;
  assign n6545 = ( n851 & n1035 ) | ( n851 & ~n6544 ) | ( n1035 & ~n6544 ) ;
  assign n6537 = ( n1486 & n2239 ) | ( n1486 & ~n2653 ) | ( n2239 & ~n2653 ) ;
  assign n6538 = n1909 | n3797 ;
  assign n6539 = n6538 ^ n995 ^ 1'b0 ;
  assign n6540 = n3971 ^ n1068 ^ 1'b0 ;
  assign n6541 = ~n6539 & n6540 ;
  assign n6542 = ( n2083 & n6537 ) | ( n2083 & ~n6541 ) | ( n6537 & ~n6541 ) ;
  assign n6543 = ( n1134 & n3120 ) | ( n1134 & n6542 ) | ( n3120 & n6542 ) ;
  assign n6536 = n6126 ^ n612 ^ n606 ;
  assign n6546 = n6545 ^ n6543 ^ n6536 ;
  assign n6548 = n6547 ^ n6546 ^ n2329 ;
  assign n6549 = n6548 ^ n897 ^ 1'b0 ;
  assign n6550 = ( ~n939 & n4244 ) | ( ~n939 & n4401 ) | ( n4244 & n4401 ) ;
  assign n6551 = n4325 ^ n1577 ^ n442 ;
  assign n6552 = n1886 & ~n5368 ;
  assign n6553 = n6551 & n6552 ;
  assign n6554 = ( n5053 & n6550 ) | ( n5053 & ~n6553 ) | ( n6550 & ~n6553 ) ;
  assign n6562 = n2747 ^ n176 ^ 1'b0 ;
  assign n6563 = n6562 ^ n3892 ^ n2331 ;
  assign n6555 = n624 ^ x22 ^ 1'b0 ;
  assign n6556 = n6555 ^ n1304 ^ 1'b0 ;
  assign n6557 = ( ~n415 & n749 ) | ( ~n415 & n3834 ) | ( n749 & n3834 ) ;
  assign n6558 = ( n901 & n2987 ) | ( n901 & n3394 ) | ( n2987 & n3394 ) ;
  assign n6559 = n6558 ^ n4062 ^ n1639 ;
  assign n6560 = ( n4328 & ~n6557 ) | ( n4328 & n6559 ) | ( ~n6557 & n6559 ) ;
  assign n6561 = ( ~n5674 & n6556 ) | ( ~n5674 & n6560 ) | ( n6556 & n6560 ) ;
  assign n6564 = n6563 ^ n6561 ^ 1'b0 ;
  assign n6565 = n514 & ~n6564 ;
  assign n6566 = ( n1684 & ~n2378 ) | ( n1684 & n2944 ) | ( ~n2378 & n2944 ) ;
  assign n6567 = n1370 ^ n1210 ^ n1165 ;
  assign n6568 = ( ~n5464 & n6566 ) | ( ~n5464 & n6567 ) | ( n6566 & n6567 ) ;
  assign n6569 = n6568 ^ n4742 ^ n4540 ;
  assign n6570 = ~n521 & n3617 ;
  assign n6571 = ( n2756 & ~n3265 ) | ( n2756 & n6570 ) | ( ~n3265 & n6570 ) ;
  assign n6572 = n4686 ^ n2121 ^ n1095 ;
  assign n6573 = ( ~n4224 & n6571 ) | ( ~n4224 & n6572 ) | ( n6571 & n6572 ) ;
  assign n6575 = ( ~n2144 & n2429 ) | ( ~n2144 & n2828 ) | ( n2429 & n2828 ) ;
  assign n6574 = n4356 | n6216 ;
  assign n6576 = n6575 ^ n6574 ^ 1'b0 ;
  assign n6577 = n1930 & n4528 ;
  assign n6578 = n6577 ^ n4003 ^ n3100 ;
  assign n6580 = n971 ^ n855 ^ 1'b0 ;
  assign n6581 = ~n4394 & n6580 ;
  assign n6579 = n5674 ^ n4546 ^ n1161 ;
  assign n6582 = n6581 ^ n6579 ^ n5690 ;
  assign n6583 = n6263 ^ n4557 ^ n904 ;
  assign n6584 = n591 & ~n3007 ;
  assign n6585 = n6583 & n6584 ;
  assign n6592 = n641 ^ n451 ^ n374 ;
  assign n6593 = n6592 ^ n4518 ^ n251 ;
  assign n6594 = ( n1842 & n3627 ) | ( n1842 & n6593 ) | ( n3627 & n6593 ) ;
  assign n6586 = ( ~n896 & n1287 ) | ( ~n896 & n3651 ) | ( n1287 & n3651 ) ;
  assign n6587 = n2910 | n6586 ;
  assign n6588 = n6587 ^ n948 ^ n668 ;
  assign n6589 = n3944 ^ n3836 ^ n1258 ;
  assign n6590 = n2539 & n6589 ;
  assign n6591 = ( n2395 & n6588 ) | ( n2395 & ~n6590 ) | ( n6588 & ~n6590 ) ;
  assign n6595 = n6594 ^ n6591 ^ n2229 ;
  assign n6596 = ( ~n781 & n1355 ) | ( ~n781 & n2417 ) | ( n1355 & n2417 ) ;
  assign n6597 = ( n565 & n972 ) | ( n565 & ~n3136 ) | ( n972 & ~n3136 ) ;
  assign n6598 = n1172 ^ n785 ^ x100 ;
  assign n6599 = n4244 | n6598 ;
  assign n6600 = n6597 & ~n6599 ;
  assign n6601 = ( x43 & n6596 ) | ( x43 & n6600 ) | ( n6596 & n6600 ) ;
  assign n6602 = n6601 ^ n1563 ^ 1'b0 ;
  assign n6603 = n676 & n1241 ;
  assign n6604 = n6603 ^ n1478 ^ 1'b0 ;
  assign n6605 = n6604 ^ n668 ^ x76 ;
  assign n6606 = ( ~n2197 & n6602 ) | ( ~n2197 & n6605 ) | ( n6602 & n6605 ) ;
  assign n6607 = n2448 ^ n1115 ^ n295 ;
  assign n6608 = n6607 ^ n6545 ^ n1934 ;
  assign n6609 = ( ~n3352 & n5892 ) | ( ~n3352 & n6608 ) | ( n5892 & n6608 ) ;
  assign n6610 = n6609 ^ n1937 ^ n1538 ;
  assign n6611 = ( n3077 & ~n6606 ) | ( n3077 & n6610 ) | ( ~n6606 & n6610 ) ;
  assign n6615 = ( n2606 & ~n4517 ) | ( n2606 & n5032 ) | ( ~n4517 & n5032 ) ;
  assign n6616 = ( n1460 & ~n2581 ) | ( n1460 & n6615 ) | ( ~n2581 & n6615 ) ;
  assign n6612 = n5918 ^ n1098 ^ n428 ;
  assign n6613 = n6612 ^ n1315 ^ n656 ;
  assign n6614 = n3970 & ~n6613 ;
  assign n6617 = n6616 ^ n6614 ^ n2024 ;
  assign n6618 = ( n214 & n647 ) | ( n214 & n1963 ) | ( n647 & n1963 ) ;
  assign n6619 = n6618 ^ n2901 ^ n1714 ;
  assign n6620 = n3206 ^ n2714 ^ n146 ;
  assign n6621 = ( n2717 & ~n6619 ) | ( n2717 & n6620 ) | ( ~n6619 & n6620 ) ;
  assign n6622 = n6621 ^ n4994 ^ n226 ;
  assign n6623 = n6545 ^ n5974 ^ n688 ;
  assign n6624 = ( n1055 & n1786 ) | ( n1055 & ~n6623 ) | ( n1786 & ~n6623 ) ;
  assign n6625 = ( n270 & n4393 ) | ( n270 & ~n6624 ) | ( n4393 & ~n6624 ) ;
  assign n6626 = n6625 ^ n6445 ^ n1349 ;
  assign n6627 = n2876 ^ n864 ^ x95 ;
  assign n6628 = n557 & n6627 ;
  assign n6629 = n6628 ^ n1479 ^ 1'b0 ;
  assign n6630 = n2209 ^ n627 ^ n330 ;
  assign n6631 = ( n1041 & ~n4108 ) | ( n1041 & n6630 ) | ( ~n4108 & n6630 ) ;
  assign n6632 = ( n1374 & ~n6629 ) | ( n1374 & n6631 ) | ( ~n6629 & n6631 ) ;
  assign n6633 = n6393 ^ n2107 ^ 1'b0 ;
  assign n6634 = n3328 & ~n6633 ;
  assign n6638 = ( n764 & n3314 ) | ( n764 & n4559 ) | ( n3314 & n4559 ) ;
  assign n6635 = ( n3581 & ~n3865 ) | ( n3581 & n5115 ) | ( ~n3865 & n5115 ) ;
  assign n6636 = n6635 ^ n4840 ^ n4392 ;
  assign n6637 = n6636 ^ n6586 ^ n259 ;
  assign n6639 = n6638 ^ n6637 ^ n3551 ;
  assign n6640 = ~n3577 & n4465 ;
  assign n6641 = ( n934 & n4098 ) | ( n934 & ~n6640 ) | ( n4098 & ~n6640 ) ;
  assign n6647 = n3287 ^ n230 ^ 1'b0 ;
  assign n6648 = ~n1753 & n6647 ;
  assign n6649 = ( ~n1154 & n6455 ) | ( ~n1154 & n6648 ) | ( n6455 & n6648 ) ;
  assign n6646 = n4920 ^ n1682 ^ n688 ;
  assign n6643 = n2753 & ~n4045 ;
  assign n6644 = n1920 & ~n6643 ;
  assign n6645 = n1785 & n6644 ;
  assign n6650 = n6649 ^ n6646 ^ n6645 ;
  assign n6642 = ( ~n160 & n4750 ) | ( ~n160 & n5540 ) | ( n4750 & n5540 ) ;
  assign n6651 = n6650 ^ n6645 ^ n6642 ;
  assign n6652 = ( n5899 & n6553 ) | ( n5899 & n6651 ) | ( n6553 & n6651 ) ;
  assign n6653 = ( n1237 & n2074 ) | ( n1237 & ~n3149 ) | ( n2074 & ~n3149 ) ;
  assign n6654 = n6653 ^ n4658 ^ n1706 ;
  assign n6660 = n3628 ^ n2760 ^ n1871 ;
  assign n6658 = n765 ^ x32 ^ 1'b0 ;
  assign n6659 = n6658 ^ n3319 ^ x42 ;
  assign n6655 = ( n4420 & n4958 ) | ( n4420 & n5032 ) | ( n4958 & n5032 ) ;
  assign n6656 = n6339 & n6655 ;
  assign n6657 = n6656 ^ n997 ^ 1'b0 ;
  assign n6661 = n6660 ^ n6659 ^ n6657 ;
  assign n6662 = n1978 ^ n1906 ^ n193 ;
  assign n6663 = n4696 | n6600 ;
  assign n6664 = ( ~n3559 & n6662 ) | ( ~n3559 & n6663 ) | ( n6662 & n6663 ) ;
  assign n6674 = n1374 ^ n666 ^ x77 ;
  assign n6665 = n2274 ^ n1954 ^ 1'b0 ;
  assign n6666 = n6665 ^ n4120 ^ n3105 ;
  assign n6667 = n3261 | n6666 ;
  assign n6668 = n6667 ^ n710 ^ n364 ;
  assign n6669 = n5133 ^ n3841 ^ n1262 ;
  assign n6670 = n6669 ^ n1140 ^ n937 ;
  assign n6671 = n6668 & n6670 ;
  assign n6672 = n6671 ^ n589 ^ 1'b0 ;
  assign n6673 = ~n5811 & n6672 ;
  assign n6675 = n6674 ^ n6673 ^ n898 ;
  assign n6676 = n5656 ^ n2021 ^ n258 ;
  assign n6677 = n6676 ^ n2205 ^ n1461 ;
  assign n6678 = ( ~n1123 & n6675 ) | ( ~n1123 & n6677 ) | ( n6675 & n6677 ) ;
  assign n6679 = n4117 ^ n1735 ^ x127 ;
  assign n6680 = n6679 ^ n4382 ^ n4094 ;
  assign n6681 = n4617 ^ n891 ^ n698 ;
  assign n6682 = ( n4751 & ~n6596 ) | ( n4751 & n6681 ) | ( ~n6596 & n6681 ) ;
  assign n6683 = n3530 ^ n2941 ^ 1'b0 ;
  assign n6684 = ~n1706 & n6683 ;
  assign n6690 = n297 & n840 ;
  assign n6688 = ( n603 & n947 ) | ( n603 & ~n6620 ) | ( n947 & ~n6620 ) ;
  assign n6689 = n6688 ^ n4379 ^ n787 ;
  assign n6686 = ( ~n558 & n1929 ) | ( ~n558 & n5064 ) | ( n1929 & n5064 ) ;
  assign n6685 = n1028 & ~n4199 ;
  assign n6687 = n6686 ^ n6685 ^ n2373 ;
  assign n6691 = n6690 ^ n6689 ^ n6687 ;
  assign n6692 = n2214 & n5157 ;
  assign n6693 = ~n6691 & n6692 ;
  assign n6698 = ( n175 & ~n315 ) | ( n175 & n2250 ) | ( ~n315 & n2250 ) ;
  assign n6696 = ( ~n449 & n1543 ) | ( ~n449 & n3419 ) | ( n1543 & n3419 ) ;
  assign n6697 = ( n1850 & ~n1911 ) | ( n1850 & n6696 ) | ( ~n1911 & n6696 ) ;
  assign n6694 = n3173 ^ n1943 ^ n1381 ;
  assign n6695 = n6694 ^ n6328 ^ n758 ;
  assign n6699 = n6698 ^ n6697 ^ n6695 ;
  assign n6705 = x116 | n337 ;
  assign n6706 = n6705 ^ n511 ^ n227 ;
  assign n6707 = n1847 & n3776 ;
  assign n6708 = ~n6706 & n6707 ;
  assign n6700 = n4775 ^ n2890 ^ n1417 ;
  assign n6701 = ( n404 & ~n3357 ) | ( n404 & n6700 ) | ( ~n3357 & n6700 ) ;
  assign n6702 = n6701 ^ n4953 ^ n2815 ;
  assign n6703 = n6702 ^ n2489 ^ n319 ;
  assign n6704 = n6703 ^ n5683 ^ n962 ;
  assign n6709 = n6708 ^ n6704 ^ n3865 ;
  assign n6710 = ( n2205 & n3159 ) | ( n2205 & n4812 ) | ( n3159 & n4812 ) ;
  assign n6711 = ( n659 & n3390 ) | ( n659 & n6710 ) | ( n3390 & n6710 ) ;
  assign n6713 = ( n445 & n2204 ) | ( n445 & ~n6369 ) | ( n2204 & ~n6369 ) ;
  assign n6712 = ( ~x67 & n1349 ) | ( ~x67 & n3847 ) | ( n1349 & n3847 ) ;
  assign n6714 = n6713 ^ n6712 ^ n1362 ;
  assign n6715 = n1014 & ~n4451 ;
  assign n6716 = n6715 ^ n2595 ^ 1'b0 ;
  assign n6717 = n6716 ^ n1715 ^ x51 ;
  assign n6718 = ( n256 & n2217 ) | ( n256 & n6717 ) | ( n2217 & n6717 ) ;
  assign n6720 = ( n1352 & ~n2386 ) | ( n1352 & n5997 ) | ( ~n2386 & n5997 ) ;
  assign n6719 = n3652 ^ n3061 ^ n1984 ;
  assign n6721 = n6720 ^ n6719 ^ n403 ;
  assign n6722 = n4281 ^ n3564 ^ n2016 ;
  assign n6723 = n5902 ^ n3761 ^ n1165 ;
  assign n6724 = n1556 ^ x101 ^ 1'b0 ;
  assign n6725 = n4846 & n6724 ;
  assign n6726 = ( n578 & n694 ) | ( n578 & ~n1192 ) | ( n694 & ~n1192 ) ;
  assign n6727 = ( ~n3400 & n4931 ) | ( ~n3400 & n6726 ) | ( n4931 & n6726 ) ;
  assign n6728 = n6725 & n6727 ;
  assign n6729 = n6723 & n6728 ;
  assign n6730 = ( n2861 & n6722 ) | ( n2861 & ~n6729 ) | ( n6722 & ~n6729 ) ;
  assign n6731 = n6157 ^ n3791 ^ n1957 ;
  assign n6732 = ~n4372 & n6731 ;
  assign n6733 = n6732 ^ n4285 ^ 1'b0 ;
  assign n6734 = n6733 ^ n4808 ^ 1'b0 ;
  assign n6735 = ~n2726 & n4054 ;
  assign n6736 = n1056 & n6735 ;
  assign n6737 = n6736 ^ n254 ^ 1'b0 ;
  assign n6738 = n4074 & ~n6737 ;
  assign n6739 = n4127 ^ n2770 ^ n494 ;
  assign n6740 = ( ~n1624 & n5716 ) | ( ~n1624 & n6705 ) | ( n5716 & n6705 ) ;
  assign n6741 = ( ~n3622 & n6739 ) | ( ~n3622 & n6740 ) | ( n6739 & n6740 ) ;
  assign n6742 = ( n4722 & ~n6738 ) | ( n4722 & n6741 ) | ( ~n6738 & n6741 ) ;
  assign n6743 = n2656 ^ n1778 ^ n915 ;
  assign n6744 = ( n2265 & n3269 ) | ( n2265 & ~n6743 ) | ( n3269 & ~n6743 ) ;
  assign n6745 = ( n1672 & n4258 ) | ( n1672 & n4546 ) | ( n4258 & n4546 ) ;
  assign n6746 = n3154 ^ n2569 ^ 1'b0 ;
  assign n6747 = n5206 & ~n6746 ;
  assign n6748 = ( n829 & ~n1728 ) | ( n829 & n3248 ) | ( ~n1728 & n3248 ) ;
  assign n6749 = n6748 ^ n5428 ^ n3080 ;
  assign n6750 = ( ~n859 & n6747 ) | ( ~n859 & n6749 ) | ( n6747 & n6749 ) ;
  assign n6752 = ( n761 & n1368 ) | ( n761 & n2773 ) | ( n1368 & n2773 ) ;
  assign n6751 = ( n943 & n2315 ) | ( n943 & n4204 ) | ( n2315 & n4204 ) ;
  assign n6753 = n6752 ^ n6751 ^ n1027 ;
  assign n6756 = ( n740 & n1566 ) | ( n740 & ~n1668 ) | ( n1566 & ~n1668 ) ;
  assign n6757 = n6756 ^ n810 ^ n399 ;
  assign n6754 = ( n1133 & ~n1178 ) | ( n1133 & n3412 ) | ( ~n1178 & n3412 ) ;
  assign n6755 = ~n4049 & n6754 ;
  assign n6758 = n6757 ^ n6755 ^ 1'b0 ;
  assign n6759 = n6758 ^ n6556 ^ x122 ;
  assign n6760 = ( n265 & n329 ) | ( n265 & ~n444 ) | ( n329 & ~n444 ) ;
  assign n6761 = n6760 ^ n3208 ^ n1113 ;
  assign n6766 = n4733 ^ n1241 ^ 1'b0 ;
  assign n6767 = ~n488 & n6766 ;
  assign n6763 = n3066 ^ n2558 ^ n482 ;
  assign n6764 = ( n840 & ~n2649 ) | ( n840 & n6763 ) | ( ~n2649 & n6763 ) ;
  assign n6762 = n1929 & n2813 ;
  assign n6765 = n6764 ^ n6762 ^ n3971 ;
  assign n6768 = n6767 ^ n6765 ^ n2082 ;
  assign n6769 = n6761 | n6768 ;
  assign n6770 = ( n345 & n1788 ) | ( n345 & ~n2083 ) | ( n1788 & ~n2083 ) ;
  assign n6771 = n3635 & ~n6770 ;
  assign n6772 = n4243 ^ n3188 ^ n617 ;
  assign n6773 = n6772 ^ n6274 ^ n6086 ;
  assign n6776 = x21 & n1167 ;
  assign n6777 = ~n547 & n6776 ;
  assign n6774 = n4511 ^ n187 ^ 1'b0 ;
  assign n6775 = n6774 ^ n4829 ^ 1'b0 ;
  assign n6778 = n6777 ^ n6775 ^ n1400 ;
  assign n6779 = n6283 ^ n4148 ^ 1'b0 ;
  assign n6780 = n1254 & n6779 ;
  assign n6781 = n5416 ^ n2959 ^ 1'b0 ;
  assign n6782 = ( n234 & n621 ) | ( n234 & ~n5484 ) | ( n621 & ~n5484 ) ;
  assign n6783 = ( n612 & ~n2522 ) | ( n612 & n6782 ) | ( ~n2522 & n6782 ) ;
  assign n6788 = n2976 ^ n2730 ^ n1263 ;
  assign n6784 = n1866 ^ n1668 ^ x17 ;
  assign n6785 = ( n415 & ~n2964 ) | ( n415 & n4914 ) | ( ~n2964 & n4914 ) ;
  assign n6786 = n4155 & ~n6785 ;
  assign n6787 = n6784 & n6786 ;
  assign n6789 = n6788 ^ n6787 ^ n1447 ;
  assign n6790 = ( n6781 & n6783 ) | ( n6781 & ~n6789 ) | ( n6783 & ~n6789 ) ;
  assign n6793 = ( n481 & n1125 ) | ( n481 & ~n1452 ) | ( n1125 & ~n1452 ) ;
  assign n6794 = n6793 ^ n1202 ^ n220 ;
  assign n6795 = ( n656 & n805 ) | ( n656 & n6794 ) | ( n805 & n6794 ) ;
  assign n6796 = n6795 ^ n6450 ^ 1'b0 ;
  assign n6791 = n5980 ^ n4836 ^ 1'b0 ;
  assign n6792 = ~n3738 & n6791 ;
  assign n6797 = n6796 ^ n6792 ^ n1139 ;
  assign n6801 = n3893 ^ n2381 ^ n1571 ;
  assign n6802 = ( x120 & n6587 ) | ( x120 & n6801 ) | ( n6587 & n6801 ) ;
  assign n6799 = ( ~x119 & n1521 ) | ( ~x119 & n2189 ) | ( n1521 & n2189 ) ;
  assign n6798 = ( n981 & n1883 ) | ( n981 & n4527 ) | ( n1883 & n4527 ) ;
  assign n6800 = n6799 ^ n6798 ^ n2547 ;
  assign n6803 = n6802 ^ n6800 ^ n4155 ;
  assign n6812 = ~n653 & n2723 ;
  assign n6808 = ( n1616 & ~n2032 ) | ( n1616 & n5189 ) | ( ~n2032 & n5189 ) ;
  assign n6807 = ( n366 & n3057 ) | ( n366 & ~n4905 ) | ( n3057 & ~n4905 ) ;
  assign n6804 = n6506 ^ n3311 ^ x5 ;
  assign n6805 = n6504 & ~n6804 ;
  assign n6806 = ( n1783 & ~n1959 ) | ( n1783 & n6805 ) | ( ~n1959 & n6805 ) ;
  assign n6809 = n6808 ^ n6807 ^ n6806 ;
  assign n6810 = n4692 & ~n6809 ;
  assign n6811 = n6810 ^ n3020 ^ 1'b0 ;
  assign n6813 = n6812 ^ n6811 ^ n466 ;
  assign n6814 = ~n1475 & n3212 ;
  assign n6815 = ~n6813 & n6814 ;
  assign n6816 = n2309 & ~n4136 ;
  assign n6817 = n6816 ^ n1848 ^ n1586 ;
  assign n6820 = n380 & n5724 ;
  assign n6821 = ~n6686 & n6820 ;
  assign n6818 = ( n382 & ~n1044 ) | ( n382 & n1301 ) | ( ~n1044 & n1301 ) ;
  assign n6819 = ( ~n788 & n4175 ) | ( ~n788 & n6818 ) | ( n4175 & n6818 ) ;
  assign n6822 = n6821 ^ n6819 ^ n1234 ;
  assign n6823 = ( n3914 & n4693 ) | ( n3914 & ~n6822 ) | ( n4693 & ~n6822 ) ;
  assign n6824 = n6823 ^ n5273 ^ 1'b0 ;
  assign n6825 = ( ~n1308 & n6817 ) | ( ~n1308 & n6824 ) | ( n6817 & n6824 ) ;
  assign n6826 = ~n2060 & n5068 ;
  assign n6827 = n6826 ^ n3159 ^ 1'b0 ;
  assign n6828 = n6076 ^ n3064 ^ n2652 ;
  assign n6829 = n6828 ^ n3493 ^ x63 ;
  assign n6830 = ( n1202 & n5597 ) | ( n1202 & ~n6829 ) | ( n5597 & ~n6829 ) ;
  assign n6831 = n2824 ^ n437 ^ 1'b0 ;
  assign n6841 = n583 & ~n1018 ;
  assign n6842 = n1730 & n6841 ;
  assign n6837 = ( ~x81 & n759 ) | ( ~x81 & n867 ) | ( n759 & n867 ) ;
  assign n6838 = n6837 ^ n2952 ^ n2749 ;
  assign n6839 = ( n810 & ~n1023 ) | ( n810 & n6838 ) | ( ~n1023 & n6838 ) ;
  assign n6832 = n5965 ^ n1308 ^ n1077 ;
  assign n6833 = n6832 ^ n918 ^ x105 ;
  assign n6834 = n6833 ^ x0 ^ 1'b0 ;
  assign n6835 = ~n1304 & n6834 ;
  assign n6836 = ~n1306 & n6835 ;
  assign n6840 = n6839 ^ n6836 ^ 1'b0 ;
  assign n6843 = n6842 ^ n6840 ^ n5978 ;
  assign n6844 = ( ~n636 & n4985 ) | ( ~n636 & n5425 ) | ( n4985 & n5425 ) ;
  assign n6845 = n819 ^ n221 ^ x23 ;
  assign n6846 = n3746 ^ n1386 ^ n1241 ;
  assign n6847 = ( n4002 & n6845 ) | ( n4002 & n6846 ) | ( n6845 & n6846 ) ;
  assign n6848 = n6847 ^ n4521 ^ 1'b0 ;
  assign n6849 = ( n1578 & ~n1673 ) | ( n1578 & n6848 ) | ( ~n1673 & n6848 ) ;
  assign n6850 = ( x119 & n1959 ) | ( x119 & n4747 ) | ( n1959 & n4747 ) ;
  assign n6851 = ( n2062 & ~n3502 ) | ( n2062 & n4058 ) | ( ~n3502 & n4058 ) ;
  assign n6852 = n1511 & n2888 ;
  assign n6853 = ~n4756 & n6852 ;
  assign n6858 = ( n683 & n1867 ) | ( n683 & n2610 ) | ( n1867 & n2610 ) ;
  assign n6854 = n449 ^ n201 ^ 1'b0 ;
  assign n6855 = n1369 & n6854 ;
  assign n6856 = n926 ^ n803 ^ 1'b0 ;
  assign n6857 = n6855 & n6856 ;
  assign n6859 = n6858 ^ n6857 ^ n6227 ;
  assign n6860 = n6859 ^ n3306 ^ 1'b0 ;
  assign n6861 = ( n6407 & n6853 ) | ( n6407 & ~n6860 ) | ( n6853 & ~n6860 ) ;
  assign n6862 = n3197 ^ n2138 ^ n1061 ;
  assign n6863 = ( n1392 & n4825 ) | ( n1392 & n6862 ) | ( n4825 & n6862 ) ;
  assign n6864 = n6863 ^ n2844 ^ n1603 ;
  assign n6865 = n6864 ^ n6040 ^ x59 ;
  assign n6866 = ( n1265 & ~n1706 ) | ( n1265 & n6106 ) | ( ~n1706 & n6106 ) ;
  assign n6867 = ( x122 & n1647 ) | ( x122 & n6866 ) | ( n1647 & n6866 ) ;
  assign n6871 = ( n905 & ~n1778 ) | ( n905 & n2576 ) | ( ~n1778 & n2576 ) ;
  assign n6872 = n6871 ^ n780 ^ n539 ;
  assign n6870 = n4329 ^ n799 ^ x62 ;
  assign n6873 = n6872 ^ n6870 ^ n6795 ;
  assign n6874 = n6873 ^ n2538 ^ 1'b0 ;
  assign n6868 = n2144 ^ n708 ^ 1'b0 ;
  assign n6869 = n4742 & ~n6868 ;
  assign n6875 = n6874 ^ n6869 ^ n5822 ;
  assign n6876 = ( n293 & n350 ) | ( n293 & ~n3249 ) | ( n350 & ~n3249 ) ;
  assign n6877 = ( n1215 & n4841 ) | ( n1215 & n6876 ) | ( n4841 & n6876 ) ;
  assign n6878 = n6877 ^ n6331 ^ n5063 ;
  assign n6879 = n6878 ^ n3718 ^ 1'b0 ;
  assign n6880 = ~n2141 & n6879 ;
  assign n6881 = ( ~n4972 & n6875 ) | ( ~n4972 & n6880 ) | ( n6875 & n6880 ) ;
  assign n6882 = ( n1133 & n1505 ) | ( n1133 & n2678 ) | ( n1505 & n2678 ) ;
  assign n6883 = ( n188 & ~n2830 ) | ( n188 & n2953 ) | ( ~n2830 & n2953 ) ;
  assign n6884 = n6883 ^ n3611 ^ x65 ;
  assign n6885 = n6733 ^ n4738 ^ n3821 ;
  assign n6886 = ( n349 & n6884 ) | ( n349 & ~n6885 ) | ( n6884 & ~n6885 ) ;
  assign n6887 = ( ~n539 & n6882 ) | ( ~n539 & n6886 ) | ( n6882 & n6886 ) ;
  assign n6896 = n5098 ^ n4204 ^ n3357 ;
  assign n6895 = n3860 ^ n1446 ^ n971 ;
  assign n6897 = n6896 ^ n6895 ^ n3558 ;
  assign n6898 = n3374 & n6897 ;
  assign n6899 = ~n609 & n6898 ;
  assign n6892 = n5957 ^ n3225 ^ 1'b0 ;
  assign n6893 = n6566 | n6892 ;
  assign n6890 = ( n602 & ~n1273 ) | ( n602 & n3893 ) | ( ~n1273 & n3893 ) ;
  assign n6891 = ( n1883 & n3499 ) | ( n1883 & ~n6890 ) | ( n3499 & ~n6890 ) ;
  assign n6889 = ( ~n755 & n4356 ) | ( ~n755 & n5505 ) | ( n4356 & n5505 ) ;
  assign n6894 = n6893 ^ n6891 ^ n6889 ;
  assign n6888 = ~n3253 & n6587 ;
  assign n6900 = n6899 ^ n6894 ^ n6888 ;
  assign n6901 = ( n4756 & n6307 ) | ( n4756 & ~n6900 ) | ( n6307 & ~n6900 ) ;
  assign n6902 = n6482 ^ n2963 ^ n1565 ;
  assign n6903 = n5725 ^ n4771 ^ n2523 ;
  assign n6904 = n6708 ^ n6119 ^ n4541 ;
  assign n6905 = n6904 ^ n4530 ^ n4473 ;
  assign n6906 = ( ~n5407 & n6903 ) | ( ~n5407 & n6905 ) | ( n6903 & n6905 ) ;
  assign n6907 = ( n4686 & n6902 ) | ( n4686 & n6906 ) | ( n6902 & n6906 ) ;
  assign n6908 = n6907 ^ n4350 ^ n3822 ;
  assign n6912 = n2843 ^ n2575 ^ 1'b0 ;
  assign n6913 = n599 | n6912 ;
  assign n6911 = ~n3859 & n5879 ;
  assign n6909 = n4395 ^ n2718 ^ x93 ;
  assign n6910 = n6909 ^ n5679 ^ n3741 ;
  assign n6914 = n6913 ^ n6911 ^ n6910 ;
  assign n6919 = n3841 ^ n2781 ^ n1645 ;
  assign n6916 = n3670 ^ n684 ^ x83 ;
  assign n6917 = n6604 ^ n2214 ^ n1154 ;
  assign n6918 = n6916 | n6917 ;
  assign n6915 = n5576 ^ n1732 ^ n728 ;
  assign n6920 = n6919 ^ n6918 ^ n6915 ;
  assign n6925 = n5041 ^ n942 ^ 1'b0 ;
  assign n6926 = ~n6306 & n6925 ;
  assign n6927 = n6926 ^ n1201 ^ 1'b0 ;
  assign n6928 = n715 & ~n6927 ;
  assign n6921 = n5554 ^ n3698 ^ n2678 ;
  assign n6922 = ( n1223 & n3964 ) | ( n1223 & ~n6921 ) | ( n3964 & ~n6921 ) ;
  assign n6923 = n5680 ^ n3581 ^ n1685 ;
  assign n6924 = ( n1696 & n6922 ) | ( n1696 & ~n6923 ) | ( n6922 & ~n6923 ) ;
  assign n6929 = n6928 ^ n6924 ^ n6832 ;
  assign n6931 = n4843 ^ n3002 ^ n2927 ;
  assign n6930 = n1918 & n3163 ;
  assign n6932 = n6931 ^ n6930 ^ 1'b0 ;
  assign n6933 = n6932 ^ n2910 ^ n967 ;
  assign n6940 = n917 & n4262 ;
  assign n6941 = ~n4566 & n6940 ;
  assign n6936 = n1192 & n3408 ;
  assign n6937 = n1270 & n6936 ;
  assign n6938 = n620 | n6937 ;
  assign n6939 = n6938 ^ n3382 ^ 1'b0 ;
  assign n6934 = x39 & ~n858 ;
  assign n6935 = ~n2881 & n6934 ;
  assign n6942 = n6941 ^ n6939 ^ n6935 ;
  assign n6943 = ( n1725 & ~n3483 ) | ( n1725 & n3515 ) | ( ~n3483 & n3515 ) ;
  assign n6944 = n6943 ^ n6361 ^ n1706 ;
  assign n6968 = n6587 ^ n6265 ^ n3820 ;
  assign n6969 = n5245 ^ n3776 ^ 1'b0 ;
  assign n6970 = ~n6968 & n6969 ;
  assign n6951 = n3916 ^ n1289 ^ n841 ;
  assign n6952 = ( n1756 & n4010 ) | ( n1756 & ~n6951 ) | ( n4010 & ~n6951 ) ;
  assign n6950 = n1383 | n5069 ;
  assign n6953 = n6952 ^ n6950 ^ 1'b0 ;
  assign n6954 = ( n354 & n1501 ) | ( n354 & ~n6953 ) | ( n1501 & ~n6953 ) ;
  assign n6947 = ( ~n280 & n2167 ) | ( ~n280 & n3229 ) | ( n2167 & n3229 ) ;
  assign n6948 = ( n170 & n2608 ) | ( n170 & n6588 ) | ( n2608 & n6588 ) ;
  assign n6949 = ( n2695 & ~n6947 ) | ( n2695 & n6948 ) | ( ~n6947 & n6948 ) ;
  assign n6945 = n311 & ~n698 ;
  assign n6946 = ~n1028 & n6945 ;
  assign n6955 = n6954 ^ n6949 ^ n6946 ;
  assign n6956 = ~n278 & n856 ;
  assign n6957 = n6956 ^ n2393 ^ n2165 ;
  assign n6958 = n6957 ^ n6623 ^ n5949 ;
  assign n6964 = ( n1158 & n3007 ) | ( n1158 & n4669 ) | ( n3007 & n4669 ) ;
  assign n6959 = n6740 ^ n1931 ^ n391 ;
  assign n6960 = ( x106 & n420 ) | ( x106 & ~n1297 ) | ( n420 & ~n1297 ) ;
  assign n6961 = n2250 ^ n2095 ^ n1612 ;
  assign n6962 = ( n379 & n6960 ) | ( n379 & n6961 ) | ( n6960 & n6961 ) ;
  assign n6963 = ( ~n717 & n6959 ) | ( ~n717 & n6962 ) | ( n6959 & n6962 ) ;
  assign n6965 = n6964 ^ n6963 ^ n4085 ;
  assign n6966 = ( n4551 & ~n6958 ) | ( n4551 & n6965 ) | ( ~n6958 & n6965 ) ;
  assign n6967 = ~n6955 & n6966 ;
  assign n6971 = n6970 ^ n6967 ^ 1'b0 ;
  assign n6972 = ( ~n3133 & n5510 ) | ( ~n3133 & n6971 ) | ( n5510 & n6971 ) ;
  assign n6973 = n6972 ^ n6469 ^ n4926 ;
  assign n6974 = ( n2718 & n2952 ) | ( n2718 & n3406 ) | ( n2952 & n3406 ) ;
  assign n6975 = n6271 ^ n4431 ^ 1'b0 ;
  assign n6976 = n2863 & ~n6975 ;
  assign n6977 = ( n6206 & ~n6974 ) | ( n6206 & n6976 ) | ( ~n6974 & n6976 ) ;
  assign n6978 = n4061 ^ n3046 ^ n1095 ;
  assign n6979 = n6978 ^ n3002 ^ n522 ;
  assign n6980 = n6979 ^ n6175 ^ n4790 ;
  assign n6981 = n6895 ^ n4327 ^ n702 ;
  assign n6982 = n6981 ^ n6354 ^ n4589 ;
  assign n6983 = n6982 ^ n6423 ^ n3657 ;
  assign n6984 = n4391 ^ n3930 ^ n2963 ;
  assign n6985 = ( ~n4038 & n4175 ) | ( ~n4038 & n4605 ) | ( n4175 & n4605 ) ;
  assign n6986 = ( n274 & n5841 ) | ( n274 & n6985 ) | ( n5841 & n6985 ) ;
  assign n6987 = ( ~n5111 & n6984 ) | ( ~n5111 & n6986 ) | ( n6984 & n6986 ) ;
  assign n6988 = ( n258 & n698 ) | ( n258 & n6301 ) | ( n698 & n6301 ) ;
  assign n6989 = n532 & ~n6988 ;
  assign n6990 = n6989 ^ n3324 ^ 1'b0 ;
  assign n6995 = n5962 ^ n4055 ^ 1'b0 ;
  assign n6996 = n3480 & ~n6995 ;
  assign n6991 = n3144 ^ n2029 ^ n881 ;
  assign n6992 = n5888 ^ n4206 ^ n3013 ;
  assign n6993 = ( n1662 & n6991 ) | ( n1662 & n6992 ) | ( n6991 & n6992 ) ;
  assign n6994 = ( n3568 & n5874 ) | ( n3568 & ~n6993 ) | ( n5874 & ~n6993 ) ;
  assign n6997 = n6996 ^ n6994 ^ n2309 ;
  assign n6998 = n5003 ^ n1204 ^ n329 ;
  assign n6999 = n6998 ^ n6690 ^ n6535 ;
  assign n7001 = n3387 ^ n1654 ^ n714 ;
  assign n7000 = n2708 ^ n2111 ^ n601 ;
  assign n7002 = n7001 ^ n7000 ^ n2045 ;
  assign n7003 = n4167 ^ n3524 ^ 1'b0 ;
  assign n7009 = ( ~n751 & n1115 ) | ( ~n751 & n6960 ) | ( n1115 & n6960 ) ;
  assign n7007 = x82 & n1655 ;
  assign n7008 = ~n4143 & n7007 ;
  assign n7004 = n2127 ^ n2050 ^ n1476 ;
  assign n7005 = n971 & ~n2803 ;
  assign n7006 = ( n1204 & n7004 ) | ( n1204 & n7005 ) | ( n7004 & n7005 ) ;
  assign n7010 = n7009 ^ n7008 ^ n7006 ;
  assign n7011 = ( ~n676 & n4157 ) | ( ~n676 & n4867 ) | ( n4157 & n4867 ) ;
  assign n7012 = ( ~n2708 & n6492 ) | ( ~n2708 & n7011 ) | ( n6492 & n7011 ) ;
  assign n7013 = n7012 ^ n4610 ^ n2031 ;
  assign n7014 = n7013 ^ n5489 ^ x87 ;
  assign n7016 = ( n955 & n4161 ) | ( n955 & n4748 ) | ( n4161 & n4748 ) ;
  assign n7015 = ( n1097 & ~n4651 ) | ( n1097 & n5060 ) | ( ~n4651 & n5060 ) ;
  assign n7017 = n7016 ^ n7015 ^ n5067 ;
  assign n7018 = n7014 & n7017 ;
  assign n7019 = n4910 ^ n1599 ^ n426 ;
  assign n7020 = n3106 ^ n2373 ^ 1'b0 ;
  assign n7021 = n5196 ^ n1932 ^ x51 ;
  assign n7022 = n6426 | n7021 ;
  assign n7023 = ( n3843 & n7020 ) | ( n3843 & n7022 ) | ( n7020 & n7022 ) ;
  assign n7024 = n1228 | n7015 ;
  assign n7025 = n1971 | n7024 ;
  assign n7026 = ( n307 & ~n1470 ) | ( n307 & n3353 ) | ( ~n1470 & n3353 ) ;
  assign n7027 = ( ~n426 & n1109 ) | ( ~n426 & n2642 ) | ( n1109 & n2642 ) ;
  assign n7028 = ( n4555 & n4692 ) | ( n4555 & n5838 ) | ( n4692 & n5838 ) ;
  assign n7029 = n7028 ^ n3832 ^ n3022 ;
  assign n7030 = ( n1662 & n7027 ) | ( n1662 & n7029 ) | ( n7027 & n7029 ) ;
  assign n7031 = ( n2960 & n7026 ) | ( n2960 & ~n7030 ) | ( n7026 & ~n7030 ) ;
  assign n7032 = n5939 ^ n1544 ^ n302 ;
  assign n7033 = ( n2634 & n5745 ) | ( n2634 & n7032 ) | ( n5745 & n7032 ) ;
  assign n7034 = n7033 ^ n5611 ^ n1784 ;
  assign n7035 = ( ~n1834 & n2899 ) | ( ~n1834 & n3855 ) | ( n2899 & n3855 ) ;
  assign n7036 = n7035 ^ n4052 ^ 1'b0 ;
  assign n7037 = n263 & n2959 ;
  assign n7038 = ~n6697 & n7037 ;
  assign n7039 = ( n4303 & n6982 ) | ( n4303 & ~n7038 ) | ( n6982 & ~n7038 ) ;
  assign n7040 = ( n1771 & n1812 ) | ( n1771 & ~n3002 ) | ( n1812 & ~n3002 ) ;
  assign n7041 = ( ~n4895 & n6655 ) | ( ~n4895 & n7040 ) | ( n6655 & n7040 ) ;
  assign n7042 = n7041 ^ n6485 ^ n1100 ;
  assign n7043 = n7042 ^ n6842 ^ n4032 ;
  assign n7044 = n3510 ^ n2310 ^ n1080 ;
  assign n7045 = n1227 | n7044 ;
  assign n7046 = n260 & ~n7045 ;
  assign n7047 = n5505 | n7046 ;
  assign n7048 = ( n818 & n1106 ) | ( n818 & ~n3429 ) | ( n1106 & ~n3429 ) ;
  assign n7049 = n5076 | n7048 ;
  assign n7050 = n2134 | n7049 ;
  assign n7051 = n393 & ~n5090 ;
  assign n7052 = n7051 ^ n3833 ^ n2100 ;
  assign n7053 = ( ~n1725 & n5635 ) | ( ~n1725 & n6229 ) | ( n5635 & n6229 ) ;
  assign n7054 = n1633 ^ n604 ^ n260 ;
  assign n7055 = n7054 ^ n1331 ^ n1169 ;
  assign n7056 = n7055 ^ n4184 ^ n1206 ;
  assign n7057 = n7056 ^ n5936 ^ n309 ;
  assign n7058 = ( ~n4623 & n7053 ) | ( ~n4623 & n7057 ) | ( n7053 & n7057 ) ;
  assign n7059 = ( n7050 & ~n7052 ) | ( n7050 & n7058 ) | ( ~n7052 & n7058 ) ;
  assign n7060 = n7059 ^ n5818 ^ n1760 ;
  assign n7061 = ( ~n330 & n410 ) | ( ~n330 & n789 ) | ( n410 & n789 ) ;
  assign n7062 = ( ~n479 & n2721 ) | ( ~n479 & n2780 ) | ( n2721 & n2780 ) ;
  assign n7063 = ( n1912 & ~n4641 ) | ( n1912 & n7062 ) | ( ~n4641 & n7062 ) ;
  assign n7064 = ( x11 & n2429 ) | ( x11 & n5369 ) | ( n2429 & n5369 ) ;
  assign n7065 = ( ~x113 & n6528 ) | ( ~x113 & n7064 ) | ( n6528 & n7064 ) ;
  assign n7066 = n6845 & n7065 ;
  assign n7067 = ( n7061 & n7063 ) | ( n7061 & n7066 ) | ( n7063 & n7066 ) ;
  assign n7068 = ( ~n2092 & n2195 ) | ( ~n2092 & n3982 ) | ( n2195 & n3982 ) ;
  assign n7069 = ( ~n2133 & n4969 ) | ( ~n2133 & n7068 ) | ( n4969 & n7068 ) ;
  assign n7070 = ( ~n1489 & n2794 ) | ( ~n1489 & n7069 ) | ( n2794 & n7069 ) ;
  assign n7071 = n2237 ^ n1548 ^ n1114 ;
  assign n7072 = ( ~n2706 & n6354 ) | ( ~n2706 & n7071 ) | ( n6354 & n7071 ) ;
  assign n7073 = n6057 ^ n1394 ^ 1'b0 ;
  assign n7074 = ( n3073 & n7072 ) | ( n3073 & n7073 ) | ( n7072 & n7073 ) ;
  assign n7075 = n6376 | n7074 ;
  assign n7076 = n7075 ^ x75 ^ 1'b0 ;
  assign n7077 = n3545 ^ n2703 ^ n1896 ;
  assign n7078 = n4552 ^ x33 ^ 1'b0 ;
  assign n7079 = ( n1927 & n3734 ) | ( n1927 & ~n5886 ) | ( n3734 & ~n5886 ) ;
  assign n7081 = n2331 ^ n1407 ^ 1'b0 ;
  assign n7080 = n6598 ^ n6307 ^ n1885 ;
  assign n7082 = n7081 ^ n7080 ^ 1'b0 ;
  assign n7083 = n7079 | n7082 ;
  assign n7084 = ( n6431 & n7078 ) | ( n6431 & ~n7083 ) | ( n7078 & ~n7083 ) ;
  assign n7085 = ~n1288 & n7084 ;
  assign n7086 = n7085 ^ n5697 ^ 1'b0 ;
  assign n7087 = ( n1393 & ~n3961 ) | ( n1393 & n4610 ) | ( ~n3961 & n4610 ) ;
  assign n7088 = n7087 ^ n3779 ^ n2171 ;
  assign n7089 = n7088 ^ n1846 ^ n1089 ;
  assign n7090 = ~n2462 & n5230 ;
  assign n7091 = ( ~x110 & n140 ) | ( ~x110 & n1400 ) | ( n140 & n1400 ) ;
  assign n7092 = ( ~n3047 & n4569 ) | ( ~n3047 & n7091 ) | ( n4569 & n7091 ) ;
  assign n7096 = n4977 ^ n4487 ^ n1281 ;
  assign n7093 = n1877 & n4108 ;
  assign n7094 = n7093 ^ n5126 ^ n641 ;
  assign n7095 = n1546 & n7094 ;
  assign n7097 = n7096 ^ n7095 ^ 1'b0 ;
  assign n7098 = n7092 & ~n7097 ;
  assign n7099 = ~n7090 & n7098 ;
  assign n7100 = n2222 ^ n1804 ^ x32 ;
  assign n7101 = n7100 ^ n3720 ^ n1718 ;
  assign n7102 = n4101 & ~n7101 ;
  assign n7103 = n6139 & n7102 ;
  assign n7105 = n3114 ^ n3049 ^ n354 ;
  assign n7106 = n7105 ^ n1589 ^ n586 ;
  assign n7104 = n6216 ^ n2149 ^ 1'b0 ;
  assign n7107 = n7106 ^ n7104 ^ n4660 ;
  assign n7108 = n4231 & ~n4281 ;
  assign n7109 = n7108 ^ n5351 ^ n4034 ;
  assign n7110 = ( ~n2272 & n7107 ) | ( ~n2272 & n7109 ) | ( n7107 & n7109 ) ;
  assign n7111 = n224 & ~n7110 ;
  assign n7112 = n5175 ^ n2015 ^ 1'b0 ;
  assign n7113 = ~n694 & n7112 ;
  assign n7114 = ~n2413 & n7113 ;
  assign n7115 = n2669 ^ n1199 ^ n1009 ;
  assign n7116 = n4004 ^ n1353 ^ 1'b0 ;
  assign n7117 = n7116 ^ n3120 ^ n490 ;
  assign n7118 = ( n4397 & n6228 ) | ( n4397 & n7117 ) | ( n6228 & n7117 ) ;
  assign n7119 = ( n2454 & n7115 ) | ( n2454 & ~n7118 ) | ( n7115 & ~n7118 ) ;
  assign n7120 = ( n1442 & ~n2315 ) | ( n1442 & n5607 ) | ( ~n2315 & n5607 ) ;
  assign n7122 = n5566 ^ n4120 ^ n1755 ;
  assign n7121 = n4774 | n6453 ;
  assign n7123 = n7122 ^ n7121 ^ n6176 ;
  assign n7124 = n5646 ^ n1998 ^ n1745 ;
  assign n7125 = ( n5547 & n7123 ) | ( n5547 & n7124 ) | ( n7123 & n7124 ) ;
  assign n7126 = ( ~x115 & n3802 ) | ( ~x115 & n6978 ) | ( n3802 & n6978 ) ;
  assign n7127 = n7126 ^ n5251 ^ n4258 ;
  assign n7134 = n1238 ^ n1102 ^ n765 ;
  assign n7128 = n4187 ^ n3420 ^ 1'b0 ;
  assign n7129 = n2600 & ~n7128 ;
  assign n7130 = ( n1695 & n3063 ) | ( n1695 & ~n7129 ) | ( n3063 & ~n7129 ) ;
  assign n7131 = n4452 | n7130 ;
  assign n7132 = n3950 & ~n7131 ;
  assign n7133 = ( ~x42 & n6686 ) | ( ~x42 & n7132 ) | ( n6686 & n7132 ) ;
  assign n7135 = n7134 ^ n7133 ^ n1256 ;
  assign n7137 = ( n687 & n2441 ) | ( n687 & n6991 ) | ( n2441 & n6991 ) ;
  assign n7136 = n5466 ^ n237 ^ 1'b0 ;
  assign n7138 = n7137 ^ n7136 ^ n3748 ;
  assign n7139 = n7138 ^ n5817 ^ n2224 ;
  assign n7140 = n7139 ^ n6497 ^ n781 ;
  assign n7141 = n3260 ^ n1910 ^ 1'b0 ;
  assign n7142 = n7140 & n7141 ;
  assign n7143 = n7142 ^ n3582 ^ 1'b0 ;
  assign n7144 = n4962 ^ n1812 ^ x24 ;
  assign n7145 = n4248 | n7144 ;
  assign n7146 = n7145 ^ n3826 ^ 1'b0 ;
  assign n7147 = n7146 ^ n5599 ^ n5501 ;
  assign n7153 = n4416 ^ n2108 ^ n1708 ;
  assign n7151 = n2310 ^ n1743 ^ n595 ;
  assign n7149 = n6537 ^ n5942 ^ n1442 ;
  assign n7148 = ~n1115 & n4714 ;
  assign n7150 = n7149 ^ n7148 ^ n4959 ;
  assign n7152 = n7151 ^ n7150 ^ n4983 ;
  assign n7154 = n7153 ^ n7152 ^ n3898 ;
  assign n7155 = ( n2468 & ~n4767 ) | ( n2468 & n4949 ) | ( ~n4767 & n4949 ) ;
  assign n7156 = ( ~n1712 & n1826 ) | ( ~n1712 & n4226 ) | ( n1826 & n4226 ) ;
  assign n7157 = ( n2024 & ~n2835 ) | ( n2024 & n7156 ) | ( ~n2835 & n7156 ) ;
  assign n7158 = n7157 ^ n5191 ^ n383 ;
  assign n7159 = ( n6535 & n7155 ) | ( n6535 & n7158 ) | ( n7155 & n7158 ) ;
  assign n7160 = ~n4014 & n5462 ;
  assign n7161 = n5027 & n7160 ;
  assign n7162 = ( n315 & n4066 ) | ( n315 & ~n7161 ) | ( n4066 & ~n7161 ) ;
  assign n7175 = n5932 ^ n5779 ^ n620 ;
  assign n7167 = n2959 ^ n258 ^ 1'b0 ;
  assign n7168 = n3462 & n7167 ;
  assign n7169 = n723 & n7168 ;
  assign n7170 = ~n1456 & n7169 ;
  assign n7171 = ( ~n1478 & n5364 ) | ( ~n1478 & n7170 ) | ( n5364 & n7170 ) ;
  assign n7172 = ( ~n1120 & n4575 ) | ( ~n1120 & n7171 ) | ( n4575 & n7171 ) ;
  assign n7173 = n7172 ^ n5695 ^ n5378 ;
  assign n7174 = n7173 ^ n1391 ^ n1316 ;
  assign n7176 = n7175 ^ n7174 ^ n377 ;
  assign n7163 = n2752 ^ n289 ^ 1'b0 ;
  assign n7164 = n1203 & ~n7163 ;
  assign n7165 = n545 & n7164 ;
  assign n7166 = n7165 ^ n1213 ^ n304 ;
  assign n7177 = n7176 ^ n7166 ^ n2175 ;
  assign n7178 = n4787 ^ n3401 ^ n1696 ;
  assign n7179 = ( ~n611 & n6367 ) | ( ~n611 & n7178 ) | ( n6367 & n7178 ) ;
  assign n7184 = ( n908 & n3471 ) | ( n908 & ~n4178 ) | ( n3471 & ~n4178 ) ;
  assign n7185 = n6192 ^ n4420 ^ n1124 ;
  assign n7186 = ( ~n2288 & n7184 ) | ( ~n2288 & n7185 ) | ( n7184 & n7185 ) ;
  assign n7187 = n7186 ^ n2166 ^ n209 ;
  assign n7180 = n6808 ^ n2678 ^ n2479 ;
  assign n7181 = n5531 ^ n1994 ^ n1621 ;
  assign n7182 = ( n977 & n3555 ) | ( n977 & ~n7181 ) | ( n3555 & ~n7181 ) ;
  assign n7183 = ( ~n1103 & n7180 ) | ( ~n1103 & n7182 ) | ( n7180 & n7182 ) ;
  assign n7188 = n7187 ^ n7183 ^ n6655 ;
  assign n7192 = ~n1600 & n1663 ;
  assign n7189 = ( n4436 & n5227 ) | ( n4436 & n6485 ) | ( n5227 & n6485 ) ;
  assign n7190 = n3768 ^ n2941 ^ n1406 ;
  assign n7191 = n7189 & n7190 ;
  assign n7193 = n7192 ^ n7191 ^ 1'b0 ;
  assign n7194 = n5159 ^ n3167 ^ n1664 ;
  assign n7195 = ( n484 & ~n3461 ) | ( n484 & n3566 ) | ( ~n3461 & n3566 ) ;
  assign n7196 = ( n187 & n6607 ) | ( n187 & ~n7195 ) | ( n6607 & ~n7195 ) ;
  assign n7197 = n658 & n4099 ;
  assign n7198 = n7197 ^ n1075 ^ n199 ;
  assign n7199 = ( ~n7194 & n7196 ) | ( ~n7194 & n7198 ) | ( n7196 & n7198 ) ;
  assign n7205 = n5230 ^ n2853 ^ 1'b0 ;
  assign n7206 = n2228 & n7205 ;
  assign n7200 = ( ~x74 & n1697 ) | ( ~x74 & n5930 ) | ( n1697 & n5930 ) ;
  assign n7201 = ( n1979 & n5837 ) | ( n1979 & n7200 ) | ( n5837 & n7200 ) ;
  assign n7202 = n1116 | n7201 ;
  assign n7203 = n7202 ^ n5695 ^ n349 ;
  assign n7204 = ( n341 & n6180 ) | ( n341 & n7203 ) | ( n6180 & n7203 ) ;
  assign n7207 = n7206 ^ n7204 ^ n4087 ;
  assign n7208 = ( x46 & n292 ) | ( x46 & ~n2797 ) | ( n292 & ~n2797 ) ;
  assign n7209 = n7208 ^ n6473 ^ n6421 ;
  assign n7210 = ( n345 & ~n6757 ) | ( n345 & n7209 ) | ( ~n6757 & n7209 ) ;
  assign n7211 = n6842 ^ n2184 ^ 1'b0 ;
  assign n7212 = ( n4072 & n4718 ) | ( n4072 & n7211 ) | ( n4718 & n7211 ) ;
  assign n7213 = n2940 & ~n7202 ;
  assign n7214 = ~n7212 & n7213 ;
  assign n7215 = ( n399 & n7210 ) | ( n399 & n7214 ) | ( n7210 & n7214 ) ;
  assign n7216 = ( n887 & ~n992 ) | ( n887 & n1465 ) | ( ~n992 & n1465 ) ;
  assign n7217 = n6921 ^ n6646 ^ n3165 ;
  assign n7218 = ( ~n555 & n3767 ) | ( ~n555 & n7217 ) | ( n3767 & n7217 ) ;
  assign n7219 = ( n1820 & ~n7216 ) | ( n1820 & n7218 ) | ( ~n7216 & n7218 ) ;
  assign n7220 = n4480 & ~n4612 ;
  assign n7221 = ~n2322 & n7220 ;
  assign n7222 = ( n1742 & n1801 ) | ( n1742 & ~n4518 ) | ( n1801 & ~n4518 ) ;
  assign n7223 = n7222 ^ n164 ^ 1'b0 ;
  assign n7224 = n2026 & ~n7223 ;
  assign n7225 = n7224 ^ n5906 ^ n4154 ;
  assign n7226 = n5405 ^ n3828 ^ n1832 ;
  assign n7227 = n7226 ^ n4132 ^ n4076 ;
  assign n7229 = n933 ^ n779 ^ n528 ;
  assign n7228 = ( n334 & ~n817 ) | ( n334 & n2710 ) | ( ~n817 & n2710 ) ;
  assign n7230 = n7229 ^ n7228 ^ n2138 ;
  assign n7231 = ( ~n7225 & n7227 ) | ( ~n7225 & n7230 ) | ( n7227 & n7230 ) ;
  assign n7232 = ( n198 & n1615 ) | ( n198 & n3642 ) | ( n1615 & n3642 ) ;
  assign n7233 = ( x9 & ~n1079 ) | ( x9 & n6726 ) | ( ~n1079 & n6726 ) ;
  assign n7234 = ( n1141 & n1326 ) | ( n1141 & n7233 ) | ( n1326 & n7233 ) ;
  assign n7235 = ( ~n2274 & n7232 ) | ( ~n2274 & n7234 ) | ( n7232 & n7234 ) ;
  assign n7237 = ( x12 & ~n490 ) | ( x12 & n3465 ) | ( ~n490 & n3465 ) ;
  assign n7236 = n5499 ^ n2155 ^ 1'b0 ;
  assign n7238 = n7237 ^ n7236 ^ n4552 ;
  assign n7239 = ~n2722 & n6845 ;
  assign n7240 = n6988 & n7239 ;
  assign n7241 = ( n318 & n7076 ) | ( n318 & ~n7240 ) | ( n7076 & ~n7240 ) ;
  assign n7242 = ( ~n1300 & n1505 ) | ( ~n1300 & n6517 ) | ( n1505 & n6517 ) ;
  assign n7243 = ( n4003 & ~n4660 ) | ( n4003 & n7242 ) | ( ~n4660 & n7242 ) ;
  assign n7244 = n7243 ^ n2763 ^ n1935 ;
  assign n7245 = ( n567 & n2964 ) | ( n567 & ~n7244 ) | ( n2964 & ~n7244 ) ;
  assign n7246 = ( n1295 & n2254 ) | ( n1295 & n4013 ) | ( n2254 & n4013 ) ;
  assign n7247 = ( n575 & n4352 ) | ( n575 & n7246 ) | ( n4352 & n7246 ) ;
  assign n7248 = n4807 ^ n1764 ^ n1026 ;
  assign n7249 = n1390 ^ n491 ^ n437 ;
  assign n7250 = n1015 | n1138 ;
  assign n7251 = n7250 ^ n3263 ^ 1'b0 ;
  assign n7252 = x17 & n3403 ;
  assign n7253 = n7252 ^ n1306 ^ 1'b0 ;
  assign n7254 = ( n383 & n7251 ) | ( n383 & ~n7253 ) | ( n7251 & ~n7253 ) ;
  assign n7255 = ( n7248 & n7249 ) | ( n7248 & n7254 ) | ( n7249 & n7254 ) ;
  assign n7256 = ( n4258 & n6276 ) | ( n4258 & n7255 ) | ( n6276 & n7255 ) ;
  assign n7258 = ( n1702 & n3731 ) | ( n1702 & n6598 ) | ( n3731 & n6598 ) ;
  assign n7257 = n5405 ^ n4231 ^ n2836 ;
  assign n7259 = n7258 ^ n7257 ^ 1'b0 ;
  assign n7260 = n5530 ^ n1337 ^ n834 ;
  assign n7261 = ( ~n1083 & n7255 ) | ( ~n1083 & n7260 ) | ( n7255 & n7260 ) ;
  assign n7262 = ( n1886 & n2537 ) | ( n1886 & n6475 ) | ( n2537 & n6475 ) ;
  assign n7263 = ( n1507 & n2014 ) | ( n1507 & ~n5262 ) | ( n2014 & ~n5262 ) ;
  assign n7264 = ( n1124 & n5763 ) | ( n1124 & ~n7263 ) | ( n5763 & ~n7263 ) ;
  assign n7265 = n4858 ^ n2172 ^ n868 ;
  assign n7266 = n5359 ^ n1361 ^ n759 ;
  assign n7267 = ( n1091 & n7265 ) | ( n1091 & n7266 ) | ( n7265 & n7266 ) ;
  assign n7268 = ( n7262 & n7264 ) | ( n7262 & ~n7267 ) | ( n7264 & ~n7267 ) ;
  assign n7269 = n556 & n4569 ;
  assign n7270 = ~n2335 & n7269 ;
  assign n7271 = ( n1918 & n2146 ) | ( n1918 & n3378 ) | ( n2146 & n3378 ) ;
  assign n7272 = n6725 & n7271 ;
  assign n7273 = n7272 ^ n4158 ^ 1'b0 ;
  assign n7274 = n1708 | n6394 ;
  assign n7275 = ( n7270 & n7273 ) | ( n7270 & n7274 ) | ( n7273 & n7274 ) ;
  assign n7276 = ( n1169 & n2338 ) | ( n1169 & ~n6571 ) | ( n2338 & ~n6571 ) ;
  assign n7277 = ( ~n3012 & n4009 ) | ( ~n3012 & n4279 ) | ( n4009 & n4279 ) ;
  assign n7283 = n5016 ^ n3505 ^ n1713 ;
  assign n7278 = n3053 ^ n337 ^ x91 ;
  assign n7279 = n7278 ^ n5771 ^ n588 ;
  assign n7280 = n7279 ^ n4424 ^ 1'b0 ;
  assign n7281 = n7280 ^ n6444 ^ n1945 ;
  assign n7282 = n7281 ^ n2356 ^ n1915 ;
  assign n7284 = n7283 ^ n7282 ^ n2419 ;
  assign n7286 = n1955 ^ n1500 ^ 1'b0 ;
  assign n7287 = ~n961 & n7286 ;
  assign n7288 = n5191 & n7287 ;
  assign n7285 = n5564 ^ n1143 ^ 1'b0 ;
  assign n7289 = n7288 ^ n7285 ^ 1'b0 ;
  assign n7290 = n7284 | n7289 ;
  assign n7291 = n2017 & n6011 ;
  assign n7292 = ~n5022 & n7291 ;
  assign n7293 = n5158 ^ n4640 ^ n625 ;
  assign n7294 = n7293 ^ n5416 ^ 1'b0 ;
  assign n7295 = ( n373 & n7292 ) | ( n373 & ~n7294 ) | ( n7292 & ~n7294 ) ;
  assign n7296 = ( n302 & n3063 ) | ( n302 & ~n6505 ) | ( n3063 & ~n6505 ) ;
  assign n7304 = ( n1803 & ~n1999 ) | ( n1803 & n4546 ) | ( ~n1999 & n4546 ) ;
  assign n7301 = n1587 ^ n992 ^ n975 ;
  assign n7302 = ( n2470 & n4153 ) | ( n2470 & n7301 ) | ( n4153 & n7301 ) ;
  assign n7298 = n1380 ^ x64 ^ 1'b0 ;
  assign n7299 = x47 & ~n7298 ;
  assign n7300 = n7299 ^ n4784 ^ n1030 ;
  assign n7297 = n3767 ^ n2757 ^ n220 ;
  assign n7303 = n7302 ^ n7300 ^ n7297 ;
  assign n7305 = n7304 ^ n7303 ^ 1'b0 ;
  assign n7306 = n7305 ^ n2938 ^ 1'b0 ;
  assign n7324 = ( x55 & n987 ) | ( x55 & ~n1830 ) | ( n987 & ~n1830 ) ;
  assign n7325 = ( n1565 & ~n1874 ) | ( n1565 & n7324 ) | ( ~n1874 & n7324 ) ;
  assign n7326 = n7325 ^ n4822 ^ n1239 ;
  assign n7322 = n6793 ^ n5735 ^ n5549 ;
  assign n7323 = ( n2043 & ~n2698 ) | ( n2043 & n7322 ) | ( ~n2698 & n7322 ) ;
  assign n7327 = n7326 ^ n7323 ^ n349 ;
  assign n7328 = ( n564 & ~n4042 ) | ( n564 & n7327 ) | ( ~n4042 & n7327 ) ;
  assign n7307 = ( n2372 & n4279 ) | ( n2372 & n4685 ) | ( n4279 & n4685 ) ;
  assign n7308 = n3893 ^ n3795 ^ n1533 ;
  assign n7309 = ( n1089 & n2537 ) | ( n1089 & n7308 ) | ( n2537 & n7308 ) ;
  assign n7310 = n7309 ^ n3206 ^ n1158 ;
  assign n7311 = n7310 ^ n2168 ^ n2035 ;
  assign n7312 = n1522 | n4121 ;
  assign n7313 = n7312 ^ n1976 ^ 1'b0 ;
  assign n7314 = ( ~n243 & n2226 ) | ( ~n243 & n4682 ) | ( n2226 & n4682 ) ;
  assign n7315 = n6752 ^ n3841 ^ n282 ;
  assign n7316 = n7315 ^ n5126 ^ 1'b0 ;
  assign n7317 = n7314 & n7316 ;
  assign n7318 = ( n6429 & n7313 ) | ( n6429 & n7317 ) | ( n7313 & n7317 ) ;
  assign n7319 = ~n5005 & n7318 ;
  assign n7320 = n3297 & n7319 ;
  assign n7321 = ( n7307 & n7311 ) | ( n7307 & ~n7320 ) | ( n7311 & ~n7320 ) ;
  assign n7329 = n7328 ^ n7321 ^ x19 ;
  assign n7337 = n1199 & n1445 ;
  assign n7338 = n7337 ^ n3514 ^ n1080 ;
  assign n7330 = ( n566 & ~n5816 ) | ( n566 & n5913 ) | ( ~n5816 & n5913 ) ;
  assign n7331 = n7330 ^ n4638 ^ n2066 ;
  assign n7332 = n4530 ^ n2937 ^ n130 ;
  assign n7333 = ( x20 & ~n3004 ) | ( x20 & n7332 ) | ( ~n3004 & n7332 ) ;
  assign n7334 = n2550 | n7333 ;
  assign n7335 = n7334 ^ n4013 ^ n788 ;
  assign n7336 = ( ~n5135 & n7331 ) | ( ~n5135 & n7335 ) | ( n7331 & n7335 ) ;
  assign n7339 = n7338 ^ n7336 ^ n757 ;
  assign n7341 = ( ~x102 & n484 ) | ( ~x102 & n1700 ) | ( n484 & n1700 ) ;
  assign n7342 = n5233 ^ n2906 ^ n313 ;
  assign n7343 = n635 & ~n1615 ;
  assign n7344 = n7342 & n7343 ;
  assign n7345 = ( n1715 & n7341 ) | ( n1715 & n7344 ) | ( n7341 & n7344 ) ;
  assign n7346 = ( ~n3688 & n5088 ) | ( ~n3688 & n7345 ) | ( n5088 & n7345 ) ;
  assign n7347 = ( n1456 & ~n2076 ) | ( n1456 & n7346 ) | ( ~n2076 & n7346 ) ;
  assign n7340 = n1986 & ~n4595 ;
  assign n7348 = n7347 ^ n7340 ^ 1'b0 ;
  assign n7349 = ~x18 & n2665 ;
  assign n7350 = n7349 ^ n5323 ^ n5288 ;
  assign n7351 = ( n362 & n5389 ) | ( n362 & n7350 ) | ( n5389 & n7350 ) ;
  assign n7352 = ( n365 & n2316 ) | ( n365 & ~n7351 ) | ( n2316 & ~n7351 ) ;
  assign n7353 = ( n1831 & n2476 ) | ( n1831 & n7352 ) | ( n2476 & n7352 ) ;
  assign n7354 = ( x52 & n1421 ) | ( x52 & n4152 ) | ( n1421 & n4152 ) ;
  assign n7362 = n3931 ^ n729 ^ n608 ;
  assign n7363 = ( n1824 & ~n1930 ) | ( n1824 & n7362 ) | ( ~n1930 & n7362 ) ;
  assign n7364 = n7363 ^ n3841 ^ n2265 ;
  assign n7365 = ( ~n2562 & n3617 ) | ( ~n2562 & n7364 ) | ( n3617 & n7364 ) ;
  assign n7355 = ( n237 & n3792 ) | ( n237 & n4793 ) | ( n3792 & n4793 ) ;
  assign n7356 = n1532 ^ n800 ^ n534 ;
  assign n7357 = ( n4808 & n7355 ) | ( n4808 & ~n7356 ) | ( n7355 & ~n7356 ) ;
  assign n7358 = ( n1080 & n1502 ) | ( n1080 & ~n7357 ) | ( n1502 & ~n7357 ) ;
  assign n7359 = n7358 ^ n5407 ^ n908 ;
  assign n7360 = n7359 ^ n4137 ^ n949 ;
  assign n7361 = n7360 ^ n6364 ^ n3744 ;
  assign n7366 = n7365 ^ n7361 ^ n3302 ;
  assign n7367 = n7366 ^ n4042 ^ n3120 ;
  assign n7382 = n7090 ^ n744 ^ x30 ;
  assign n7381 = ( n740 & n1686 ) | ( n740 & ~n3367 ) | ( n1686 & ~n3367 ) ;
  assign n7383 = n7382 ^ n7381 ^ n910 ;
  assign n7374 = n3254 ^ n2039 ^ n1922 ;
  assign n7375 = ( n2656 & n4733 ) | ( n2656 & ~n7374 ) | ( n4733 & ~n7374 ) ;
  assign n7376 = x93 & ~n4878 ;
  assign n7377 = n7376 ^ n1620 ^ 1'b0 ;
  assign n7378 = ( ~n6421 & n6846 ) | ( ~n6421 & n7377 ) | ( n6846 & n7377 ) ;
  assign n7379 = n3280 ^ n2773 ^ x113 ;
  assign n7380 = ( ~n7375 & n7378 ) | ( ~n7375 & n7379 ) | ( n7378 & n7379 ) ;
  assign n7369 = n529 & ~n4500 ;
  assign n7368 = n1616 & n7299 ;
  assign n7370 = n7369 ^ n7368 ^ n5724 ;
  assign n7371 = ( n2749 & ~n4236 ) | ( n2749 & n6031 ) | ( ~n4236 & n6031 ) ;
  assign n7372 = n1925 | n7371 ;
  assign n7373 = ( ~n3567 & n7370 ) | ( ~n3567 & n7372 ) | ( n7370 & n7372 ) ;
  assign n7384 = n7383 ^ n7380 ^ n7373 ;
  assign n7385 = ( x82 & ~n2811 ) | ( x82 & n3931 ) | ( ~n2811 & n3931 ) ;
  assign n7392 = n3141 ^ n2081 ^ n175 ;
  assign n7388 = n3581 ^ n2620 ^ n283 ;
  assign n7387 = ( n1059 & ~n5962 ) | ( n1059 & n7009 ) | ( ~n5962 & n7009 ) ;
  assign n7389 = n7388 ^ n7387 ^ 1'b0 ;
  assign n7390 = n7389 ^ n5207 ^ n1986 ;
  assign n7391 = ( ~n3150 & n7305 ) | ( ~n3150 & n7390 ) | ( n7305 & n7390 ) ;
  assign n7386 = n6307 ^ n3752 ^ 1'b0 ;
  assign n7393 = n7392 ^ n7391 ^ n7386 ;
  assign n7394 = ( n2203 & ~n7385 ) | ( n2203 & n7393 ) | ( ~n7385 & n7393 ) ;
  assign n7395 = n4303 ^ n1211 ^ n700 ;
  assign n7396 = n5407 ^ n3315 ^ n2395 ;
  assign n7397 = ( n342 & n7395 ) | ( n342 & n7396 ) | ( n7395 & n7396 ) ;
  assign n7398 = n3319 ^ n1868 ^ n1833 ;
  assign n7399 = n7398 ^ n1554 ^ 1'b0 ;
  assign n7406 = n2396 & n4775 ;
  assign n7407 = ( n2104 & n2528 ) | ( n2104 & ~n5284 ) | ( n2528 & ~n5284 ) ;
  assign n7408 = ( n4290 & ~n7322 ) | ( n4290 & n7407 ) | ( ~n7322 & n7407 ) ;
  assign n7409 = ( ~n903 & n7406 ) | ( ~n903 & n7408 ) | ( n7406 & n7408 ) ;
  assign n7400 = ( n529 & ~n686 ) | ( n529 & n2958 ) | ( ~n686 & n2958 ) ;
  assign n7401 = ( ~n1747 & n3181 ) | ( ~n1747 & n7400 ) | ( n3181 & n7400 ) ;
  assign n7402 = ( n2964 & n6095 ) | ( n2964 & ~n7401 ) | ( n6095 & ~n7401 ) ;
  assign n7403 = n1517 ^ n1324 ^ n708 ;
  assign n7404 = n7403 ^ n5706 ^ n775 ;
  assign n7405 = ( n1475 & ~n7402 ) | ( n1475 & n7404 ) | ( ~n7402 & n7404 ) ;
  assign n7410 = n7409 ^ n7405 ^ n4730 ;
  assign n7412 = n7187 ^ n5339 ^ n2881 ;
  assign n7413 = ( n1653 & ~n2773 ) | ( n1653 & n7412 ) | ( ~n2773 & n7412 ) ;
  assign n7411 = ( n729 & ~n3912 ) | ( n729 & n5505 ) | ( ~n3912 & n5505 ) ;
  assign n7414 = n7413 ^ n7411 ^ n1379 ;
  assign n7415 = ( n2253 & n2749 ) | ( n2253 & ~n6926 ) | ( n2749 & ~n6926 ) ;
  assign n7416 = ( n734 & n4258 ) | ( n734 & n7415 ) | ( n4258 & n7415 ) ;
  assign n7417 = ( n4865 & ~n7414 ) | ( n4865 & n7416 ) | ( ~n7414 & n7416 ) ;
  assign n7418 = n1717 ^ n1164 ^ n772 ;
  assign n7419 = ( n1176 & ~n6338 ) | ( n1176 & n7418 ) | ( ~n6338 & n7418 ) ;
  assign n7420 = n4669 ^ n3548 ^ n2108 ;
  assign n7421 = n2039 | n7420 ;
  assign n7422 = n7419 | n7421 ;
  assign n7423 = n6519 ^ n4886 ^ n1902 ;
  assign n7424 = ( ~n3770 & n7422 ) | ( ~n3770 & n7423 ) | ( n7422 & n7423 ) ;
  assign n7425 = n6314 ^ n1237 ^ 1'b0 ;
  assign n7426 = ~n4254 & n7425 ;
  assign n7427 = n4684 & n7426 ;
  assign n7428 = n5799 ^ n3575 ^ n1321 ;
  assign n7431 = ( x29 & n3156 ) | ( x29 & ~n4304 ) | ( n3156 & ~n4304 ) ;
  assign n7429 = ( ~n5006 & n6092 ) | ( ~n5006 & n7051 ) | ( n6092 & n7051 ) ;
  assign n7430 = x90 & ~n7429 ;
  assign n7432 = n7431 ^ n7430 ^ 1'b0 ;
  assign n7433 = ( n1973 & n6658 ) | ( n1973 & ~n7432 ) | ( n6658 & ~n7432 ) ;
  assign n7434 = ( n1399 & n3763 ) | ( n1399 & n5417 ) | ( n3763 & n5417 ) ;
  assign n7435 = n7434 ^ n6612 ^ n6425 ;
  assign n7436 = ( ~n827 & n7393 ) | ( ~n827 & n7435 ) | ( n7393 & n7435 ) ;
  assign n7443 = ( n1004 & ~n1430 ) | ( n1004 & n3088 ) | ( ~n1430 & n3088 ) ;
  assign n7442 = ( n2379 & n4908 ) | ( n2379 & n6457 ) | ( n4908 & n6457 ) ;
  assign n7440 = n4775 ^ n4066 ^ n1977 ;
  assign n7437 = n6372 ^ n1832 ^ 1'b0 ;
  assign n7438 = ~n3142 & n7437 ;
  assign n7439 = ( n2879 & n4213 ) | ( n2879 & ~n7438 ) | ( n4213 & ~n7438 ) ;
  assign n7441 = n7440 ^ n7439 ^ n2830 ;
  assign n7444 = n7443 ^ n7442 ^ n7441 ;
  assign n7445 = ( ~n2521 & n3703 ) | ( ~n2521 & n5313 ) | ( n3703 & n5313 ) ;
  assign n7446 = n7445 ^ n5890 ^ n5708 ;
  assign n7447 = n6802 ^ n1172 ^ n292 ;
  assign n7448 = n7447 ^ n6397 ^ n2830 ;
  assign n7449 = n1787 | n6476 ;
  assign n7450 = n4892 | n7449 ;
  assign n7451 = ~n4853 & n7450 ;
  assign n7452 = ( x32 & n2014 ) | ( x32 & n2912 ) | ( n2014 & n2912 ) ;
  assign n7453 = n4309 | n7452 ;
  assign n7454 = n7453 ^ n3714 ^ 1'b0 ;
  assign n7455 = n7454 ^ n4483 ^ n4156 ;
  assign n7456 = n5794 ^ n2774 ^ n2744 ;
  assign n7457 = n2104 & n2335 ;
  assign n7458 = n7457 ^ n2734 ^ 1'b0 ;
  assign n7459 = n3898 ^ n3325 ^ 1'b0 ;
  assign n7460 = ( n2598 & n5669 ) | ( n2598 & ~n7459 ) | ( n5669 & ~n7459 ) ;
  assign n7461 = ( ~n2998 & n7458 ) | ( ~n2998 & n7460 ) | ( n7458 & n7460 ) ;
  assign n7462 = ( n6948 & ~n7456 ) | ( n6948 & n7461 ) | ( ~n7456 & n7461 ) ;
  assign n7463 = ~n7455 & n7462 ;
  assign n7464 = n7463 ^ n4683 ^ 1'b0 ;
  assign n7465 = ( n2952 & n3330 ) | ( n2952 & n3951 ) | ( n3330 & n3951 ) ;
  assign n7466 = ( n4079 & n4143 ) | ( n4079 & n7465 ) | ( n4143 & n7465 ) ;
  assign n7467 = n1819 ^ n1285 ^ n608 ;
  assign n7468 = ( n377 & ~n582 ) | ( n377 & n1979 ) | ( ~n582 & n1979 ) ;
  assign n7469 = ( n5110 & n7467 ) | ( n5110 & n7468 ) | ( n7467 & n7468 ) ;
  assign n7470 = n2514 ^ n2339 ^ n1245 ;
  assign n7471 = n4410 ^ n2113 ^ n986 ;
  assign n7472 = ( n1391 & n4196 ) | ( n1391 & n7471 ) | ( n4196 & n7471 ) ;
  assign n7473 = ( ~x109 & n7470 ) | ( ~x109 & n7472 ) | ( n7470 & n7472 ) ;
  assign n7474 = ( n1295 & n1576 ) | ( n1295 & n2239 ) | ( n1576 & n2239 ) ;
  assign n7475 = n7474 ^ n5532 ^ n370 ;
  assign n7476 = ( n1838 & n6889 ) | ( n1838 & ~n7475 ) | ( n6889 & ~n7475 ) ;
  assign n7480 = n5125 ^ n4696 ^ n1143 ;
  assign n7481 = ( n5634 & n6593 ) | ( n5634 & n7480 ) | ( n6593 & n7480 ) ;
  assign n7477 = n1953 ^ n1866 ^ n952 ;
  assign n7478 = ( n494 & ~n6801 ) | ( n494 & n7477 ) | ( ~n6801 & n7477 ) ;
  assign n7479 = ( n417 & n6738 ) | ( n417 & n7478 ) | ( n6738 & n7478 ) ;
  assign n7482 = n7481 ^ n7479 ^ 1'b0 ;
  assign n7483 = ~n7476 & n7482 ;
  assign n7484 = ~n4423 & n5011 ;
  assign n7485 = n2063 & ~n4754 ;
  assign n7486 = n7485 ^ n1559 ^ n863 ;
  assign n7488 = n6485 ^ n3851 ^ n2017 ;
  assign n7487 = ( n788 & n1771 ) | ( n788 & n3638 ) | ( n1771 & n3638 ) ;
  assign n7489 = n7488 ^ n7487 ^ n6126 ;
  assign n7490 = n4878 ^ n2194 ^ n1917 ;
  assign n7491 = n7490 ^ n581 ^ 1'b0 ;
  assign n7492 = ( n7486 & n7489 ) | ( n7486 & ~n7491 ) | ( n7489 & ~n7491 ) ;
  assign n7493 = ( n661 & n2534 ) | ( n661 & ~n2821 ) | ( n2534 & ~n2821 ) ;
  assign n7494 = n4223 ^ n3901 ^ n1724 ;
  assign n7495 = n7494 ^ n4742 ^ 1'b0 ;
  assign n7496 = ( n6004 & n7493 ) | ( n6004 & n7495 ) | ( n7493 & n7495 ) ;
  assign n7497 = ( n1902 & n3905 ) | ( n1902 & n6336 ) | ( n3905 & n6336 ) ;
  assign n7498 = ( x37 & n835 ) | ( x37 & n2204 ) | ( n835 & n2204 ) ;
  assign n7499 = ( n230 & n1012 ) | ( n230 & ~n7498 ) | ( n1012 & ~n7498 ) ;
  assign n7500 = ( n2211 & n3412 ) | ( n2211 & n7499 ) | ( n3412 & n7499 ) ;
  assign n7501 = ( n2316 & n3064 ) | ( n2316 & ~n7500 ) | ( n3064 & ~n7500 ) ;
  assign n7502 = ( n129 & n516 ) | ( n129 & ~n2232 ) | ( n516 & ~n2232 ) ;
  assign n7503 = n2108 ^ n1800 ^ 1'b0 ;
  assign n7504 = n7502 & n7503 ;
  assign n7505 = n2963 ^ n2316 ^ n1140 ;
  assign n7506 = n7505 ^ n1921 ^ n1846 ;
  assign n7507 = n7506 ^ n5504 ^ n3275 ;
  assign n7508 = ( n2891 & n7504 ) | ( n2891 & ~n7507 ) | ( n7504 & ~n7507 ) ;
  assign n7509 = n7501 | n7508 ;
  assign n7510 = n2042 & ~n7509 ;
  assign n7511 = n4841 ^ n2279 ^ n689 ;
  assign n7512 = n2085 | n7511 ;
  assign n7513 = ( n1175 & n4666 ) | ( n1175 & n7512 ) | ( n4666 & n7512 ) ;
  assign n7514 = n7513 ^ n5660 ^ 1'b0 ;
  assign n7517 = ( n2428 & ~n3770 ) | ( n2428 & n5718 ) | ( ~n3770 & n5718 ) ;
  assign n7518 = n7517 ^ n640 ^ x99 ;
  assign n7515 = x73 | n962 ;
  assign n7516 = ( n2347 & n7442 ) | ( n2347 & n7515 ) | ( n7442 & n7515 ) ;
  assign n7519 = n7518 ^ n7516 ^ n4135 ;
  assign n7520 = ( ~n6558 & n7514 ) | ( ~n6558 & n7519 ) | ( n7514 & n7519 ) ;
  assign n7521 = n7068 ^ n1303 ^ 1'b0 ;
  assign n7522 = x44 & ~n7521 ;
  assign n7523 = n5428 | n7522 ;
  assign n7524 = ( n2367 & n5692 ) | ( n2367 & n7253 ) | ( n5692 & n7253 ) ;
  assign n7531 = ( ~x96 & n212 ) | ( ~x96 & n2724 ) | ( n212 & n2724 ) ;
  assign n7532 = ( x28 & n331 ) | ( x28 & n7531 ) | ( n331 & n7531 ) ;
  assign n7533 = n7532 ^ n5145 ^ n138 ;
  assign n7529 = ( n888 & n4129 ) | ( n888 & n6543 ) | ( n4129 & n6543 ) ;
  assign n7530 = ( ~n2296 & n7325 ) | ( ~n2296 & n7529 ) | ( n7325 & n7529 ) ;
  assign n7525 = ( n2265 & n2969 ) | ( n2265 & n4281 ) | ( n2969 & n4281 ) ;
  assign n7526 = ( n2021 & n3374 ) | ( n2021 & ~n7525 ) | ( n3374 & ~n7525 ) ;
  assign n7527 = n7526 ^ n1765 ^ n1377 ;
  assign n7528 = ( ~n848 & n6804 ) | ( ~n848 & n7527 ) | ( n6804 & n7527 ) ;
  assign n7534 = n7533 ^ n7530 ^ n7528 ;
  assign n7536 = ( ~n2054 & n2539 ) | ( ~n2054 & n2609 ) | ( n2539 & n2609 ) ;
  assign n7537 = ( n624 & ~n4057 ) | ( n624 & n4966 ) | ( ~n4057 & n4966 ) ;
  assign n7538 = ~n7536 & n7537 ;
  assign n7535 = n6455 ^ n1854 ^ n1035 ;
  assign n7539 = n7538 ^ n7535 ^ 1'b0 ;
  assign n7540 = x4 | n1557 ;
  assign n7541 = n7540 ^ n1820 ^ 1'b0 ;
  assign n7542 = n7541 ^ n4996 ^ 1'b0 ;
  assign n7543 = ~n3473 & n7542 ;
  assign n7544 = ( n824 & ~n1710 ) | ( n824 & n7543 ) | ( ~n1710 & n7543 ) ;
  assign n7545 = ( x81 & n2779 ) | ( x81 & ~n3744 ) | ( n2779 & ~n3744 ) ;
  assign n7546 = n7545 ^ n4384 ^ n589 ;
  assign n7547 = n7546 ^ n6059 ^ n4302 ;
  assign n7548 = n7547 ^ n4824 ^ n479 ;
  assign n7549 = ( n7539 & ~n7544 ) | ( n7539 & n7548 ) | ( ~n7544 & n7548 ) ;
  assign n7550 = ( x95 & ~n2281 ) | ( x95 & n3466 ) | ( ~n2281 & n3466 ) ;
  assign n7551 = ( n3729 & n4229 ) | ( n3729 & ~n7550 ) | ( n4229 & ~n7550 ) ;
  assign n7552 = n5114 ^ n4694 ^ n2309 ;
  assign n7556 = n1801 ^ n1707 ^ n1363 ;
  assign n7557 = n7556 ^ n1704 ^ n818 ;
  assign n7558 = n1365 & n5389 ;
  assign n7559 = ( n1907 & ~n7557 ) | ( n1907 & n7558 ) | ( ~n7557 & n7558 ) ;
  assign n7553 = ( n203 & ~n803 ) | ( n203 & n2139 ) | ( ~n803 & n2139 ) ;
  assign n7554 = n6437 & ~n7553 ;
  assign n7555 = n4116 & n7554 ;
  assign n7560 = n7559 ^ n7555 ^ n4387 ;
  assign n7561 = ~n5268 & n7560 ;
  assign n7562 = n7561 ^ n904 ^ 1'b0 ;
  assign n7563 = ( ~n344 & n1121 ) | ( ~n344 & n1475 ) | ( n1121 & n1475 ) ;
  assign n7564 = ( n477 & n3260 ) | ( n477 & n4145 ) | ( n3260 & n4145 ) ;
  assign n7565 = ( ~n6079 & n6816 ) | ( ~n6079 & n7564 ) | ( n6816 & n7564 ) ;
  assign n7566 = ( n2254 & n7563 ) | ( n2254 & n7565 ) | ( n7563 & n7565 ) ;
  assign n7586 = n7537 ^ n6877 ^ n5512 ;
  assign n7584 = n1723 | n2535 ;
  assign n7585 = n1502 | n7584 ;
  assign n7587 = n7586 ^ n7585 ^ n6253 ;
  assign n7567 = n5777 ^ n4661 ^ n1603 ;
  assign n7568 = n7567 ^ n1490 ^ n1151 ;
  assign n7569 = ( n2015 & n6494 ) | ( n2015 & n7568 ) | ( n6494 & n7568 ) ;
  assign n7579 = n2082 ^ n1253 ^ 1'b0 ;
  assign n7580 = ( ~n1839 & n2558 ) | ( ~n1839 & n7579 ) | ( n2558 & n7579 ) ;
  assign n7575 = n867 & n1686 ;
  assign n7576 = n7575 ^ n932 ^ 1'b0 ;
  assign n7577 = n7576 ^ n2211 ^ n1921 ;
  assign n7573 = ( n988 & n1377 ) | ( n988 & ~n1447 ) | ( n1377 & ~n1447 ) ;
  assign n7574 = n7573 ^ n6627 ^ n1779 ;
  assign n7571 = n2834 ^ n2819 ^ n544 ;
  assign n7570 = n3544 ^ n1638 ^ n1502 ;
  assign n7572 = n7571 ^ n7570 ^ n2121 ;
  assign n7578 = n7577 ^ n7574 ^ n7572 ;
  assign n7581 = n7580 ^ n7578 ^ n4800 ;
  assign n7582 = ( n3438 & n7569 ) | ( n3438 & n7581 ) | ( n7569 & n7581 ) ;
  assign n7583 = ( n2402 & n2785 ) | ( n2402 & n7582 ) | ( n2785 & n7582 ) ;
  assign n7588 = n7587 ^ n7583 ^ 1'b0 ;
  assign n7589 = n7567 ^ n2964 ^ n2895 ;
  assign n7590 = n7589 ^ n7038 ^ n2858 ;
  assign n7591 = ( ~n3813 & n7434 ) | ( ~n3813 & n7590 ) | ( n7434 & n7590 ) ;
  assign n7592 = n6492 ^ n5706 ^ n5412 ;
  assign n7593 = ( x46 & ~n1992 ) | ( x46 & n2018 ) | ( ~n1992 & n2018 ) ;
  assign n7595 = n4607 ^ n2339 ^ n2179 ;
  assign n7594 = ( n1100 & ~n2462 ) | ( n1100 & n3764 ) | ( ~n2462 & n3764 ) ;
  assign n7596 = n7595 ^ n7594 ^ n3853 ;
  assign n7597 = ( ~n189 & n3446 ) | ( ~n189 & n7596 ) | ( n3446 & n7596 ) ;
  assign n7598 = ( n7592 & ~n7593 ) | ( n7592 & n7597 ) | ( ~n7593 & n7597 ) ;
  assign n7599 = ( n463 & n2385 ) | ( n463 & ~n3514 ) | ( n2385 & ~n3514 ) ;
  assign n7600 = n7599 ^ n3086 ^ 1'b0 ;
  assign n7601 = n6078 ^ n5287 ^ 1'b0 ;
  assign n7602 = n571 | n597 ;
  assign n7603 = ( ~n5575 & n7601 ) | ( ~n5575 & n7602 ) | ( n7601 & n7602 ) ;
  assign n7604 = n6845 ^ n1682 ^ n296 ;
  assign n7605 = n4868 ^ n710 ^ n661 ;
  assign n7606 = ( n2245 & n7604 ) | ( n2245 & ~n7605 ) | ( n7604 & ~n7605 ) ;
  assign n7607 = ( n1723 & n5257 ) | ( n1723 & ~n7606 ) | ( n5257 & ~n7606 ) ;
  assign n7608 = ( n701 & n4105 ) | ( n701 & n7607 ) | ( n4105 & n7607 ) ;
  assign n7609 = ( ~n7600 & n7603 ) | ( ~n7600 & n7608 ) | ( n7603 & n7608 ) ;
  assign n7610 = ( n1911 & n4864 ) | ( n1911 & ~n7609 ) | ( n4864 & ~n7609 ) ;
  assign n7611 = n3975 ^ n1880 ^ n471 ;
  assign n7612 = ( ~n2823 & n5234 ) | ( ~n2823 & n7611 ) | ( n5234 & n7611 ) ;
  assign n7613 = n7612 ^ n2573 ^ n200 ;
  assign n7618 = n1084 ^ n539 ^ x110 ;
  assign n7619 = ( n1499 & ~n3430 ) | ( n1499 & n7618 ) | ( ~n3430 & n7618 ) ;
  assign n7620 = ( n996 & ~n2116 ) | ( n996 & n5775 ) | ( ~n2116 & n5775 ) ;
  assign n7621 = n7620 ^ n5457 ^ n4228 ;
  assign n7622 = n7621 ^ n6118 ^ n4422 ;
  assign n7623 = ( n5065 & n7619 ) | ( n5065 & ~n7622 ) | ( n7619 & ~n7622 ) ;
  assign n7616 = ( n968 & ~n3186 ) | ( n968 & n4101 ) | ( ~n3186 & n4101 ) ;
  assign n7617 = ( n3259 & n4381 ) | ( n3259 & n7616 ) | ( n4381 & n7616 ) ;
  assign n7614 = ~n799 & n5610 ;
  assign n7615 = ( n3467 & n4944 ) | ( n3467 & ~n7614 ) | ( n4944 & ~n7614 ) ;
  assign n7624 = n7623 ^ n7617 ^ n7615 ;
  assign n7625 = ( ~n445 & n2392 ) | ( ~n445 & n2971 ) | ( n2392 & n2971 ) ;
  assign n7626 = n6648 ^ n861 ^ 1'b0 ;
  assign n7627 = ( n773 & n779 ) | ( n773 & n6317 ) | ( n779 & n6317 ) ;
  assign n7628 = ( ~n4661 & n7626 ) | ( ~n4661 & n7627 ) | ( n7626 & n7627 ) ;
  assign n7629 = n3133 | n7628 ;
  assign n7630 = n2609 ^ n209 ^ 1'b0 ;
  assign n7631 = n7629 | n7630 ;
  assign n7632 = ( n1690 & n7625 ) | ( n1690 & n7631 ) | ( n7625 & n7631 ) ;
  assign n7633 = ( n497 & n3742 ) | ( n497 & n5323 ) | ( n3742 & n5323 ) ;
  assign n7634 = ( x63 & n1094 ) | ( x63 & ~n7633 ) | ( n1094 & ~n7633 ) ;
  assign n7635 = n7558 ^ n2795 ^ n2509 ;
  assign n7636 = n449 & ~n7635 ;
  assign n7637 = n6897 & ~n7203 ;
  assign n7638 = n1244 & n7637 ;
  assign n7639 = ( n2881 & n3408 ) | ( n2881 & n7601 ) | ( n3408 & n7601 ) ;
  assign n7640 = ( n1689 & ~n7638 ) | ( n1689 & n7639 ) | ( ~n7638 & n7639 ) ;
  assign n7641 = n7640 ^ n5220 ^ n297 ;
  assign n7642 = n4168 ^ n3638 ^ n1336 ;
  assign n7643 = x81 & ~n7642 ;
  assign n7644 = n1514 & n7643 ;
  assign n7645 = n2824 ^ n2131 ^ n2062 ;
  assign n7646 = n7645 ^ n6324 ^ n2683 ;
  assign n7648 = n1733 ^ n681 ^ n199 ;
  assign n7649 = n7648 ^ n255 ^ 1'b0 ;
  assign n7647 = ( n2610 & n2784 ) | ( n2610 & ~n7356 ) | ( n2784 & ~n7356 ) ;
  assign n7650 = n7649 ^ n7647 ^ n5412 ;
  assign n7651 = n6587 ^ n1568 ^ 1'b0 ;
  assign n7652 = n6233 ^ n3349 ^ n1169 ;
  assign n7653 = n5041 & n7652 ;
  assign n7654 = ~n7651 & n7653 ;
  assign n7655 = n7654 ^ n3030 ^ n1692 ;
  assign n7656 = ( n5900 & n7650 ) | ( n5900 & ~n7655 ) | ( n7650 & ~n7655 ) ;
  assign n7657 = n7001 ^ n6216 ^ n2219 ;
  assign n7658 = ( x12 & n7184 ) | ( x12 & n7657 ) | ( n7184 & n7657 ) ;
  assign n7659 = n7658 ^ n2893 ^ n2757 ;
  assign n7660 = n2204 ^ n1958 ^ 1'b0 ;
  assign n7661 = n7660 ^ n1314 ^ n669 ;
  assign n7662 = n4720 & n7661 ;
  assign n7663 = n2340 ^ n801 ^ n562 ;
  assign n7664 = n5285 ^ n3225 ^ 1'b0 ;
  assign n7665 = n7663 & ~n7664 ;
  assign n7668 = ( n169 & n3404 ) | ( n169 & n6301 ) | ( n3404 & n6301 ) ;
  assign n7666 = ( n924 & n1274 ) | ( n924 & ~n5376 ) | ( n1274 & ~n5376 ) ;
  assign n7667 = n7666 ^ n7625 ^ n6383 ;
  assign n7669 = n7668 ^ n7667 ^ n5033 ;
  assign n7670 = ( n2415 & n7665 ) | ( n2415 & n7669 ) | ( n7665 & n7669 ) ;
  assign n7671 = ( ~n921 & n2141 ) | ( ~n921 & n4430 ) | ( n2141 & n4430 ) ;
  assign n7672 = ( ~n906 & n7670 ) | ( ~n906 & n7671 ) | ( n7670 & n7671 ) ;
  assign n7673 = n7672 ^ n6465 ^ 1'b0 ;
  assign n7674 = n4772 & n7673 ;
  assign n7680 = n1558 | n3789 ;
  assign n7681 = n7680 ^ n2947 ^ n2041 ;
  assign n7678 = ( n1442 & ~n2015 ) | ( n1442 & n2896 ) | ( ~n2015 & n2896 ) ;
  assign n7675 = ~n2339 & n2466 ;
  assign n7676 = ~x49 & n7675 ;
  assign n7677 = n4527 & ~n7676 ;
  assign n7679 = n7678 ^ n7677 ^ 1'b0 ;
  assign n7682 = n7681 ^ n7679 ^ n7206 ;
  assign n7683 = ( n2393 & ~n5249 ) | ( n2393 & n7001 ) | ( ~n5249 & n7001 ) ;
  assign n7684 = ( ~n1877 & n5703 ) | ( ~n1877 & n7683 ) | ( n5703 & n7683 ) ;
  assign n7685 = n4257 ^ n2354 ^ n228 ;
  assign n7686 = n3249 ^ n2953 ^ n1499 ;
  assign n7687 = ( ~n1499 & n2169 ) | ( ~n1499 & n7686 ) | ( n2169 & n7686 ) ;
  assign n7688 = n7687 ^ n6059 ^ n3063 ;
  assign n7689 = ~n7685 & n7688 ;
  assign n7690 = ~n1357 & n7689 ;
  assign n7691 = ~n956 & n7690 ;
  assign n7692 = ( n2228 & n2416 ) | ( n2228 & ~n2761 ) | ( n2416 & ~n2761 ) ;
  assign n7693 = n7692 ^ n280 ^ 1'b0 ;
  assign n7694 = ( ~x17 & n2156 ) | ( ~x17 & n7693 ) | ( n2156 & n7693 ) ;
  assign n7698 = n955 | n5530 ;
  assign n7695 = n173 | n2494 ;
  assign n7696 = ( n5177 & ~n5793 ) | ( n5177 & n6749 ) | ( ~n5793 & n6749 ) ;
  assign n7697 = ( n5685 & ~n7695 ) | ( n5685 & n7696 ) | ( ~n7695 & n7696 ) ;
  assign n7699 = n7698 ^ n7697 ^ n1780 ;
  assign n7700 = ( n7527 & n7694 ) | ( n7527 & n7699 ) | ( n7694 & n7699 ) ;
  assign n7701 = n5765 ^ n1436 ^ 1'b0 ;
  assign n7702 = ( x48 & n2825 ) | ( x48 & n6002 ) | ( n2825 & n6002 ) ;
  assign n7703 = n7702 ^ n4746 ^ 1'b0 ;
  assign n7704 = n4983 | n7703 ;
  assign n7709 = ( ~n1360 & n3047 ) | ( ~n1360 & n3828 ) | ( n3047 & n3828 ) ;
  assign n7710 = ( n1485 & n5823 ) | ( n1485 & ~n7709 ) | ( n5823 & ~n7709 ) ;
  assign n7706 = n1852 & n1865 ;
  assign n7707 = ( n3624 & n5719 ) | ( n3624 & ~n7706 ) | ( n5719 & ~n7706 ) ;
  assign n7708 = ( n986 & n6804 ) | ( n986 & n7707 ) | ( n6804 & n7707 ) ;
  assign n7711 = n7710 ^ n7708 ^ n3245 ;
  assign n7705 = n733 & n6098 ;
  assign n7712 = n7711 ^ n7705 ^ 1'b0 ;
  assign n7713 = ( ~n1816 & n2213 ) | ( ~n1816 & n6809 ) | ( n2213 & n6809 ) ;
  assign n7714 = n7713 ^ n3244 ^ 1'b0 ;
  assign n7717 = n4939 ^ n4395 ^ n3318 ;
  assign n7715 = ( n3381 & n5109 ) | ( n3381 & ~n6602 ) | ( n5109 & ~n6602 ) ;
  assign n7716 = n7715 ^ n7511 ^ n606 ;
  assign n7718 = n7717 ^ n7716 ^ n614 ;
  assign n7720 = n1654 ^ n470 ^ 1'b0 ;
  assign n7721 = n4017 & n7720 ;
  assign n7719 = n784 & ~n3922 ;
  assign n7722 = n7721 ^ n7719 ^ 1'b0 ;
  assign n7723 = ( n1162 & ~n3463 ) | ( n1162 & n4144 ) | ( ~n3463 & n4144 ) ;
  assign n7726 = n4487 ^ n3520 ^ n982 ;
  assign n7724 = n3104 ^ n858 ^ n819 ;
  assign n7725 = n7724 ^ n2620 ^ n2064 ;
  assign n7727 = n7726 ^ n7725 ^ n2762 ;
  assign n7728 = ( n7722 & n7723 ) | ( n7722 & ~n7727 ) | ( n7723 & ~n7727 ) ;
  assign n7730 = n197 & ~n5998 ;
  assign n7729 = n6600 ^ n2246 ^ n2176 ;
  assign n7731 = n7730 ^ n7729 ^ n5269 ;
  assign n7732 = n2826 | n7731 ;
  assign n7733 = n256 & n3572 ;
  assign n7734 = ( n2478 & ~n6781 ) | ( n2478 & n7733 ) | ( ~n6781 & n7733 ) ;
  assign n7735 = n424 & n7734 ;
  assign n7736 = n7735 ^ n963 ^ 1'b0 ;
  assign n7737 = n7041 ^ n5555 ^ n3201 ;
  assign n7738 = ( n280 & n348 ) | ( n280 & ~n1830 ) | ( n348 & ~n1830 ) ;
  assign n7739 = n3447 ^ n1879 ^ n714 ;
  assign n7740 = ( ~n6816 & n7738 ) | ( ~n6816 & n7739 ) | ( n7738 & n7739 ) ;
  assign n7741 = n7740 ^ n1972 ^ 1'b0 ;
  assign n7742 = n7737 | n7741 ;
  assign n7743 = ( n3716 & n3934 ) | ( n3716 & n4517 ) | ( n3934 & n4517 ) ;
  assign n7746 = ( n1506 & n2076 ) | ( n1506 & n5367 ) | ( n2076 & n5367 ) ;
  assign n7747 = n4487 ^ n3120 ^ 1'b0 ;
  assign n7748 = n7746 & ~n7747 ;
  assign n7744 = n5745 ^ n3318 ^ n1771 ;
  assign n7745 = ( ~n1319 & n3822 ) | ( ~n1319 & n7744 ) | ( n3822 & n7744 ) ;
  assign n7749 = n7748 ^ n7745 ^ 1'b0 ;
  assign n7750 = ( n3800 & ~n4500 ) | ( n3800 & n7749 ) | ( ~n4500 & n7749 ) ;
  assign n7751 = n479 | n1406 ;
  assign n7752 = ( n1596 & n2417 ) | ( n1596 & ~n7751 ) | ( n2417 & ~n7751 ) ;
  assign n7756 = n3673 ^ n2654 ^ x79 ;
  assign n7753 = ( n172 & n3701 ) | ( n172 & ~n4274 ) | ( n3701 & ~n4274 ) ;
  assign n7754 = n3039 | n3473 ;
  assign n7755 = n7753 & ~n7754 ;
  assign n7757 = n7756 ^ n7755 ^ n4877 ;
  assign n7758 = ( ~n2321 & n3821 ) | ( ~n2321 & n7757 ) | ( n3821 & n7757 ) ;
  assign n7759 = n3467 ^ n3286 ^ n983 ;
  assign n7760 = ( n7029 & ~n7758 ) | ( n7029 & n7759 ) | ( ~n7758 & n7759 ) ;
  assign n7761 = ( ~n1755 & n2009 ) | ( ~n1755 & n7760 ) | ( n2009 & n7760 ) ;
  assign n7762 = n7761 ^ n7628 ^ 1'b0 ;
  assign n7763 = n2082 | n3572 ;
  assign n7764 = n7198 ^ n4203 ^ n2189 ;
  assign n7767 = ( ~n2556 & n3452 ) | ( ~n2556 & n5448 ) | ( n3452 & n5448 ) ;
  assign n7766 = n4511 ^ n2345 ^ n285 ;
  assign n7765 = n2580 & ~n2992 ;
  assign n7768 = n7767 ^ n7766 ^ n7765 ;
  assign n7769 = ( n1863 & n5319 ) | ( n1863 & n5976 ) | ( n5319 & n5976 ) ;
  assign n7770 = x39 & n7769 ;
  assign n7771 = ~n6316 & n7770 ;
  assign n7772 = n3164 & ~n7601 ;
  assign n7773 = n7771 & n7772 ;
  assign n7774 = n7773 ^ n5826 ^ n563 ;
  assign n7775 = n3564 ^ x118 ^ 1'b0 ;
  assign n7776 = n7774 & ~n7775 ;
  assign n7784 = n1370 ^ n435 ^ x32 ;
  assign n7785 = ( n146 & n1788 ) | ( n146 & n2228 ) | ( n1788 & n2228 ) ;
  assign n7786 = ( n1566 & n7784 ) | ( n1566 & ~n7785 ) | ( n7784 & ~n7785 ) ;
  assign n7787 = n7786 ^ n7507 ^ n4251 ;
  assign n7783 = n6326 ^ n5332 ^ n2525 ;
  assign n7781 = n1524 ^ n617 ^ 1'b0 ;
  assign n7777 = n5456 ^ n2058 ^ n716 ;
  assign n7778 = n7777 ^ n4050 ^ n837 ;
  assign n7779 = ~n736 & n7778 ;
  assign n7780 = n7779 ^ n4426 ^ 1'b0 ;
  assign n7782 = n7781 ^ n7780 ^ n1757 ;
  assign n7788 = n7787 ^ n7783 ^ n7782 ;
  assign n7789 = n1630 | n7402 ;
  assign n7790 = n3170 | n7789 ;
  assign n7791 = ( n4067 & ~n5872 ) | ( n4067 & n7790 ) | ( ~n5872 & n7790 ) ;
  assign n7805 = n6819 ^ n3365 ^ n596 ;
  assign n7799 = ( n1707 & ~n2083 ) | ( n1707 & n4874 ) | ( ~n2083 & n4874 ) ;
  assign n7800 = n7317 ^ n6921 ^ n1153 ;
  assign n7801 = n7800 ^ n6152 ^ n1472 ;
  assign n7802 = n7801 ^ n7514 ^ n6672 ;
  assign n7803 = n7802 ^ n7158 ^ n147 ;
  assign n7804 = ( n5026 & ~n7799 ) | ( n5026 & n7803 ) | ( ~n7799 & n7803 ) ;
  assign n7797 = n2902 ^ n2581 ^ n575 ;
  assign n7792 = n4624 ^ n408 ^ n256 ;
  assign n7794 = n5051 ^ n3447 ^ n1314 ;
  assign n7793 = ( n1024 & n3234 ) | ( n1024 & ~n6143 ) | ( n3234 & ~n6143 ) ;
  assign n7795 = n7794 ^ n7793 ^ n2286 ;
  assign n7796 = ( n602 & ~n7792 ) | ( n602 & n7795 ) | ( ~n7792 & n7795 ) ;
  assign n7798 = n7797 ^ n7796 ^ n2610 ;
  assign n7806 = n7805 ^ n7804 ^ n7798 ;
  assign n7807 = n4539 ^ n3085 ^ n451 ;
  assign n7808 = ( n4053 & n7726 ) | ( n4053 & n7807 ) | ( n7726 & n7807 ) ;
  assign n7809 = ( n1700 & n6812 ) | ( n1700 & ~n7808 ) | ( n6812 & ~n7808 ) ;
  assign n7813 = n4704 ^ n2850 ^ n1112 ;
  assign n7814 = n7813 ^ n3533 ^ 1'b0 ;
  assign n7815 = ~n2731 & n7814 ;
  assign n7810 = n4178 ^ n692 ^ 1'b0 ;
  assign n7811 = n874 & ~n1257 ;
  assign n7812 = n7810 & n7811 ;
  assign n7816 = n7815 ^ n7812 ^ n6838 ;
  assign n7817 = n4695 & ~n6119 ;
  assign n7818 = ( n2637 & n3369 ) | ( n2637 & ~n7817 ) | ( n3369 & ~n7817 ) ;
  assign n7819 = n7818 ^ n1173 ^ 1'b0 ;
  assign n7820 = n7816 & n7819 ;
  assign n7821 = ( x99 & n3148 ) | ( x99 & n6175 ) | ( n3148 & n6175 ) ;
  assign n7822 = n2175 ^ n1934 ^ 1'b0 ;
  assign n7823 = n7822 ^ n7001 ^ n6062 ;
  assign n7824 = ( ~n881 & n2101 ) | ( ~n881 & n5301 ) | ( n2101 & n5301 ) ;
  assign n7825 = ( ~n4306 & n4327 ) | ( ~n4306 & n5062 ) | ( n4327 & n5062 ) ;
  assign n7826 = n7825 ^ n7237 ^ n1525 ;
  assign n7827 = n7826 ^ n7395 ^ n2653 ;
  assign n7828 = ( n6544 & ~n7606 ) | ( n6544 & n7827 ) | ( ~n7606 & n7827 ) ;
  assign n7829 = ( n4875 & ~n7824 ) | ( n4875 & n7828 ) | ( ~n7824 & n7828 ) ;
  assign n7830 = ( n6263 & n7823 ) | ( n6263 & n7829 ) | ( n7823 & n7829 ) ;
  assign n7832 = n3115 ^ n1935 ^ n749 ;
  assign n7833 = ( n134 & ~n364 ) | ( n134 & n7832 ) | ( ~n364 & n7832 ) ;
  assign n7831 = n1144 | n4800 ;
  assign n7834 = n7833 ^ n7831 ^ 1'b0 ;
  assign n7835 = ( n4138 & ~n6209 ) | ( n4138 & n7358 ) | ( ~n6209 & n7358 ) ;
  assign n7839 = n3777 ^ n2374 ^ n543 ;
  assign n7836 = ( n1203 & n2641 ) | ( n1203 & ~n4888 ) | ( n2641 & ~n4888 ) ;
  assign n7837 = n7836 ^ n6098 ^ n617 ;
  assign n7838 = ( ~n1544 & n4778 ) | ( ~n1544 & n7837 ) | ( n4778 & n7837 ) ;
  assign n7840 = n7839 ^ n7838 ^ n1467 ;
  assign n7841 = n4795 ^ n3588 ^ n804 ;
  assign n7842 = n239 & n7841 ;
  assign n7843 = ( ~n4178 & n5124 ) | ( ~n4178 & n5530 ) | ( n5124 & n5530 ) ;
  assign n7844 = n7843 ^ n6152 ^ n3944 ;
  assign n7845 = ( n3624 & n6143 ) | ( n3624 & n7403 ) | ( n6143 & n7403 ) ;
  assign n7846 = n6443 ^ x95 ^ 1'b0 ;
  assign n7847 = n1408 & ~n7846 ;
  assign n7848 = ( ~n1350 & n2676 ) | ( ~n1350 & n7365 ) | ( n2676 & n7365 ) ;
  assign n7849 = ( n2326 & n7847 ) | ( n2326 & ~n7848 ) | ( n7847 & ~n7848 ) ;
  assign n7854 = ( n2068 & n4064 ) | ( n2068 & ~n5858 ) | ( n4064 & ~n5858 ) ;
  assign n7850 = n6666 ^ n3232 ^ n2987 ;
  assign n7851 = n3716 ^ n2653 ^ n1315 ;
  assign n7852 = n7851 ^ n7391 ^ n4897 ;
  assign n7853 = ( n974 & n7850 ) | ( n974 & n7852 ) | ( n7850 & n7852 ) ;
  assign n7855 = n7854 ^ n7853 ^ n337 ;
  assign n7856 = n2117 ^ n984 ^ n625 ;
  assign n7866 = ( ~n417 & n1895 ) | ( ~n417 & n2472 ) | ( n1895 & n2472 ) ;
  assign n7865 = n6362 ^ n6315 ^ n3449 ;
  assign n7867 = n7866 ^ n7865 ^ n5896 ;
  assign n7857 = n5257 ^ n3635 ^ 1'b0 ;
  assign n7859 = n5254 ^ n3090 ^ n2923 ;
  assign n7858 = ( n2354 & ~n6146 ) | ( n2354 & n6643 ) | ( ~n6146 & n6643 ) ;
  assign n7860 = n7859 ^ n7858 ^ n6583 ;
  assign n7861 = n1211 & ~n1230 ;
  assign n7862 = n7860 & n7861 ;
  assign n7863 = ( n453 & n3836 ) | ( n453 & n5091 ) | ( n3836 & n5091 ) ;
  assign n7864 = ( n7857 & n7862 ) | ( n7857 & n7863 ) | ( n7862 & n7863 ) ;
  assign n7868 = n7867 ^ n7864 ^ n2716 ;
  assign n7877 = ( n3575 & ~n4413 ) | ( n3575 & n5076 ) | ( ~n4413 & n5076 ) ;
  assign n7870 = n5999 | n7287 ;
  assign n7871 = n7870 ^ n2079 ^ n1337 ;
  assign n7872 = n4728 ^ n4153 ^ 1'b0 ;
  assign n7873 = ~n7028 & n7872 ;
  assign n7874 = ( n6253 & n7871 ) | ( n6253 & ~n7873 ) | ( n7871 & ~n7873 ) ;
  assign n7875 = ( n2614 & ~n4694 ) | ( n2614 & n7874 ) | ( ~n4694 & n7874 ) ;
  assign n7869 = ( ~n226 & n931 ) | ( ~n226 & n6520 ) | ( n931 & n6520 ) ;
  assign n7876 = n7875 ^ n7869 ^ n201 ;
  assign n7878 = n7877 ^ n7876 ^ n3103 ;
  assign n7884 = n5224 ^ n3504 ^ n2048 ;
  assign n7882 = n4475 | n6547 ;
  assign n7883 = n447 | n7882 ;
  assign n7885 = n7884 ^ n7883 ^ n737 ;
  assign n7879 = n6812 ^ n2657 ^ n2467 ;
  assign n7880 = n7879 ^ n7638 ^ n2838 ;
  assign n7881 = n5779 & n7880 ;
  assign n7886 = n7885 ^ n7881 ^ 1'b0 ;
  assign n7887 = n401 | n5480 ;
  assign n7888 = n7887 ^ n7182 ^ n915 ;
  assign n7889 = n1839 & ~n4916 ;
  assign n7890 = n7889 ^ n642 ^ 1'b0 ;
  assign n7891 = ( n6338 & n7888 ) | ( n6338 & ~n7890 ) | ( n7888 & ~n7890 ) ;
  assign n7892 = n7891 ^ n2117 ^ n796 ;
  assign n7893 = n2228 ^ n2062 ^ n1024 ;
  assign n7894 = ( n3964 & ~n5475 ) | ( n3964 & n7893 ) | ( ~n5475 & n7893 ) ;
  assign n7895 = ( x73 & ~n606 ) | ( x73 & n2550 ) | ( ~n606 & n2550 ) ;
  assign n7896 = n7895 ^ n2181 ^ n1724 ;
  assign n7897 = ( ~n2587 & n4387 ) | ( ~n2587 & n6271 ) | ( n4387 & n6271 ) ;
  assign n7898 = n7897 ^ n2745 ^ 1'b0 ;
  assign n7899 = n7898 ^ n7854 ^ n3930 ;
  assign n7900 = n6158 ^ n2731 ^ 1'b0 ;
  assign n7901 = n7899 | n7900 ;
  assign n7902 = ( n832 & n1601 ) | ( n832 & n4711 ) | ( n1601 & n4711 ) ;
  assign n7903 = n7611 ^ n3390 ^ n2119 ;
  assign n7904 = n3113 ^ n2338 ^ n1226 ;
  assign n7905 = ( n7648 & n7903 ) | ( n7648 & n7904 ) | ( n7903 & n7904 ) ;
  assign n7906 = ~n2201 & n3682 ;
  assign n7907 = ( ~n1128 & n7905 ) | ( ~n1128 & n7906 ) | ( n7905 & n7906 ) ;
  assign n7908 = ( n847 & n2140 ) | ( n847 & ~n3645 ) | ( n2140 & ~n3645 ) ;
  assign n7909 = n7908 ^ n2887 ^ n673 ;
  assign n7916 = n1254 ^ n984 ^ n498 ;
  assign n7910 = n1716 ^ n683 ^ n632 ;
  assign n7911 = n7887 ^ n2775 ^ 1'b0 ;
  assign n7912 = n5857 ^ n1684 ^ n1427 ;
  assign n7913 = n7912 ^ n3060 ^ 1'b0 ;
  assign n7914 = ~n2928 & n7913 ;
  assign n7915 = ( n7910 & n7911 ) | ( n7910 & ~n7914 ) | ( n7911 & ~n7914 ) ;
  assign n7917 = n7916 ^ n7915 ^ n3897 ;
  assign n7918 = n7917 ^ n2537 ^ n2393 ;
  assign n7919 = ( n4176 & n7909 ) | ( n4176 & ~n7918 ) | ( n7909 & ~n7918 ) ;
  assign n7920 = n4541 ^ n2073 ^ n366 ;
  assign n7921 = ( n2565 & ~n7635 ) | ( n2565 & n7920 ) | ( ~n7635 & n7920 ) ;
  assign n7923 = n3633 ^ n2441 ^ n2127 ;
  assign n7924 = n7923 ^ n2360 ^ 1'b0 ;
  assign n7922 = ( ~n1335 & n3709 ) | ( ~n1335 & n7813 ) | ( n3709 & n7813 ) ;
  assign n7925 = n7924 ^ n7922 ^ n4197 ;
  assign n7926 = n7925 ^ n3121 ^ n880 ;
  assign n7927 = ( ~n6283 & n7465 ) | ( ~n6283 & n7926 ) | ( n7465 & n7926 ) ;
  assign n7928 = ( n2575 & n7921 ) | ( n2575 & n7927 ) | ( n7921 & n7927 ) ;
  assign n7929 = n7388 ^ n2940 ^ n547 ;
  assign n7930 = n5785 ^ n4380 ^ n2141 ;
  assign n7931 = n7317 ^ n4274 ^ n1415 ;
  assign n7932 = n7931 ^ n5459 ^ n2596 ;
  assign n7933 = ( x76 & ~n7930 ) | ( x76 & n7932 ) | ( ~n7930 & n7932 ) ;
  assign n7934 = ( n1670 & n2317 ) | ( n1670 & n7933 ) | ( n2317 & n7933 ) ;
  assign n7935 = n4644 ^ n4298 ^ n697 ;
  assign n7936 = ( n7929 & ~n7934 ) | ( n7929 & n7935 ) | ( ~n7934 & n7935 ) ;
  assign n7938 = n6774 ^ n2917 ^ n1378 ;
  assign n7939 = n7938 ^ n2612 ^ n1712 ;
  assign n7940 = ( ~n1685 & n5904 ) | ( ~n1685 & n7939 ) | ( n5904 & n7939 ) ;
  assign n7937 = ( n2748 & n4528 ) | ( n2748 & n7378 ) | ( n4528 & n7378 ) ;
  assign n7941 = n7940 ^ n7937 ^ n1429 ;
  assign n7942 = ( n353 & n1137 ) | ( n353 & n3829 ) | ( n1137 & n3829 ) ;
  assign n7943 = n7942 ^ n7148 ^ n2908 ;
  assign n7944 = n6200 ^ n3558 ^ n1988 ;
  assign n7945 = n7944 ^ n2869 ^ x48 ;
  assign n7946 = ( n994 & ~n2260 ) | ( n994 & n7945 ) | ( ~n2260 & n7945 ) ;
  assign n7947 = n1520 ^ n1280 ^ n317 ;
  assign n7948 = n7947 ^ n6428 ^ n3964 ;
  assign n7949 = n7948 ^ n3069 ^ n1184 ;
  assign n7950 = ( n2608 & n3935 ) | ( n2608 & n7949 ) | ( n3935 & n7949 ) ;
  assign n7951 = ( ~n1321 & n3369 ) | ( ~n1321 & n4546 ) | ( n3369 & n4546 ) ;
  assign n7952 = ( n5847 & n7604 ) | ( n5847 & n7951 ) | ( n7604 & n7951 ) ;
  assign n7953 = ( ~n1609 & n4433 ) | ( ~n1609 & n7952 ) | ( n4433 & n7952 ) ;
  assign n7954 = ( n4650 & ~n7950 ) | ( n4650 & n7953 ) | ( ~n7950 & n7953 ) ;
  assign n7955 = n6213 ^ n3668 ^ 1'b0 ;
  assign n7956 = n3930 & ~n7955 ;
  assign n7958 = n4475 | n5900 ;
  assign n7957 = n2718 | n7104 ;
  assign n7959 = n7958 ^ n7957 ^ n3733 ;
  assign n7960 = ( ~n3672 & n7956 ) | ( ~n3672 & n7959 ) | ( n7956 & n7959 ) ;
  assign n7961 = ( n2213 & n5836 ) | ( n2213 & n6763 ) | ( n5836 & n6763 ) ;
  assign n7962 = n7961 ^ n7081 ^ n1413 ;
  assign n7963 = n3234 ^ n3158 ^ n1085 ;
  assign n7964 = ( n1811 & ~n5456 ) | ( n1811 & n7963 ) | ( ~n5456 & n7963 ) ;
  assign n7965 = ( n893 & n3778 ) | ( n893 & n7964 ) | ( n3778 & n7964 ) ;
  assign n7966 = n6486 ^ n2083 ^ n1572 ;
  assign n7967 = ( n3236 & n3904 ) | ( n3236 & n5167 ) | ( n3904 & n5167 ) ;
  assign n7968 = ( n882 & ~n7201 ) | ( n882 & n7967 ) | ( ~n7201 & n7967 ) ;
  assign n7969 = ( n145 & ~n7966 ) | ( n145 & n7968 ) | ( ~n7966 & n7968 ) ;
  assign n7970 = ( ~n4525 & n7965 ) | ( ~n4525 & n7969 ) | ( n7965 & n7969 ) ;
  assign n7971 = ( n1169 & ~n4474 ) | ( n1169 & n7967 ) | ( ~n4474 & n7967 ) ;
  assign n7972 = n1032 | n7971 ;
  assign n7973 = n2563 & n7972 ;
  assign n7974 = ~n1049 & n7973 ;
  assign n7975 = ~n3153 & n5316 ;
  assign n7976 = n7975 ^ n5056 ^ 1'b0 ;
  assign n7977 = n7976 ^ n7925 ^ n6335 ;
  assign n7978 = n3138 ^ n2330 ^ n1473 ;
  assign n7979 = n2470 ^ n995 ^ 1'b0 ;
  assign n7980 = n7979 ^ n4120 ^ n2349 ;
  assign n7981 = n7980 ^ n7594 ^ n2060 ;
  assign n7982 = n7978 & ~n7981 ;
  assign n7983 = ~n4424 & n7982 ;
  assign n7984 = ( ~n3105 & n6705 ) | ( ~n3105 & n7983 ) | ( n6705 & n7983 ) ;
  assign n7985 = ( n796 & n1741 ) | ( n796 & ~n2015 ) | ( n1741 & ~n2015 ) ;
  assign n7986 = n7985 ^ n4371 ^ n2536 ;
  assign n7988 = n957 ^ n839 ^ n563 ;
  assign n7987 = n1979 ^ n749 ^ 1'b0 ;
  assign n7989 = n7988 ^ n7987 ^ x97 ;
  assign n7990 = n6042 ^ n2390 ^ n2123 ;
  assign n7991 = n7990 ^ n2696 ^ n1760 ;
  assign n7992 = ( n381 & n1207 ) | ( n381 & ~n7991 ) | ( n1207 & ~n7991 ) ;
  assign n7993 = ( n7826 & ~n7989 ) | ( n7826 & n7992 ) | ( ~n7989 & n7992 ) ;
  assign n8006 = n4867 ^ n1099 ^ x25 ;
  assign n8001 = x96 & n5846 ;
  assign n8002 = n8001 ^ n1827 ^ 1'b0 ;
  assign n8003 = n6911 ^ n5149 ^ n2770 ;
  assign n8004 = n8003 ^ n4570 ^ n2152 ;
  assign n8005 = ( ~n3431 & n8002 ) | ( ~n3431 & n8004 ) | ( n8002 & n8004 ) ;
  assign n7996 = n4120 | n5077 ;
  assign n7997 = n883 | n7996 ;
  assign n7998 = ( ~n3285 & n4876 ) | ( ~n3285 & n7997 ) | ( n4876 & n7997 ) ;
  assign n7995 = n1831 ^ n235 ^ 1'b0 ;
  assign n7999 = n7998 ^ n7995 ^ 1'b0 ;
  assign n7994 = n3937 ^ n1330 ^ n1204 ;
  assign n8000 = n7999 ^ n7994 ^ n3888 ;
  assign n8007 = n8006 ^ n8005 ^ n8000 ;
  assign n8019 = n6833 ^ n3930 ^ n582 ;
  assign n8020 = ( n2101 & n5496 ) | ( n2101 & ~n8019 ) | ( n5496 & ~n8019 ) ;
  assign n8011 = n3424 ^ n3304 ^ n1239 ;
  assign n8008 = ( n2154 & n3272 ) | ( n2154 & ~n4487 ) | ( n3272 & ~n4487 ) ;
  assign n8012 = n3677 | n7477 ;
  assign n8013 = n3170 | n8012 ;
  assign n8014 = n689 & n8013 ;
  assign n8015 = ~n8008 & n8014 ;
  assign n8016 = n7545 ^ n2112 ^ n1270 ;
  assign n8017 = ( n8011 & ~n8015 ) | ( n8011 & n8016 ) | ( ~n8015 & n8016 ) ;
  assign n8009 = n6909 & n8008 ;
  assign n8010 = n8009 ^ n3460 ^ n1486 ;
  assign n8018 = n8017 ^ n8010 ^ n1341 ;
  assign n8021 = n8020 ^ n8018 ^ n3693 ;
  assign n8028 = ( n274 & n1041 ) | ( n274 & n4954 ) | ( n1041 & n4954 ) ;
  assign n8029 = n8028 ^ n3304 ^ n3239 ;
  assign n8026 = ( n4576 & n5791 ) | ( n4576 & ~n7308 ) | ( n5791 & ~n7308 ) ;
  assign n8027 = ~n1680 & n8026 ;
  assign n8030 = n8029 ^ n8027 ^ 1'b0 ;
  assign n8025 = n7363 ^ n1770 ^ n1586 ;
  assign n8023 = ( ~n2326 & n2369 ) | ( ~n2326 & n3318 ) | ( n2369 & n3318 ) ;
  assign n8022 = n1091 & ~n1457 ;
  assign n8024 = n8023 ^ n8022 ^ 1'b0 ;
  assign n8031 = n8030 ^ n8025 ^ n8024 ;
  assign n8032 = ( x15 & n6011 ) | ( x15 & n8031 ) | ( n6011 & n8031 ) ;
  assign n8035 = n2993 ^ n1116 ^ n474 ;
  assign n8034 = ( n1008 & n4624 ) | ( n1008 & n6434 ) | ( n4624 & n6434 ) ;
  assign n8036 = n8035 ^ n8034 ^ n6315 ;
  assign n8033 = ( n1372 & ~n4148 ) | ( n1372 & n5934 ) | ( ~n4148 & n5934 ) ;
  assign n8037 = n8036 ^ n8033 ^ n5055 ;
  assign n8038 = n1354 | n7910 ;
  assign n8039 = n5020 ^ n3947 ^ n1609 ;
  assign n8040 = ( n3543 & n3905 ) | ( n3543 & ~n8039 ) | ( n3905 & ~n8039 ) ;
  assign n8041 = ( n868 & n7687 ) | ( n868 & ~n8040 ) | ( n7687 & ~n8040 ) ;
  assign n8042 = ( n517 & n6130 ) | ( n517 & n8041 ) | ( n6130 & n8041 ) ;
  assign n8043 = n806 ^ n385 ^ n206 ;
  assign n8044 = n8043 ^ n7698 ^ n1702 ;
  assign n8045 = ( x16 & ~n7871 ) | ( x16 & n8044 ) | ( ~n7871 & n8044 ) ;
  assign n8046 = n2536 ^ n1799 ^ n1757 ;
  assign n8047 = n2649 ^ n621 ^ n497 ;
  assign n8048 = n8047 ^ n6320 ^ n1090 ;
  assign n8049 = n8048 ^ n7287 ^ 1'b0 ;
  assign n8050 = ~n6458 & n8049 ;
  assign n8051 = ( ~n4038 & n8046 ) | ( ~n4038 & n8050 ) | ( n8046 & n8050 ) ;
  assign n8053 = n3996 ^ n1321 ^ n951 ;
  assign n8054 = n8053 ^ n3377 ^ x95 ;
  assign n8055 = ( ~x97 & n5754 ) | ( ~x97 & n5846 ) | ( n5754 & n5846 ) ;
  assign n8056 = n8055 ^ n3961 ^ n198 ;
  assign n8057 = ( n2887 & ~n4608 ) | ( n2887 & n8056 ) | ( ~n4608 & n8056 ) ;
  assign n8058 = n7625 | n8057 ;
  assign n8059 = n8058 ^ n1444 ^ 1'b0 ;
  assign n8060 = n8059 ^ n7317 ^ n1772 ;
  assign n8061 = n8060 ^ n5805 ^ n4964 ;
  assign n8062 = ( ~n408 & n8054 ) | ( ~n408 & n8061 ) | ( n8054 & n8061 ) ;
  assign n8052 = n2269 ^ n616 ^ x22 ;
  assign n8063 = n8062 ^ n8052 ^ n6971 ;
  assign n8064 = ( n435 & n2680 ) | ( n435 & ~n3349 ) | ( n2680 & ~n3349 ) ;
  assign n8065 = ( x99 & ~n685 ) | ( x99 & n2080 ) | ( ~n685 & n2080 ) ;
  assign n8066 = n8064 | n8065 ;
  assign n8067 = n7342 ^ n6797 ^ n5495 ;
  assign n8068 = ( x7 & ~n4682 ) | ( x7 & n5398 ) | ( ~n4682 & n5398 ) ;
  assign n8069 = n1717 ^ n990 ^ 1'b0 ;
  assign n8070 = n8068 | n8069 ;
  assign n8071 = ( n5035 & ~n6536 ) | ( n5035 & n8070 ) | ( ~n6536 & n8070 ) ;
  assign n8072 = n8071 ^ n7005 ^ n5699 ;
  assign n8073 = ~n1474 & n3230 ;
  assign n8074 = n767 ^ n240 ^ n164 ;
  assign n8075 = ( ~n1263 & n8073 ) | ( ~n1263 & n8074 ) | ( n8073 & n8074 ) ;
  assign n8076 = n8075 ^ n7119 ^ n5512 ;
  assign n8083 = n3361 ^ n2332 ^ n517 ;
  assign n8084 = n8083 ^ n735 ^ n254 ;
  assign n8082 = n5092 ^ n2997 ^ n2701 ;
  assign n8078 = n1383 ^ n644 ^ n475 ;
  assign n8077 = n2259 & ~n5808 ;
  assign n8079 = n8078 ^ n8077 ^ 1'b0 ;
  assign n8080 = n4359 ^ n3822 ^ 1'b0 ;
  assign n8081 = n8079 | n8080 ;
  assign n8085 = n8084 ^ n8082 ^ n8081 ;
  assign n8091 = n3882 ^ n1032 ^ n637 ;
  assign n8090 = ( n1703 & n2833 ) | ( n1703 & ~n6492 ) | ( n2833 & ~n6492 ) ;
  assign n8092 = n8091 ^ n8090 ^ n6054 ;
  assign n8093 = ( ~n676 & n1087 ) | ( ~n676 & n8092 ) | ( n1087 & n8092 ) ;
  assign n8086 = ( n2505 & n3788 ) | ( n2505 & n5245 ) | ( n3788 & n5245 ) ;
  assign n8087 = ( ~n469 & n740 ) | ( ~n469 & n8086 ) | ( n740 & n8086 ) ;
  assign n8088 = n8087 ^ n4443 ^ 1'b0 ;
  assign n8089 = n7558 | n8088 ;
  assign n8094 = n8093 ^ n8089 ^ n6629 ;
  assign n8095 = n6076 ^ n4142 ^ n603 ;
  assign n8096 = n8095 ^ n2642 ^ x69 ;
  assign n8097 = n7676 ^ n6846 ^ n2530 ;
  assign n8098 = n8097 ^ n882 ^ 1'b0 ;
  assign n8099 = ( n3102 & ~n8096 ) | ( n3102 & n8098 ) | ( ~n8096 & n8098 ) ;
  assign n8100 = ( n1801 & ~n2290 ) | ( n1801 & n3035 ) | ( ~n2290 & n3035 ) ;
  assign n8101 = ( n3865 & n6922 ) | ( n3865 & ~n8100 ) | ( n6922 & ~n8100 ) ;
  assign n8102 = ( n723 & n3751 ) | ( n723 & ~n8101 ) | ( n3751 & ~n8101 ) ;
  assign n8103 = ( n1558 & n3012 ) | ( n1558 & n4023 ) | ( n3012 & n4023 ) ;
  assign n8104 = ( n622 & ~n3930 ) | ( n622 & n8103 ) | ( ~n3930 & n8103 ) ;
  assign n8105 = n3040 & ~n4646 ;
  assign n8106 = n8105 ^ n7619 ^ 1'b0 ;
  assign n8107 = ( n3809 & ~n5997 ) | ( n3809 & n8106 ) | ( ~n5997 & n8106 ) ;
  assign n8108 = n8107 ^ n2328 ^ 1'b0 ;
  assign n8109 = n8104 & ~n8108 ;
  assign n8110 = ( n2610 & n8102 ) | ( n2610 & ~n8109 ) | ( n8102 & ~n8109 ) ;
  assign n8111 = n4038 ^ n3488 ^ 1'b0 ;
  assign n8112 = n5180 & ~n8111 ;
  assign n8113 = ( n5291 & n6567 ) | ( n5291 & ~n8112 ) | ( n6567 & ~n8112 ) ;
  assign n8122 = n1710 ^ n582 ^ 1'b0 ;
  assign n8119 = ( n1717 & n1979 ) | ( n1717 & n2487 ) | ( n1979 & n2487 ) ;
  assign n8116 = n3220 & ~n6602 ;
  assign n8117 = n8116 ^ n5834 ^ 1'b0 ;
  assign n8114 = ( n803 & n973 ) | ( n803 & n1823 ) | ( n973 & n1823 ) ;
  assign n8115 = ( ~n191 & n771 ) | ( ~n191 & n8114 ) | ( n771 & n8114 ) ;
  assign n8118 = n8117 ^ n8115 ^ x37 ;
  assign n8120 = n8119 ^ n8118 ^ n3241 ;
  assign n8121 = n2452 & ~n8120 ;
  assign n8123 = n8122 ^ n8121 ^ 1'b0 ;
  assign n8125 = n521 | n3138 ;
  assign n8126 = n8125 ^ n1247 ^ 1'b0 ;
  assign n8124 = n1861 & n7470 ;
  assign n8127 = n8126 ^ n8124 ^ n3223 ;
  assign n8128 = n762 ^ n566 ^ 1'b0 ;
  assign n8129 = n3561 & ~n8128 ;
  assign n8130 = n8129 ^ n198 ^ 1'b0 ;
  assign n8131 = n7479 ^ n3963 ^ n1271 ;
  assign n8132 = n219 & n662 ;
  assign n8133 = ~n8131 & n8132 ;
  assign n8134 = n4002 ^ n3719 ^ n1629 ;
  assign n8135 = n8134 ^ n4916 ^ n2326 ;
  assign n8136 = ~n4985 & n8135 ;
  assign n8137 = ~n4238 & n8136 ;
  assign n8138 = ( n1295 & n2450 ) | ( n1295 & ~n3234 ) | ( n2450 & ~n3234 ) ;
  assign n8139 = ( ~n653 & n780 ) | ( ~n653 & n8138 ) | ( n780 & n8138 ) ;
  assign n8140 = n8139 ^ n4199 ^ n3748 ;
  assign n8141 = n2124 & ~n8140 ;
  assign n8142 = ( n1012 & n2048 ) | ( n1012 & ~n7683 ) | ( n2048 & ~n7683 ) ;
  assign n8143 = n6509 & ~n8142 ;
  assign n8144 = n8026 ^ n4742 ^ n2142 ;
  assign n8145 = ( n728 & n3566 ) | ( n728 & n8144 ) | ( n3566 & n8144 ) ;
  assign n8146 = n5795 ^ n1333 ^ 1'b0 ;
  assign n8147 = n7594 & ~n8146 ;
  assign n8149 = n2200 ^ n286 ^ n249 ;
  assign n8148 = n6031 ^ n3414 ^ n1260 ;
  assign n8150 = n8149 ^ n8148 ^ n4102 ;
  assign n8151 = ( n429 & n3509 ) | ( n429 & ~n3759 ) | ( n3509 & ~n3759 ) ;
  assign n8154 = n6109 ^ n4620 ^ n3514 ;
  assign n8152 = n238 | n319 ;
  assign n8153 = n1625 | n8152 ;
  assign n8155 = n8154 ^ n8153 ^ n7390 ;
  assign n8156 = ( n8092 & ~n8151 ) | ( n8092 & n8155 ) | ( ~n8151 & n8155 ) ;
  assign n8157 = ( n8147 & ~n8150 ) | ( n8147 & n8156 ) | ( ~n8150 & n8156 ) ;
  assign n8167 = n333 ^ x17 ^ 1'b0 ;
  assign n8168 = n3499 & n8167 ;
  assign n8164 = ~n5004 & n7419 ;
  assign n8165 = ~n3920 & n8164 ;
  assign n8162 = n6065 ^ n589 ^ n132 ;
  assign n8163 = ( n3411 & n5718 ) | ( n3411 & n8162 ) | ( n5718 & n8162 ) ;
  assign n8166 = n8165 ^ n8163 ^ n967 ;
  assign n8158 = n1400 ^ n1358 ^ 1'b0 ;
  assign n8159 = n924 & ~n8158 ;
  assign n8160 = n8159 ^ n3558 ^ n1179 ;
  assign n8161 = ( n5761 & ~n5788 ) | ( n5761 & n8160 ) | ( ~n5788 & n8160 ) ;
  assign n8169 = n8168 ^ n8166 ^ n8161 ;
  assign n8170 = n2396 ^ n651 ^ 1'b0 ;
  assign n8171 = n6437 ^ n2041 ^ 1'b0 ;
  assign n8172 = ( ~n1158 & n1285 ) | ( ~n1158 & n1860 ) | ( n1285 & n1860 ) ;
  assign n8173 = n8172 ^ n7786 ^ 1'b0 ;
  assign n8174 = ~n6713 & n8173 ;
  assign n8175 = n6021 ^ n1522 ^ 1'b0 ;
  assign n8176 = ( n2657 & ~n8135 ) | ( n2657 & n8175 ) | ( ~n8135 & n8175 ) ;
  assign n8177 = ( n1217 & n3070 ) | ( n1217 & n4404 ) | ( n3070 & n4404 ) ;
  assign n8181 = n5599 ^ n5065 ^ 1'b0 ;
  assign n8182 = ~n1164 & n8181 ;
  assign n8178 = ( n239 & ~n3122 ) | ( n239 & n5803 ) | ( ~n3122 & n5803 ) ;
  assign n8179 = ~n994 & n8178 ;
  assign n8180 = n8179 ^ n4346 ^ 1'b0 ;
  assign n8183 = n8182 ^ n8180 ^ n5079 ;
  assign n8184 = ~n787 & n2551 ;
  assign n8185 = n6065 ^ n4224 ^ n2236 ;
  assign n8196 = ( n2000 & ~n2374 ) | ( n2000 & n2390 ) | ( ~n2374 & n2390 ) ;
  assign n8197 = n8196 ^ n1527 ^ n900 ;
  assign n8198 = ( ~n932 & n1446 ) | ( ~n932 & n8197 ) | ( n1446 & n8197 ) ;
  assign n8188 = n704 & ~n1638 ;
  assign n8189 = n8188 ^ n1093 ^ 1'b0 ;
  assign n8190 = n8189 ^ n4739 ^ n658 ;
  assign n8191 = ( ~x22 & n2079 ) | ( ~x22 & n3681 ) | ( n2079 & n3681 ) ;
  assign n8192 = x61 & n1093 ;
  assign n8193 = ( ~n2577 & n3256 ) | ( ~n2577 & n8192 ) | ( n3256 & n8192 ) ;
  assign n8194 = ( ~x126 & n8191 ) | ( ~x126 & n8193 ) | ( n8191 & n8193 ) ;
  assign n8195 = ( n1423 & n8190 ) | ( n1423 & n8194 ) | ( n8190 & n8194 ) ;
  assign n8186 = n1837 & n6986 ;
  assign n8187 = n8186 ^ n1593 ^ 1'b0 ;
  assign n8199 = n8198 ^ n8195 ^ n8187 ;
  assign n8200 = ( n8184 & n8185 ) | ( n8184 & n8199 ) | ( n8185 & n8199 ) ;
  assign n8201 = ( n1240 & ~n1362 ) | ( n1240 & n3650 ) | ( ~n1362 & n3650 ) ;
  assign n8202 = ( n2434 & ~n3855 ) | ( n2434 & n8201 ) | ( ~n3855 & n8201 ) ;
  assign n8203 = n8202 ^ n5379 ^ x31 ;
  assign n8204 = n8203 ^ n5617 ^ n5537 ;
  assign n8205 = n1442 ^ n952 ^ n283 ;
  assign n8206 = ( n2598 & n3264 ) | ( n2598 & n8205 ) | ( n3264 & n8205 ) ;
  assign n8207 = ( n4107 & ~n5719 ) | ( n4107 & n8206 ) | ( ~n5719 & n8206 ) ;
  assign n8208 = ( ~n5389 & n6701 ) | ( ~n5389 & n8207 ) | ( n6701 & n8207 ) ;
  assign n8209 = ( n1860 & n4142 ) | ( n1860 & ~n8208 ) | ( n4142 & ~n8208 ) ;
  assign n8210 = ( ~n905 & n2374 ) | ( ~n905 & n8209 ) | ( n2374 & n8209 ) ;
  assign n8212 = ( ~n314 & n1140 ) | ( ~n314 & n2890 ) | ( n1140 & n2890 ) ;
  assign n8211 = ( n2690 & n3514 ) | ( n2690 & ~n6713 ) | ( n3514 & ~n6713 ) ;
  assign n8213 = n8212 ^ n8211 ^ 1'b0 ;
  assign n8214 = n2513 ^ n1614 ^ 1'b0 ;
  assign n8215 = x8 & n8214 ;
  assign n8216 = n706 | n1884 ;
  assign n8217 = n8216 ^ n1409 ^ 1'b0 ;
  assign n8218 = ( ~n1184 & n2127 ) | ( ~n1184 & n8217 ) | ( n2127 & n8217 ) ;
  assign n8219 = n5629 ^ n5160 ^ 1'b0 ;
  assign n8224 = n2745 ^ n2708 ^ n926 ;
  assign n8225 = ( ~n4964 & n6120 ) | ( ~n4964 & n8224 ) | ( n6120 & n8224 ) ;
  assign n8220 = ~n521 & n2398 ;
  assign n8221 = ( ~n497 & n3662 ) | ( ~n497 & n5716 ) | ( n3662 & n5716 ) ;
  assign n8222 = ( ~x49 & n8220 ) | ( ~x49 & n8221 ) | ( n8220 & n8221 ) ;
  assign n8223 = ( ~n201 & n2728 ) | ( ~n201 & n8222 ) | ( n2728 & n8222 ) ;
  assign n8226 = n8225 ^ n8223 ^ n5113 ;
  assign n8227 = ( ~n1868 & n2439 ) | ( ~n1868 & n8226 ) | ( n2439 & n8226 ) ;
  assign n8228 = ( n2726 & n3479 ) | ( n2726 & ~n3791 ) | ( n3479 & ~n3791 ) ;
  assign n8229 = n5605 ^ n4144 ^ n3103 ;
  assign n8230 = ( n387 & ~n4673 ) | ( n387 & n8229 ) | ( ~n4673 & n8229 ) ;
  assign n8231 = ( ~n1979 & n8228 ) | ( ~n1979 & n8230 ) | ( n8228 & n8230 ) ;
  assign n8232 = n4830 ^ n2941 ^ n1006 ;
  assign n8233 = ( n1893 & n7573 ) | ( n1893 & n8232 ) | ( n7573 & n8232 ) ;
  assign n8234 = n8233 ^ n4713 ^ n1003 ;
  assign n8235 = n906 | n8234 ;
  assign n8236 = n8235 ^ n3325 ^ 1'b0 ;
  assign n8237 = n8236 ^ n7864 ^ n4814 ;
  assign n8241 = n3397 | n3710 ;
  assign n8238 = n3264 ^ n215 ^ 1'b0 ;
  assign n8239 = n740 & ~n8238 ;
  assign n8240 = n8239 ^ n5723 ^ 1'b0 ;
  assign n8242 = n8241 ^ n8240 ^ n498 ;
  assign n8249 = ( n266 & n2553 ) | ( n266 & ~n6757 ) | ( n2553 & ~n6757 ) ;
  assign n8243 = ( n3447 & ~n4385 ) | ( n3447 & n4400 ) | ( ~n4385 & n4400 ) ;
  assign n8244 = ~n640 & n8243 ;
  assign n8245 = ( ~n2160 & n3778 ) | ( ~n2160 & n4887 ) | ( n3778 & n4887 ) ;
  assign n8246 = ~n8244 & n8245 ;
  assign n8247 = ~n3683 & n8246 ;
  assign n8248 = n8247 ^ n5296 ^ n4818 ;
  assign n8250 = n8249 ^ n8248 ^ n2420 ;
  assign n8251 = n8250 ^ n3253 ^ 1'b0 ;
  assign n8252 = ( n2453 & ~n8190 ) | ( n2453 & n8251 ) | ( ~n8190 & n8251 ) ;
  assign n8253 = n3822 ^ n3442 ^ n2159 ;
  assign n8254 = n2132 | n3041 ;
  assign n8255 = ( n7786 & n8253 ) | ( n7786 & n8254 ) | ( n8253 & n8254 ) ;
  assign n8256 = ( n220 & n1558 ) | ( n220 & ~n7652 ) | ( n1558 & ~n7652 ) ;
  assign n8257 = n8256 ^ n1898 ^ 1'b0 ;
  assign n8258 = n8255 | n8257 ;
  assign n8259 = ( n382 & n1277 ) | ( n382 & ~n1644 ) | ( n1277 & ~n1644 ) ;
  assign n8260 = n7951 ^ n5339 ^ n3241 ;
  assign n8261 = n8260 ^ n1853 ^ n748 ;
  assign n8262 = n8259 & n8261 ;
  assign n8263 = n7681 ^ n2069 ^ 1'b0 ;
  assign n8264 = ~n3874 & n8263 ;
  assign n8265 = n527 | n1366 ;
  assign n8269 = n794 ^ n428 ^ n175 ;
  assign n8270 = ( x108 & n3528 ) | ( x108 & ~n8269 ) | ( n3528 & ~n8269 ) ;
  assign n8266 = ( ~n1060 & n2507 ) | ( ~n1060 & n4045 ) | ( n2507 & n4045 ) ;
  assign n8267 = ( ~n439 & n7287 ) | ( ~n439 & n8266 ) | ( n7287 & n8266 ) ;
  assign n8268 = n8267 ^ n3999 ^ n3068 ;
  assign n8271 = n8270 ^ n8268 ^ n7062 ;
  assign n8272 = n8253 ^ n3724 ^ n3064 ;
  assign n8273 = n8272 ^ n7688 ^ n1808 ;
  assign n8274 = ( n536 & ~n5007 ) | ( n536 & n8273 ) | ( ~n5007 & n8273 ) ;
  assign n8275 = ( n3704 & n5560 ) | ( n3704 & n8274 ) | ( n5560 & n8274 ) ;
  assign n8276 = ( n276 & n8271 ) | ( n276 & ~n8275 ) | ( n8271 & ~n8275 ) ;
  assign n8277 = ( ~n417 & n3171 ) | ( ~n417 & n5592 ) | ( n3171 & n5592 ) ;
  assign n8294 = n8035 ^ n4241 ^ n1577 ;
  assign n8295 = ( n6042 & ~n7679 ) | ( n6042 & n8294 ) | ( ~n7679 & n8294 ) ;
  assign n8292 = n3171 | n6482 ;
  assign n8293 = n8292 ^ n4064 ^ 1'b0 ;
  assign n8279 = n751 & ~n5405 ;
  assign n8278 = ( n1336 & n1932 ) | ( n1336 & n4027 ) | ( n1932 & n4027 ) ;
  assign n8280 = n8279 ^ n8278 ^ n4723 ;
  assign n8281 = ( n578 & n1273 ) | ( n578 & ~n4626 ) | ( n1273 & ~n4626 ) ;
  assign n8287 = n5530 ^ n836 ^ n461 ;
  assign n8284 = n7924 ^ n5654 ^ n966 ;
  assign n8285 = ( n4447 & n7196 ) | ( n4447 & ~n8284 ) | ( n7196 & ~n8284 ) ;
  assign n8286 = ( ~n368 & n6028 ) | ( ~n368 & n8285 ) | ( n6028 & n8285 ) ;
  assign n8282 = n4725 ^ n2793 ^ 1'b0 ;
  assign n8283 = ( n596 & ~n4349 ) | ( n596 & n8282 ) | ( ~n4349 & n8282 ) ;
  assign n8288 = n8287 ^ n8286 ^ n8283 ;
  assign n8289 = ~n8281 & n8288 ;
  assign n8290 = n8289 ^ n5931 ^ 1'b0 ;
  assign n8291 = ( n5661 & ~n8280 ) | ( n5661 & n8290 ) | ( ~n8280 & n8290 ) ;
  assign n8296 = n8295 ^ n8293 ^ n8291 ;
  assign n8302 = n5411 ^ n4374 ^ n4091 ;
  assign n8300 = ( ~n173 & n376 ) | ( ~n173 & n2436 ) | ( n376 & n2436 ) ;
  assign n8301 = ( n915 & n4550 ) | ( n915 & ~n8300 ) | ( n4550 & ~n8300 ) ;
  assign n8297 = n1265 ^ n277 ^ 1'b0 ;
  assign n8298 = n8297 ^ n2396 ^ n286 ;
  assign n8299 = ( n699 & n7858 ) | ( n699 & ~n8298 ) | ( n7858 & ~n8298 ) ;
  assign n8303 = n8302 ^ n8301 ^ n8299 ;
  assign n8304 = ( n4789 & ~n6475 ) | ( n4789 & n8303 ) | ( ~n6475 & n8303 ) ;
  assign n8305 = ( n2308 & n6051 ) | ( n2308 & n6467 ) | ( n6051 & n6467 ) ;
  assign n8306 = ( ~n6691 & n7483 ) | ( ~n6691 & n8305 ) | ( n7483 & n8305 ) ;
  assign n8307 = n6848 ^ n2318 ^ n839 ;
  assign n8308 = n2733 ^ n674 ^ 1'b0 ;
  assign n8309 = ( x56 & n8307 ) | ( x56 & ~n8308 ) | ( n8307 & ~n8308 ) ;
  assign n8311 = n5190 ^ n3513 ^ n1666 ;
  assign n8312 = n8311 ^ n2174 ^ 1'b0 ;
  assign n8313 = n4997 & ~n8312 ;
  assign n8314 = n8313 ^ n4954 ^ n1684 ;
  assign n8310 = ( n4901 & ~n5619 ) | ( n4901 & n6406 ) | ( ~n5619 & n6406 ) ;
  assign n8315 = n8314 ^ n8310 ^ n986 ;
  assign n8316 = n8315 ^ n4744 ^ n1583 ;
  assign n8317 = n5643 ^ n4871 ^ n714 ;
  assign n8318 = ~n962 & n8317 ;
  assign n8319 = n8318 ^ n2833 ^ 1'b0 ;
  assign n8320 = ( n414 & n3266 ) | ( n414 & n4052 ) | ( n3266 & n4052 ) ;
  assign n8321 = n5303 ^ n5026 ^ n742 ;
  assign n8322 = ~n8320 & n8321 ;
  assign n8323 = n8322 ^ n2629 ^ 1'b0 ;
  assign n8325 = n3063 ^ n2534 ^ n507 ;
  assign n8324 = ( n294 & n3286 ) | ( n294 & n7207 ) | ( n3286 & n7207 ) ;
  assign n8326 = n8325 ^ n8324 ^ 1'b0 ;
  assign n8327 = ( n2807 & ~n3124 ) | ( n2807 & n7866 ) | ( ~n3124 & n7866 ) ;
  assign n8328 = n8327 ^ n6838 ^ n4510 ;
  assign n8329 = n2455 & n7113 ;
  assign n8330 = ~n7793 & n8329 ;
  assign n8331 = n8328 | n8330 ;
  assign n8332 = n8331 ^ n6594 ^ n5066 ;
  assign n8333 = n6635 ^ n4977 ^ n3184 ;
  assign n8334 = n3736 & n8333 ;
  assign n8335 = n8334 ^ n2521 ^ 1'b0 ;
  assign n8336 = n1205 | n2962 ;
  assign n8337 = ( ~n1549 & n4173 ) | ( ~n1549 & n4587 ) | ( n4173 & n4587 ) ;
  assign n8338 = n8337 ^ n3720 ^ n1039 ;
  assign n8339 = ( n614 & n1352 ) | ( n614 & n2853 ) | ( n1352 & n2853 ) ;
  assign n8340 = n8339 ^ n6184 ^ n5583 ;
  assign n8341 = n8340 ^ n2232 ^ n711 ;
  assign n8342 = ( n989 & ~n8338 ) | ( n989 & n8341 ) | ( ~n8338 & n8341 ) ;
  assign n8344 = ( n1614 & n2664 ) | ( n1614 & ~n6669 ) | ( n2664 & ~n6669 ) ;
  assign n8343 = n7498 ^ n3722 ^ n940 ;
  assign n8345 = n8344 ^ n8343 ^ n6955 ;
  assign n8346 = n8345 ^ n248 ^ 1'b0 ;
  assign n8347 = n4574 | n8346 ;
  assign n8348 = ( n2342 & n4626 ) | ( n2342 & n4910 ) | ( n4626 & n4910 ) ;
  assign n8349 = ( ~n6477 & n8138 ) | ( ~n6477 & n8348 ) | ( n8138 & n8348 ) ;
  assign n8350 = ( ~n524 & n636 ) | ( ~n524 & n4484 ) | ( n636 & n4484 ) ;
  assign n8351 = n8350 ^ n6107 ^ n664 ;
  assign n8358 = n6890 ^ n4105 ^ n4048 ;
  assign n8352 = ( n3688 & n4519 ) | ( n3688 & n5269 ) | ( n4519 & n5269 ) ;
  assign n8353 = n4220 ^ n2438 ^ 1'b0 ;
  assign n8354 = n329 | n8353 ;
  assign n8355 = ( n2046 & n8352 ) | ( n2046 & n8354 ) | ( n8352 & n8354 ) ;
  assign n8356 = ( n3779 & n5828 ) | ( n3779 & n8355 ) | ( n5828 & n8355 ) ;
  assign n8357 = n8356 ^ n2340 ^ n1633 ;
  assign n8359 = n8358 ^ n8357 ^ n2227 ;
  assign n8360 = n8359 ^ n7989 ^ n4213 ;
  assign n8361 = ~n492 & n2174 ;
  assign n8362 = n8361 ^ n2377 ^ 1'b0 ;
  assign n8363 = x21 & n8362 ;
  assign n8365 = ~x23 & n5703 ;
  assign n8364 = n5539 ^ n5044 ^ n624 ;
  assign n8366 = n8365 ^ n8364 ^ n1110 ;
  assign n8367 = ( ~x81 & n8363 ) | ( ~x81 & n8366 ) | ( n8363 & n8366 ) ;
  assign n8368 = ( ~n5781 & n8360 ) | ( ~n5781 & n8367 ) | ( n8360 & n8367 ) ;
  assign n8369 = n4158 ^ n3159 ^ n2263 ;
  assign n8370 = ~n2594 & n8369 ;
  assign n8371 = n4722 ^ n4262 ^ n3776 ;
  assign n8372 = n8371 ^ n3677 ^ x28 ;
  assign n8373 = n8370 | n8372 ;
  assign n8387 = ( n1410 & ~n3012 ) | ( n1410 & n3517 ) | ( ~n3012 & n3517 ) ;
  assign n8382 = n1853 | n5936 ;
  assign n8383 = n3305 ^ n3272 ^ n906 ;
  assign n8384 = n8383 ^ n460 ^ n261 ;
  assign n8385 = ( n626 & n5088 ) | ( n626 & ~n8384 ) | ( n5088 & ~n8384 ) ;
  assign n8386 = ( ~n4003 & n8382 ) | ( ~n4003 & n8385 ) | ( n8382 & n8385 ) ;
  assign n8378 = n6442 ^ n4296 ^ n2125 ;
  assign n8377 = n7078 ^ n5520 ^ n1400 ;
  assign n8376 = n4779 | n6812 ;
  assign n8379 = n8378 ^ n8377 ^ n8376 ;
  assign n8380 = n8379 ^ n7914 ^ n2733 ;
  assign n8374 = n3820 ^ n3395 ^ 1'b0 ;
  assign n8375 = n8374 ^ n8286 ^ n3026 ;
  assign n8381 = n8380 ^ n8375 ^ n8044 ;
  assign n8388 = n8387 ^ n8386 ^ n8381 ;
  assign n8389 = ( n259 & n2253 ) | ( n259 & ~n3184 ) | ( n2253 & ~n3184 ) ;
  assign n8390 = n4583 ^ n730 ^ 1'b0 ;
  assign n8391 = n8389 | n8390 ;
  assign n8393 = ( x11 & n232 ) | ( x11 & n1489 ) | ( n232 & n1489 ) ;
  assign n8392 = ( x91 & ~n969 ) | ( x91 & n4288 ) | ( ~n969 & n4288 ) ;
  assign n8394 = n8393 ^ n8392 ^ n6743 ;
  assign n8395 = ( n1018 & n1030 ) | ( n1018 & ~n2434 ) | ( n1030 & ~n2434 ) ;
  assign n8396 = ( n2117 & n4250 ) | ( n2117 & n8395 ) | ( n4250 & n8395 ) ;
  assign n8397 = n8396 ^ n6028 ^ n3131 ;
  assign n8398 = ( n2255 & n8394 ) | ( n2255 & n8397 ) | ( n8394 & n8397 ) ;
  assign n8399 = n5351 ^ n4772 ^ n881 ;
  assign n8400 = ( n2443 & n2656 ) | ( n2443 & n2947 ) | ( n2656 & n2947 ) ;
  assign n8401 = n8400 ^ n1695 ^ n469 ;
  assign n8402 = n1155 & n8401 ;
  assign n8403 = n8402 ^ n2554 ^ 1'b0 ;
  assign n8404 = ( ~n5410 & n8399 ) | ( ~n5410 & n8403 ) | ( n8399 & n8403 ) ;
  assign n8412 = ( n738 & n1386 ) | ( n738 & n2727 ) | ( n1386 & n2727 ) ;
  assign n8409 = n7810 ^ n5933 ^ 1'b0 ;
  assign n8410 = n136 & ~n8409 ;
  assign n8405 = ( ~n992 & n2063 ) | ( ~n992 & n4044 ) | ( n2063 & n4044 ) ;
  assign n8406 = n8405 ^ n4939 ^ n1748 ;
  assign n8407 = n8406 ^ n2277 ^ n1009 ;
  assign n8408 = n7545 & ~n8407 ;
  assign n8411 = n8410 ^ n8408 ^ n1413 ;
  assign n8413 = n8412 ^ n8411 ^ n1593 ;
  assign n8414 = ( n138 & n2378 ) | ( n138 & ~n4059 ) | ( n2378 & ~n4059 ) ;
  assign n8418 = ( n1894 & ~n3704 ) | ( n1894 & n5700 ) | ( ~n3704 & n5700 ) ;
  assign n8419 = n4135 & n8418 ;
  assign n8420 = ~n5338 & n8419 ;
  assign n8415 = n2449 & n5081 ;
  assign n8416 = ( n5293 & n5792 ) | ( n5293 & n6583 ) | ( n5792 & n6583 ) ;
  assign n8417 = n8415 | n8416 ;
  assign n8421 = n8420 ^ n8417 ^ 1'b0 ;
  assign n8422 = ( n1157 & n1686 ) | ( n1157 & n2534 ) | ( n1686 & n2534 ) ;
  assign n8423 = ~n4097 & n8422 ;
  assign n8424 = n8423 ^ n4530 ^ 1'b0 ;
  assign n8425 = n6112 ^ n3330 ^ x28 ;
  assign n8426 = n8425 ^ n8285 ^ n4907 ;
  assign n8427 = n8424 | n8426 ;
  assign n8428 = n7873 | n8427 ;
  assign n8429 = n2879 & n7173 ;
  assign n8430 = n8429 ^ n4250 ^ 1'b0 ;
  assign n8431 = n8430 ^ n5246 ^ 1'b0 ;
  assign n8432 = ~n3095 & n8431 ;
  assign n8434 = n2314 ^ n2213 ^ 1'b0 ;
  assign n8435 = n6665 & ~n8434 ;
  assign n8440 = n1964 | n7195 ;
  assign n8441 = n1606 | n8440 ;
  assign n8436 = n2098 ^ n388 ^ 1'b0 ;
  assign n8437 = n1861 & ~n8436 ;
  assign n8438 = ( n2294 & n3356 ) | ( n2294 & n8437 ) | ( n3356 & n8437 ) ;
  assign n8439 = ( n3290 & n3969 ) | ( n3290 & n8438 ) | ( n3969 & n8438 ) ;
  assign n8442 = n8441 ^ n8439 ^ n1270 ;
  assign n8443 = ( n6882 & ~n8435 ) | ( n6882 & n8442 ) | ( ~n8435 & n8442 ) ;
  assign n8433 = n1992 & n6148 ;
  assign n8444 = n8443 ^ n8433 ^ 1'b0 ;
  assign n8445 = ( n950 & n1327 ) | ( n950 & ~n3449 ) | ( n1327 & ~n3449 ) ;
  assign n8447 = ( n678 & n1076 ) | ( n678 & n1211 ) | ( n1076 & n1211 ) ;
  assign n8446 = n7841 ^ n4608 ^ x16 ;
  assign n8448 = n8447 ^ n8446 ^ n1503 ;
  assign n8449 = n3483 ^ n974 ^ 1'b0 ;
  assign n8450 = ~n7786 & n8449 ;
  assign n8451 = ( n8445 & n8448 ) | ( n8445 & n8450 ) | ( n8448 & n8450 ) ;
  assign n8452 = n1716 & ~n8451 ;
  assign n8453 = n3143 ^ n2296 ^ n1138 ;
  assign n8454 = n5151 ^ n2433 ^ n1431 ;
  assign n8455 = ( n165 & n888 ) | ( n165 & ~n8454 ) | ( n888 & ~n8454 ) ;
  assign n8456 = n8455 ^ n6883 ^ n2550 ;
  assign n8457 = n7692 ^ x93 ^ x43 ;
  assign n8458 = n8457 ^ n6956 ^ n3516 ;
  assign n8459 = ~n983 & n5643 ;
  assign n8460 = n8458 & n8459 ;
  assign n8461 = n206 & ~n8460 ;
  assign n8462 = n2617 ^ n487 ^ n392 ;
  assign n8463 = ( n642 & n2063 ) | ( n642 & ~n8462 ) | ( n2063 & ~n8462 ) ;
  assign n8464 = n5360 | n8463 ;
  assign n8465 = n1462 & ~n8464 ;
  assign n8466 = ( n3781 & n8461 ) | ( n3781 & n8465 ) | ( n8461 & n8465 ) ;
  assign n8467 = ( ~n8453 & n8456 ) | ( ~n8453 & n8466 ) | ( n8456 & n8466 ) ;
  assign n8492 = ( n910 & n1226 ) | ( n910 & n5389 ) | ( n1226 & n5389 ) ;
  assign n8493 = ( n1799 & n3504 ) | ( n1799 & n8492 ) | ( n3504 & n8492 ) ;
  assign n8488 = n2069 | n2831 ;
  assign n8489 = n145 & ~n8488 ;
  assign n8490 = n6743 ^ n2322 ^ n795 ;
  assign n8491 = ( n2752 & ~n8489 ) | ( n2752 & n8490 ) | ( ~n8489 & n8490 ) ;
  assign n8481 = n6957 ^ n4651 ^ n1998 ;
  assign n8482 = ( n2060 & n2996 ) | ( n2060 & ~n4016 ) | ( n2996 & ~n4016 ) ;
  assign n8483 = n8482 ^ n7307 ^ 1'b0 ;
  assign n8484 = n8481 | n8483 ;
  assign n8475 = ( ~n3465 & n7879 ) | ( ~n3465 & n8100 ) | ( n7879 & n8100 ) ;
  assign n8476 = ( n2976 & n6787 ) | ( n2976 & n8475 ) | ( n6787 & n8475 ) ;
  assign n8477 = n3114 | n8383 ;
  assign n8478 = n8476 & ~n8477 ;
  assign n8479 = n8478 ^ n4762 ^ n3089 ;
  assign n8472 = n5376 ^ n4183 ^ n3702 ;
  assign n8473 = ( n2402 & n8211 ) | ( n2402 & n8472 ) | ( n8211 & n8472 ) ;
  assign n8474 = ( n2270 & ~n4023 ) | ( n2270 & n8473 ) | ( ~n4023 & n8473 ) ;
  assign n8469 = n6627 ^ n3176 ^ n683 ;
  assign n8468 = n2766 & n3137 ;
  assign n8470 = n8469 ^ n8468 ^ 1'b0 ;
  assign n8471 = ( n2662 & n7288 ) | ( n2662 & n8470 ) | ( n7288 & n8470 ) ;
  assign n8480 = n8479 ^ n8474 ^ n8471 ;
  assign n8485 = n8484 ^ n8480 ^ n6287 ;
  assign n8486 = n8485 ^ n7143 ^ n5636 ;
  assign n8487 = n8486 ^ n641 ^ 1'b0 ;
  assign n8494 = n8493 ^ n8491 ^ n8487 ;
  assign n8496 = n3749 & ~n7200 ;
  assign n8495 = n5316 ^ n251 ^ 1'b0 ;
  assign n8497 = n8496 ^ n8495 ^ 1'b0 ;
  assign n8498 = n8497 ^ n7321 ^ n7176 ;
  assign n8499 = n4434 ^ n1975 ^ n1826 ;
  assign n8500 = ( n314 & n7869 ) | ( n314 & n8499 ) | ( n7869 & n8499 ) ;
  assign n8503 = n1121 ^ x68 ^ 1'b0 ;
  assign n8504 = n8503 ^ n7211 ^ 1'b0 ;
  assign n8505 = ~n2127 & n8504 ;
  assign n8506 = n8505 ^ n3840 ^ n3235 ;
  assign n8501 = ( n2370 & ~n3342 ) | ( n2370 & n7216 ) | ( ~n3342 & n7216 ) ;
  assign n8502 = ( n4100 & n6691 ) | ( n4100 & n8501 ) | ( n6691 & n8501 ) ;
  assign n8507 = n8506 ^ n8502 ^ 1'b0 ;
  assign n8508 = n7888 ^ n4391 ^ n1897 ;
  assign n8510 = n4342 ^ n1522 ^ n1138 ;
  assign n8509 = n4906 ^ n3131 ^ n294 ;
  assign n8511 = n8510 ^ n8509 ^ n961 ;
  assign n8512 = n3671 ^ n1130 ^ 1'b0 ;
  assign n8513 = n7730 & n8512 ;
  assign n8514 = n7505 ^ n3466 ^ n2694 ;
  assign n8515 = ( ~n608 & n4196 ) | ( ~n608 & n5070 ) | ( n4196 & n5070 ) ;
  assign n8518 = ( n211 & n437 ) | ( n211 & ~n6896 ) | ( n437 & ~n6896 ) ;
  assign n8519 = ( n994 & ~n1198 ) | ( n994 & n8518 ) | ( ~n1198 & n8518 ) ;
  assign n8517 = n2170 | n2942 ;
  assign n8520 = n8519 ^ n8517 ^ 1'b0 ;
  assign n8516 = n7592 ^ n6618 ^ n1286 ;
  assign n8521 = n8520 ^ n8516 ^ n1218 ;
  assign n8522 = ( n8514 & n8515 ) | ( n8514 & ~n8521 ) | ( n8515 & ~n8521 ) ;
  assign n8524 = ( n3964 & ~n4493 ) | ( n3964 & n6525 ) | ( ~n4493 & n6525 ) ;
  assign n8525 = ( n930 & ~n3075 ) | ( n930 & n8524 ) | ( ~n3075 & n8524 ) ;
  assign n8523 = n6868 | n7608 ;
  assign n8526 = n8525 ^ n8523 ^ 1'b0 ;
  assign n8527 = ( ~n2823 & n6336 ) | ( ~n2823 & n8526 ) | ( n6336 & n8526 ) ;
  assign n8528 = n7134 ^ n1579 ^ n806 ;
  assign n8529 = n8528 ^ n4354 ^ n1533 ;
  assign n8530 = n8529 ^ n4393 ^ n1663 ;
  assign n8531 = ( n1146 & n6636 ) | ( n1146 & ~n8530 ) | ( n6636 & ~n8530 ) ;
  assign n8532 = ( ~n164 & n4074 ) | ( ~n164 & n6449 ) | ( n4074 & n6449 ) ;
  assign n8533 = n8165 ^ n474 ^ 1'b0 ;
  assign n8534 = ( n1172 & n5224 ) | ( n1172 & ~n5516 ) | ( n5224 & ~n5516 ) ;
  assign n8535 = ( ~n617 & n791 ) | ( ~n617 & n8534 ) | ( n791 & n8534 ) ;
  assign n8536 = ( x120 & n5496 ) | ( x120 & n8225 ) | ( n5496 & n8225 ) ;
  assign n8537 = n8492 ^ n7243 ^ n2862 ;
  assign n8538 = n8537 ^ n7695 ^ n3168 ;
  assign n8539 = ( n1068 & n7506 ) | ( n1068 & n8211 ) | ( n7506 & n8211 ) ;
  assign n8540 = ( n2659 & n2927 ) | ( n2659 & n8510 ) | ( n2927 & n8510 ) ;
  assign n8541 = ( n756 & ~n3098 ) | ( n756 & n8528 ) | ( ~n3098 & n8528 ) ;
  assign n8542 = n8541 ^ n2728 ^ n1122 ;
  assign n8543 = n8542 ^ n6555 ^ 1'b0 ;
  assign n8544 = n2532 & n8543 ;
  assign n8545 = ( n5643 & ~n8540 ) | ( n5643 & n8544 ) | ( ~n8540 & n8544 ) ;
  assign n8546 = ( n8538 & n8539 ) | ( n8538 & n8545 ) | ( n8539 & n8545 ) ;
  assign n8547 = ( n8535 & ~n8536 ) | ( n8535 & n8546 ) | ( ~n8536 & n8546 ) ;
  assign n8548 = ( n1311 & n1859 ) | ( n1311 & ~n7590 ) | ( n1859 & ~n7590 ) ;
  assign n8549 = ( n166 & n662 ) | ( n166 & n1059 ) | ( n662 & n1059 ) ;
  assign n8550 = n8437 ^ n2534 ^ n1086 ;
  assign n8551 = n8550 ^ n5551 ^ n4533 ;
  assign n8552 = n4614 & ~n8551 ;
  assign n8553 = n7985 ^ n2463 ^ n1801 ;
  assign n8554 = n8553 ^ n7151 ^ n2658 ;
  assign n8559 = ~n6449 & n8288 ;
  assign n8556 = n1678 ^ n1363 ^ n1154 ;
  assign n8555 = n5895 ^ n2354 ^ n1813 ;
  assign n8557 = n8556 ^ n8555 ^ n5743 ;
  assign n8558 = n2089 & n8557 ;
  assign n8560 = n8559 ^ n8558 ^ 1'b0 ;
  assign n8561 = n4127 ^ n3738 ^ 1'b0 ;
  assign n8562 = n1888 | n8561 ;
  assign n8563 = ( x63 & n1044 ) | ( x63 & n1748 ) | ( n1044 & n1748 ) ;
  assign n8564 = ( n1167 & n3127 ) | ( n1167 & n4605 ) | ( n3127 & n4605 ) ;
  assign n8565 = ( n8562 & n8563 ) | ( n8562 & ~n8564 ) | ( n8563 & ~n8564 ) ;
  assign n8566 = n2455 ^ n1447 ^ n921 ;
  assign n8567 = ( n1690 & ~n2862 ) | ( n1690 & n8566 ) | ( ~n2862 & n8566 ) ;
  assign n8568 = n4473 ^ n1847 ^ n1579 ;
  assign n8569 = ( n5182 & n7553 ) | ( n5182 & ~n8568 ) | ( n7553 & ~n8568 ) ;
  assign n8570 = ( ~n3964 & n6774 ) | ( ~n3964 & n8569 ) | ( n6774 & n8569 ) ;
  assign n8571 = ( ~n8565 & n8567 ) | ( ~n8565 & n8570 ) | ( n8567 & n8570 ) ;
  assign n8572 = n8571 ^ n4234 ^ n1730 ;
  assign n8573 = ( n713 & ~n1148 ) | ( n713 & n5602 ) | ( ~n1148 & n5602 ) ;
  assign n8574 = ( n1128 & n2135 ) | ( n1128 & n3489 ) | ( n2135 & n3489 ) ;
  assign n8575 = n1806 & n8574 ;
  assign n8576 = ( n1165 & n3371 ) | ( n1165 & n5249 ) | ( n3371 & n5249 ) ;
  assign n8577 = n8576 ^ n3114 ^ 1'b0 ;
  assign n8578 = ( n4850 & n8575 ) | ( n4850 & n8577 ) | ( n8575 & n8577 ) ;
  assign n8579 = ( ~n325 & n8573 ) | ( ~n325 & n8578 ) | ( n8573 & n8578 ) ;
  assign n8580 = n8579 ^ n7419 ^ n3861 ;
  assign n8581 = ( n3391 & n4436 ) | ( n3391 & ~n8580 ) | ( n4436 & ~n8580 ) ;
  assign n8582 = ( n753 & n2874 ) | ( n753 & n8581 ) | ( n2874 & n8581 ) ;
  assign n8583 = n8582 ^ n7104 ^ n4199 ;
  assign n8584 = ( n1610 & n1902 ) | ( n1610 & n2779 ) | ( n1902 & n2779 ) ;
  assign n8585 = ( n1064 & n7186 ) | ( n1064 & n8584 ) | ( n7186 & n8584 ) ;
  assign n8586 = ( n1789 & n3417 ) | ( n1789 & n8585 ) | ( n3417 & n8585 ) ;
  assign n8587 = n1623 ^ n1574 ^ 1'b0 ;
  assign n8588 = n8587 ^ n5821 ^ n3098 ;
  assign n8589 = ~n5077 & n8588 ;
  assign n8590 = n8589 ^ n4102 ^ 1'b0 ;
  assign n8594 = ( n1461 & ~n1559 ) | ( n1461 & n3274 ) | ( ~n1559 & n3274 ) ;
  assign n8593 = x26 & ~n5357 ;
  assign n8595 = n8594 ^ n8593 ^ 1'b0 ;
  assign n8591 = n5723 ^ n5517 ^ n1895 ;
  assign n8592 = n4068 & n8591 ;
  assign n8596 = n8595 ^ n8592 ^ 1'b0 ;
  assign n8598 = n7116 ^ n3138 ^ n704 ;
  assign n8597 = ( n1958 & n2641 ) | ( n1958 & n6205 ) | ( n2641 & n6205 ) ;
  assign n8599 = n8598 ^ n8597 ^ n6511 ;
  assign n8601 = n7799 ^ n2750 ^ n2678 ;
  assign n8600 = n4057 & ~n7308 ;
  assign n8602 = n8601 ^ n8600 ^ 1'b0 ;
  assign n8604 = ( ~n410 & n7302 ) | ( ~n410 & n7825 ) | ( n7302 & n7825 ) ;
  assign n8603 = n6871 ^ n6542 ^ n452 ;
  assign n8605 = n8604 ^ n8603 ^ n7681 ;
  assign n8606 = n6530 ^ n4132 ^ n1526 ;
  assign n8615 = n7729 ^ n4032 ^ n984 ;
  assign n8613 = ( n983 & ~n1004 ) | ( n983 & n1034 ) | ( ~n1004 & n1034 ) ;
  assign n8611 = ( ~n2322 & n4198 ) | ( ~n2322 & n4359 ) | ( n4198 & n4359 ) ;
  assign n8612 = ( n3524 & n6149 ) | ( n3524 & ~n8611 ) | ( n6149 & ~n8611 ) ;
  assign n8607 = ( x62 & n1521 ) | ( x62 & ~n7777 ) | ( n1521 & ~n7777 ) ;
  assign n8608 = ( n555 & n3335 ) | ( n555 & n3865 ) | ( n3335 & n3865 ) ;
  assign n8609 = n6627 ^ n4387 ^ n2214 ;
  assign n8610 = ( n8607 & n8608 ) | ( n8607 & n8609 ) | ( n8608 & n8609 ) ;
  assign n8614 = n8613 ^ n8612 ^ n8610 ;
  assign n8616 = n8615 ^ n8614 ^ n4883 ;
  assign n8617 = ( n4110 & n8606 ) | ( n4110 & n8616 ) | ( n8606 & n8616 ) ;
  assign n8618 = ( n8602 & n8605 ) | ( n8602 & n8617 ) | ( n8605 & n8617 ) ;
  assign n8623 = n3663 ^ n1986 ^ n1161 ;
  assign n8624 = n8623 ^ n7442 ^ n153 ;
  assign n8619 = n8074 ^ n3103 ^ n1060 ;
  assign n8620 = n1899 ^ n193 ^ x83 ;
  assign n8621 = n8620 ^ n2538 ^ n1322 ;
  assign n8622 = ( n4801 & n8619 ) | ( n4801 & n8621 ) | ( n8619 & n8621 ) ;
  assign n8625 = n8624 ^ n8622 ^ n2703 ;
  assign n8629 = ( n331 & n2759 ) | ( n331 & ~n4722 ) | ( n2759 & ~n4722 ) ;
  assign n8627 = n4188 ^ n4054 ^ n2754 ;
  assign n8628 = ( n827 & n1411 ) | ( n827 & ~n8627 ) | ( n1411 & ~n8627 ) ;
  assign n8626 = ( n1886 & n4241 ) | ( n1886 & ~n4944 ) | ( n4241 & ~n4944 ) ;
  assign n8630 = n8629 ^ n8628 ^ n8626 ;
  assign n8631 = n8630 ^ n7077 ^ n3092 ;
  assign n8635 = n2390 ^ n1617 ^ n710 ;
  assign n8634 = n7107 ^ n4501 ^ 1'b0 ;
  assign n8632 = ( ~n2549 & n2935 ) | ( ~n2549 & n7836 ) | ( n2935 & n7836 ) ;
  assign n8633 = n8632 ^ n3867 ^ 1'b0 ;
  assign n8636 = n8635 ^ n8634 ^ n8633 ;
  assign n8637 = n7776 ^ n3128 ^ n895 ;
  assign n8638 = n5014 ^ n2153 ^ n178 ;
  assign n8639 = n5206 ^ n4520 ^ n1215 ;
  assign n8640 = ( n196 & n8462 ) | ( n196 & n8639 ) | ( n8462 & n8639 ) ;
  assign n8641 = n3728 & ~n8640 ;
  assign n8642 = ( n4838 & ~n7431 ) | ( n4838 & n7966 ) | ( ~n7431 & n7966 ) ;
  assign n8643 = n8642 ^ n2045 ^ x97 ;
  assign n8644 = n2414 ^ n1207 ^ n785 ;
  assign n8645 = n6616 ^ n2760 ^ n1918 ;
  assign n8646 = ( n4551 & n8644 ) | ( n4551 & n8645 ) | ( n8644 & n8645 ) ;
  assign n8647 = ( ~n6412 & n8643 ) | ( ~n6412 & n8646 ) | ( n8643 & n8646 ) ;
  assign n8648 = ( ~x96 & n8641 ) | ( ~x96 & n8647 ) | ( n8641 & n8647 ) ;
  assign n8649 = ( n1022 & n8638 ) | ( n1022 & ~n8648 ) | ( n8638 & ~n8648 ) ;
  assign n8656 = ( n4780 & ~n5242 ) | ( n4780 & n6921 ) | ( ~n5242 & n6921 ) ;
  assign n8650 = ( ~n2422 & n3531 ) | ( ~n2422 & n6566 ) | ( n3531 & n6566 ) ;
  assign n8651 = ( n990 & ~n4945 ) | ( n990 & n8650 ) | ( ~n4945 & n8650 ) ;
  assign n8652 = ( ~x115 & n1826 ) | ( ~x115 & n7037 ) | ( n1826 & n7037 ) ;
  assign n8653 = n8652 ^ n8642 ^ n7324 ;
  assign n8654 = ( n192 & n8651 ) | ( n192 & ~n8653 ) | ( n8651 & ~n8653 ) ;
  assign n8655 = ( ~n3224 & n8096 ) | ( ~n3224 & n8654 ) | ( n8096 & n8654 ) ;
  assign n8657 = n8656 ^ n8655 ^ n3312 ;
  assign n8658 = n6070 ^ n5930 ^ n2974 ;
  assign n8659 = n4434 ^ n4309 ^ n3131 ;
  assign n8660 = ( n2268 & n3143 ) | ( n2268 & ~n8659 ) | ( n3143 & ~n8659 ) ;
  assign n8664 = n6457 ^ n980 ^ n530 ;
  assign n8661 = ( n372 & n971 ) | ( n372 & n3580 ) | ( n971 & n3580 ) ;
  assign n8662 = ( ~x30 & n305 ) | ( ~x30 & n8661 ) | ( n305 & n8661 ) ;
  assign n8663 = n8662 ^ n760 ^ n735 ;
  assign n8665 = n8664 ^ n8663 ^ n3669 ;
  assign n8666 = ( ~n400 & n1255 ) | ( ~n400 & n2706 ) | ( n1255 & n2706 ) ;
  assign n8667 = ( n5281 & n7342 ) | ( n5281 & ~n7995 ) | ( n7342 & ~n7995 ) ;
  assign n8668 = ( n3127 & ~n8666 ) | ( n3127 & n8667 ) | ( ~n8666 & n8667 ) ;
  assign n8669 = n6630 ^ n4352 ^ n3117 ;
  assign n8670 = ( n1232 & n2901 ) | ( n1232 & ~n8669 ) | ( n2901 & ~n8669 ) ;
  assign n8672 = n6751 ^ n3122 ^ n1845 ;
  assign n8671 = ( ~n780 & n891 ) | ( ~n780 & n1898 ) | ( n891 & n1898 ) ;
  assign n8673 = n8672 ^ n8671 ^ n4943 ;
  assign n8674 = n8673 ^ n4197 ^ x92 ;
  assign n8675 = ~n4790 & n8674 ;
  assign n8676 = n8675 ^ n7694 ^ 1'b0 ;
  assign n8677 = n2121 ^ n1972 ^ n203 ;
  assign n8694 = ( n912 & ~n1309 ) | ( n912 & n2175 ) | ( ~n1309 & n2175 ) ;
  assign n8695 = n2100 ^ n1913 ^ 1'b0 ;
  assign n8696 = n8694 | n8695 ;
  assign n8697 = n8696 ^ n7138 ^ n1753 ;
  assign n8686 = n475 & ~n885 ;
  assign n8687 = ( n3430 & n7725 ) | ( n3430 & ~n8686 ) | ( n7725 & ~n8686 ) ;
  assign n8688 = n8475 ^ n3227 ^ n2372 ;
  assign n8689 = ( n1390 & n2151 ) | ( n1390 & n2843 ) | ( n2151 & n2843 ) ;
  assign n8690 = n8689 ^ n6903 ^ n1589 ;
  assign n8691 = ( n3985 & n8688 ) | ( n3985 & n8690 ) | ( n8688 & n8690 ) ;
  assign n8692 = n8687 & n8691 ;
  assign n8693 = ~n1395 & n8692 ;
  assign n8680 = n2088 & ~n2882 ;
  assign n8681 = n7851 & n8680 ;
  assign n8682 = n8681 ^ n4665 ^ n2392 ;
  assign n8683 = n8682 ^ n8356 ^ 1'b0 ;
  assign n8684 = n4634 | n8683 ;
  assign n8678 = n469 & ~n4045 ;
  assign n8679 = ~n4655 & n8678 ;
  assign n8685 = n8684 ^ n8679 ^ n4890 ;
  assign n8698 = n8697 ^ n8693 ^ n8685 ;
  assign n8699 = ( n6129 & n8677 ) | ( n6129 & ~n8698 ) | ( n8677 & ~n8698 ) ;
  assign n8707 = n8301 ^ n8100 ^ n2878 ;
  assign n8705 = ~n3172 & n4655 ;
  assign n8706 = n6809 & n8705 ;
  assign n8701 = x7 & x89 ;
  assign n8702 = ~n1692 & n8701 ;
  assign n8703 = n8702 ^ n4045 ^ 1'b0 ;
  assign n8700 = n671 | n7698 ;
  assign n8704 = n8703 ^ n8700 ^ n5528 ;
  assign n8708 = n8707 ^ n8706 ^ n8704 ;
  assign n8713 = ( x43 & n1191 ) | ( x43 & n1766 ) | ( n1191 & n1766 ) ;
  assign n8709 = n6961 ^ n627 ^ 1'b0 ;
  assign n8710 = n1000 & n8709 ;
  assign n8711 = n5098 ^ n5009 ^ n1392 ;
  assign n8712 = ( ~n142 & n8710 ) | ( ~n142 & n8711 ) | ( n8710 & n8711 ) ;
  assign n8714 = n8713 ^ n8712 ^ n4266 ;
  assign n8715 = ( n3231 & n3440 ) | ( n3231 & n6121 ) | ( n3440 & n6121 ) ;
  assign n8716 = ~n3372 & n8715 ;
  assign n8717 = n3669 ^ n2095 ^ n411 ;
  assign n8718 = n5802 ^ n223 ^ 1'b0 ;
  assign n8719 = ( n2349 & n4643 ) | ( n2349 & ~n7573 ) | ( n4643 & ~n7573 ) ;
  assign n8720 = ( n5325 & ~n8718 ) | ( n5325 & n8719 ) | ( ~n8718 & n8719 ) ;
  assign n8721 = ( n6725 & ~n8717 ) | ( n6725 & n8720 ) | ( ~n8717 & n8720 ) ;
  assign n8722 = n4285 & ~n8721 ;
  assign n8723 = n4895 & n8722 ;
  assign n8724 = n7987 & ~n8723 ;
  assign n8725 = n8724 ^ n4530 ^ 1'b0 ;
  assign n8726 = ( n6051 & n8716 ) | ( n6051 & ~n8725 ) | ( n8716 & ~n8725 ) ;
  assign n8727 = ( x79 & ~n713 ) | ( x79 & n2461 ) | ( ~n713 & n2461 ) ;
  assign n8728 = ~n1692 & n8727 ;
  assign n8729 = n8343 ^ n3676 ^ n2245 ;
  assign n8730 = ( n1173 & n8728 ) | ( n1173 & n8729 ) | ( n8728 & n8729 ) ;
  assign n8731 = ( n1258 & n3105 ) | ( n1258 & ~n8730 ) | ( n3105 & ~n8730 ) ;
  assign n8732 = n238 | n8731 ;
  assign n8733 = ( ~n784 & n2204 ) | ( ~n784 & n4610 ) | ( n2204 & n4610 ) ;
  assign n8734 = n8093 & ~n8733 ;
  assign n8739 = ( n794 & n2309 ) | ( n794 & n2622 ) | ( n2309 & n2622 ) ;
  assign n8740 = n8739 ^ n7287 ^ n3662 ;
  assign n8736 = n6818 ^ n6514 ^ n4898 ;
  assign n8737 = n4688 | n8736 ;
  assign n8738 = n8737 ^ n4914 ^ 1'b0 ;
  assign n8735 = n5197 ^ n3803 ^ n303 ;
  assign n8741 = n8740 ^ n8738 ^ n8735 ;
  assign n8742 = n3247 ^ n1645 ^ n479 ;
  assign n8743 = n6206 ^ n4129 ^ n3095 ;
  assign n8744 = ( ~n7476 & n8742 ) | ( ~n7476 & n8743 ) | ( n8742 & n8743 ) ;
  assign n8745 = n8744 ^ n4400 ^ n1128 ;
  assign n8746 = n8745 ^ n6031 ^ n5275 ;
  assign n8747 = n2348 ^ n1068 ^ 1'b0 ;
  assign n8748 = ( n252 & n2924 ) | ( n252 & n8747 ) | ( n2924 & n8747 ) ;
  assign n8749 = n757 | n8748 ;
  assign n8750 = ( ~n870 & n3635 ) | ( ~n870 & n8749 ) | ( n3635 & n8749 ) ;
  assign n8751 = n8750 ^ n3933 ^ 1'b0 ;
  assign n8752 = n4785 ^ n4122 ^ n317 ;
  assign n8758 = n7134 ^ n2082 ^ 1'b0 ;
  assign n8753 = ( x58 & n2406 ) | ( x58 & n2521 ) | ( n2406 & n2521 ) ;
  assign n8754 = n8753 ^ n8623 ^ n4054 ;
  assign n8755 = n2135 ^ n545 ^ n363 ;
  assign n8756 = n8755 ^ n3599 ^ 1'b0 ;
  assign n8757 = n8754 & ~n8756 ;
  assign n8759 = n8758 ^ n8757 ^ n3568 ;
  assign n8760 = ( n610 & n5143 ) | ( n610 & n8759 ) | ( n5143 & n8759 ) ;
  assign n8761 = n8760 ^ n5379 ^ n383 ;
  assign n8762 = ~n3845 & n5776 ;
  assign n8763 = ( n401 & ~n7608 ) | ( n401 & n8535 ) | ( ~n7608 & n8535 ) ;
  assign n8764 = n2941 ^ n1817 ^ n855 ;
  assign n8765 = n5134 & ~n8764 ;
  assign n8766 = n8765 ^ n7679 ^ n539 ;
  assign n8767 = ~n6163 & n8017 ;
  assign n8768 = ( n771 & n1878 ) | ( n771 & ~n6449 ) | ( n1878 & ~n6449 ) ;
  assign n8769 = n8768 ^ n6964 ^ 1'b0 ;
  assign n8778 = ( x64 & n2135 ) | ( x64 & n2813 ) | ( n2135 & n2813 ) ;
  assign n8777 = n4830 ^ n926 ^ 1'b0 ;
  assign n8779 = n8778 ^ n8777 ^ n5052 ;
  assign n8770 = ( ~n329 & n612 ) | ( ~n329 & n2172 ) | ( n612 & n2172 ) ;
  assign n8771 = n8770 ^ n2667 ^ x73 ;
  assign n8772 = ( n2178 & n6210 ) | ( n2178 & ~n8771 ) | ( n6210 & ~n8771 ) ;
  assign n8773 = n5984 ^ n2638 ^ n354 ;
  assign n8774 = n1508 & ~n4944 ;
  assign n8775 = ( n1735 & n3352 ) | ( n1735 & n8774 ) | ( n3352 & n8774 ) ;
  assign n8776 = ( n8772 & n8773 ) | ( n8772 & ~n8775 ) | ( n8773 & ~n8775 ) ;
  assign n8780 = n8779 ^ n8776 ^ n1110 ;
  assign n8781 = n7681 ^ n1752 ^ n256 ;
  assign n8782 = n3182 ^ n2329 ^ n1973 ;
  assign n8783 = n4209 ^ n2906 ^ n1570 ;
  assign n8784 = ( n5204 & n6310 ) | ( n5204 & n8783 ) | ( n6310 & n8783 ) ;
  assign n8785 = ( n343 & ~n8782 ) | ( n343 & n8784 ) | ( ~n8782 & n8784 ) ;
  assign n8786 = n5362 ^ n3901 ^ 1'b0 ;
  assign n8787 = n2132 & ~n8786 ;
  assign n8788 = ( ~n5826 & n6462 ) | ( ~n5826 & n8787 ) | ( n6462 & n8787 ) ;
  assign n8789 = ( n8781 & n8785 ) | ( n8781 & ~n8788 ) | ( n8785 & ~n8788 ) ;
  assign n8790 = n5225 ^ n337 ^ 1'b0 ;
  assign n8792 = ( n1069 & n1446 ) | ( n1069 & n7706 ) | ( n1446 & n7706 ) ;
  assign n8791 = n6832 ^ n5829 ^ n2837 ;
  assign n8793 = n8792 ^ n8791 ^ n2558 ;
  assign n8794 = n1823 ^ n1808 ^ n771 ;
  assign n8795 = ( n760 & ~n4920 ) | ( n760 & n8739 ) | ( ~n4920 & n8739 ) ;
  assign n8796 = n8795 ^ n3609 ^ n3325 ;
  assign n8797 = ( ~n245 & n2173 ) | ( ~n245 & n4380 ) | ( n2173 & n4380 ) ;
  assign n8798 = n8797 ^ n6926 ^ n812 ;
  assign n8799 = ( ~n8794 & n8796 ) | ( ~n8794 & n8798 ) | ( n8796 & n8798 ) ;
  assign n8800 = ( n2083 & n8793 ) | ( n2083 & n8799 ) | ( n8793 & n8799 ) ;
  assign n8801 = ( n1014 & ~n1206 ) | ( n1014 & n1470 ) | ( ~n1206 & n1470 ) ;
  assign n8802 = ( ~n3064 & n3940 ) | ( ~n3064 & n8159 ) | ( n3940 & n8159 ) ;
  assign n8803 = n8802 ^ n5940 ^ n5790 ;
  assign n8804 = ( n241 & n2556 ) | ( n241 & ~n8803 ) | ( n2556 & ~n8803 ) ;
  assign n8805 = n8801 | n8804 ;
  assign n8806 = ( n1059 & n1558 ) | ( n1059 & n3942 ) | ( n1558 & n3942 ) ;
  assign n8807 = ( n2641 & n5998 ) | ( n2641 & ~n8806 ) | ( n5998 & ~n8806 ) ;
  assign n8808 = n8807 ^ n8594 ^ n7257 ;
  assign n8809 = ( x37 & ~n654 ) | ( x37 & n4298 ) | ( ~n654 & n4298 ) ;
  assign n8810 = n8809 ^ n6688 ^ n3735 ;
  assign n8811 = n8810 ^ n3763 ^ n2459 ;
  assign n8812 = ~n5361 & n8811 ;
  assign n8813 = n6649 ^ n3510 ^ n486 ;
  assign n8814 = n8813 ^ n2295 ^ 1'b0 ;
  assign n8815 = ( n7706 & n8165 ) | ( n7706 & n8814 ) | ( n8165 & n8814 ) ;
  assign n8816 = ( n3711 & n5038 ) | ( n3711 & ~n5180 ) | ( n5038 & ~n5180 ) ;
  assign n8817 = ( ~n4089 & n4807 ) | ( ~n4089 & n8816 ) | ( n4807 & n8816 ) ;
  assign n8818 = ~n8815 & n8817 ;
  assign n8819 = n502 & n8818 ;
  assign n8820 = n6458 ^ n5237 ^ n3401 ;
  assign n8821 = ( n3521 & n6136 ) | ( n3521 & n8820 ) | ( n6136 & n8820 ) ;
  assign n8822 = n7164 ^ n1278 ^ 1'b0 ;
  assign n8823 = n8821 & ~n8822 ;
  assign n8824 = n6059 & n8823 ;
  assign n8825 = ~n7689 & n8824 ;
  assign n8826 = n7476 ^ n2353 ^ n1843 ;
  assign n8831 = ( n1342 & n1752 ) | ( n1342 & ~n3998 ) | ( n1752 & ~n3998 ) ;
  assign n8832 = ( n170 & ~n2266 ) | ( n170 & n6893 ) | ( ~n2266 & n6893 ) ;
  assign n8834 = ( n3215 & n3400 ) | ( n3215 & n4348 ) | ( n3400 & n4348 ) ;
  assign n8833 = ( x20 & ~n2357 ) | ( x20 & n3300 ) | ( ~n2357 & n3300 ) ;
  assign n8835 = n8834 ^ n8833 ^ n4947 ;
  assign n8836 = ( n8831 & n8832 ) | ( n8831 & n8835 ) | ( n8832 & n8835 ) ;
  assign n8829 = ( n681 & n1161 ) | ( n681 & n3635 ) | ( n1161 & n3635 ) ;
  assign n8827 = ( n1305 & n5111 ) | ( n1305 & n7400 ) | ( n5111 & n7400 ) ;
  assign n8828 = ( n5441 & n6453 ) | ( n5441 & n8827 ) | ( n6453 & n8827 ) ;
  assign n8830 = n8829 ^ n8828 ^ n6275 ;
  assign n8837 = n8836 ^ n8830 ^ n7350 ;
  assign n8839 = n1494 ^ n343 ^ 1'b0 ;
  assign n8838 = n8626 ^ n7450 ^ n3357 ;
  assign n8840 = n8839 ^ n8838 ^ n5021 ;
  assign n8841 = n917 & ~n8840 ;
  assign n8842 = n4153 & n8841 ;
  assign n8843 = n8842 ^ n8295 ^ n2389 ;
  assign n8844 = n4530 ^ n4515 ^ n2035 ;
  assign n8845 = n8844 ^ n2905 ^ n1362 ;
  assign n8846 = n8101 ^ n6432 ^ 1'b0 ;
  assign n8847 = n8845 & ~n8846 ;
  assign n8848 = ( n1385 & ~n2574 ) | ( n1385 & n4058 ) | ( ~n2574 & n4058 ) ;
  assign n8849 = ( n1282 & n1802 ) | ( n1282 & n3589 ) | ( n1802 & n3589 ) ;
  assign n8850 = ( n260 & ~n8848 ) | ( n260 & n8849 ) | ( ~n8848 & n8849 ) ;
  assign n8851 = n8850 ^ n2551 ^ n1293 ;
  assign n8852 = n5639 & n8851 ;
  assign n8853 = n8852 ^ n3628 ^ n542 ;
  assign n8854 = ( n6095 & n7827 ) | ( n6095 & ~n8853 ) | ( n7827 & ~n8853 ) ;
  assign n8855 = ( ~n8131 & n8847 ) | ( ~n8131 & n8854 ) | ( n8847 & n8854 ) ;
  assign n8856 = ( n1913 & n2266 ) | ( n1913 & n2931 ) | ( n2266 & n2931 ) ;
  assign n8857 = n8856 ^ n4757 ^ n2106 ;
  assign n8858 = ( ~n2003 & n5723 ) | ( ~n2003 & n5775 ) | ( n5723 & n5775 ) ;
  assign n8859 = n8858 ^ n6158 ^ 1'b0 ;
  assign n8860 = n8857 | n8859 ;
  assign n8861 = n1122 | n8860 ;
  assign n8863 = n7363 ^ n6984 ^ n788 ;
  assign n8862 = n8530 ^ n6537 ^ n5564 ;
  assign n8864 = n8863 ^ n8862 ^ n386 ;
  assign n8865 = ( n8035 & n8861 ) | ( n8035 & n8864 ) | ( n8861 & n8864 ) ;
  assign n8866 = n5457 ^ n1095 ^ 1'b0 ;
  assign n8868 = n4126 | n8623 ;
  assign n8869 = n8868 ^ n8153 ^ 1'b0 ;
  assign n8867 = ( n6521 & n8352 ) | ( n6521 & n8608 ) | ( n8352 & n8608 ) ;
  assign n8870 = n8869 ^ n8867 ^ n1135 ;
  assign n8871 = ( n8865 & ~n8866 ) | ( n8865 & n8870 ) | ( ~n8866 & n8870 ) ;
  assign n8877 = n5379 ^ n1863 ^ n1288 ;
  assign n8874 = n2399 ^ n362 ^ 1'b0 ;
  assign n8875 = ( n3351 & n5765 ) | ( n3351 & ~n8874 ) | ( n5765 & ~n8874 ) ;
  assign n8876 = ~n922 & n8875 ;
  assign n8878 = n8877 ^ n8876 ^ 1'b0 ;
  assign n8872 = ( ~n1774 & n2014 ) | ( ~n1774 & n3158 ) | ( n2014 & n3158 ) ;
  assign n8873 = ( n2843 & n7803 ) | ( n2843 & n8872 ) | ( n7803 & n8872 ) ;
  assign n8879 = n8878 ^ n8873 ^ 1'b0 ;
  assign n8880 = n450 & ~n4064 ;
  assign n8881 = n4896 & n8880 ;
  assign n8882 = ( ~n5063 & n6028 ) | ( ~n5063 & n8881 ) | ( n6028 & n8881 ) ;
  assign n8886 = n5791 ^ n3555 ^ n2833 ;
  assign n8885 = n5128 ^ n4505 ^ n1587 ;
  assign n8887 = n8886 ^ n8885 ^ 1'b0 ;
  assign n8883 = n6542 ^ n3103 ^ n2150 ;
  assign n8884 = n2072 & n8883 ;
  assign n8888 = n8887 ^ n8884 ^ n376 ;
  assign n8889 = ( n3728 & ~n4685 ) | ( n3728 & n8294 ) | ( ~n4685 & n8294 ) ;
  assign n8890 = n8889 ^ n8463 ^ n5758 ;
  assign n8891 = n6569 & n8890 ;
  assign n8892 = n2039 & n8891 ;
  assign n8894 = n967 & n1822 ;
  assign n8895 = n8894 ^ n5930 ^ 1'b0 ;
  assign n8896 = n8895 ^ n5411 ^ n3951 ;
  assign n8893 = ~n187 & n2775 ;
  assign n8897 = n8896 ^ n8893 ^ 1'b0 ;
  assign n8898 = ( n6283 & ~n8486 ) | ( n6283 & n8897 ) | ( ~n8486 & n8897 ) ;
  assign n8899 = n3253 ^ n2615 ^ n2575 ;
  assign n8900 = n1099 | n6012 ;
  assign n8901 = ( ~n619 & n3101 ) | ( ~n619 & n7647 ) | ( n3101 & n7647 ) ;
  assign n8902 = n480 & ~n2040 ;
  assign n8903 = ( n3470 & ~n8901 ) | ( n3470 & n8902 ) | ( ~n8901 & n8902 ) ;
  assign n8904 = ( ~n2975 & n4334 ) | ( ~n2975 & n8903 ) | ( n4334 & n8903 ) ;
  assign n8905 = n8904 ^ n8653 ^ n2143 ;
  assign n8906 = n3276 ^ n2839 ^ n1522 ;
  assign n8907 = n7349 | n8906 ;
  assign n8908 = ( ~n8900 & n8905 ) | ( ~n8900 & n8907 ) | ( n8905 & n8907 ) ;
  assign n8909 = ( ~n4020 & n8899 ) | ( ~n4020 & n8908 ) | ( n8899 & n8908 ) ;
  assign n8910 = n7137 ^ n3759 ^ 1'b0 ;
  assign n8913 = n6299 ^ n2378 ^ 1'b0 ;
  assign n8914 = n8913 ^ n4512 ^ n2411 ;
  assign n8912 = n8778 ^ n3039 ^ n767 ;
  assign n8911 = ( n454 & n1094 ) | ( n454 & ~n5066 ) | ( n1094 & ~n5066 ) ;
  assign n8915 = n8914 ^ n8912 ^ n8911 ;
  assign n8916 = ( ~n5500 & n8910 ) | ( ~n5500 & n8915 ) | ( n8910 & n8915 ) ;
  assign n8917 = n7767 ^ n4798 ^ n4265 ;
  assign n8918 = n8917 ^ n3007 ^ 1'b0 ;
  assign n8919 = n5385 & n8918 ;
  assign n8929 = n3119 ^ n2219 ^ n351 ;
  assign n8920 = ( n943 & ~n2931 ) | ( n943 & n4979 ) | ( ~n2931 & n4979 ) ;
  assign n8921 = ( n779 & n2195 ) | ( n779 & n8920 ) | ( n2195 & n8920 ) ;
  assign n8922 = ( n1113 & n1965 ) | ( n1113 & ~n2460 ) | ( n1965 & ~n2460 ) ;
  assign n8923 = n8922 ^ n5227 ^ n3736 ;
  assign n8924 = ( n196 & n838 ) | ( n196 & ~n1119 ) | ( n838 & ~n1119 ) ;
  assign n8925 = n8924 ^ n1734 ^ 1'b0 ;
  assign n8926 = n8925 ^ n5258 ^ n1600 ;
  assign n8927 = n8926 ^ n8225 ^ n4265 ;
  assign n8928 = ( n8921 & n8923 ) | ( n8921 & ~n8927 ) | ( n8923 & ~n8927 ) ;
  assign n8930 = n8929 ^ n8928 ^ n8799 ;
  assign n8931 = n740 & ~n2518 ;
  assign n8932 = n8931 ^ n283 ^ 1'b0 ;
  assign n8933 = n8932 ^ n6289 ^ n3841 ;
  assign n8934 = n4840 ^ n1286 ^ n586 ;
  assign n8935 = n1927 ^ n659 ^ n469 ;
  assign n8936 = ( n8653 & n8934 ) | ( n8653 & n8935 ) | ( n8934 & n8935 ) ;
  assign n8937 = ( n6638 & ~n8933 ) | ( n6638 & n8936 ) | ( ~n8933 & n8936 ) ;
  assign n8942 = n3535 ^ n2140 ^ n2011 ;
  assign n8943 = n8942 ^ n6099 ^ n3071 ;
  assign n8938 = n1661 ^ n909 ^ n788 ;
  assign n8939 = n8938 ^ n3519 ^ n1113 ;
  assign n8940 = ( n1104 & n1436 ) | ( n1104 & ~n8939 ) | ( n1436 & ~n8939 ) ;
  assign n8941 = n8940 ^ n8059 ^ n4589 ;
  assign n8944 = n8943 ^ n8941 ^ x32 ;
  assign n8945 = n8622 ^ n3518 ^ n2021 ;
  assign n8947 = n4099 ^ n575 ^ n300 ;
  assign n8946 = n1032 & ~n7137 ;
  assign n8948 = n8947 ^ n8946 ^ n4269 ;
  assign n8949 = n6132 & n6821 ;
  assign n8950 = ( n898 & n3126 ) | ( n898 & n7389 ) | ( n3126 & n7389 ) ;
  assign n8951 = n2759 ^ x83 ^ 1'b0 ;
  assign n8952 = ( n826 & ~n1602 ) | ( n826 & n8951 ) | ( ~n1602 & n8951 ) ;
  assign n8953 = ( n4669 & n8422 ) | ( n4669 & n8952 ) | ( n8422 & n8952 ) ;
  assign n8954 = ( n1492 & ~n3827 ) | ( n1492 & n7229 ) | ( ~n3827 & n7229 ) ;
  assign n8955 = ( n1802 & n8953 ) | ( n1802 & n8954 ) | ( n8953 & n8954 ) ;
  assign n8956 = ( ~n1283 & n8950 ) | ( ~n1283 & n8955 ) | ( n8950 & n8955 ) ;
  assign n8957 = n8191 | n8956 ;
  assign n8958 = n6234 ^ n2722 ^ n1138 ;
  assign n8959 = n8958 ^ n5741 ^ n5027 ;
  assign n8960 = ( n1044 & n2204 ) | ( n1044 & ~n5917 ) | ( n2204 & ~n5917 ) ;
  assign n8961 = n2905 & n3244 ;
  assign n8962 = ~n8960 & n8961 ;
  assign n8963 = ~n7737 & n8962 ;
  assign n8964 = ( n8460 & n8959 ) | ( n8460 & n8963 ) | ( n8959 & n8963 ) ;
  assign n8970 = n289 & ~n880 ;
  assign n8971 = ~x96 & n8970 ;
  assign n8972 = ( x20 & n5159 ) | ( x20 & n8971 ) | ( n5159 & n8971 ) ;
  assign n8965 = ( n1823 & n2665 ) | ( n1823 & n6828 ) | ( n2665 & n6828 ) ;
  assign n8966 = n8965 ^ n2890 ^ n834 ;
  assign n8967 = ~n5578 & n6959 ;
  assign n8968 = ( n2187 & ~n6566 ) | ( n2187 & n8967 ) | ( ~n6566 & n8967 ) ;
  assign n8969 = ~n8966 & n8968 ;
  assign n8973 = n8972 ^ n8969 ^ n7656 ;
  assign n8974 = ( ~n2596 & n3600 ) | ( ~n2596 & n7371 ) | ( n3600 & n7371 ) ;
  assign n8975 = n2881 & ~n8974 ;
  assign n8976 = n8975 ^ n6621 ^ 1'b0 ;
  assign n8977 = ( n997 & n4425 ) | ( n997 & ~n4868 ) | ( n4425 & ~n4868 ) ;
  assign n8978 = n7504 ^ n1466 ^ n307 ;
  assign n8980 = ( n2507 & ~n3289 ) | ( n2507 & n4221 ) | ( ~n3289 & n4221 ) ;
  assign n8979 = n6249 ^ n3471 ^ n2055 ;
  assign n8981 = n8980 ^ n8979 ^ n7407 ;
  assign n8982 = n4183 ^ n2960 ^ n255 ;
  assign n8983 = ( ~n8405 & n8981 ) | ( ~n8405 & n8982 ) | ( n8981 & n8982 ) ;
  assign n8984 = n8983 ^ n8627 ^ n7432 ;
  assign n8985 = ( n7906 & n8978 ) | ( n7906 & n8984 ) | ( n8978 & n8984 ) ;
  assign n8990 = n6998 ^ n3970 ^ n166 ;
  assign n8991 = ( n3553 & n5363 ) | ( n3553 & ~n8990 ) | ( n5363 & ~n8990 ) ;
  assign n8992 = n8991 ^ n748 ^ n474 ;
  assign n8986 = n4015 ^ n2253 ^ n144 ;
  assign n8987 = n1810 ^ n822 ^ n793 ;
  assign n8988 = ( n4693 & n4800 ) | ( n4693 & n8987 ) | ( n4800 & n8987 ) ;
  assign n8989 = n8986 & n8988 ;
  assign n8993 = n8992 ^ n8989 ^ 1'b0 ;
  assign n8994 = n8993 ^ n5590 ^ n2771 ;
  assign n8995 = ( n1446 & ~n2756 ) | ( n1446 & n8537 ) | ( ~n2756 & n8537 ) ;
  assign n8996 = n2594 ^ n2019 ^ n1441 ;
  assign n8997 = n8996 ^ n8354 ^ n7356 ;
  assign n8998 = ( ~n359 & n8995 ) | ( ~n359 & n8997 ) | ( n8995 & n8997 ) ;
  assign n8999 = n5566 ^ n1638 ^ n1207 ;
  assign n9001 = ( x12 & n815 ) | ( x12 & n1195 ) | ( n815 & n1195 ) ;
  assign n9002 = n4342 ^ n1223 ^ 1'b0 ;
  assign n9003 = ~n9001 & n9002 ;
  assign n9004 = ( n1240 & n5898 ) | ( n1240 & ~n6504 ) | ( n5898 & ~n6504 ) ;
  assign n9005 = n9004 ^ n4676 ^ n3576 ;
  assign n9006 = ( n1915 & n9003 ) | ( n1915 & n9005 ) | ( n9003 & n9005 ) ;
  assign n9000 = ( n679 & n2290 ) | ( n679 & ~n8361 ) | ( n2290 & ~n8361 ) ;
  assign n9007 = n9006 ^ n9000 ^ n514 ;
  assign n9008 = n9007 ^ n6172 ^ n1852 ;
  assign n9009 = ( n6840 & ~n8999 ) | ( n6840 & n9008 ) | ( ~n8999 & n9008 ) ;
  assign n9010 = ( n1074 & ~n8998 ) | ( n1074 & n9009 ) | ( ~n8998 & n9009 ) ;
  assign n9016 = ( ~n1988 & n4055 ) | ( ~n1988 & n4797 ) | ( n4055 & n4797 ) ;
  assign n9017 = n9016 ^ n4258 ^ x52 ;
  assign n9011 = n1521 & n5063 ;
  assign n9012 = ~n1044 & n9011 ;
  assign n9013 = ( n856 & n1384 ) | ( n856 & ~n3821 ) | ( n1384 & ~n3821 ) ;
  assign n9014 = ( n7845 & n9012 ) | ( n7845 & n9013 ) | ( n9012 & n9013 ) ;
  assign n9015 = ( n2338 & n6194 ) | ( n2338 & ~n9014 ) | ( n6194 & ~n9014 ) ;
  assign n9018 = n9017 ^ n9015 ^ n4050 ;
  assign n9021 = n5503 ^ n2491 ^ 1'b0 ;
  assign n9022 = ~n1238 & n9021 ;
  assign n9020 = ( ~n3803 & n5365 ) | ( ~n3803 & n7266 ) | ( n5365 & n7266 ) ;
  assign n9023 = n9022 ^ n9020 ^ 1'b0 ;
  assign n9024 = n2298 & ~n9023 ;
  assign n9025 = n9024 ^ n7618 ^ n2922 ;
  assign n9019 = ( n1099 & ~n1909 ) | ( n1099 & n3713 ) | ( ~n1909 & n3713 ) ;
  assign n9026 = n9025 ^ n9019 ^ n8473 ;
  assign n9027 = ( n540 & n2583 ) | ( n540 & n3725 ) | ( n2583 & n3725 ) ;
  assign n9028 = n9027 ^ n7374 ^ n2257 ;
  assign n9029 = ( ~n2151 & n5745 ) | ( ~n2151 & n9028 ) | ( n5745 & n9028 ) ;
  assign n9030 = ~n5378 & n6336 ;
  assign n9031 = ( ~n1009 & n9029 ) | ( ~n1009 & n9030 ) | ( n9029 & n9030 ) ;
  assign n9032 = n1259 & ~n9014 ;
  assign n9033 = n3267 & ~n8086 ;
  assign n9034 = n7021 ^ n5667 ^ n4838 ;
  assign n9035 = n3111 ^ n1978 ^ 1'b0 ;
  assign n9036 = n2941 ^ n2906 ^ n1362 ;
  assign n9037 = ( n549 & n9035 ) | ( n549 & n9036 ) | ( n9035 & n9036 ) ;
  assign n9038 = ( n1774 & n9034 ) | ( n1774 & n9037 ) | ( n9034 & n9037 ) ;
  assign n9039 = n9038 ^ n8518 ^ n8366 ;
  assign n9040 = n4789 ^ n137 ^ x65 ;
  assign n9041 = ( n2684 & n3431 ) | ( n2684 & n9040 ) | ( n3431 & n9040 ) ;
  assign n9042 = n2756 ^ n146 ^ 1'b0 ;
  assign n9043 = n9042 ^ n2216 ^ n1261 ;
  assign n9044 = n9043 ^ n8807 ^ 1'b0 ;
  assign n9045 = n9044 ^ n7718 ^ n203 ;
  assign n9046 = n5003 ^ n1034 ^ 1'b0 ;
  assign n9047 = n907 & ~n4582 ;
  assign n9048 = n9046 & n9047 ;
  assign n9049 = n9048 ^ n4796 ^ n4018 ;
  assign n9050 = ( n2612 & n5005 ) | ( n2612 & n6157 ) | ( n5005 & n6157 ) ;
  assign n9051 = n9050 ^ n5069 ^ n1750 ;
  assign n9052 = ( n1048 & n3268 ) | ( n1048 & ~n9051 ) | ( n3268 & ~n9051 ) ;
  assign n9053 = ( n1113 & n5833 ) | ( n1113 & n9052 ) | ( n5833 & n9052 ) ;
  assign n9054 = n3798 ^ n3369 ^ n2917 ;
  assign n9055 = n2496 & ~n9054 ;
  assign n9056 = n9055 ^ n8009 ^ 1'b0 ;
  assign n9057 = n9056 ^ x102 ^ 1'b0 ;
  assign n9058 = n1394 & n9057 ;
  assign n9059 = n9058 ^ n3570 ^ x22 ;
  assign n9060 = n7548 ^ n5476 ^ n1067 ;
  assign n9068 = n2605 & n3658 ;
  assign n9069 = n563 & ~n9068 ;
  assign n9061 = n8934 ^ n6600 ^ n1920 ;
  assign n9064 = ( ~n2146 & n2344 ) | ( ~n2146 & n7274 ) | ( n2344 & n7274 ) ;
  assign n9062 = n7929 ^ n6455 ^ n852 ;
  assign n9063 = n3709 | n9062 ;
  assign n9065 = n9064 ^ n9063 ^ 1'b0 ;
  assign n9066 = ( n3294 & n8702 ) | ( n3294 & ~n9065 ) | ( n8702 & ~n9065 ) ;
  assign n9067 = ( ~n6874 & n9061 ) | ( ~n6874 & n9066 ) | ( n9061 & n9066 ) ;
  assign n9070 = n9069 ^ n9067 ^ n7441 ;
  assign n9071 = n9070 ^ n2218 ^ x124 ;
  assign n9072 = n5043 ^ n2537 ^ 1'b0 ;
  assign n9073 = n3023 & n9072 ;
  assign n9075 = n3053 | n3814 ;
  assign n9076 = ( ~n314 & n3747 ) | ( ~n314 & n9075 ) | ( n3747 & n9075 ) ;
  assign n9074 = ( ~n2889 & n2954 ) | ( ~n2889 & n6475 ) | ( n2954 & n6475 ) ;
  assign n9077 = n9076 ^ n9074 ^ 1'b0 ;
  assign n9078 = ( n7190 & ~n9073 ) | ( n7190 & n9077 ) | ( ~n9073 & n9077 ) ;
  assign n9079 = ( x113 & n3139 ) | ( x113 & ~n4739 ) | ( n3139 & ~n4739 ) ;
  assign n9081 = ~n2011 & n2015 ;
  assign n9082 = n9081 ^ n848 ^ 1'b0 ;
  assign n9080 = ( n4032 & ~n6411 ) | ( n4032 & n7903 ) | ( ~n6411 & n7903 ) ;
  assign n9083 = n9082 ^ n9080 ^ 1'b0 ;
  assign n9084 = n6922 & n9083 ;
  assign n9085 = ( n7934 & ~n9079 ) | ( n7934 & n9084 ) | ( ~n9079 & n9084 ) ;
  assign n9090 = n7037 ^ n3597 ^ n1856 ;
  assign n9091 = ( n187 & ~n7389 ) | ( n187 & n9090 ) | ( ~n7389 & n9090 ) ;
  assign n9086 = n5398 ^ n2687 ^ 1'b0 ;
  assign n9087 = n2148 & ~n9086 ;
  assign n9088 = n9087 ^ n2649 ^ 1'b0 ;
  assign n9089 = n1988 & n9088 ;
  assign n9092 = n9091 ^ n9089 ^ n5840 ;
  assign n9093 = n5403 ^ n4629 ^ 1'b0 ;
  assign n9094 = n2490 & ~n9093 ;
  assign n9095 = n2976 ^ n2431 ^ 1'b0 ;
  assign n9096 = n9095 ^ n7322 ^ n135 ;
  assign n9097 = ( ~n1037 & n1135 ) | ( ~n1037 & n9096 ) | ( n1135 & n9096 ) ;
  assign n9098 = ( n3186 & n9094 ) | ( n3186 & ~n9097 ) | ( n9094 & ~n9097 ) ;
  assign n9099 = ~n3619 & n9098 ;
  assign n9100 = n9092 & n9099 ;
  assign n9101 = n3602 ^ n3560 ^ 1'b0 ;
  assign n9102 = ~n1075 & n9101 ;
  assign n9103 = n5658 & n9102 ;
  assign n9104 = n9103 ^ n6541 ^ n705 ;
  assign n9105 = n7029 ^ n6729 ^ n2923 ;
  assign n9106 = ( n8595 & n8666 ) | ( n8595 & ~n9105 ) | ( n8666 & ~n9105 ) ;
  assign n9107 = ( n309 & ~n7570 ) | ( n309 & n8454 ) | ( ~n7570 & n8454 ) ;
  assign n9108 = ( n630 & ~n7921 ) | ( n630 & n9107 ) | ( ~n7921 & n9107 ) ;
  assign n9109 = n5233 ^ n1743 ^ n547 ;
  assign n9110 = n9109 ^ n7817 ^ n6880 ;
  assign n9112 = ( n2742 & ~n5060 ) | ( n2742 & n7866 ) | ( ~n5060 & n7866 ) ;
  assign n9111 = n2275 | n7978 ;
  assign n9113 = n9112 ^ n9111 ^ n6935 ;
  assign n9114 = ( n752 & ~n2595 ) | ( n752 & n3762 ) | ( ~n2595 & n3762 ) ;
  assign n9115 = ( n1968 & ~n8624 ) | ( n1968 & n8713 ) | ( ~n8624 & n8713 ) ;
  assign n9116 = ( ~n3890 & n9114 ) | ( ~n3890 & n9115 ) | ( n9114 & n9115 ) ;
  assign n9117 = n4213 & n6697 ;
  assign n9120 = ~n1457 & n1738 ;
  assign n9121 = n9120 ^ n2372 ^ 1'b0 ;
  assign n9122 = n9121 ^ n8748 ^ n4184 ;
  assign n9118 = ( x21 & ~n191 ) | ( x21 & n1573 ) | ( ~n191 & n1573 ) ;
  assign n9119 = ( n199 & n7140 ) | ( n199 & n9118 ) | ( n7140 & n9118 ) ;
  assign n9123 = n9122 ^ n9119 ^ n7944 ;
  assign n9130 = ( n227 & n2144 ) | ( n227 & ~n8642 ) | ( n2144 & ~n8642 ) ;
  assign n9126 = n1545 & ~n2660 ;
  assign n9127 = n9126 ^ n1255 ^ 1'b0 ;
  assign n9128 = n9127 ^ n7299 ^ n2188 ;
  assign n9124 = ( x112 & n3609 ) | ( x112 & ~n5649 ) | ( n3609 & ~n5649 ) ;
  assign n9125 = ( n2286 & n3708 ) | ( n2286 & ~n9124 ) | ( n3708 & ~n9124 ) ;
  assign n9129 = n9128 ^ n9125 ^ n2387 ;
  assign n9131 = n9130 ^ n9129 ^ n3111 ;
  assign n9132 = n9131 ^ n2490 ^ 1'b0 ;
  assign n9133 = n8458 ^ n6697 ^ n6435 ;
  assign n9134 = ~n6922 & n9046 ;
  assign n9135 = n9134 ^ n5339 ^ n3438 ;
  assign n9136 = n9135 ^ n3688 ^ n657 ;
  assign n9137 = ( ~n4945 & n5860 ) | ( ~n4945 & n7184 ) | ( n5860 & n7184 ) ;
  assign n9138 = ( ~n7311 & n9136 ) | ( ~n7311 & n9137 ) | ( n9136 & n9137 ) ;
  assign n9139 = ( n5079 & ~n9133 ) | ( n5079 & n9138 ) | ( ~n9133 & n9138 ) ;
  assign n9146 = ( n826 & n3573 ) | ( n826 & ~n4157 ) | ( n3573 & ~n4157 ) ;
  assign n9143 = ( n1301 & n1771 ) | ( n1301 & n5725 ) | ( n1771 & n5725 ) ;
  assign n9144 = n2129 | n9143 ;
  assign n9145 = n9144 ^ n1912 ^ 1'b0 ;
  assign n9140 = n1793 ^ n1371 ^ x57 ;
  assign n9141 = ( ~n2143 & n6586 ) | ( ~n2143 & n7753 ) | ( n6586 & n7753 ) ;
  assign n9142 = ( ~n6483 & n9140 ) | ( ~n6483 & n9141 ) | ( n9140 & n9141 ) ;
  assign n9147 = n9146 ^ n9145 ^ n9142 ;
  assign n9148 = n3578 & ~n9147 ;
  assign n9149 = n7240 & n9148 ;
  assign n9150 = n9149 ^ n7406 ^ n4775 ;
  assign n9151 = ( n3238 & n5806 ) | ( n3238 & ~n7443 ) | ( n5806 & ~n7443 ) ;
  assign n9152 = ( ~n2563 & n3224 ) | ( ~n2563 & n9151 ) | ( n3224 & n9151 ) ;
  assign n9153 = n5607 ^ n3719 ^ n1841 ;
  assign n9154 = n9153 ^ n8274 ^ n4338 ;
  assign n9157 = n644 & ~n2239 ;
  assign n9158 = n9157 ^ n3550 ^ 1'b0 ;
  assign n9159 = ( ~n781 & n7887 ) | ( ~n781 & n9158 ) | ( n7887 & n9158 ) ;
  assign n9155 = n5809 ^ n5434 ^ n3328 ;
  assign n9156 = n9155 ^ n8960 ^ n388 ;
  assign n9160 = n9159 ^ n9156 ^ n4379 ;
  assign n9161 = n7854 ^ n6974 ^ n3229 ;
  assign n9162 = ~n273 & n3083 ;
  assign n9163 = n9161 & n9162 ;
  assign n9164 = ( n3516 & ~n4498 ) | ( n3516 & n6785 ) | ( ~n4498 & n6785 ) ;
  assign n9165 = ( n5507 & ~n6553 ) | ( n5507 & n9164 ) | ( ~n6553 & n9164 ) ;
  assign n9166 = n6613 ^ n5062 ^ n2025 ;
  assign n9167 = n9166 ^ n1497 ^ n267 ;
  assign n9168 = ( n5350 & n7721 ) | ( n5350 & ~n9167 ) | ( n7721 & ~n9167 ) ;
  assign n9169 = ( n1044 & n6625 ) | ( n1044 & n9168 ) | ( n6625 & n9168 ) ;
  assign n9174 = n3601 ^ n2801 ^ n569 ;
  assign n9175 = ( n2811 & n7121 ) | ( n2811 & n9174 ) | ( n7121 & n9174 ) ;
  assign n9170 = n6701 ^ n6012 ^ n4488 ;
  assign n9171 = ( n592 & ~n792 ) | ( n592 & n3708 ) | ( ~n792 & n3708 ) ;
  assign n9172 = ( n5038 & ~n9170 ) | ( n5038 & n9171 ) | ( ~n9170 & n9171 ) ;
  assign n9173 = ( n2531 & n5792 ) | ( n2531 & ~n9172 ) | ( n5792 & ~n9172 ) ;
  assign n9176 = n9175 ^ n9173 ^ 1'b0 ;
  assign n9177 = n8327 & ~n9176 ;
  assign n9178 = ( n1023 & n2615 ) | ( n1023 & n2663 ) | ( n2615 & n2663 ) ;
  assign n9179 = n9178 ^ n4481 ^ 1'b0 ;
  assign n9180 = n7139 & ~n9179 ;
  assign n9184 = ( n3352 & n4137 ) | ( n3352 & ~n4472 ) | ( n4137 & ~n4472 ) ;
  assign n9182 = n7755 ^ n4670 ^ x113 ;
  assign n9183 = n9182 ^ n446 ^ 1'b0 ;
  assign n9181 = n7748 ^ n5274 ^ n5258 ;
  assign n9185 = n9184 ^ n9183 ^ n9181 ;
  assign n9186 = ( x57 & ~n9180 ) | ( x57 & n9185 ) | ( ~n9180 & n9185 ) ;
  assign n9189 = n8758 ^ n8378 ^ n4739 ;
  assign n9190 = ( n3099 & ~n3686 ) | ( n3099 & n9189 ) | ( ~n3686 & n9189 ) ;
  assign n9187 = ~n2958 & n6970 ;
  assign n9188 = ~n4135 & n9187 ;
  assign n9191 = n9190 ^ n9188 ^ n6292 ;
  assign n9198 = ( n1202 & n3613 ) | ( n1202 & n5281 ) | ( n3613 & n5281 ) ;
  assign n9192 = n5166 ^ n1798 ^ n730 ;
  assign n9193 = ( n3720 & n5846 ) | ( n3720 & ~n9192 ) | ( n5846 & ~n9192 ) ;
  assign n9194 = n9193 ^ n7335 ^ n1588 ;
  assign n9195 = n5180 ^ n2558 ^ n1361 ;
  assign n9196 = ~n1242 & n9195 ;
  assign n9197 = ~n9194 & n9196 ;
  assign n9199 = n9198 ^ n9197 ^ n852 ;
  assign n9200 = ( n411 & n2987 ) | ( n411 & ~n4880 ) | ( n2987 & ~n4880 ) ;
  assign n9201 = n9200 ^ n8151 ^ n5864 ;
  assign n9206 = n9173 ^ n850 ^ n319 ;
  assign n9204 = ( ~n503 & n1834 ) | ( ~n503 & n3717 ) | ( n1834 & n3717 ) ;
  assign n9202 = n1407 ^ n415 ^ 1'b0 ;
  assign n9203 = n9202 ^ n2816 ^ n1666 ;
  assign n9205 = n9204 ^ n9203 ^ n1709 ;
  assign n9207 = n9206 ^ n9205 ^ n7265 ;
  assign n9212 = n1895 ^ n1342 ^ n291 ;
  assign n9210 = n2597 ^ n2218 ^ 1'b0 ;
  assign n9211 = ~n3131 & n9210 ;
  assign n9208 = n3823 ^ n3694 ^ n3372 ;
  assign n9209 = n9208 ^ n9105 ^ n2139 ;
  assign n9213 = n9212 ^ n9211 ^ n9209 ;
  assign n9214 = n7485 ^ n4674 ^ n962 ;
  assign n9216 = n6235 ^ n660 ^ 1'b0 ;
  assign n9217 = n4399 | n9216 ;
  assign n9215 = ( n500 & ~n4493 ) | ( n500 & n8911 ) | ( ~n4493 & n8911 ) ;
  assign n9218 = n9217 ^ n9215 ^ n595 ;
  assign n9219 = ( ~n913 & n5359 ) | ( ~n913 & n5456 ) | ( n5359 & n5456 ) ;
  assign n9220 = ( ~n6502 & n8870 ) | ( ~n6502 & n9219 ) | ( n8870 & n9219 ) ;
  assign n9221 = ~n7283 & n8520 ;
  assign n9222 = n9221 ^ n4359 ^ 1'b0 ;
  assign n9223 = n9222 ^ n4361 ^ n1343 ;
  assign n9224 = ( n555 & n1586 ) | ( n555 & n4969 ) | ( n1586 & n4969 ) ;
  assign n9225 = n8074 ^ n1373 ^ x8 ;
  assign n9226 = ( n5463 & n6747 ) | ( n5463 & n9225 ) | ( n6747 & n9225 ) ;
  assign n9227 = n9224 | n9226 ;
  assign n9228 = n3461 | n9227 ;
  assign n9229 = n1681 | n7170 ;
  assign n9230 = n9229 ^ n3051 ^ n1030 ;
  assign n9231 = ( n4478 & n9228 ) | ( n4478 & ~n9230 ) | ( n9228 & ~n9230 ) ;
  assign n9232 = ( ~n844 & n5312 ) | ( ~n844 & n9231 ) | ( n5312 & n9231 ) ;
  assign n9233 = ( n5192 & n6855 ) | ( n5192 & n9232 ) | ( n6855 & n9232 ) ;
  assign n9234 = ( n4605 & n9223 ) | ( n4605 & n9233 ) | ( n9223 & n9233 ) ;
  assign n9235 = n986 & n2115 ;
  assign n9236 = ( n1233 & n1860 ) | ( n1233 & n9235 ) | ( n1860 & n9235 ) ;
  assign n9237 = ~n2232 & n8939 ;
  assign n9238 = n9237 ^ n7204 ^ n1695 ;
  assign n9247 = n4062 ^ n482 ^ 1'b0 ;
  assign n9245 = n1418 & n3905 ;
  assign n9246 = n9245 ^ n7931 ^ n1360 ;
  assign n9239 = n4945 ^ n1878 ^ x15 ;
  assign n9240 = ( ~n4618 & n5088 ) | ( ~n4618 & n5880 ) | ( n5088 & n5880 ) ;
  assign n9241 = n9240 ^ n5294 ^ n1822 ;
  assign n9242 = ( n677 & n9239 ) | ( n677 & n9241 ) | ( n9239 & n9241 ) ;
  assign n9243 = n4618 & n6097 ;
  assign n9244 = n9242 & n9243 ;
  assign n9248 = n9247 ^ n9246 ^ n9244 ;
  assign n9249 = ( n1343 & ~n1846 ) | ( n1343 & n3349 ) | ( ~n1846 & n3349 ) ;
  assign n9250 = ( n3479 & ~n5587 ) | ( n3479 & n8294 ) | ( ~n5587 & n8294 ) ;
  assign n9251 = n9249 & ~n9250 ;
  assign n9252 = ~n2630 & n9251 ;
  assign n9253 = n5064 & ~n6118 ;
  assign n9254 = ~n1445 & n9253 ;
  assign n9255 = n6754 & ~n9254 ;
  assign n9256 = ~n4024 & n9255 ;
  assign n9259 = ( ~n328 & n1239 ) | ( ~n328 & n2085 ) | ( n1239 & n2085 ) ;
  assign n9257 = n3989 ^ n2595 ^ n1635 ;
  assign n9258 = ( n5785 & n7635 ) | ( n5785 & n9257 ) | ( n7635 & n9257 ) ;
  assign n9260 = n9259 ^ n9258 ^ n1545 ;
  assign n9261 = ( n5569 & n7805 ) | ( n5569 & ~n9260 ) | ( n7805 & ~n9260 ) ;
  assign n9262 = ( n3996 & n9256 ) | ( n3996 & n9261 ) | ( n9256 & n9261 ) ;
  assign n9263 = n5217 ^ n5019 ^ n2221 ;
  assign n9264 = n4225 ^ n438 ^ n135 ;
  assign n9265 = n9264 ^ n9024 ^ n3389 ;
  assign n9268 = ( n1146 & n1548 ) | ( n1146 & n2414 ) | ( n1548 & n2414 ) ;
  assign n9269 = n9268 ^ n2925 ^ n1318 ;
  assign n9266 = ~n1114 & n2168 ;
  assign n9267 = n9266 ^ n4884 ^ 1'b0 ;
  assign n9270 = n9269 ^ n9267 ^ n658 ;
  assign n9271 = ( n4162 & n9265 ) | ( n4162 & n9270 ) | ( n9265 & n9270 ) ;
  assign n9272 = n6172 & n6792 ;
  assign n9273 = n9272 ^ n2322 ^ 1'b0 ;
  assign n9274 = ( n432 & n764 ) | ( n432 & ~n4874 ) | ( n764 & ~n4874 ) ;
  assign n9275 = ( n1008 & ~n3625 ) | ( n1008 & n8885 ) | ( ~n3625 & n8885 ) ;
  assign n9276 = ( n1171 & n9274 ) | ( n1171 & n9275 ) | ( n9274 & n9275 ) ;
  assign n9277 = ( ~n6280 & n7792 ) | ( ~n6280 & n9276 ) | ( n7792 & n9276 ) ;
  assign n9278 = ( n3149 & n7687 ) | ( n3149 & ~n9277 ) | ( n7687 & ~n9277 ) ;
  assign n9279 = ( n2475 & ~n6428 ) | ( n2475 & n8275 ) | ( ~n6428 & n8275 ) ;
  assign n9280 = ( ~n223 & n6108 ) | ( ~n223 & n9279 ) | ( n6108 & n9279 ) ;
  assign n9281 = n9280 ^ n9178 ^ n8598 ;
  assign n9282 = ( n4665 & n9278 ) | ( n4665 & n9281 ) | ( n9278 & n9281 ) ;
  assign n9283 = ( n4034 & ~n5201 ) | ( n4034 & n7572 ) | ( ~n5201 & n7572 ) ;
  assign n9284 = n9283 ^ n5647 ^ n4878 ;
  assign n9285 = ( n1553 & ~n2967 ) | ( n1553 & n9284 ) | ( ~n2967 & n9284 ) ;
  assign n9286 = ( n354 & n1503 ) | ( n354 & ~n9285 ) | ( n1503 & ~n9285 ) ;
  assign n9287 = n9286 ^ n165 ^ x19 ;
  assign n9288 = n7922 ^ n7500 ^ n1447 ;
  assign n9289 = ( ~n5639 & n6979 ) | ( ~n5639 & n9288 ) | ( n6979 & n9288 ) ;
  assign n9290 = n670 & n3202 ;
  assign n9291 = n4812 & ~n9290 ;
  assign n9292 = n9291 ^ n8355 ^ 1'b0 ;
  assign n9293 = n3347 ^ n906 ^ 1'b0 ;
  assign n9294 = ~n9292 & n9293 ;
  assign n9295 = n8212 ^ n235 ^ 1'b0 ;
  assign n9296 = n9294 & n9295 ;
  assign n9297 = n3563 ^ n1440 ^ n1275 ;
  assign n9298 = n9297 ^ n3675 ^ 1'b0 ;
  assign n9299 = n1859 | n9298 ;
  assign n9300 = n5113 ^ n3869 ^ n2194 ;
  assign n9301 = ( n3244 & n4827 ) | ( n3244 & n6616 ) | ( n4827 & n6616 ) ;
  assign n9302 = ( n609 & ~n9300 ) | ( n609 & n9301 ) | ( ~n9300 & n9301 ) ;
  assign n9303 = ( n207 & ~n861 ) | ( n207 & n1630 ) | ( ~n861 & n1630 ) ;
  assign n9304 = n7787 & n9303 ;
  assign n9305 = n8295 ^ n3800 ^ 1'b0 ;
  assign n9306 = ( ~n945 & n2380 ) | ( ~n945 & n5131 ) | ( n2380 & n5131 ) ;
  assign n9307 = ( n2019 & n2073 ) | ( n2019 & ~n6998 ) | ( n2073 & ~n6998 ) ;
  assign n9308 = n7711 ^ n2500 ^ 1'b0 ;
  assign n9309 = n9307 & ~n9308 ;
  assign n9310 = ( n1644 & ~n9306 ) | ( n1644 & n9309 ) | ( ~n9306 & n9309 ) ;
  assign n9311 = n1361 & n5610 ;
  assign n9312 = ~n7693 & n9311 ;
  assign n9313 = n4628 ^ n2426 ^ n190 ;
  assign n9314 = n9313 ^ n5914 ^ n3229 ;
  assign n9315 = ( n1976 & n9312 ) | ( n1976 & n9314 ) | ( n9312 & n9314 ) ;
  assign n9316 = n2600 ^ n2357 ^ n1172 ;
  assign n9317 = ( ~n3231 & n9315 ) | ( ~n3231 & n9316 ) | ( n9315 & n9316 ) ;
  assign n9318 = ~n684 & n823 ;
  assign n9319 = n9318 ^ n6157 ^ 1'b0 ;
  assign n9320 = ~n9109 & n9319 ;
  assign n9321 = n9317 & n9320 ;
  assign n9322 = ( ~n3323 & n8899 ) | ( ~n3323 & n9321 ) | ( n8899 & n9321 ) ;
  assign n9323 = n9322 ^ n4291 ^ x116 ;
  assign n9324 = n7333 ^ n4960 ^ n2308 ;
  assign n9325 = n9324 ^ n8537 ^ n5649 ;
  assign n9326 = ( n2509 & ~n5446 ) | ( n2509 & n9325 ) | ( ~n5446 & n9325 ) ;
  assign n9327 = n2394 ^ n1328 ^ 1'b0 ;
  assign n9328 = n9327 ^ n8325 ^ n495 ;
  assign n9329 = n7158 ^ n4614 ^ n352 ;
  assign n9330 = n9329 ^ n719 ^ n709 ;
  assign n9331 = ( ~n688 & n9151 ) | ( ~n688 & n9330 ) | ( n9151 & n9330 ) ;
  assign n9332 = ( ~n1024 & n4133 ) | ( ~n1024 & n9331 ) | ( n4133 & n9331 ) ;
  assign n9333 = ( ~n3671 & n7382 ) | ( ~n3671 & n7600 ) | ( n7382 & n7600 ) ;
  assign n9334 = n9333 ^ n9264 ^ n1973 ;
  assign n9345 = n8035 ^ n3092 ^ 1'b0 ;
  assign n9346 = n7046 | n9345 ;
  assign n9342 = n3143 ^ n2871 ^ n1012 ;
  assign n9343 = n9342 ^ n2480 ^ 1'b0 ;
  assign n9344 = n9343 ^ n4019 ^ 1'b0 ;
  assign n9340 = n1230 ^ n1072 ^ n1002 ;
  assign n9336 = n6686 ^ n5369 ^ 1'b0 ;
  assign n9337 = n2332 | n9336 ;
  assign n9338 = n9337 ^ n567 ^ n168 ;
  assign n9339 = n9338 ^ n4679 ^ n293 ;
  assign n9335 = n4896 ^ n1854 ^ n601 ;
  assign n9341 = n9340 ^ n9339 ^ n9335 ;
  assign n9347 = n9346 ^ n9344 ^ n9341 ;
  assign n9348 = ( n3261 & n9334 ) | ( n3261 & n9347 ) | ( n9334 & n9347 ) ;
  assign n9349 = ( n4906 & n7411 ) | ( n4906 & n7810 ) | ( n7411 & n7810 ) ;
  assign n9350 = ( ~n3160 & n6155 ) | ( ~n3160 & n9349 ) | ( n6155 & n9349 ) ;
  assign n9360 = n3208 ^ n2958 ^ n705 ;
  assign n9361 = n9360 ^ n2795 ^ n1937 ;
  assign n9358 = x35 & n4860 ;
  assign n9359 = ~n7168 & n9358 ;
  assign n9356 = n3391 ^ n3010 ^ n1620 ;
  assign n9357 = n9356 ^ n3639 ^ 1'b0 ;
  assign n9362 = n9361 ^ n9359 ^ n9357 ;
  assign n9352 = ( ~n3359 & n3693 ) | ( ~n3359 & n7197 ) | ( n3693 & n7197 ) ;
  assign n9351 = n2443 ^ n1378 ^ n1165 ;
  assign n9353 = n9352 ^ n9351 ^ n5840 ;
  assign n9354 = ( n3323 & ~n6535 ) | ( n3323 & n9353 ) | ( ~n6535 & n9353 ) ;
  assign n9355 = n9354 ^ n5937 ^ n4860 ;
  assign n9363 = n9362 ^ n9355 ^ n1805 ;
  assign n9365 = n1461 ^ n907 ^ n704 ;
  assign n9364 = n6752 ^ n2397 ^ x7 ;
  assign n9366 = n9365 ^ n9364 ^ n1820 ;
  assign n9367 = ( n3699 & n4683 ) | ( n3699 & n5064 ) | ( n4683 & n5064 ) ;
  assign n9368 = n9367 ^ n1809 ^ n769 ;
  assign n9369 = ( n1770 & n2825 ) | ( n1770 & n2837 ) | ( n2825 & n2837 ) ;
  assign n9370 = ( ~x92 & n2695 ) | ( ~x92 & n3175 ) | ( n2695 & n3175 ) ;
  assign n9371 = n8159 ^ n3307 ^ 1'b0 ;
  assign n9372 = ( n1313 & ~n9370 ) | ( n1313 & n9371 ) | ( ~n9370 & n9371 ) ;
  assign n9373 = n8153 ^ n7392 ^ n1878 ;
  assign n9374 = ( n3371 & n4795 ) | ( n3371 & ~n5359 ) | ( n4795 & ~n5359 ) ;
  assign n9375 = ( n294 & n2641 ) | ( n294 & n7666 ) | ( n2641 & n7666 ) ;
  assign n9376 = ( n551 & n906 ) | ( n551 & n9375 ) | ( n906 & n9375 ) ;
  assign n9377 = ( ~n2390 & n9374 ) | ( ~n2390 & n9376 ) | ( n9374 & n9376 ) ;
  assign n9378 = ( n751 & ~n1152 ) | ( n751 & n8659 ) | ( ~n1152 & n8659 ) ;
  assign n9379 = n9378 ^ n7237 ^ n5992 ;
  assign n9380 = ( x127 & ~n2023 ) | ( x127 & n5695 ) | ( ~n2023 & n5695 ) ;
  assign n9381 = n9380 ^ n2265 ^ n1205 ;
  assign n9382 = ( n9377 & n9379 ) | ( n9377 & ~n9381 ) | ( n9379 & ~n9381 ) ;
  assign n9383 = ( n2660 & n5300 ) | ( n2660 & n9382 ) | ( n5300 & n9382 ) ;
  assign n9384 = ( ~n9372 & n9373 ) | ( ~n9372 & n9383 ) | ( n9373 & n9383 ) ;
  assign n9385 = n2329 & ~n3227 ;
  assign n9386 = ( ~x69 & n1112 ) | ( ~x69 & n9090 ) | ( n1112 & n9090 ) ;
  assign n9387 = n1921 & n9386 ;
  assign n9388 = ~n8050 & n9387 ;
  assign n9389 = n9388 ^ n7853 ^ 1'b0 ;
  assign n9390 = n9385 & n9389 ;
  assign n9392 = ~n5835 & n6570 ;
  assign n9391 = n6179 ^ n3597 ^ n1414 ;
  assign n9393 = n9392 ^ n9391 ^ n1198 ;
  assign n9394 = ( n4050 & ~n4842 ) | ( n4050 & n4987 ) | ( ~n4842 & n4987 ) ;
  assign n9399 = n8239 ^ n792 ^ x12 ;
  assign n9395 = n7364 ^ n3186 ^ n2360 ;
  assign n9396 = n7596 ^ n7546 ^ n1335 ;
  assign n9397 = n9396 ^ n5782 ^ n1209 ;
  assign n9398 = ( n5695 & n9395 ) | ( n5695 & n9397 ) | ( n9395 & n9397 ) ;
  assign n9400 = n9399 ^ n9398 ^ n8541 ;
  assign n9401 = ( n2260 & n9394 ) | ( n2260 & n9400 ) | ( n9394 & n9400 ) ;
  assign n9402 = n1838 | n2447 ;
  assign n9403 = ( n5575 & n6267 ) | ( n5575 & n9402 ) | ( n6267 & n9402 ) ;
  assign n9404 = n6185 ^ n3983 ^ n984 ;
  assign n9405 = ( n5803 & n9403 ) | ( n5803 & ~n9404 ) | ( n9403 & ~n9404 ) ;
  assign n9406 = n2484 ^ n1124 ^ 1'b0 ;
  assign n9407 = n4674 ^ n2204 ^ 1'b0 ;
  assign n9408 = ~n7924 & n9407 ;
  assign n9409 = n5980 & n6668 ;
  assign n9410 = n9409 ^ n597 ^ 1'b0 ;
  assign n9418 = n3716 ^ n2875 ^ n417 ;
  assign n9419 = n9418 ^ n3160 ^ n1298 ;
  assign n9411 = n985 | n5471 ;
  assign n9412 = n799 | n9411 ;
  assign n9413 = n5327 ^ n834 ^ n408 ;
  assign n9414 = ( n563 & n3112 ) | ( n563 & n4160 ) | ( n3112 & n4160 ) ;
  assign n9415 = n9414 ^ n7556 ^ n1650 ;
  assign n9416 = ( n6589 & n9413 ) | ( n6589 & n9415 ) | ( n9413 & n9415 ) ;
  assign n9417 = ( n3352 & ~n9412 ) | ( n3352 & n9416 ) | ( ~n9412 & n9416 ) ;
  assign n9420 = n9419 ^ n9417 ^ n5737 ;
  assign n9421 = n9420 ^ n3874 ^ n3605 ;
  assign n9422 = x47 & n3724 ;
  assign n9423 = n9422 ^ n2779 ^ 1'b0 ;
  assign n9424 = ( n1411 & n2741 ) | ( n1411 & n3911 ) | ( n2741 & n3911 ) ;
  assign n9425 = n843 & n5745 ;
  assign n9426 = n9425 ^ n1262 ^ 1'b0 ;
  assign n9427 = ~n9424 & n9426 ;
  assign n9428 = ~n9423 & n9427 ;
  assign n9429 = n7334 ^ n2298 ^ 1'b0 ;
  assign n9430 = ( ~n5114 & n5220 ) | ( ~n5114 & n5886 ) | ( n5220 & n5886 ) ;
  assign n9431 = n9430 ^ n4528 ^ n584 ;
  assign n9432 = ( n422 & n2075 ) | ( n422 & ~n9431 ) | ( n2075 & ~n9431 ) ;
  assign n9433 = ( n472 & n9429 ) | ( n472 & n9432 ) | ( n9429 & n9432 ) ;
  assign n9434 = n8325 ^ n5191 ^ n3228 ;
  assign n9435 = ( n1565 & n2218 ) | ( n1565 & ~n9434 ) | ( n2218 & ~n9434 ) ;
  assign n9436 = ( n2759 & n6392 ) | ( n2759 & ~n9435 ) | ( n6392 & ~n9435 ) ;
  assign n9438 = ( n2381 & n2484 ) | ( n2381 & n9372 ) | ( n2484 & n9372 ) ;
  assign n9437 = ( n260 & n694 ) | ( n260 & ~n3825 ) | ( n694 & ~n3825 ) ;
  assign n9439 = n9438 ^ n9437 ^ n8584 ;
  assign n9440 = n3246 | n3828 ;
  assign n9441 = ( n2866 & n8912 ) | ( n2866 & n9440 ) | ( n8912 & n9440 ) ;
  assign n9442 = ( ~n9436 & n9439 ) | ( ~n9436 & n9441 ) | ( n9439 & n9441 ) ;
  assign n9443 = ( ~x126 & n1377 ) | ( ~x126 & n3498 ) | ( n1377 & n3498 ) ;
  assign n9444 = ( n3440 & n7141 ) | ( n3440 & ~n7196 ) | ( n7141 & ~n7196 ) ;
  assign n9445 = ( ~n3307 & n4728 ) | ( ~n3307 & n5515 ) | ( n4728 & n5515 ) ;
  assign n9446 = n9445 ^ n2486 ^ 1'b0 ;
  assign n9447 = n4953 & n9446 ;
  assign n9448 = ( ~n9443 & n9444 ) | ( ~n9443 & n9447 ) | ( n9444 & n9447 ) ;
  assign n9457 = n2172 & ~n7910 ;
  assign n9458 = n9457 ^ n3095 ^ 1'b0 ;
  assign n9452 = n6845 ^ n5351 ^ n3647 ;
  assign n9450 = n9264 ^ n2080 ^ n1150 ;
  assign n9449 = ( x10 & ~n2935 ) | ( x10 & n3009 ) | ( ~n2935 & n3009 ) ;
  assign n9451 = n9450 ^ n9449 ^ n7307 ;
  assign n9453 = n9452 ^ n9451 ^ 1'b0 ;
  assign n9454 = n6453 ^ n5556 ^ n2583 ;
  assign n9455 = n641 & ~n9454 ;
  assign n9456 = n9453 & n9455 ;
  assign n9459 = n9458 ^ n9456 ^ n5773 ;
  assign n9460 = n6662 ^ n1806 ^ 1'b0 ;
  assign n9461 = n6926 ^ n3676 ^ n2769 ;
  assign n9462 = n9461 ^ n8611 ^ 1'b0 ;
  assign n9463 = n1803 | n5754 ;
  assign n9464 = n2065 & ~n9463 ;
  assign n9465 = n2213 ^ n1591 ^ x16 ;
  assign n9466 = n9465 ^ n5430 ^ n965 ;
  assign n9467 = ( n1700 & n7282 ) | ( n1700 & ~n9466 ) | ( n7282 & ~n9466 ) ;
  assign n9468 = ( ~n4862 & n9464 ) | ( ~n4862 & n9467 ) | ( n9464 & n9467 ) ;
  assign n9469 = ( n319 & n9257 ) | ( n319 & ~n9468 ) | ( n9257 & ~n9468 ) ;
  assign n9470 = ( n4076 & ~n9462 ) | ( n4076 & n9469 ) | ( ~n9462 & n9469 ) ;
  assign n9471 = n6517 ^ n1767 ^ n1677 ;
  assign n9481 = ( ~n2460 & n2987 ) | ( ~n2460 & n4004 ) | ( n2987 & n4004 ) ;
  assign n9482 = n9481 ^ n1490 ^ 1'b0 ;
  assign n9479 = n1397 ^ n439 ^ 1'b0 ;
  assign n9480 = n9479 ^ n8947 ^ n6490 ;
  assign n9483 = n9482 ^ n9480 ^ n475 ;
  assign n9484 = n9483 ^ n1738 ^ 1'b0 ;
  assign n9472 = ~n3521 & n7301 ;
  assign n9473 = n3500 & n9472 ;
  assign n9474 = ( ~x6 & n5074 ) | ( ~x6 & n9473 ) | ( n5074 & n9473 ) ;
  assign n9475 = ( n300 & n2980 ) | ( n300 & ~n4115 ) | ( n2980 & ~n4115 ) ;
  assign n9476 = n5724 & ~n9475 ;
  assign n9477 = ( n651 & n9474 ) | ( n651 & n9476 ) | ( n9474 & n9476 ) ;
  assign n9478 = ( n2327 & ~n4832 ) | ( n2327 & n9477 ) | ( ~n4832 & n9477 ) ;
  assign n9485 = n9484 ^ n9478 ^ n2025 ;
  assign n9486 = n7156 ^ n4780 ^ n3813 ;
  assign n9487 = n9486 ^ n8369 ^ n3123 ;
  assign n9488 = ( ~n2093 & n7699 ) | ( ~n2093 & n9487 ) | ( n7699 & n9487 ) ;
  assign n9489 = ( n1609 & n9485 ) | ( n1609 & n9488 ) | ( n9485 & n9488 ) ;
  assign n9490 = ( n5974 & ~n9471 ) | ( n5974 & n9489 ) | ( ~n9471 & n9489 ) ;
  assign n9491 = n996 ^ n907 ^ n241 ;
  assign n9492 = n1917 | n9491 ;
  assign n9499 = n3576 ^ n2083 ^ n339 ;
  assign n9500 = n9499 ^ n7966 ^ x96 ;
  assign n9501 = ( n3463 & n6951 ) | ( n3463 & n9500 ) | ( n6951 & n9500 ) ;
  assign n9502 = n9501 ^ n7435 ^ n2232 ;
  assign n9493 = ( n2039 & n2564 ) | ( n2039 & n4482 ) | ( n2564 & n4482 ) ;
  assign n9494 = ( n2673 & n4660 ) | ( n2673 & n9493 ) | ( n4660 & n9493 ) ;
  assign n9495 = n9494 ^ n3365 ^ n1785 ;
  assign n9496 = ( n805 & n3129 ) | ( n805 & ~n9495 ) | ( n3129 & ~n9495 ) ;
  assign n9497 = ~n6884 & n9496 ;
  assign n9498 = ( n721 & n5590 ) | ( n721 & n9497 ) | ( n5590 & n9497 ) ;
  assign n9503 = n9502 ^ n9498 ^ n8619 ;
  assign n9504 = ~n351 & n6313 ;
  assign n9506 = ( n1372 & n4228 ) | ( n1372 & n6832 ) | ( n4228 & n6832 ) ;
  assign n9505 = ( n1813 & ~n2028 ) | ( n1813 & n9319 ) | ( ~n2028 & n9319 ) ;
  assign n9507 = n9506 ^ n9505 ^ n5206 ;
  assign n9508 = n3059 & ~n9507 ;
  assign n9509 = ( n7382 & ~n9504 ) | ( n7382 & n9508 ) | ( ~n9504 & n9508 ) ;
  assign n9510 = ( n222 & n2019 ) | ( n222 & n3990 ) | ( n2019 & n3990 ) ;
  assign n9511 = n2633 & n9510 ;
  assign n9512 = ~n1655 & n9511 ;
  assign n9513 = ( ~n704 & n949 ) | ( ~n704 & n9512 ) | ( n949 & n9512 ) ;
  assign n9514 = ( x55 & n3459 ) | ( x55 & n9513 ) | ( n3459 & n9513 ) ;
  assign n9515 = ( n7729 & ~n7981 ) | ( n7729 & n9514 ) | ( ~n7981 & n9514 ) ;
  assign n9521 = n2076 ^ n264 ^ 1'b0 ;
  assign n9522 = ~n584 & n9521 ;
  assign n9519 = n1860 & n9513 ;
  assign n9520 = n9519 ^ n6528 ^ x9 ;
  assign n9523 = n9522 ^ n9520 ^ n6694 ;
  assign n9516 = ~n415 & n504 ;
  assign n9517 = ~n1247 & n9516 ;
  assign n9518 = n6434 | n9517 ;
  assign n9524 = n9523 ^ n9518 ^ n729 ;
  assign n9525 = n609 & ~n2334 ;
  assign n9526 = n9525 ^ n2345 ^ 1'b0 ;
  assign n9527 = ( n7181 & n9524 ) | ( n7181 & ~n9526 ) | ( n9524 & ~n9526 ) ;
  assign n9528 = ( ~n609 & n2379 ) | ( ~n609 & n5410 ) | ( n2379 & n5410 ) ;
  assign n9529 = n9528 ^ n420 ^ n259 ;
  assign n9530 = ( n835 & ~n6520 ) | ( n835 & n9438 ) | ( ~n6520 & n9438 ) ;
  assign n9531 = ( x22 & n9529 ) | ( x22 & ~n9530 ) | ( n9529 & ~n9530 ) ;
  assign n9540 = ~n2173 & n8677 ;
  assign n9539 = ~n1347 & n2375 ;
  assign n9541 = n9540 ^ n9539 ^ 1'b0 ;
  assign n9542 = ( ~n790 & n2037 ) | ( ~n790 & n9541 ) | ( n2037 & n9541 ) ;
  assign n9537 = n7406 ^ n4009 ^ 1'b0 ;
  assign n9538 = n6629 | n9537 ;
  assign n9543 = n9542 ^ n9538 ^ 1'b0 ;
  assign n9532 = n6233 ^ n5101 ^ n1547 ;
  assign n9533 = n4618 ^ n1951 ^ n1462 ;
  assign n9534 = n9533 ^ n2173 ^ n1330 ;
  assign n9535 = n9532 | n9534 ;
  assign n9536 = n2954 & n9535 ;
  assign n9544 = n9543 ^ n9536 ^ 1'b0 ;
  assign n9549 = ( ~n546 & n734 ) | ( ~n546 & n2007 ) | ( n734 & n2007 ) ;
  assign n9550 = n7009 ^ n6233 ^ n735 ;
  assign n9551 = ( n2805 & ~n9549 ) | ( n2805 & n9550 ) | ( ~n9549 & n9550 ) ;
  assign n9552 = ( ~n532 & n2443 ) | ( ~n532 & n9551 ) | ( n2443 & n9551 ) ;
  assign n9545 = n3907 ^ n706 ^ n399 ;
  assign n9546 = n9545 ^ x45 ^ 1'b0 ;
  assign n9547 = n1447 | n9546 ;
  assign n9548 = n9547 ^ n3834 ^ n1314 ;
  assign n9553 = n9552 ^ n9548 ^ n5684 ;
  assign n9563 = ( n1052 & n5791 ) | ( n1052 & n6284 ) | ( n5791 & n6284 ) ;
  assign n9564 = ( n6911 & n7694 ) | ( n6911 & n9563 ) | ( n7694 & n9563 ) ;
  assign n9559 = n6544 ^ n3882 ^ n364 ;
  assign n9560 = n9559 ^ n5488 ^ 1'b0 ;
  assign n9561 = ~n2899 & n9560 ;
  assign n9557 = ( n1000 & n1052 ) | ( n1000 & ~n1511 ) | ( n1052 & ~n1511 ) ;
  assign n9555 = n8747 ^ n4940 ^ n4349 ;
  assign n9556 = ( ~n6217 & n6586 ) | ( ~n6217 & n9555 ) | ( n6586 & n9555 ) ;
  assign n9554 = n2152 ^ n1848 ^ n1841 ;
  assign n9558 = n9557 ^ n9556 ^ n9554 ;
  assign n9562 = n9561 ^ n9558 ^ n6019 ;
  assign n9565 = n9564 ^ n9562 ^ 1'b0 ;
  assign n9566 = n9553 & ~n9565 ;
  assign n9573 = ( ~n295 & n451 ) | ( ~n295 & n1886 ) | ( n451 & n1886 ) ;
  assign n9569 = ( ~n1226 & n2520 ) | ( ~n1226 & n5607 ) | ( n2520 & n5607 ) ;
  assign n9570 = ( n2496 & n2927 ) | ( n2496 & ~n9569 ) | ( n2927 & ~n9569 ) ;
  assign n9567 = ( n551 & n1259 ) | ( n551 & ~n5514 ) | ( n1259 & ~n5514 ) ;
  assign n9568 = n9567 ^ n1008 ^ 1'b0 ;
  assign n9571 = n9570 ^ n9568 ^ n7580 ;
  assign n9572 = n8305 & n9571 ;
  assign n9574 = n9573 ^ n9572 ^ n1751 ;
  assign n9575 = ( ~n1361 & n1373 ) | ( ~n1361 & n2259 ) | ( n1373 & n2259 ) ;
  assign n9578 = ( n4770 & ~n5216 ) | ( n4770 & n9474 ) | ( ~n5216 & n9474 ) ;
  assign n9576 = n2432 & ~n8785 ;
  assign n9577 = ~n7225 & n9576 ;
  assign n9579 = n9578 ^ n9577 ^ n8584 ;
  assign n9586 = n3833 & ~n7479 ;
  assign n9587 = ~n7532 & n9586 ;
  assign n9588 = n9587 ^ n4325 ^ n3195 ;
  assign n9583 = n1833 ^ n249 ^ 1'b0 ;
  assign n9581 = n3107 & n3433 ;
  assign n9582 = n5293 & n9581 ;
  assign n9584 = n9583 ^ n9582 ^ 1'b0 ;
  assign n9580 = x123 & n3547 ;
  assign n9585 = n9584 ^ n9580 ^ 1'b0 ;
  assign n9589 = n9588 ^ n9585 ^ n1100 ;
  assign n9590 = ( ~n484 & n1598 ) | ( ~n484 & n4160 ) | ( n1598 & n4160 ) ;
  assign n9591 = ( ~n1533 & n3386 ) | ( ~n1533 & n9590 ) | ( n3386 & n9590 ) ;
  assign n9592 = n9591 ^ n7607 ^ 1'b0 ;
  assign n9593 = n5834 & ~n9592 ;
  assign n9594 = ( n1998 & ~n4836 ) | ( n1998 & n9593 ) | ( ~n4836 & n9593 ) ;
  assign n9595 = n7465 ^ n3056 ^ n1985 ;
  assign n9596 = n9595 ^ n5807 ^ n418 ;
  assign n9597 = n9596 ^ n4319 ^ n1863 ;
  assign n9598 = ( ~n945 & n4108 ) | ( ~n945 & n4620 ) | ( n4108 & n4620 ) ;
  assign n9599 = n6210 & n9598 ;
  assign n9600 = n9599 ^ n1466 ^ 1'b0 ;
  assign n9601 = n2345 | n3532 ;
  assign n9602 = n9601 ^ x13 ^ 1'b0 ;
  assign n9603 = ( ~n3415 & n3559 ) | ( ~n3415 & n9602 ) | ( n3559 & n9602 ) ;
  assign n9604 = ( n1781 & ~n8082 ) | ( n1781 & n9222 ) | ( ~n8082 & n9222 ) ;
  assign n9605 = ~n4491 & n9604 ;
  assign n9606 = n9603 & n9605 ;
  assign n9607 = x88 & n392 ;
  assign n9608 = ( n824 & n4640 ) | ( n824 & ~n9607 ) | ( n4640 & ~n9607 ) ;
  assign n9609 = ( n1444 & n1482 ) | ( n1444 & ~n2304 ) | ( n1482 & ~n2304 ) ;
  assign n9610 = n9609 ^ n4392 ^ n3815 ;
  assign n9611 = n9610 ^ n3420 ^ 1'b0 ;
  assign n9612 = n3543 ^ n2146 ^ 1'b0 ;
  assign n9613 = n9612 ^ n8071 ^ n1802 ;
  assign n9614 = ( n9608 & n9611 ) | ( n9608 & ~n9613 ) | ( n9611 & ~n9613 ) ;
  assign n9615 = n9614 ^ n566 ^ x50 ;
  assign n9616 = n5484 ^ n4718 ^ n4444 ;
  assign n9617 = n3853 ^ x98 ^ 1'b0 ;
  assign n9618 = ( n2377 & ~n5942 ) | ( n2377 & n9617 ) | ( ~n5942 & n9617 ) ;
  assign n9619 = ( n436 & n3528 ) | ( n436 & n8856 ) | ( n3528 & n8856 ) ;
  assign n9620 = ( n8656 & n9618 ) | ( n8656 & ~n9619 ) | ( n9618 & ~n9619 ) ;
  assign n9621 = ( n1086 & ~n9616 ) | ( n1086 & n9620 ) | ( ~n9616 & n9620 ) ;
  assign n9622 = n9170 ^ n3654 ^ n2961 ;
  assign n9623 = ( ~n4701 & n8753 ) | ( ~n4701 & n9622 ) | ( n8753 & n9622 ) ;
  assign n9624 = ( n2113 & n5947 ) | ( n2113 & n9623 ) | ( n5947 & n9623 ) ;
  assign n9633 = ( ~n280 & n3776 ) | ( ~n280 & n8562 ) | ( n3776 & n8562 ) ;
  assign n9630 = n9365 ^ n2365 ^ 1'b0 ;
  assign n9631 = n9630 ^ n1671 ^ n817 ;
  assign n9627 = n1747 | n7263 ;
  assign n9628 = n9627 ^ n4954 ^ 1'b0 ;
  assign n9629 = n9628 ^ n6336 ^ n358 ;
  assign n9632 = n9631 ^ n9629 ^ n8580 ;
  assign n9634 = n9633 ^ n9632 ^ n3630 ;
  assign n9625 = n3642 ^ n2555 ^ n2375 ;
  assign n9626 = n5474 & n9625 ;
  assign n9635 = n9634 ^ n9626 ^ 1'b0 ;
  assign n9636 = n997 | n1848 ;
  assign n9637 = n9636 ^ n2250 ^ 1'b0 ;
  assign n9638 = n3173 | n9637 ;
  assign n9639 = n3037 | n9638 ;
  assign n9640 = n4085 & n7517 ;
  assign n9641 = ~n1889 & n9640 ;
  assign n9642 = ( n901 & ~n1053 ) | ( n901 & n7620 ) | ( ~n1053 & n7620 ) ;
  assign n9643 = ( n913 & n2168 ) | ( n913 & ~n9642 ) | ( n2168 & ~n9642 ) ;
  assign n9644 = n9643 ^ n5439 ^ 1'b0 ;
  assign n9645 = n6541 & ~n9644 ;
  assign n9646 = ( ~n1833 & n6895 ) | ( ~n1833 & n9645 ) | ( n6895 & n9645 ) ;
  assign n9647 = ( n4680 & n9641 ) | ( n4680 & ~n9646 ) | ( n9641 & ~n9646 ) ;
  assign n9648 = n7189 & n9647 ;
  assign n9649 = n276 & n9648 ;
  assign n9652 = n5892 ^ n5021 ^ 1'b0 ;
  assign n9650 = n4414 ^ n3773 ^ n1197 ;
  assign n9651 = n9650 ^ n4482 ^ n3657 ;
  assign n9653 = n9652 ^ n9651 ^ 1'b0 ;
  assign n9658 = n1510 ^ n1091 ^ n990 ;
  assign n9654 = n3685 & ~n9465 ;
  assign n9655 = n3139 & ~n3397 ;
  assign n9656 = n9655 ^ n4717 ^ 1'b0 ;
  assign n9657 = ( n9643 & n9654 ) | ( n9643 & ~n9656 ) | ( n9654 & ~n9656 ) ;
  assign n9659 = n9658 ^ n9657 ^ n2768 ;
  assign n9665 = n8489 ^ n3758 ^ 1'b0 ;
  assign n9660 = n5137 ^ n2622 ^ n2520 ;
  assign n9661 = ( ~n206 & n467 ) | ( ~n206 & n9660 ) | ( n467 & n9660 ) ;
  assign n9662 = ( n874 & ~n5155 ) | ( n874 & n9661 ) | ( ~n5155 & n9661 ) ;
  assign n9663 = ( n4665 & n5144 ) | ( n4665 & ~n6613 ) | ( n5144 & ~n6613 ) ;
  assign n9664 = n9662 & ~n9663 ;
  assign n9666 = n9665 ^ n9664 ^ 1'b0 ;
  assign n9667 = ( n511 & n2042 ) | ( n511 & n3550 ) | ( n2042 & n3550 ) ;
  assign n9668 = n9667 ^ n8806 ^ n7403 ;
  assign n9669 = ( ~n446 & n5871 ) | ( ~n446 & n9235 ) | ( n5871 & n9235 ) ;
  assign n9671 = n6863 ^ n1292 ^ n690 ;
  assign n9670 = ( n4852 & ~n7077 ) | ( n4852 & n7906 ) | ( ~n7077 & n7906 ) ;
  assign n9672 = n9671 ^ n9670 ^ n9585 ;
  assign n9673 = n4440 ^ n3468 ^ n1474 ;
  assign n9674 = ( n5092 & ~n5578 ) | ( n5092 & n9673 ) | ( ~n5578 & n9673 ) ;
  assign n9675 = n9674 ^ n6577 ^ n5545 ;
  assign n9676 = n1533 | n9675 ;
  assign n9677 = n9676 ^ n2153 ^ 1'b0 ;
  assign n9678 = ( n2252 & ~n4410 ) | ( n2252 & n7773 ) | ( ~n4410 & n7773 ) ;
  assign n9687 = ( n816 & n2699 ) | ( n816 & n7004 ) | ( n2699 & n7004 ) ;
  assign n9688 = ( n2379 & n5701 ) | ( n2379 & ~n9687 ) | ( n5701 & ~n9687 ) ;
  assign n9685 = n3302 ^ n336 ^ x12 ;
  assign n9683 = ( ~n287 & n611 ) | ( ~n287 & n4555 ) | ( n611 & n4555 ) ;
  assign n9682 = ( n2330 & ~n4088 ) | ( n2330 & n7168 ) | ( ~n4088 & n7168 ) ;
  assign n9679 = n4890 ^ n4120 ^ n3197 ;
  assign n9680 = n4005 & ~n9679 ;
  assign n9681 = n9680 ^ n3078 ^ 1'b0 ;
  assign n9684 = n9683 ^ n9682 ^ n9681 ;
  assign n9686 = n9685 ^ n9684 ^ n5554 ;
  assign n9689 = n9688 ^ n9686 ^ n8030 ;
  assign n9690 = n9689 ^ n3564 ^ 1'b0 ;
  assign n9691 = n3002 & ~n9690 ;
  assign n9692 = n1085 ^ n310 ^ 1'b0 ;
  assign n9693 = n283 & n9692 ;
  assign n9694 = ( n4713 & n5522 ) | ( n4713 & n9693 ) | ( n5522 & n9693 ) ;
  assign n9695 = n9694 ^ n1988 ^ n374 ;
  assign n9696 = ( n486 & ~n5095 ) | ( n486 & n9127 ) | ( ~n5095 & n9127 ) ;
  assign n9697 = ( n1506 & n9695 ) | ( n1506 & ~n9696 ) | ( n9695 & ~n9696 ) ;
  assign n9698 = n9697 ^ n7123 ^ n138 ;
  assign n9699 = ( n3593 & ~n5667 ) | ( n3593 & n8272 ) | ( ~n5667 & n8272 ) ;
  assign n9700 = ( n1335 & n9520 ) | ( n1335 & ~n9699 ) | ( n9520 & ~n9699 ) ;
  assign n9701 = ( n4683 & n8664 ) | ( n4683 & ~n9700 ) | ( n8664 & ~n9700 ) ;
  assign n9702 = ( n6065 & n9698 ) | ( n6065 & n9701 ) | ( n9698 & n9701 ) ;
  assign n9703 = ( n366 & ~n755 ) | ( n366 & n6565 ) | ( ~n755 & n6565 ) ;
  assign n9704 = n4617 ^ n4449 ^ n2901 ;
  assign n9706 = ( n1262 & n2419 ) | ( n1262 & ~n4429 ) | ( n2419 & ~n4429 ) ;
  assign n9707 = ( n1135 & ~n5331 ) | ( n1135 & n9706 ) | ( ~n5331 & n9706 ) ;
  assign n9705 = n9096 ^ n5903 ^ n4265 ;
  assign n9708 = n9707 ^ n9705 ^ n2148 ;
  assign n9709 = n4423 & n4959 ;
  assign n9710 = n3505 | n3873 ;
  assign n9711 = n9709 & ~n9710 ;
  assign n9712 = n6613 ^ n2378 ^ n1496 ;
  assign n9713 = n9712 ^ n6537 ^ n1252 ;
  assign n9714 = ( n4303 & n5618 ) | ( n4303 & n9713 ) | ( n5618 & n9713 ) ;
  assign n9715 = ( n6428 & n7080 ) | ( n6428 & ~n9714 ) | ( n7080 & ~n9714 ) ;
  assign n9717 = ( n878 & n4408 ) | ( n878 & n6665 ) | ( n4408 & n6665 ) ;
  assign n9716 = n2455 | n4328 ;
  assign n9718 = n9717 ^ n9716 ^ n4843 ;
  assign n9719 = ( ~n3357 & n3500 ) | ( ~n3357 & n4374 ) | ( n3500 & n4374 ) ;
  assign n9720 = ( n1874 & n3214 ) | ( n1874 & n9719 ) | ( n3214 & n9719 ) ;
  assign n9721 = ( n556 & n5526 ) | ( n556 & n7027 ) | ( n5526 & n7027 ) ;
  assign n9722 = ( n591 & n3813 ) | ( n591 & n5012 ) | ( n3813 & n5012 ) ;
  assign n9723 = n9722 ^ n8150 ^ n2314 ;
  assign n9724 = ( ~n8933 & n9721 ) | ( ~n8933 & n9723 ) | ( n9721 & n9723 ) ;
  assign n9725 = ( n7616 & n9720 ) | ( n7616 & n9724 ) | ( n9720 & n9724 ) ;
  assign n9726 = ( n4905 & n9718 ) | ( n4905 & n9725 ) | ( n9718 & n9725 ) ;
  assign n9727 = ( n9711 & ~n9715 ) | ( n9711 & n9726 ) | ( ~n9715 & n9726 ) ;
  assign n9728 = ( n572 & n9708 ) | ( n572 & n9727 ) | ( n9708 & n9727 ) ;
  assign n9729 = ( n1578 & n5371 ) | ( n1578 & ~n8330 ) | ( n5371 & ~n8330 ) ;
  assign n9731 = ( x27 & ~n529 ) | ( x27 & n1661 ) | ( ~n529 & n1661 ) ;
  assign n9730 = n2246 ^ n2125 ^ n2057 ;
  assign n9732 = n9731 ^ n9730 ^ n9259 ;
  assign n9733 = ( ~n5972 & n8801 ) | ( ~n5972 & n9732 ) | ( n8801 & n9732 ) ;
  assign n9735 = n398 & ~n541 ;
  assign n9736 = ( n1276 & n7799 ) | ( n1276 & n9735 ) | ( n7799 & n9735 ) ;
  assign n9737 = n9736 ^ n4188 ^ n157 ;
  assign n9734 = n5564 | n8074 ;
  assign n9738 = n9737 ^ n9734 ^ 1'b0 ;
  assign n9739 = ( n230 & ~n9733 ) | ( n230 & n9738 ) | ( ~n9733 & n9738 ) ;
  assign n9740 = ( n1726 & ~n4228 ) | ( n1726 & n5214 ) | ( ~n4228 & n5214 ) ;
  assign n9741 = n9740 ^ n1181 ^ n880 ;
  assign n9742 = n9741 ^ n3526 ^ n193 ;
  assign n9743 = ( ~n8899 & n9739 ) | ( ~n8899 & n9742 ) | ( n9739 & n9742 ) ;
  assign n9744 = ( n290 & n2063 ) | ( n290 & ~n4444 ) | ( n2063 & ~n4444 ) ;
  assign n9745 = ( n213 & n733 ) | ( n213 & ~n1233 ) | ( n733 & ~n1233 ) ;
  assign n9749 = n2426 | n8119 ;
  assign n9746 = n592 & n861 ;
  assign n9747 = n9746 ^ n2912 ^ 1'b0 ;
  assign n9748 = ~n2877 & n9747 ;
  assign n9750 = n9749 ^ n9748 ^ 1'b0 ;
  assign n9751 = n9745 & ~n9750 ;
  assign n9752 = ( n1998 & n3290 ) | ( n1998 & n3904 ) | ( n3290 & n3904 ) ;
  assign n9753 = n9436 ^ n4122 ^ 1'b0 ;
  assign n9754 = ( ~n2059 & n9274 ) | ( ~n2059 & n9753 ) | ( n9274 & n9753 ) ;
  assign n9755 = ~n1033 & n9754 ;
  assign n9756 = ~n9752 & n9755 ;
  assign n9757 = ( ~n3403 & n4759 ) | ( ~n3403 & n6601 ) | ( n4759 & n6601 ) ;
  assign n9758 = ( n4150 & ~n4860 ) | ( n4150 & n9757 ) | ( ~n4860 & n9757 ) ;
  assign n9759 = ( n326 & n5249 ) | ( n326 & n7506 ) | ( n5249 & n7506 ) ;
  assign n9760 = ( ~n510 & n2601 ) | ( ~n510 & n9759 ) | ( n2601 & n9759 ) ;
  assign n9761 = n5771 ^ n3173 ^ n1881 ;
  assign n9762 = n9761 ^ n5318 ^ n4760 ;
  assign n9763 = ( ~n3047 & n9760 ) | ( ~n3047 & n9762 ) | ( n9760 & n9762 ) ;
  assign n9764 = n9354 ^ n1785 ^ 1'b0 ;
  assign n9765 = n855 & ~n7201 ;
  assign n9766 = ~n3058 & n9765 ;
  assign n9767 = ( ~n1192 & n6415 ) | ( ~n1192 & n6454 ) | ( n6415 & n6454 ) ;
  assign n9768 = n7858 ^ n5088 ^ 1'b0 ;
  assign n9769 = n9212 & n9768 ;
  assign n9770 = ( n9766 & ~n9767 ) | ( n9766 & n9769 ) | ( ~n9767 & n9769 ) ;
  assign n9771 = ( ~n4765 & n7939 ) | ( ~n4765 & n9770 ) | ( n7939 & n9770 ) ;
  assign n9777 = ( n1755 & ~n2758 ) | ( n1755 & n7663 ) | ( ~n2758 & n7663 ) ;
  assign n9772 = ( n297 & ~n460 ) | ( n297 & n960 ) | ( ~n460 & n960 ) ;
  assign n9773 = n1386 | n2604 ;
  assign n9774 = n2065 & ~n9773 ;
  assign n9775 = ( ~n324 & n3131 ) | ( ~n324 & n9774 ) | ( n3131 & n9774 ) ;
  assign n9776 = ( n2880 & n9772 ) | ( n2880 & n9775 ) | ( n9772 & n9775 ) ;
  assign n9778 = n9777 ^ n9776 ^ 1'b0 ;
  assign n9779 = n4062 & ~n9778 ;
  assign n9780 = n2736 ^ n1037 ^ n159 ;
  assign n9781 = ( n390 & ~n824 ) | ( n390 & n9780 ) | ( ~n824 & n9780 ) ;
  assign n9782 = ( ~n6044 & n8450 ) | ( ~n6044 & n8681 ) | ( n8450 & n8681 ) ;
  assign n9783 = ( n636 & n5716 ) | ( n636 & ~n5942 ) | ( n5716 & ~n5942 ) ;
  assign n9784 = n6555 ^ n2462 ^ n706 ;
  assign n9785 = n9784 ^ n7558 ^ n3471 ;
  assign n9786 = n9785 ^ n2279 ^ n2038 ;
  assign n9787 = ( ~n774 & n3829 ) | ( ~n774 & n4275 ) | ( n3829 & n4275 ) ;
  assign n9788 = ( ~n5619 & n9786 ) | ( ~n5619 & n9787 ) | ( n9786 & n9787 ) ;
  assign n9795 = n7282 ^ n1715 ^ n568 ;
  assign n9792 = ~n1275 & n8576 ;
  assign n9793 = ~n7400 & n9792 ;
  assign n9794 = ( n1259 & n1967 ) | ( n1259 & n9793 ) | ( n1967 & n9793 ) ;
  assign n9790 = n5678 ^ n235 ^ 1'b0 ;
  assign n9789 = n5434 ^ n5284 ^ n2215 ;
  assign n9791 = n9790 ^ n9789 ^ n1017 ;
  assign n9796 = n9795 ^ n9794 ^ n9791 ;
  assign n9797 = ( ~n4732 & n5597 ) | ( ~n4732 & n5886 ) | ( n5597 & n5886 ) ;
  assign n9798 = n9797 ^ n3337 ^ n2265 ;
  assign n9799 = ( n393 & n1998 ) | ( n393 & n8206 ) | ( n1998 & n8206 ) ;
  assign n9800 = n9799 ^ n7237 ^ n4720 ;
  assign n9805 = n5230 ^ n3665 ^ n1782 ;
  assign n9806 = n9805 ^ n4257 ^ n3474 ;
  assign n9801 = ( n3067 & ~n5918 ) | ( n3067 & n8103 ) | ( ~n5918 & n8103 ) ;
  assign n9802 = ( n6913 & n7716 ) | ( n6913 & n9801 ) | ( n7716 & n9801 ) ;
  assign n9803 = n9802 ^ n4710 ^ 1'b0 ;
  assign n9804 = ~n7257 & n9803 ;
  assign n9807 = n9806 ^ n9804 ^ n736 ;
  assign n9808 = n5131 ^ n1811 ^ n166 ;
  assign n9809 = n9808 ^ n6896 ^ 1'b0 ;
  assign n9810 = ~n6118 & n9809 ;
  assign n9811 = ( n206 & ~n4608 ) | ( n206 & n5074 ) | ( ~n4608 & n5074 ) ;
  assign n9812 = n1581 & n9811 ;
  assign n9813 = ~n9810 & n9812 ;
  assign n9814 = n9813 ^ n9397 ^ n6828 ;
  assign n9815 = n357 & n1837 ;
  assign n9816 = ~n153 & n9815 ;
  assign n9817 = n4083 ^ n3834 ^ n2947 ;
  assign n9818 = ( n8209 & ~n9816 ) | ( n8209 & n9817 ) | ( ~n9816 & n9817 ) ;
  assign n9820 = n5282 ^ n1926 ^ n1143 ;
  assign n9819 = n7471 ^ n7302 ^ n7225 ;
  assign n9821 = n9820 ^ n9819 ^ n3644 ;
  assign n9822 = ( n9814 & n9818 ) | ( n9814 & n9821 ) | ( n9818 & n9821 ) ;
  assign n9823 = ( n409 & n1035 ) | ( n409 & n5169 ) | ( n1035 & n5169 ) ;
  assign n9833 = n3992 & ~n8872 ;
  assign n9831 = n2527 ^ n812 ^ 1'b0 ;
  assign n9832 = x57 & n9831 ;
  assign n9829 = n3471 ^ n1131 ^ n767 ;
  assign n9830 = n7498 & ~n9829 ;
  assign n9834 = n9833 ^ n9832 ^ n9830 ;
  assign n9827 = n7866 ^ n6764 ^ 1'b0 ;
  assign n9824 = n2849 & n9423 ;
  assign n9825 = n4020 & n9824 ;
  assign n9826 = n7206 & ~n9825 ;
  assign n9828 = n9827 ^ n9826 ^ 1'b0 ;
  assign n9835 = n9834 ^ n9828 ^ n3735 ;
  assign n9836 = n5784 ^ n5351 ^ n1198 ;
  assign n9837 = n9836 ^ n4684 ^ n336 ;
  assign n9838 = n9837 ^ n3187 ^ n1131 ;
  assign n9839 = n9838 ^ n1293 ^ n499 ;
  assign n9840 = ( n1788 & n5825 ) | ( n1788 & n7695 ) | ( n5825 & n7695 ) ;
  assign n9841 = ( n2933 & n6712 ) | ( n2933 & n9840 ) | ( n6712 & n9840 ) ;
  assign n9842 = n9167 ^ n3234 ^ n1992 ;
  assign n9843 = ( n3843 & ~n4470 ) | ( n3843 & n9842 ) | ( ~n4470 & n9842 ) ;
  assign n9844 = n3338 ^ n1161 ^ 1'b0 ;
  assign n9845 = n9843 | n9844 ;
  assign n9846 = n5567 ^ n3074 ^ n2923 ;
  assign n9847 = n9846 ^ n5416 ^ n3127 ;
  assign n9848 = ( n811 & n2326 ) | ( n811 & n9847 ) | ( n2326 & n9847 ) ;
  assign n9849 = ( n361 & n4514 ) | ( n361 & n9848 ) | ( n4514 & n9848 ) ;
  assign n9850 = n9849 ^ n6338 ^ 1'b0 ;
  assign n9851 = ( n6575 & n9845 ) | ( n6575 & ~n9850 ) | ( n9845 & ~n9850 ) ;
  assign n9854 = n5064 ^ n4452 ^ 1'b0 ;
  assign n9852 = ( n718 & n2742 ) | ( n718 & ~n7999 ) | ( n2742 & ~n7999 ) ;
  assign n9853 = n9852 ^ n4884 ^ 1'b0 ;
  assign n9855 = n9854 ^ n9853 ^ n1289 ;
  assign n9860 = n4861 ^ n2652 ^ n1403 ;
  assign n9861 = ( n1957 & n3139 ) | ( n1957 & ~n9860 ) | ( n3139 & ~n9860 ) ;
  assign n9862 = ~n4457 & n7873 ;
  assign n9863 = ~n7434 & n9862 ;
  assign n9864 = ( n8942 & n9861 ) | ( n8942 & ~n9863 ) | ( n9861 & ~n9863 ) ;
  assign n9856 = n5817 ^ n1256 ^ 1'b0 ;
  assign n9857 = n1387 & ~n9856 ;
  assign n9858 = n9857 ^ n1895 ^ n809 ;
  assign n9859 = ~n731 & n9858 ;
  assign n9865 = n9864 ^ n9859 ^ n4795 ;
  assign n9866 = ( ~n960 & n5607 ) | ( ~n960 & n7309 ) | ( n5607 & n7309 ) ;
  assign n9867 = ( n524 & ~n3100 ) | ( n524 & n4392 ) | ( ~n3100 & n4392 ) ;
  assign n9868 = ( n2104 & n6182 ) | ( n2104 & n9867 ) | ( n6182 & n9867 ) ;
  assign n9869 = ( ~n481 & n581 ) | ( ~n481 & n5398 ) | ( n581 & n5398 ) ;
  assign n9870 = ( n883 & ~n1114 ) | ( n883 & n9869 ) | ( ~n1114 & n9869 ) ;
  assign n9871 = n9870 ^ n4633 ^ 1'b0 ;
  assign n9872 = ( ~n1608 & n5115 ) | ( ~n1608 & n9871 ) | ( n5115 & n9871 ) ;
  assign n9873 = ( n2490 & n3946 ) | ( n2490 & n4511 ) | ( n3946 & n4511 ) ;
  assign n9874 = n9873 ^ n3892 ^ n968 ;
  assign n9875 = n8028 ^ n2944 ^ 1'b0 ;
  assign n9876 = n8856 | n9875 ;
  assign n9877 = n7459 & ~n9876 ;
  assign n9878 = n9877 ^ n6957 ^ n3494 ;
  assign n9879 = n9874 | n9878 ;
  assign n9880 = n9872 | n9879 ;
  assign n9881 = n5768 ^ n4285 ^ n2446 ;
  assign n9884 = n4161 ^ n1774 ^ 1'b0 ;
  assign n9882 = n5522 ^ n4741 ^ n3285 ;
  assign n9883 = ( n196 & n7379 ) | ( n196 & ~n9882 ) | ( n7379 & ~n9882 ) ;
  assign n9885 = n9884 ^ n9883 ^ 1'b0 ;
  assign n9886 = n9885 ^ n4868 ^ 1'b0 ;
  assign n9887 = ( n3666 & n9881 ) | ( n3666 & n9886 ) | ( n9881 & n9886 ) ;
  assign n9889 = ( n6609 & n7346 ) | ( n6609 & ~n9706 ) | ( n7346 & ~n9706 ) ;
  assign n9888 = ( n4385 & n4863 ) | ( n4385 & n6509 ) | ( n4863 & n6509 ) ;
  assign n9890 = n9889 ^ n9888 ^ n1450 ;
  assign n9892 = ( n2648 & ~n6318 ) | ( n2648 & n6821 ) | ( ~n6318 & n6821 ) ;
  assign n9893 = ( n1597 & n7730 ) | ( n1597 & ~n9892 ) | ( n7730 & ~n9892 ) ;
  assign n9894 = ~n6808 & n9893 ;
  assign n9895 = ( n2664 & n5637 ) | ( n2664 & ~n9894 ) | ( n5637 & ~n9894 ) ;
  assign n9891 = n5999 ^ n3751 ^ n2876 ;
  assign n9896 = n9895 ^ n9891 ^ n494 ;
  assign n9897 = ( n4189 & ~n7512 ) | ( n4189 & n8742 ) | ( ~n7512 & n8742 ) ;
  assign n9898 = ( ~n7616 & n8582 ) | ( ~n7616 & n9897 ) | ( n8582 & n9897 ) ;
  assign n9906 = n7989 ^ n3861 ^ n2470 ;
  assign n9905 = n9568 ^ n8947 ^ n2828 ;
  assign n9903 = ( ~n964 & n5142 ) | ( ~n964 & n5294 ) | ( n5142 & n5294 ) ;
  assign n9901 = n4759 ^ n4118 ^ n1629 ;
  assign n9899 = n7799 ^ n2963 ^ n2881 ;
  assign n9900 = ( n1556 & ~n6122 ) | ( n1556 & n9899 ) | ( ~n6122 & n9899 ) ;
  assign n9902 = n9901 ^ n9900 ^ 1'b0 ;
  assign n9904 = n9903 ^ n9902 ^ n6991 ;
  assign n9907 = n9906 ^ n9905 ^ n9904 ;
  assign n9910 = ( n1559 & n7408 ) | ( n1559 & ~n7756 ) | ( n7408 & ~n7756 ) ;
  assign n9908 = n4577 ^ n2697 ^ 1'b0 ;
  assign n9909 = n6685 & n9908 ;
  assign n9911 = n9910 ^ n9909 ^ n7330 ;
  assign n9912 = n9911 ^ n6795 ^ n5076 ;
  assign n9915 = n4633 ^ n2028 ^ n745 ;
  assign n9914 = n3509 ^ n1620 ^ n465 ;
  assign n9913 = ( n627 & n3506 ) | ( n627 & ~n9278 ) | ( n3506 & ~n9278 ) ;
  assign n9916 = n9915 ^ n9914 ^ n9913 ;
  assign n9917 = n5683 ^ n1198 ^ n707 ;
  assign n9918 = n8652 & n9917 ;
  assign n9919 = n9918 ^ n3359 ^ 1'b0 ;
  assign n9920 = n9876 ^ n7825 ^ n335 ;
  assign n9921 = n6666 & n9920 ;
  assign n9922 = ( n455 & ~n608 ) | ( n455 & n5398 ) | ( ~n608 & n5398 ) ;
  assign n9923 = n7574 ^ n539 ^ 1'b0 ;
  assign n9924 = n9923 ^ n6362 ^ n4287 ;
  assign n9925 = ( n9129 & ~n9922 ) | ( n9129 & n9924 ) | ( ~n9922 & n9924 ) ;
  assign n9926 = n2206 ^ n1711 ^ 1'b0 ;
  assign n9927 = ( n403 & n7158 ) | ( n403 & ~n9926 ) | ( n7158 & ~n9926 ) ;
  assign n9928 = n1977 | n2449 ;
  assign n9929 = n9928 ^ n7356 ^ 1'b0 ;
  assign n9930 = ( n8348 & ~n9927 ) | ( n8348 & n9929 ) | ( ~n9927 & n9929 ) ;
  assign n9931 = n1173 & n9930 ;
  assign n9932 = n9339 & n9931 ;
  assign n9933 = ( x115 & n726 ) | ( x115 & ~n1298 ) | ( n726 & ~n1298 ) ;
  assign n9934 = n9933 ^ n3597 ^ n2066 ;
  assign n9935 = ( n1760 & n3992 ) | ( n1760 & ~n9934 ) | ( n3992 & ~n9934 ) ;
  assign n9936 = n8857 ^ n4336 ^ n3601 ;
  assign n9937 = n9936 ^ n8997 ^ 1'b0 ;
  assign n9938 = n9937 ^ n4594 ^ n3809 ;
  assign n9939 = n9938 ^ n7924 ^ n4796 ;
  assign n9940 = ( n1918 & n7130 ) | ( n1918 & ~n9939 ) | ( n7130 & ~n9939 ) ;
  assign n9941 = ( n1474 & n4358 ) | ( n1474 & ~n9359 ) | ( n4358 & ~n9359 ) ;
  assign n9942 = n7197 ^ n6715 ^ n3819 ;
  assign n9943 = n6565 & ~n9942 ;
  assign n9944 = ~n9941 & n9943 ;
  assign n9946 = n3989 ^ n2498 ^ 1'b0 ;
  assign n9947 = n1294 & ~n9946 ;
  assign n9948 = n9947 ^ n2178 ^ n1192 ;
  assign n9949 = n9948 ^ n7240 ^ n1626 ;
  assign n9945 = ( ~n2330 & n3892 ) | ( ~n2330 & n5639 ) | ( n3892 & n5639 ) ;
  assign n9950 = n9949 ^ n9945 ^ n6479 ;
  assign n9951 = ( n1094 & n6069 ) | ( n1094 & ~n7201 ) | ( n6069 & ~n7201 ) ;
  assign n9952 = n9951 ^ n4790 ^ n334 ;
  assign n9953 = n2470 ^ n1375 ^ n1067 ;
  assign n9954 = n565 | n9953 ;
  assign n9956 = ( ~n1602 & n7278 ) | ( ~n1602 & n7531 ) | ( n7278 & n7531 ) ;
  assign n9955 = n7211 ^ n6893 ^ n2983 ;
  assign n9957 = n9956 ^ n9955 ^ n581 ;
  assign n9963 = n6078 ^ n377 ^ 1'b0 ;
  assign n9964 = n6864 & ~n9963 ;
  assign n9965 = ( n2637 & n8240 ) | ( n2637 & ~n8659 ) | ( n8240 & ~n8659 ) ;
  assign n9966 = n9965 ^ n2314 ^ 1'b0 ;
  assign n9967 = ~n9964 & n9966 ;
  assign n9961 = ( ~n2924 & n4038 ) | ( ~n2924 & n4767 ) | ( n4038 & n4767 ) ;
  assign n9958 = n3702 ^ n286 ^ 1'b0 ;
  assign n9959 = ~n423 & n9958 ;
  assign n9960 = n9959 ^ n5840 ^ n2073 ;
  assign n9962 = n9961 ^ n9960 ^ n7858 ;
  assign n9968 = n9967 ^ n9962 ^ n7419 ;
  assign n9969 = ( n9954 & n9957 ) | ( n9954 & ~n9968 ) | ( n9957 & ~n9968 ) ;
  assign n9970 = n6398 ^ n4517 ^ n2389 ;
  assign n9971 = ( ~n292 & n1130 ) | ( ~n292 & n9970 ) | ( n1130 & n9970 ) ;
  assign n9972 = ( n1684 & n5083 ) | ( n1684 & n8039 ) | ( n5083 & n8039 ) ;
  assign n9973 = ( ~n1679 & n1965 ) | ( ~n1679 & n4459 ) | ( n1965 & n4459 ) ;
  assign n9974 = ( n5098 & ~n9972 ) | ( n5098 & n9973 ) | ( ~n9972 & n9973 ) ;
  assign n9975 = n4485 ^ n4098 ^ n1984 ;
  assign n9977 = n9465 ^ n3105 ^ 1'b0 ;
  assign n9976 = n2181 ^ n1554 ^ n265 ;
  assign n9978 = n9977 ^ n9976 ^ n6855 ;
  assign n9979 = n3942 & n9978 ;
  assign n9980 = ~n9975 & n9979 ;
  assign n9981 = n9980 ^ n5753 ^ n444 ;
  assign n9982 = n5864 & n9981 ;
  assign n9983 = n1855 & ~n9658 ;
  assign n9984 = ( x47 & n2949 ) | ( x47 & ~n7106 ) | ( n2949 & ~n7106 ) ;
  assign n9985 = ( n3172 & n5581 ) | ( n3172 & n9884 ) | ( n5581 & n9884 ) ;
  assign n9986 = ( n5740 & n8187 ) | ( n5740 & ~n9985 ) | ( n8187 & ~n9985 ) ;
  assign n9987 = n9986 ^ n1049 ^ n783 ;
  assign n9988 = n7042 ^ n6801 ^ 1'b0 ;
  assign n9989 = ~n9987 & n9988 ;
  assign n9990 = n3784 ^ n512 ^ 1'b0 ;
  assign n9991 = n9990 ^ n4848 ^ n1645 ;
  assign n9992 = n9991 ^ n1580 ^ 1'b0 ;
  assign n9993 = n8674 ^ n7989 ^ n5296 ;
  assign n9995 = n5823 ^ n4445 ^ x11 ;
  assign n9994 = n9484 ^ n2673 ^ n532 ;
  assign n9996 = n9995 ^ n9994 ^ n281 ;
  assign n9997 = n3258 & n8154 ;
  assign n9998 = n7652 ^ n5430 ^ n4591 ;
  assign n9999 = ( n135 & n7545 ) | ( n135 & ~n9998 ) | ( n7545 & ~n9998 ) ;
  assign n10000 = ( n8356 & ~n9997 ) | ( n8356 & n9999 ) | ( ~n9997 & n9999 ) ;
  assign n10008 = n841 & n3075 ;
  assign n10001 = n7032 ^ n5630 ^ n2657 ;
  assign n10002 = ( ~n1262 & n2138 ) | ( ~n1262 & n3697 ) | ( n2138 & n3697 ) ;
  assign n10003 = ( ~n1374 & n2560 ) | ( ~n1374 & n10002 ) | ( n2560 & n10002 ) ;
  assign n10004 = n270 & n10003 ;
  assign n10005 = ~n2110 & n10004 ;
  assign n10006 = ( n1777 & ~n9759 ) | ( n1777 & n10005 ) | ( ~n9759 & n10005 ) ;
  assign n10007 = n10001 & ~n10006 ;
  assign n10009 = n10008 ^ n10007 ^ 1'b0 ;
  assign n10016 = n8795 ^ n4856 ^ n2409 ;
  assign n10017 = n10016 ^ n2262 ^ n2156 ;
  assign n10010 = n8770 ^ n3206 ^ n584 ;
  assign n10011 = ( ~n334 & n5914 ) | ( ~n334 & n6011 ) | ( n5914 & n6011 ) ;
  assign n10012 = ( n2722 & ~n7815 ) | ( n2722 & n10011 ) | ( ~n7815 & n10011 ) ;
  assign n10013 = n10012 ^ n9275 ^ n7480 ;
  assign n10014 = ( n6204 & n10010 ) | ( n6204 & n10013 ) | ( n10010 & n10013 ) ;
  assign n10015 = n10014 ^ n2825 ^ n289 ;
  assign n10018 = n10017 ^ n10015 ^ n287 ;
  assign n10019 = ( ~x37 & n482 ) | ( ~x37 & n1926 ) | ( n482 & n1926 ) ;
  assign n10020 = ( n6450 & n8039 ) | ( n6450 & ~n10019 ) | ( n8039 & ~n10019 ) ;
  assign n10021 = n7026 ^ n3550 ^ x116 ;
  assign n10022 = n2823 | n10021 ;
  assign n10023 = n10020 | n10022 ;
  assign n10024 = ( x57 & n7281 ) | ( x57 & n10023 ) | ( n7281 & n10023 ) ;
  assign n10026 = n180 & n2354 ;
  assign n10025 = n7755 ^ n2402 ^ n1913 ;
  assign n10027 = n10026 ^ n10025 ^ n7377 ;
  assign n10028 = ( x106 & n1289 ) | ( x106 & n9020 ) | ( n1289 & n9020 ) ;
  assign n10029 = ( n905 & n6557 ) | ( n905 & ~n6858 ) | ( n6557 & ~n6858 ) ;
  assign n10030 = ( n864 & ~n7940 ) | ( n864 & n10029 ) | ( ~n7940 & n10029 ) ;
  assign n10031 = n3206 & ~n4153 ;
  assign n10032 = n8297 & n10031 ;
  assign n10033 = ( n756 & n3116 ) | ( n756 & ~n10032 ) | ( n3116 & ~n10032 ) ;
  assign n10034 = n10033 ^ n7278 ^ n2291 ;
  assign n10035 = n4770 & ~n6957 ;
  assign n10036 = n10035 ^ n3615 ^ 1'b0 ;
  assign n10038 = n8354 ^ n6044 ^ 1'b0 ;
  assign n10039 = ( n982 & n2649 ) | ( n982 & ~n10038 ) | ( n2649 & ~n10038 ) ;
  assign n10037 = n4761 ^ n4730 ^ n2659 ;
  assign n10040 = n10039 ^ n10037 ^ n7689 ;
  assign n10041 = n5697 & n10040 ;
  assign n10042 = n10041 ^ n3120 ^ 1'b0 ;
  assign n10043 = n10042 ^ n9642 ^ n6206 ;
  assign n10044 = ( n1927 & n2462 ) | ( n1927 & ~n7987 ) | ( n2462 & ~n7987 ) ;
  assign n10045 = ( n2318 & n4329 ) | ( n2318 & n10044 ) | ( n4329 & n10044 ) ;
  assign n10046 = n2698 | n10045 ;
  assign n10047 = ( n5090 & n6523 ) | ( n5090 & ~n10046 ) | ( n6523 & ~n10046 ) ;
  assign n10048 = n10047 ^ n7258 ^ n2471 ;
  assign n10049 = n10048 ^ n9861 ^ n9578 ;
  assign n10050 = n829 & n6228 ;
  assign n10051 = n3030 ^ n467 ^ 1'b0 ;
  assign n10052 = n10051 ^ n8920 ^ 1'b0 ;
  assign n10053 = n10052 ^ n6895 ^ x57 ;
  assign n10054 = n4422 & ~n10053 ;
  assign n10055 = ( n1738 & n10050 ) | ( n1738 & n10054 ) | ( n10050 & n10054 ) ;
  assign n10056 = ~n908 & n10055 ;
  assign n10062 = n370 | n2854 ;
  assign n10063 = n5999 & ~n10062 ;
  assign n10057 = n4682 ^ n3653 ^ n817 ;
  assign n10058 = n10057 ^ n2358 ^ 1'b0 ;
  assign n10059 = n9147 | n10058 ;
  assign n10060 = n10059 ^ n6676 ^ n3825 ;
  assign n10061 = n10060 ^ n8844 ^ n1594 ;
  assign n10064 = n10063 ^ n10061 ^ n2353 ;
  assign n10073 = ( n1463 & n3153 ) | ( n1463 & ~n5779 ) | ( n3153 & ~n5779 ) ;
  assign n10065 = ( n3630 & n5008 ) | ( n3630 & n9801 ) | ( n5008 & n9801 ) ;
  assign n10068 = ( n410 & n1079 ) | ( n410 & n1863 ) | ( n1079 & n1863 ) ;
  assign n10067 = ( x50 & n503 ) | ( x50 & ~n3517 ) | ( n503 & ~n3517 ) ;
  assign n10066 = n5294 ^ n3142 ^ x36 ;
  assign n10069 = n10068 ^ n10067 ^ n10066 ;
  assign n10070 = n10069 ^ n6096 ^ 1'b0 ;
  assign n10071 = n8222 ^ n3997 ^ n1664 ;
  assign n10072 = ( n10065 & ~n10070 ) | ( n10065 & n10071 ) | ( ~n10070 & n10071 ) ;
  assign n10074 = n10073 ^ n10072 ^ n674 ;
  assign n10079 = n4770 ^ n4532 ^ n192 ;
  assign n10077 = n9259 ^ n6698 ^ n4141 ;
  assign n10078 = n10077 ^ n8356 ^ n4162 ;
  assign n10075 = ( x61 & ~n2234 ) | ( x61 & n6099 ) | ( ~n2234 & n6099 ) ;
  assign n10076 = n10075 ^ n9450 ^ n8412 ;
  assign n10080 = n10079 ^ n10078 ^ n10076 ;
  assign n10081 = n10074 & ~n10080 ;
  assign n10082 = n6713 ^ n1783 ^ 1'b0 ;
  assign n10083 = n2255 & ~n10082 ;
  assign n10084 = n10083 ^ n1869 ^ n674 ;
  assign n10085 = n4931 ^ n801 ^ 1'b0 ;
  assign n10086 = n5173 ^ n3073 ^ 1'b0 ;
  assign n10087 = n4610 & ~n10086 ;
  assign n10088 = ( n2476 & ~n3488 ) | ( n2476 & n3672 ) | ( ~n3488 & n3672 ) ;
  assign n10089 = ( ~x73 & n10087 ) | ( ~x73 & n10088 ) | ( n10087 & n10088 ) ;
  assign n10090 = ( ~n543 & n1421 ) | ( ~n543 & n2407 ) | ( n1421 & n2407 ) ;
  assign n10091 = n10090 ^ n4167 ^ n1247 ;
  assign n10092 = ( ~n10085 & n10089 ) | ( ~n10085 & n10091 ) | ( n10089 & n10091 ) ;
  assign n10099 = ( n791 & n2924 ) | ( n791 & ~n3575 ) | ( n2924 & ~n3575 ) ;
  assign n10098 = ~n1705 & n2884 ;
  assign n10093 = n3797 & n9573 ;
  assign n10094 = n8534 ^ n8273 ^ n965 ;
  assign n10095 = ( ~n3308 & n10093 ) | ( ~n3308 & n10094 ) | ( n10093 & n10094 ) ;
  assign n10096 = ~n8219 & n10095 ;
  assign n10097 = n10096 ^ n8580 ^ 1'b0 ;
  assign n10100 = n10099 ^ n10098 ^ n10097 ;
  assign n10101 = n6515 ^ n3219 ^ n3028 ;
  assign n10102 = ( n5722 & n7341 ) | ( n5722 & n10101 ) | ( n7341 & n10101 ) ;
  assign n10103 = n2178 ^ n853 ^ n210 ;
  assign n10104 = n10103 ^ n6210 ^ n1890 ;
  assign n10105 = ( n1757 & ~n3165 ) | ( n1757 & n8913 ) | ( ~n3165 & n8913 ) ;
  assign n10106 = ( x56 & n1179 ) | ( x56 & ~n4779 ) | ( n1179 & ~n4779 ) ;
  assign n10107 = ( n6446 & n9462 ) | ( n6446 & n10106 ) | ( n9462 & n10106 ) ;
  assign n10108 = ( ~n276 & n10105 ) | ( ~n276 & n10107 ) | ( n10105 & n10107 ) ;
  assign n10109 = ( x112 & n4328 ) | ( x112 & ~n7273 ) | ( n4328 & ~n7273 ) ;
  assign n10110 = n10109 ^ n2253 ^ n1436 ;
  assign n10111 = n9165 ^ n8302 ^ n1170 ;
  assign n10115 = n942 ^ n881 ^ n586 ;
  assign n10112 = ( ~n1052 & n1775 ) | ( ~n1052 & n4233 ) | ( n1775 & n4233 ) ;
  assign n10113 = n211 & ~n10112 ;
  assign n10114 = n9118 & n10113 ;
  assign n10116 = n10115 ^ n10114 ^ n9683 ;
  assign n10117 = ( n6271 & n8862 ) | ( n6271 & n8956 ) | ( n8862 & n8956 ) ;
  assign n10118 = ( n1753 & n8598 ) | ( n1753 & n10117 ) | ( n8598 & n10117 ) ;
  assign n10119 = n573 & ~n1951 ;
  assign n10120 = n1451 & n10119 ;
  assign n10121 = n10120 ^ n5969 ^ n4608 ;
  assign n10122 = ( n7292 & n9742 ) | ( n7292 & n10121 ) | ( n9742 & n10121 ) ;
  assign n10127 = n1588 ^ n1315 ^ n358 ;
  assign n10123 = n1764 & n8869 ;
  assign n10124 = n1984 & n10123 ;
  assign n10125 = n10124 ^ n5924 ^ n5630 ;
  assign n10126 = ( n278 & ~n8832 ) | ( n278 & n10125 ) | ( ~n8832 & n10125 ) ;
  assign n10128 = n10127 ^ n10126 ^ n9025 ;
  assign n10134 = n7663 ^ n6135 ^ n2438 ;
  assign n10135 = ~n816 & n10134 ;
  assign n10136 = n10135 ^ n2520 ^ 1'b0 ;
  assign n10131 = n5284 ^ n1525 ^ n986 ;
  assign n10132 = n10131 ^ n3148 ^ n1492 ;
  assign n10129 = n7284 ^ n2826 ^ n274 ;
  assign n10130 = n10129 ^ n6781 ^ n3726 ;
  assign n10133 = n10132 ^ n10130 ^ n3564 ;
  assign n10137 = n10136 ^ n10133 ^ n5195 ;
  assign n10138 = n9512 ^ n1801 ^ 1'b0 ;
  assign n10139 = n9573 ^ n298 ^ 1'b0 ;
  assign n10140 = n10139 ^ n2080 ^ n1744 ;
  assign n10141 = ~n2570 & n10140 ;
  assign n10142 = n10141 ^ n8099 ^ 1'b0 ;
  assign n10143 = n4094 ^ n3976 ^ n1958 ;
  assign n10144 = n10143 ^ n10033 ^ n7297 ;
  assign n10145 = ( n9600 & ~n10142 ) | ( n9600 & n10144 ) | ( ~n10142 & n10144 ) ;
  assign n10146 = ( n1599 & ~n3830 ) | ( n1599 & n4328 ) | ( ~n3830 & n4328 ) ;
  assign n10147 = n10146 ^ n3506 ^ n2106 ;
  assign n10148 = ( n448 & n1345 ) | ( n448 & n1367 ) | ( n1345 & n1367 ) ;
  assign n10149 = n10148 ^ n8565 ^ n1601 ;
  assign n10150 = ( n2151 & n3861 ) | ( n2151 & ~n9933 ) | ( n3861 & ~n9933 ) ;
  assign n10151 = ( n8588 & n10149 ) | ( n8588 & n10150 ) | ( n10149 & n10150 ) ;
  assign n10152 = ( n1024 & n1837 ) | ( n1024 & ~n8470 ) | ( n1837 & ~n8470 ) ;
  assign n10153 = ~n2135 & n10152 ;
  assign n10154 = n938 & ~n10153 ;
  assign n10155 = n10154 ^ n4721 ^ n2580 ;
  assign n10156 = ( n915 & n2297 ) | ( n915 & n4446 ) | ( n2297 & n4446 ) ;
  assign n10157 = ( ~n2830 & n6088 ) | ( ~n2830 & n10156 ) | ( n6088 & n10156 ) ;
  assign n10158 = ~n2615 & n6148 ;
  assign n10159 = n10157 & n10158 ;
  assign n10160 = n7498 ^ n6767 ^ 1'b0 ;
  assign n10161 = ~n10159 & n10160 ;
  assign n10162 = ( x40 & n5556 ) | ( x40 & ~n5818 ) | ( n5556 & ~n5818 ) ;
  assign n10163 = n7157 ^ n3170 ^ 1'b0 ;
  assign n10164 = n8048 & ~n10163 ;
  assign n10165 = n10164 ^ x66 ^ 1'b0 ;
  assign n10166 = ( ~n3465 & n10162 ) | ( ~n3465 & n10165 ) | ( n10162 & n10165 ) ;
  assign n10167 = n10166 ^ n9342 ^ n1427 ;
  assign n10170 = ~n609 & n3219 ;
  assign n10168 = n5486 ^ n5014 ^ n2785 ;
  assign n10169 = n10168 ^ n9109 ^ n4251 ;
  assign n10171 = n10170 ^ n10169 ^ n3489 ;
  assign n10172 = ( n1366 & n7810 ) | ( n1366 & n9683 ) | ( n7810 & n9683 ) ;
  assign n10173 = n10172 ^ n3409 ^ 1'b0 ;
  assign n10174 = n3207 ^ n1039 ^ 1'b0 ;
  assign n10175 = ( ~x98 & n5622 ) | ( ~x98 & n6086 ) | ( n5622 & n6086 ) ;
  assign n10176 = n10175 ^ n1849 ^ 1'b0 ;
  assign n10177 = ( n152 & n10174 ) | ( n152 & n10176 ) | ( n10174 & n10176 ) ;
  assign n10178 = n4635 ^ n3489 ^ n337 ;
  assign n10179 = n2663 ^ n2285 ^ n1367 ;
  assign n10180 = n10179 ^ n1632 ^ 1'b0 ;
  assign n10181 = n10180 ^ n4717 ^ n4140 ;
  assign n10182 = n10181 ^ n2446 ^ n1144 ;
  assign n10183 = ( ~n8784 & n10178 ) | ( ~n8784 & n10182 ) | ( n10178 & n10182 ) ;
  assign n10184 = ( n8339 & n10177 ) | ( n8339 & n10183 ) | ( n10177 & n10183 ) ;
  assign n10185 = n10184 ^ n4553 ^ n3287 ;
  assign n10186 = ( ~n1449 & n1510 ) | ( ~n1449 & n1881 ) | ( n1510 & n1881 ) ;
  assign n10187 = ( n5177 & n5695 ) | ( n5177 & n10186 ) | ( n5695 & n10186 ) ;
  assign n10188 = n10187 ^ n7033 ^ 1'b0 ;
  assign n10189 = ( n1946 & n2277 ) | ( n1946 & ~n2991 ) | ( n2277 & ~n2991 ) ;
  assign n10190 = n10189 ^ n9075 ^ n6790 ;
  assign n10191 = ( n799 & n3557 ) | ( n799 & ~n4875 ) | ( n3557 & ~n4875 ) ;
  assign n10194 = n3419 ^ n2465 ^ n1393 ;
  assign n10195 = n1780 & ~n10194 ;
  assign n10196 = n10195 ^ n3215 ^ 1'b0 ;
  assign n10192 = n2148 ^ n1937 ^ 1'b0 ;
  assign n10193 = n586 & ~n10192 ;
  assign n10197 = n10196 ^ n10193 ^ n5718 ;
  assign n10198 = n10197 ^ n6130 ^ 1'b0 ;
  assign n10199 = n9235 | n10198 ;
  assign n10200 = ( n9069 & n9663 ) | ( n9069 & ~n10199 ) | ( n9663 & ~n10199 ) ;
  assign n10201 = ~n10191 & n10200 ;
  assign n10202 = n10190 & n10201 ;
  assign n10203 = n6443 ^ n6439 ^ n3307 ;
  assign n10204 = ( ~n2339 & n4416 ) | ( ~n2339 & n4704 ) | ( n4416 & n4704 ) ;
  assign n10205 = n10204 ^ n7375 ^ n4032 ;
  assign n10206 = n10205 ^ n1439 ^ 1'b0 ;
  assign n10210 = n530 | n1257 ;
  assign n10207 = ( x76 & n1254 ) | ( x76 & ~n7037 ) | ( n1254 & ~n7037 ) ;
  assign n10208 = n3524 & n10207 ;
  assign n10209 = n10208 ^ n6932 ^ 1'b0 ;
  assign n10211 = n10210 ^ n10209 ^ n9487 ;
  assign n10212 = ( n10203 & n10206 ) | ( n10203 & n10211 ) | ( n10206 & n10211 ) ;
  assign n10213 = n785 & n9399 ;
  assign n10214 = n2815 & n4448 ;
  assign n10215 = n10213 & n10214 ;
  assign n10216 = n5846 ^ n5009 ^ n767 ;
  assign n10217 = n9732 | n10216 ;
  assign n10218 = n10217 ^ n293 ^ 1'b0 ;
  assign n10219 = ( n999 & n1566 ) | ( n999 & ~n4974 ) | ( n1566 & ~n4974 ) ;
  assign n10220 = ( n10215 & ~n10218 ) | ( n10215 & n10219 ) | ( ~n10218 & n10219 ) ;
  assign n10224 = ( n2989 & n3717 ) | ( n2989 & n4206 ) | ( n3717 & n4206 ) ;
  assign n10223 = ( n5466 & n6705 ) | ( n5466 & n6888 ) | ( n6705 & n6888 ) ;
  assign n10221 = x102 & n1286 ;
  assign n10222 = n9224 & n10221 ;
  assign n10225 = n10224 ^ n10223 ^ n10222 ;
  assign n10226 = ( n2767 & ~n7015 ) | ( n2767 & n10225 ) | ( ~n7015 & n10225 ) ;
  assign n10227 = n2751 & n5893 ;
  assign n10228 = n10227 ^ n4225 ^ 1'b0 ;
  assign n10229 = n10228 ^ n3830 ^ n2703 ;
  assign n10237 = ( n6357 & ~n7156 ) | ( n6357 & n7979 ) | ( ~n7156 & n7979 ) ;
  assign n10234 = ( n832 & n1808 ) | ( n832 & n2930 ) | ( n1808 & n2930 ) ;
  assign n10235 = n10234 ^ n1751 ^ n591 ;
  assign n10232 = ( n3861 & n5661 ) | ( n3861 & ~n10066 ) | ( n5661 & ~n10066 ) ;
  assign n10233 = n10232 ^ n1148 ^ n133 ;
  assign n10236 = n10235 ^ n10233 ^ 1'b0 ;
  assign n10238 = n10237 ^ n10236 ^ n1341 ;
  assign n10239 = n10238 ^ n10011 ^ n3793 ;
  assign n10230 = ( n745 & n1608 ) | ( n745 & ~n2305 ) | ( n1608 & ~n2305 ) ;
  assign n10231 = n10230 ^ n3479 ^ n1181 ;
  assign n10240 = n10239 ^ n10231 ^ n7317 ;
  assign n10241 = ( n5420 & n6307 ) | ( n5420 & ~n10240 ) | ( n6307 & ~n10240 ) ;
  assign n10242 = n6233 ^ n3611 ^ n1737 ;
  assign n10244 = n8476 ^ n7404 ^ n4678 ;
  assign n10243 = ( n187 & n4116 ) | ( n187 & ~n8248 ) | ( n4116 & ~n8248 ) ;
  assign n10245 = n10244 ^ n10243 ^ n9195 ;
  assign n10246 = ( ~n8394 & n10242 ) | ( ~n8394 & n10245 ) | ( n10242 & n10245 ) ;
  assign n10247 = n7621 ^ n4257 ^ n1430 ;
  assign n10248 = n10247 ^ n3768 ^ 1'b0 ;
  assign n10249 = ( n4039 & ~n4516 ) | ( n4039 & n6409 ) | ( ~n4516 & n6409 ) ;
  assign n10250 = n10249 ^ n8980 ^ 1'b0 ;
  assign n10251 = ( n2226 & ~n4896 ) | ( n2226 & n7933 ) | ( ~n4896 & n7933 ) ;
  assign n10252 = ( n5619 & n6539 ) | ( n5619 & n10251 ) | ( n6539 & n10251 ) ;
  assign n10253 = ( n8195 & ~n9699 ) | ( n8195 & n10252 ) | ( ~n9699 & n10252 ) ;
  assign n10254 = n1917 ^ n1442 ^ n982 ;
  assign n10255 = ( n6860 & n8458 ) | ( n6860 & ~n10254 ) | ( n8458 & ~n10254 ) ;
  assign n10256 = ( x36 & ~n641 ) | ( x36 & n7512 ) | ( ~n641 & n7512 ) ;
  assign n10257 = n4299 & n6313 ;
  assign n10258 = ( ~n405 & n3627 ) | ( ~n405 & n9174 ) | ( n3627 & n9174 ) ;
  assign n10259 = ( n8551 & n10257 ) | ( n8551 & ~n10258 ) | ( n10257 & ~n10258 ) ;
  assign n10263 = ( n2801 & ~n3331 ) | ( n2801 & n8294 ) | ( ~n3331 & n8294 ) ;
  assign n10264 = ( n206 & ~n1795 ) | ( n206 & n10263 ) | ( ~n1795 & n10263 ) ;
  assign n10260 = n6373 ^ n249 ^ 1'b0 ;
  assign n10261 = ~n864 & n10260 ;
  assign n10262 = n10261 ^ n6157 ^ n1135 ;
  assign n10265 = n10264 ^ n10262 ^ n8983 ;
  assign n10266 = n10265 ^ n6396 ^ n3691 ;
  assign n10267 = n1684 | n1739 ;
  assign n10268 = n10267 ^ n7493 ^ 1'b0 ;
  assign n10269 = n10268 ^ n6023 ^ n536 ;
  assign n10270 = n4722 ^ n3189 ^ n2010 ;
  assign n10271 = n1902 | n7577 ;
  assign n10272 = n5418 ^ n4842 ^ n818 ;
  assign n10273 = ( n1565 & n1825 ) | ( n1565 & n2398 ) | ( n1825 & n2398 ) ;
  assign n10274 = ( ~n2129 & n10272 ) | ( ~n2129 & n10273 ) | ( n10272 & n10273 ) ;
  assign n10275 = ( n446 & n982 ) | ( n446 & ~n10274 ) | ( n982 & ~n10274 ) ;
  assign n10276 = ( n2235 & ~n4283 ) | ( n2235 & n6896 ) | ( ~n4283 & n6896 ) ;
  assign n10277 = n2345 ^ n2165 ^ n1293 ;
  assign n10278 = ( ~n5284 & n10276 ) | ( ~n5284 & n10277 ) | ( n10276 & n10277 ) ;
  assign n10279 = n10278 ^ n7824 ^ 1'b0 ;
  assign n10280 = ~n8481 & n10279 ;
  assign n10281 = ( n8148 & n9584 ) | ( n8148 & n10280 ) | ( n9584 & n10280 ) ;
  assign n10282 = n10281 ^ n8981 ^ n7264 ;
  assign n10283 = ( ~n10271 & n10275 ) | ( ~n10271 & n10282 ) | ( n10275 & n10282 ) ;
  assign n10284 = n2078 | n9585 ;
  assign n10285 = n5660 | n10284 ;
  assign n10286 = n10285 ^ n9341 ^ n3596 ;
  assign n10287 = n9094 ^ n6700 ^ n5312 ;
  assign n10288 = ( ~n2397 & n4013 ) | ( ~n2397 & n10287 ) | ( n4013 & n10287 ) ;
  assign n10289 = n9603 | n10288 ;
  assign n10290 = n1636 | n10289 ;
  assign n10291 = n5110 ^ n4816 ^ n3099 ;
  assign n10292 = ( n5617 & n9596 ) | ( n5617 & ~n10291 ) | ( n9596 & ~n10291 ) ;
  assign n10293 = ( n1262 & ~n10290 ) | ( n1262 & n10292 ) | ( ~n10290 & n10292 ) ;
  assign n10298 = ( n4328 & ~n8969 ) | ( n4328 & n9732 ) | ( ~n8969 & n9732 ) ;
  assign n10295 = n8877 ^ n1913 ^ x37 ;
  assign n10296 = n10295 ^ n7945 ^ 1'b0 ;
  assign n10294 = n3365 & ~n9770 ;
  assign n10297 = n10296 ^ n10294 ^ 1'b0 ;
  assign n10299 = n10298 ^ n10297 ^ 1'b0 ;
  assign n10300 = n7196 ^ n5020 ^ n996 ;
  assign n10301 = n1133 & ~n6598 ;
  assign n10302 = n10301 ^ n6189 ^ 1'b0 ;
  assign n10303 = ( n466 & n967 ) | ( n466 & n10302 ) | ( n967 & n10302 ) ;
  assign n10306 = n7726 ^ n4605 ^ n1394 ;
  assign n10304 = n2055 ^ n1633 ^ n1185 ;
  assign n10305 = n10304 ^ n3734 ^ n524 ;
  assign n10307 = n10306 ^ n10305 ^ x41 ;
  assign n10308 = n4805 & n6596 ;
  assign n10309 = n8515 & n10308 ;
  assign n10310 = ( ~n1244 & n4066 ) | ( ~n1244 & n10309 ) | ( n4066 & n10309 ) ;
  assign n10311 = ( ~n4758 & n10307 ) | ( ~n4758 & n10310 ) | ( n10307 & n10310 ) ;
  assign n10312 = ( ~n5250 & n10303 ) | ( ~n5250 & n10311 ) | ( n10303 & n10311 ) ;
  assign n10313 = n205 & ~n2686 ;
  assign n10314 = n1341 & n10313 ;
  assign n10315 = n10314 ^ n4685 ^ n1750 ;
  assign n10316 = n10315 ^ n5878 ^ n3145 ;
  assign n10317 = n10246 ^ n305 ^ 1'b0 ;
  assign n10318 = n3422 ^ n3111 ^ 1'b0 ;
  assign n10319 = n390 & ~n5625 ;
  assign n10320 = n10319 ^ n4311 ^ n3493 ;
  assign n10323 = n6806 ^ n6100 ^ n1736 ;
  assign n10321 = ( n1380 & n7476 ) | ( n1380 & n8821 ) | ( n7476 & n8821 ) ;
  assign n10322 = n10321 ^ n4058 ^ n3993 ;
  assign n10324 = n10323 ^ n10322 ^ n6137 ;
  assign n10325 = ( x40 & ~n10050 ) | ( x40 & n10324 ) | ( ~n10050 & n10324 ) ;
  assign n10326 = n5060 ^ n2781 ^ n1569 ;
  assign n10327 = ( n1936 & n8135 ) | ( n1936 & ~n10326 ) | ( n8135 & ~n10326 ) ;
  assign n10328 = n6613 ^ n1859 ^ n1689 ;
  assign n10329 = n180 ^ x101 ^ 1'b0 ;
  assign n10330 = n284 & n10329 ;
  assign n10331 = ( x92 & n898 ) | ( x92 & ~n904 ) | ( n898 & ~n904 ) ;
  assign n10332 = ( n1715 & n10330 ) | ( n1715 & ~n10331 ) | ( n10330 & ~n10331 ) ;
  assign n10333 = ( n1649 & n7151 ) | ( n1649 & n10332 ) | ( n7151 & n10332 ) ;
  assign n10334 = ( n418 & n1016 ) | ( n418 & ~n4906 ) | ( n1016 & ~n4906 ) ;
  assign n10335 = ( n10328 & n10333 ) | ( n10328 & n10334 ) | ( n10333 & n10334 ) ;
  assign n10337 = n6251 & n9257 ;
  assign n10338 = ~x34 & n10337 ;
  assign n10336 = ( ~n983 & n1037 ) | ( ~n983 & n5153 ) | ( n1037 & n5153 ) ;
  assign n10339 = n10338 ^ n10336 ^ 1'b0 ;
  assign n10340 = ( n1050 & n7192 ) | ( n1050 & ~n10339 ) | ( n7192 & ~n10339 ) ;
  assign n10341 = ~n3720 & n3846 ;
  assign n10342 = n10341 ^ n4386 ^ 1'b0 ;
  assign n10343 = n3023 ^ n1836 ^ 1'b0 ;
  assign n10344 = n954 | n10343 ;
  assign n10345 = ( n1150 & ~n6648 ) | ( n1150 & n10344 ) | ( ~n6648 & n10344 ) ;
  assign n10346 = n1342 | n10345 ;
  assign n10347 = n4874 & ~n10346 ;
  assign n10348 = ( n1549 & ~n4746 ) | ( n1549 & n10347 ) | ( ~n4746 & n10347 ) ;
  assign n10349 = ( ~n6875 & n10342 ) | ( ~n6875 & n10348 ) | ( n10342 & n10348 ) ;
  assign n10350 = n9830 & n10349 ;
  assign n10351 = n10350 ^ n502 ^ 1'b0 ;
  assign n10352 = ( ~n7837 & n10088 ) | ( ~n7837 & n10351 ) | ( n10088 & n10351 ) ;
  assign n10353 = n8684 ^ n1685 ^ n1619 ;
  assign n10354 = n10353 ^ n3998 ^ n2596 ;
  assign n10355 = n8829 ^ n5008 ^ n2013 ;
  assign n10356 = n10355 ^ n3310 ^ n794 ;
  assign n10357 = n3931 ^ n3865 ^ n1553 ;
  assign n10358 = ( n1465 & n1510 ) | ( n1465 & n6454 ) | ( n1510 & n6454 ) ;
  assign n10359 = ( n6819 & n10357 ) | ( n6819 & ~n10358 ) | ( n10357 & ~n10358 ) ;
  assign n10360 = ( n8645 & n10356 ) | ( n8645 & n10359 ) | ( n10356 & n10359 ) ;
  assign n10361 = n375 ^ n147 ^ x109 ;
  assign n10362 = ~n8651 & n10361 ;
  assign n10363 = n10362 ^ n7132 ^ 1'b0 ;
  assign n10364 = ( ~n2988 & n7429 ) | ( ~n2988 & n10363 ) | ( n7429 & n10363 ) ;
  assign n10365 = ( n6200 & n10360 ) | ( n6200 & n10364 ) | ( n10360 & n10364 ) ;
  assign n10366 = n10365 ^ n1093 ^ n478 ;
  assign n10367 = n3715 & n10366 ;
  assign n10368 = ~n6867 & n10367 ;
  assign n10373 = n9225 ^ n5777 ^ n4919 ;
  assign n10371 = n8754 ^ n2747 ^ n211 ;
  assign n10369 = n9510 ^ n1562 ^ n1386 ;
  assign n10370 = n8101 | n10369 ;
  assign n10372 = n10371 ^ n10370 ^ 1'b0 ;
  assign n10374 = n10373 ^ n10372 ^ n1771 ;
  assign n10375 = ( ~n1653 & n1910 ) | ( ~n1653 & n4556 ) | ( n1910 & n4556 ) ;
  assign n10376 = n10375 ^ n6423 ^ n133 ;
  assign n10377 = n3082 & n10376 ;
  assign n10378 = ~n4403 & n6562 ;
  assign n10379 = n10378 ^ n2013 ^ 1'b0 ;
  assign n10383 = n2771 | n4419 ;
  assign n10384 = n10383 ^ n5129 ^ 1'b0 ;
  assign n10388 = n5382 & n7890 ;
  assign n10389 = ( x8 & n4066 ) | ( x8 & ~n10388 ) | ( n4066 & ~n10388 ) ;
  assign n10387 = n4554 & ~n7447 ;
  assign n10390 = n10389 ^ n10387 ^ 1'b0 ;
  assign n10391 = n10390 ^ n10178 ^ n1289 ;
  assign n10385 = ( n491 & n577 ) | ( n491 & n3547 ) | ( n577 & n3547 ) ;
  assign n10386 = n10385 ^ n460 ^ 1'b0 ;
  assign n10392 = n10391 ^ n10386 ^ n6607 ;
  assign n10395 = n6332 ^ n4774 ^ n3217 ;
  assign n10393 = n1391 | n8758 ;
  assign n10394 = ( n1420 & n4850 ) | ( n1420 & ~n10393 ) | ( n4850 & ~n10393 ) ;
  assign n10396 = n10395 ^ n10394 ^ n2000 ;
  assign n10397 = n10392 & n10396 ;
  assign n10398 = n10384 & ~n10397 ;
  assign n10380 = ( n1915 & n2328 ) | ( n1915 & ~n3939 ) | ( n2328 & ~n3939 ) ;
  assign n10381 = ( n3122 & n3271 ) | ( n3122 & n10380 ) | ( n3271 & n10380 ) ;
  assign n10382 = n10381 ^ n5168 ^ n1426 ;
  assign n10399 = n10398 ^ n10382 ^ 1'b0 ;
  assign n10401 = ( n2454 & ~n6164 ) | ( n2454 & n8566 ) | ( ~n6164 & n8566 ) ;
  assign n10400 = ( n1089 & ~n1798 ) | ( n1089 & n4294 ) | ( ~n1798 & n4294 ) ;
  assign n10402 = n10401 ^ n10400 ^ n5420 ;
  assign n10403 = n10402 ^ n1158 ^ n945 ;
  assign n10404 = ( n187 & n440 ) | ( n187 & ~n2844 ) | ( n440 & ~n2844 ) ;
  assign n10405 = n8247 ^ n5464 ^ 1'b0 ;
  assign n10406 = ~n10404 & n10405 ;
  assign n10413 = ( n2148 & ~n2400 ) | ( n2148 & n6655 ) | ( ~n2400 & n6655 ) ;
  assign n10411 = n9054 ^ n2404 ^ n699 ;
  assign n10412 = ( ~n3182 & n5088 ) | ( ~n3182 & n10411 ) | ( n5088 & n10411 ) ;
  assign n10407 = ( n2452 & n3616 ) | ( n2452 & ~n4725 ) | ( n3616 & ~n4725 ) ;
  assign n10408 = n7096 ^ n6981 ^ n620 ;
  assign n10409 = ( ~n6040 & n10407 ) | ( ~n6040 & n10408 ) | ( n10407 & n10408 ) ;
  assign n10410 = n10409 ^ n3272 ^ n1443 ;
  assign n10414 = n10413 ^ n10412 ^ n10410 ;
  assign n10416 = n9889 ^ n3275 ^ n1728 ;
  assign n10415 = ( n1617 & n7413 ) | ( n1617 & ~n8187 ) | ( n7413 & ~n8187 ) ;
  assign n10417 = n10416 ^ n10415 ^ n7043 ;
  assign n10418 = n3673 ^ n2137 ^ n908 ;
  assign n10419 = n10418 ^ n172 ^ 1'b0 ;
  assign n10420 = n3737 & n10419 ;
  assign n10421 = ~n7366 & n10420 ;
  assign n10423 = n1595 ^ n1055 ^ n442 ;
  assign n10422 = n3515 | n9118 ;
  assign n10424 = n10423 ^ n10422 ^ 1'b0 ;
  assign n10431 = n5194 ^ n228 ^ 1'b0 ;
  assign n10428 = n5919 ^ n5788 ^ 1'b0 ;
  assign n10429 = ~n452 & n10428 ;
  assign n10425 = ( n1883 & n3048 ) | ( n1883 & ~n4335 ) | ( n3048 & ~n4335 ) ;
  assign n10426 = ( ~n4640 & n4785 ) | ( ~n4640 & n8896 ) | ( n4785 & n8896 ) ;
  assign n10427 = ( n3652 & n10425 ) | ( n3652 & n10426 ) | ( n10425 & n10426 ) ;
  assign n10430 = n10429 ^ n10427 ^ n6410 ;
  assign n10432 = n10431 ^ n10430 ^ n6079 ;
  assign n10433 = ~n3432 & n5386 ;
  assign n10434 = n10433 ^ n2472 ^ 1'b0 ;
  assign n10435 = n5418 ^ n140 ^ 1'b0 ;
  assign n10436 = n2274 & n10435 ;
  assign n10437 = ( n7404 & ~n10434 ) | ( n7404 & n10436 ) | ( ~n10434 & n10436 ) ;
  assign n10438 = n6127 ^ n1578 ^ n1076 ;
  assign n10439 = n5258 & ~n10112 ;
  assign n10440 = n10439 ^ n2942 ^ n631 ;
  assign n10447 = n2981 ^ n907 ^ x62 ;
  assign n10448 = n294 & ~n10447 ;
  assign n10449 = n6812 & n10448 ;
  assign n10441 = n5262 ^ n2892 ^ n445 ;
  assign n10442 = n10441 ^ n5912 ^ 1'b0 ;
  assign n10443 = n5576 ^ n4279 ^ n398 ;
  assign n10444 = ( ~n2805 & n10442 ) | ( ~n2805 & n10443 ) | ( n10442 & n10443 ) ;
  assign n10445 = n10444 ^ n3740 ^ n3026 ;
  assign n10446 = ( n2948 & ~n5414 ) | ( n2948 & n10445 ) | ( ~n5414 & n10445 ) ;
  assign n10450 = n10449 ^ n10446 ^ n1794 ;
  assign n10451 = n7833 ^ n4944 ^ 1'b0 ;
  assign n10459 = n9964 ^ n2481 ^ 1'b0 ;
  assign n10457 = ( ~n260 & n1362 ) | ( ~n260 & n4235 ) | ( n1362 & n4235 ) ;
  assign n10458 = ( ~n827 & n6310 ) | ( ~n827 & n10457 ) | ( n6310 & n10457 ) ;
  assign n10452 = ( n1165 & n2208 ) | ( n1165 & n2797 ) | ( n2208 & n2797 ) ;
  assign n10453 = ~n5162 & n10452 ;
  assign n10454 = n10037 & n10453 ;
  assign n10455 = n10454 ^ n4604 ^ n4004 ;
  assign n10456 = n10455 ^ n8615 ^ n5533 ;
  assign n10460 = n10459 ^ n10458 ^ n10456 ;
  assign n10461 = ( n2814 & n5472 ) | ( n2814 & n8080 ) | ( n5472 & n8080 ) ;
  assign n10462 = ( n5530 & n7229 ) | ( n5530 & ~n10461 ) | ( n7229 & ~n10461 ) ;
  assign n10465 = n2314 ^ n1849 ^ n1592 ;
  assign n10466 = ( ~n1994 & n8906 ) | ( ~n1994 & n10465 ) | ( n8906 & n10465 ) ;
  assign n10467 = ( ~n6194 & n6903 ) | ( ~n6194 & n10466 ) | ( n6903 & n10466 ) ;
  assign n10468 = n2234 | n10467 ;
  assign n10463 = n4925 ^ n3438 ^ n2462 ;
  assign n10464 = ( n8415 & ~n10002 ) | ( n8415 & n10463 ) | ( ~n10002 & n10463 ) ;
  assign n10469 = n10468 ^ n10464 ^ n5551 ;
  assign n10470 = n10469 ^ n9152 ^ n5055 ;
  assign n10472 = n2527 ^ n1270 ^ n627 ;
  assign n10473 = n10472 ^ n3782 ^ x2 ;
  assign n10474 = ( n1391 & n5210 ) | ( n1391 & n10473 ) | ( n5210 & n10473 ) ;
  assign n10471 = n10005 ^ n9661 ^ n6135 ;
  assign n10475 = n10474 ^ n10471 ^ 1'b0 ;
  assign n10477 = ~n1749 & n2751 ;
  assign n10478 = n2651 & n10477 ;
  assign n10479 = ( n2149 & n4370 ) | ( n2149 & n10478 ) | ( n4370 & n10478 ) ;
  assign n10476 = ( n4501 & n5731 ) | ( n4501 & n10181 ) | ( n5731 & n10181 ) ;
  assign n10480 = n10479 ^ n10476 ^ n303 ;
  assign n10482 = ( n3257 & n3984 ) | ( n3257 & ~n6076 ) | ( n3984 & ~n6076 ) ;
  assign n10483 = ~n5535 & n8601 ;
  assign n10484 = n10483 ^ n9805 ^ 1'b0 ;
  assign n10485 = ( n2765 & n10482 ) | ( n2765 & n10484 ) | ( n10482 & n10484 ) ;
  assign n10481 = n4150 ^ n3954 ^ n165 ;
  assign n10486 = n10485 ^ n10481 ^ 1'b0 ;
  assign n10487 = n3633 & ~n10486 ;
  assign n10488 = n7905 ^ n7595 ^ n2594 ;
  assign n10489 = n10488 ^ n10060 ^ n5083 ;
  assign n10490 = ( n10480 & n10487 ) | ( n10480 & n10489 ) | ( n10487 & n10489 ) ;
  assign n10495 = n5429 ^ n4471 ^ n293 ;
  assign n10491 = ( n2014 & ~n2409 ) | ( n2014 & n6615 ) | ( ~n2409 & n6615 ) ;
  assign n10492 = n8256 ^ n5599 ^ n3289 ;
  assign n10493 = ( n868 & n1871 ) | ( n868 & ~n10492 ) | ( n1871 & ~n10492 ) ;
  assign n10494 = n10491 | n10493 ;
  assign n10496 = n10495 ^ n10494 ^ 1'b0 ;
  assign n10497 = n3414 | n10496 ;
  assign n10498 = n10497 ^ n7251 ^ 1'b0 ;
  assign n10499 = n9022 ^ n3895 ^ n1442 ;
  assign n10500 = ( n502 & ~n4188 ) | ( n502 & n10396 ) | ( ~n4188 & n10396 ) ;
  assign n10501 = ( n8323 & n9981 ) | ( n8323 & ~n10500 ) | ( n9981 & ~n10500 ) ;
  assign n10502 = n3937 ^ n439 ^ 1'b0 ;
  assign n10514 = n1494 & ~n6354 ;
  assign n10515 = ( n2240 & n5233 ) | ( n2240 & n9482 ) | ( n5233 & n9482 ) ;
  assign n10516 = ( n1522 & n10514 ) | ( n1522 & ~n10515 ) | ( n10514 & ~n10515 ) ;
  assign n10505 = ( n1517 & n1971 ) | ( n1517 & n3867 ) | ( n1971 & n3867 ) ;
  assign n10506 = n10505 ^ n7325 ^ n6292 ;
  assign n10507 = n9257 ^ n4078 ^ 1'b0 ;
  assign n10508 = n793 & n10507 ;
  assign n10511 = n4650 ^ n2525 ^ x14 ;
  assign n10509 = ~n2029 & n9846 ;
  assign n10510 = n2425 & n10509 ;
  assign n10512 = n10511 ^ n10510 ^ n8044 ;
  assign n10513 = ( n10506 & n10508 ) | ( n10506 & n10512 ) | ( n10508 & n10512 ) ;
  assign n10504 = ( n751 & n2383 ) | ( n751 & ~n4387 ) | ( n2383 & ~n4387 ) ;
  assign n10517 = n10516 ^ n10513 ^ n10504 ;
  assign n10503 = n606 ^ n260 ^ 1'b0 ;
  assign n10518 = n10517 ^ n10503 ^ n563 ;
  assign n10522 = n5276 ^ n1482 ^ n329 ;
  assign n10523 = n10522 ^ n9247 ^ n6806 ;
  assign n10524 = n10523 ^ n7153 ^ n681 ;
  assign n10521 = ( n1137 & n1586 ) | ( n1137 & ~n5784 ) | ( n1586 & ~n5784 ) ;
  assign n10519 = n978 ^ x4 ^ 1'b0 ;
  assign n10520 = ( n1366 & ~n3853 ) | ( n1366 & n10519 ) | ( ~n3853 & n10519 ) ;
  assign n10525 = n10524 ^ n10521 ^ n10520 ;
  assign n10526 = n1635 | n9462 ;
  assign n10527 = n5423 & ~n10526 ;
  assign n10528 = ( n3984 & n8187 ) | ( n3984 & ~n10527 ) | ( n8187 & ~n10527 ) ;
  assign n10529 = ( n309 & n2149 ) | ( n309 & n4355 ) | ( n2149 & n4355 ) ;
  assign n10530 = ( n201 & n10380 ) | ( n201 & ~n10529 ) | ( n10380 & ~n10529 ) ;
  assign n10534 = ( ~n3175 & n4152 ) | ( ~n3175 & n4998 ) | ( n4152 & n4998 ) ;
  assign n10531 = ~n2856 & n7642 ;
  assign n10532 = n10531 ^ n6163 ^ 1'b0 ;
  assign n10533 = n7836 | n10532 ;
  assign n10535 = n10534 ^ n10533 ^ 1'b0 ;
  assign n10536 = n2060 & ~n7365 ;
  assign n10537 = n10536 ^ n9810 ^ 1'b0 ;
  assign n10538 = ~n5359 & n10537 ;
  assign n10539 = n10538 ^ n7733 ^ 1'b0 ;
  assign n10540 = n7686 ^ n1494 ^ 1'b0 ;
  assign n10541 = ~n5484 & n10540 ;
  assign n10542 = ( n3271 & n10539 ) | ( n3271 & ~n10541 ) | ( n10539 & ~n10541 ) ;
  assign n10545 = ( n834 & n921 ) | ( n834 & ~n981 ) | ( n921 & ~n981 ) ;
  assign n10546 = ( n6583 & n10326 ) | ( n6583 & ~n10545 ) | ( n10326 & ~n10545 ) ;
  assign n10543 = n222 & n1590 ;
  assign n10544 = n10543 ^ n8667 ^ 1'b0 ;
  assign n10547 = n10546 ^ n10544 ^ n5096 ;
  assign n10548 = ~n966 & n4178 ;
  assign n10549 = ~n8783 & n10548 ;
  assign n10550 = ( n157 & ~n688 ) | ( n157 & n2352 ) | ( ~n688 & n2352 ) ;
  assign n10551 = ( n3713 & ~n5733 ) | ( n3713 & n8026 ) | ( ~n5733 & n8026 ) ;
  assign n10552 = n10223 & ~n10551 ;
  assign n10553 = ( ~n1789 & n5520 ) | ( ~n1789 & n10552 ) | ( n5520 & n10552 ) ;
  assign n10554 = ( n3018 & ~n10550 ) | ( n3018 & n10553 ) | ( ~n10550 & n10553 ) ;
  assign n10555 = ~n10549 & n10554 ;
  assign n10556 = ~n3893 & n4757 ;
  assign n10557 = ( n592 & n1923 ) | ( n592 & ~n5131 ) | ( n1923 & ~n5131 ) ;
  assign n10558 = n7586 ^ n6072 ^ n2850 ;
  assign n10559 = n9482 | n10558 ;
  assign n10560 = n10559 ^ n8142 ^ 1'b0 ;
  assign n10561 = ( n3966 & n6833 ) | ( n3966 & ~n9337 ) | ( n6833 & ~n9337 ) ;
  assign n10562 = n659 & n10561 ;
  assign n10563 = ( n10557 & n10560 ) | ( n10557 & n10562 ) | ( n10560 & n10562 ) ;
  assign n10564 = n5912 ^ n5101 ^ n3788 ;
  assign n10565 = n10564 ^ n4771 ^ 1'b0 ;
  assign n10572 = ( ~n8447 & n9146 ) | ( ~n8447 & n10052 ) | ( n9146 & n10052 ) ;
  assign n10573 = n10572 ^ n5083 ^ n4486 ;
  assign n10570 = n2938 ^ n2890 ^ n983 ;
  assign n10569 = ( ~n342 & n525 ) | ( ~n342 & n7777 ) | ( n525 & n7777 ) ;
  assign n10571 = n10570 ^ n10569 ^ n4335 ;
  assign n10566 = n5629 ^ n2023 ^ n870 ;
  assign n10567 = ( n4028 & ~n7054 ) | ( n4028 & n10566 ) | ( ~n7054 & n10566 ) ;
  assign n10568 = n10567 ^ n8095 ^ n462 ;
  assign n10574 = n10573 ^ n10571 ^ n10568 ;
  assign n10577 = n4021 & ~n4298 ;
  assign n10578 = ( n2303 & n9877 ) | ( n2303 & n10577 ) | ( n9877 & n10577 ) ;
  assign n10575 = ~n456 & n844 ;
  assign n10576 = n10575 ^ n1004 ^ 1'b0 ;
  assign n10579 = n10578 ^ n10576 ^ n8606 ;
  assign n10583 = ( n2427 & ~n6231 ) | ( n2427 & n8134 ) | ( ~n6231 & n8134 ) ;
  assign n10580 = n4512 & ~n4964 ;
  assign n10581 = n10580 ^ n6332 ^ n322 ;
  assign n10582 = ~n2031 & n10581 ;
  assign n10584 = n10583 ^ n10582 ^ n639 ;
  assign n10586 = ( n511 & n3683 ) | ( n511 & n7893 ) | ( n3683 & n7893 ) ;
  assign n10585 = n4508 ^ n4090 ^ n2547 ;
  assign n10587 = n10586 ^ n10585 ^ n1351 ;
  assign n10588 = n6666 ^ n6446 ^ n4587 ;
  assign n10591 = ( n3837 & n4744 ) | ( n3837 & ~n9786 ) | ( n4744 & ~n9786 ) ;
  assign n10589 = n8162 ^ n1820 ^ 1'b0 ;
  assign n10590 = ~n834 & n10589 ;
  assign n10592 = n10591 ^ n10590 ^ n4457 ;
  assign n10593 = n10588 & n10592 ;
  assign n10594 = ~n10587 & n10593 ;
  assign n10601 = ( n1454 & n2786 ) | ( n1454 & n5782 ) | ( n2786 & n5782 ) ;
  assign n10595 = ( n6454 & ~n7905 ) | ( n6454 & n10032 ) | ( ~n7905 & n10032 ) ;
  assign n10596 = n10595 ^ n5572 ^ n1556 ;
  assign n10597 = ( n4066 & n7115 ) | ( n4066 & ~n10596 ) | ( n7115 & ~n10596 ) ;
  assign n10598 = n3828 | n6935 ;
  assign n10599 = n10598 ^ n6199 ^ n309 ;
  assign n10600 = ( ~n6209 & n10597 ) | ( ~n6209 & n10599 ) | ( n10597 & n10599 ) ;
  assign n10602 = n10601 ^ n10600 ^ 1'b0 ;
  assign n10603 = n9014 ^ n6140 ^ 1'b0 ;
  assign n10604 = n3136 ^ n1371 ^ n1240 ;
  assign n10605 = n6715 | n10604 ;
  assign n10606 = n5213 | n10605 ;
  assign n10607 = n4890 & n10606 ;
  assign n10608 = n10607 ^ n10361 ^ 1'b0 ;
  assign n10609 = n5545 ^ n2850 ^ n138 ;
  assign n10610 = n10609 ^ n700 ^ n522 ;
  assign n10611 = ( ~x90 & n4994 ) | ( ~x90 & n10610 ) | ( n4994 & n10610 ) ;
  assign n10612 = n8407 ^ n6669 ^ 1'b0 ;
  assign n10613 = ( n332 & ~n1666 ) | ( n332 & n3173 ) | ( ~n1666 & n3173 ) ;
  assign n10614 = n10612 & n10613 ;
  assign n10615 = n2420 ^ n1802 ^ n993 ;
  assign n10616 = n10615 ^ n8149 ^ n3181 ;
  assign n10617 = n10616 ^ n8685 ^ 1'b0 ;
  assign n10624 = n919 | n2365 ;
  assign n10623 = n7032 ^ n2869 ^ n166 ;
  assign n10618 = n8509 ^ n7342 ^ n4132 ;
  assign n10619 = n9480 ^ n1732 ^ n1444 ;
  assign n10620 = ( n5381 & n8207 ) | ( n5381 & ~n10619 ) | ( n8207 & ~n10619 ) ;
  assign n10621 = n5285 & ~n10620 ;
  assign n10622 = ( ~n4443 & n10618 ) | ( ~n4443 & n10621 ) | ( n10618 & n10621 ) ;
  assign n10625 = n10624 ^ n10623 ^ n10622 ;
  assign n10626 = n1801 ^ n1555 ^ x21 ;
  assign n10627 = ( n2576 & n5658 ) | ( n2576 & n9882 ) | ( n5658 & n9882 ) ;
  assign n10628 = n10627 ^ n8206 ^ x6 ;
  assign n10629 = ( n1339 & n7172 ) | ( n1339 & n10628 ) | ( n7172 & n10628 ) ;
  assign n10630 = ( n512 & n2823 ) | ( n512 & ~n3716 ) | ( n2823 & ~n3716 ) ;
  assign n10631 = n10630 ^ n3709 ^ 1'b0 ;
  assign n10632 = ( n10626 & n10629 ) | ( n10626 & ~n10631 ) | ( n10629 & ~n10631 ) ;
  assign n10633 = ( n858 & n6041 ) | ( n858 & n10632 ) | ( n6041 & n10632 ) ;
  assign n10634 = n4897 & n7113 ;
  assign n10635 = n1940 ^ n1921 ^ 1'b0 ;
  assign n10636 = ( n5327 & n5535 ) | ( n5327 & n10635 ) | ( n5535 & n10635 ) ;
  assign n10637 = n10636 ^ n6957 ^ n6821 ;
  assign n10650 = n972 | n6098 ;
  assign n10648 = ~n1265 & n9376 ;
  assign n10649 = n10648 ^ n10136 ^ 1'b0 ;
  assign n10638 = n2648 & n6960 ;
  assign n10639 = n6446 & n10638 ;
  assign n10640 = ( ~n5727 & n10179 ) | ( ~n5727 & n10639 ) | ( n10179 & n10639 ) ;
  assign n10641 = n2042 | n2726 ;
  assign n10642 = n4840 & ~n10641 ;
  assign n10643 = ( n1840 & n8933 ) | ( n1840 & n10642 ) | ( n8933 & n10642 ) ;
  assign n10644 = ( ~x50 & n383 ) | ( ~x50 & n8245 ) | ( n383 & n8245 ) ;
  assign n10645 = ( n4195 & n7174 ) | ( n4195 & n10644 ) | ( n7174 & n10644 ) ;
  assign n10646 = ~n10643 & n10645 ;
  assign n10647 = n10640 & n10646 ;
  assign n10651 = n10650 ^ n10649 ^ n10647 ;
  assign n10663 = ( n265 & ~n1444 ) | ( n265 & n2556 ) | ( ~n1444 & n2556 ) ;
  assign n10662 = ( n1163 & n5211 ) | ( n1163 & n6872 ) | ( n5211 & n6872 ) ;
  assign n10664 = n10663 ^ n10662 ^ n7837 ;
  assign n10652 = n3908 | n5083 ;
  assign n10653 = ( ~n7341 & n8126 ) | ( ~n7341 & n10652 ) | ( n8126 & n10652 ) ;
  assign n10655 = n10598 ^ n8489 ^ n6335 ;
  assign n10654 = ( n256 & n3046 ) | ( n256 & n9873 ) | ( n3046 & n9873 ) ;
  assign n10656 = n10655 ^ n10654 ^ n2296 ;
  assign n10657 = n4036 & ~n8261 ;
  assign n10658 = ( ~n2943 & n10656 ) | ( ~n2943 & n10657 ) | ( n10656 & n10657 ) ;
  assign n10659 = n10658 ^ n9976 ^ n1372 ;
  assign n10660 = n10659 ^ n6668 ^ n5777 ;
  assign n10661 = n10653 & n10660 ;
  assign n10665 = n10664 ^ n10661 ^ 1'b0 ;
  assign n10666 = n10665 ^ n4739 ^ n167 ;
  assign n10667 = n4454 ^ n2427 ^ 1'b0 ;
  assign n10668 = ( ~n2590 & n7394 ) | ( ~n2590 & n10667 ) | ( n7394 & n10667 ) ;
  assign n10676 = n6767 ^ n4404 ^ n3640 ;
  assign n10677 = n1391 & ~n10676 ;
  assign n10674 = ( ~n2443 & n3147 ) | ( ~n2443 & n7792 ) | ( n3147 & n7792 ) ;
  assign n10669 = ( n1086 & n1215 ) | ( n1086 & ~n8650 ) | ( n1215 & ~n8650 ) ;
  assign n10670 = n5749 ^ n4326 ^ n3741 ;
  assign n10671 = n10670 ^ n7709 ^ n6985 ;
  assign n10672 = ( ~n1238 & n10669 ) | ( ~n1238 & n10671 ) | ( n10669 & n10671 ) ;
  assign n10673 = ( n1148 & n9434 ) | ( n1148 & n10672 ) | ( n9434 & n10672 ) ;
  assign n10675 = n10674 ^ n10673 ^ n5495 ;
  assign n10678 = n10677 ^ n10675 ^ n9373 ;
  assign n10679 = ( ~n280 & n10668 ) | ( ~n280 & n10678 ) | ( n10668 & n10678 ) ;
  assign n10680 = n837 | n9643 ;
  assign n10681 = ( n3570 & n7879 ) | ( n3570 & n10680 ) | ( n7879 & n10680 ) ;
  assign n10682 = n6435 ^ n4799 ^ n2907 ;
  assign n10683 = n10682 ^ n10393 ^ n2904 ;
  assign n10684 = ( n1174 & ~n10681 ) | ( n1174 & n10683 ) | ( ~n10681 & n10683 ) ;
  assign n10685 = n7568 ^ n5487 ^ n569 ;
  assign n10686 = ( ~n2432 & n6862 ) | ( ~n2432 & n10685 ) | ( n6862 & n10685 ) ;
  assign n10687 = n3334 & n3539 ;
  assign n10688 = n10686 & n10687 ;
  assign n10689 = ( ~n537 & n3605 ) | ( ~n537 & n7270 ) | ( n3605 & n7270 ) ;
  assign n10690 = n2851 | n10689 ;
  assign n10691 = n5353 & ~n10690 ;
  assign n10692 = ( n8499 & n9876 ) | ( n8499 & ~n10691 ) | ( n9876 & ~n10691 ) ;
  assign n10693 = ( ~n1335 & n10688 ) | ( ~n1335 & n10692 ) | ( n10688 & n10692 ) ;
  assign n10694 = n9860 ^ n8162 ^ 1'b0 ;
  assign n10695 = ( ~n1368 & n1753 ) | ( ~n1368 & n1905 ) | ( n1753 & n1905 ) ;
  assign n10696 = n10695 ^ n9851 ^ n2320 ;
  assign n10697 = n6530 ^ n6458 ^ n2021 ;
  assign n10698 = x95 & ~n557 ;
  assign n10699 = n5467 ^ n5441 ^ n5194 ;
  assign n10700 = n10699 ^ n6770 ^ n3891 ;
  assign n10701 = n10698 | n10700 ;
  assign n10702 = n9646 & ~n10701 ;
  assign n10703 = ( n10219 & n10697 ) | ( n10219 & n10702 ) | ( n10697 & n10702 ) ;
  assign n10704 = n4342 ^ n2336 ^ n214 ;
  assign n10705 = ( n1095 & ~n1512 ) | ( n1095 & n10704 ) | ( ~n1512 & n10704 ) ;
  assign n10706 = n9847 ^ n6256 ^ 1'b0 ;
  assign n10707 = ( ~n3827 & n3976 ) | ( ~n3827 & n10706 ) | ( n3976 & n10706 ) ;
  assign n10708 = ( ~n1365 & n7196 ) | ( ~n1365 & n10447 ) | ( n7196 & n10447 ) ;
  assign n10709 = n5024 & ~n6643 ;
  assign n10710 = n10709 ^ n1720 ^ 1'b0 ;
  assign n10711 = n3529 ^ n1455 ^ 1'b0 ;
  assign n10712 = n10626 | n10711 ;
  assign n10713 = n557 & n10712 ;
  assign n10715 = n4030 & n4725 ;
  assign n10716 = n4413 & n10715 ;
  assign n10714 = ( n2469 & n2965 ) | ( n2469 & n3232 ) | ( n2965 & n3232 ) ;
  assign n10717 = n10716 ^ n10714 ^ 1'b0 ;
  assign n10718 = ( n10710 & ~n10713 ) | ( n10710 & n10717 ) | ( ~n10713 & n10717 ) ;
  assign n10719 = ( ~n6242 & n10708 ) | ( ~n6242 & n10718 ) | ( n10708 & n10718 ) ;
  assign n10720 = n3366 ^ n2572 ^ n1601 ;
  assign n10721 = n10720 ^ n630 ^ n484 ;
  assign n10722 = n10721 ^ n966 ^ n134 ;
  assign n10723 = n10622 ^ n9873 ^ n1109 ;
  assign n10724 = n10723 ^ n376 ^ 1'b0 ;
  assign n10725 = n7784 ^ n2238 ^ 1'b0 ;
  assign n10726 = ( n239 & ~n1625 ) | ( n239 & n1735 ) | ( ~n1625 & n1735 ) ;
  assign n10727 = n930 ^ n816 ^ 1'b0 ;
  assign n10728 = ~n10726 & n10727 ;
  assign n10729 = n10728 ^ n9602 ^ n2965 ;
  assign n10730 = ( n1121 & n10725 ) | ( n1121 & ~n10729 ) | ( n10725 & ~n10729 ) ;
  assign n10731 = n1010 & n1410 ;
  assign n10732 = n10731 ^ n3270 ^ 1'b0 ;
  assign n10733 = ( n644 & n1824 ) | ( n644 & ~n2000 ) | ( n1824 & ~n2000 ) ;
  assign n10735 = ( n3311 & ~n6592 ) | ( n3311 & n7531 ) | ( ~n6592 & n7531 ) ;
  assign n10736 = n10735 ^ n3441 ^ n2816 ;
  assign n10734 = n10721 ^ n4655 ^ n225 ;
  assign n10737 = n10736 ^ n10734 ^ n7050 ;
  assign n10738 = n10737 ^ n6806 ^ x74 ;
  assign n10739 = n9662 ^ n7528 ^ 1'b0 ;
  assign n10753 = n5553 ^ n4439 ^ n427 ;
  assign n10750 = ( ~n3797 & n5639 ) | ( ~n3797 & n6434 ) | ( n5639 & n6434 ) ;
  assign n10749 = n4943 ^ n1696 ^ n1487 ;
  assign n10751 = n10750 ^ n10749 ^ n2147 ;
  assign n10740 = ( n678 & ~n1500 ) | ( n678 & n3586 ) | ( ~n1500 & n3586 ) ;
  assign n10741 = ( n8740 & ~n10178 ) | ( n8740 & n10740 ) | ( ~n10178 & n10740 ) ;
  assign n10742 = n2849 ^ n2367 ^ n995 ;
  assign n10743 = n10742 ^ n4706 ^ n4513 ;
  assign n10744 = n5802 ^ n748 ^ n211 ;
  assign n10745 = ( n574 & ~n7531 ) | ( n574 & n10744 ) | ( ~n7531 & n10744 ) ;
  assign n10746 = ( n10741 & ~n10743 ) | ( n10741 & n10745 ) | ( ~n10743 & n10745 ) ;
  assign n10747 = n5058 ^ n2700 ^ n1323 ;
  assign n10748 = ( n5658 & n10746 ) | ( n5658 & n10747 ) | ( n10746 & n10747 ) ;
  assign n10752 = n10751 ^ n10748 ^ n6637 ;
  assign n10754 = n10753 ^ n10752 ^ n746 ;
  assign n10755 = ( n1964 & ~n10739 ) | ( n1964 & n10754 ) | ( ~n10739 & n10754 ) ;
  assign n10756 = n10755 ^ n10067 ^ n1401 ;
  assign n10757 = ( ~n3609 & n10738 ) | ( ~n3609 & n10756 ) | ( n10738 & n10756 ) ;
  assign n10758 = n5796 ^ n4281 ^ n4076 ;
  assign n10770 = n1348 ^ n240 ^ 1'b0 ;
  assign n10763 = ~n767 & n8639 ;
  assign n10764 = n10763 ^ n4962 ^ 1'b0 ;
  assign n10762 = n484 | n3095 ;
  assign n10765 = n10764 ^ n10762 ^ 1'b0 ;
  assign n10766 = ( n1620 & n3575 ) | ( n1620 & ~n5911 ) | ( n3575 & ~n5911 ) ;
  assign n10767 = ( n5496 & n6102 ) | ( n5496 & ~n8687 ) | ( n6102 & ~n8687 ) ;
  assign n10768 = n10766 | n10767 ;
  assign n10769 = n10765 & ~n10768 ;
  assign n10759 = ( n4361 & ~n4963 ) | ( n4361 & n7870 ) | ( ~n4963 & n7870 ) ;
  assign n10760 = ( ~n528 & n10182 ) | ( ~n528 & n10759 ) | ( n10182 & n10759 ) ;
  assign n10761 = n10760 ^ n6133 ^ n3889 ;
  assign n10771 = n10770 ^ n10769 ^ n10761 ;
  assign n10772 = ~n812 & n834 ;
  assign n10773 = ( ~n1817 & n8620 ) | ( ~n1817 & n10772 ) | ( n8620 & n10772 ) ;
  assign n10774 = ( n1614 & n8510 ) | ( n1614 & n10773 ) | ( n8510 & n10773 ) ;
  assign n10775 = n10774 ^ n9817 ^ n3242 ;
  assign n10776 = n10775 ^ n5559 ^ n2298 ;
  assign n10777 = n10776 ^ n3930 ^ n3443 ;
  assign n10779 = ( ~n2674 & n10207 ) | ( ~n2674 & n10557 ) | ( n10207 & n10557 ) ;
  assign n10778 = ( n514 & n5389 ) | ( n514 & n5672 ) | ( n5389 & n5672 ) ;
  assign n10780 = n10779 ^ n10778 ^ n6888 ;
  assign n10781 = ( n4362 & n4458 ) | ( n4362 & n10780 ) | ( n4458 & n10780 ) ;
  assign n10782 = ( n731 & ~n6804 ) | ( n731 & n8371 ) | ( ~n6804 & n8371 ) ;
  assign n10783 = n7107 ^ n3187 ^ 1'b0 ;
  assign n10784 = ( n4201 & ~n5754 ) | ( n4201 & n10783 ) | ( ~n5754 & n10783 ) ;
  assign n10788 = n3665 | n9224 ;
  assign n10787 = n9016 ^ n5743 ^ n955 ;
  assign n10785 = n7822 ^ n760 ^ 1'b0 ;
  assign n10786 = ( n4577 & ~n10078 ) | ( n4577 & n10785 ) | ( ~n10078 & n10785 ) ;
  assign n10789 = n10788 ^ n10787 ^ n10786 ;
  assign n10790 = n9350 ^ n8836 ^ n7887 ;
  assign n10791 = n8503 ^ n5269 ^ n4556 ;
  assign n10792 = ( n530 & ~n7924 ) | ( n530 & n10791 ) | ( ~n7924 & n10791 ) ;
  assign n10793 = ( n1982 & ~n6329 ) | ( n1982 & n8247 ) | ( ~n6329 & n8247 ) ;
  assign n10794 = ( n8641 & n10792 ) | ( n8641 & ~n10793 ) | ( n10792 & ~n10793 ) ;
  assign n10795 = ( ~n3359 & n3837 ) | ( ~n3359 & n6299 ) | ( n3837 & n6299 ) ;
  assign n10796 = n3887 & ~n10795 ;
  assign n10797 = ( n1590 & ~n3037 ) | ( n1590 & n5635 ) | ( ~n3037 & n5635 ) ;
  assign n10798 = n10797 ^ n5462 ^ n3488 ;
  assign n10799 = ( n2714 & n3431 ) | ( n2714 & n10798 ) | ( n3431 & n10798 ) ;
  assign n10800 = n3519 ^ n2762 ^ n1870 ;
  assign n10801 = n10800 ^ n3367 ^ 1'b0 ;
  assign n10802 = n7903 & n10801 ;
  assign n10803 = n1639 ^ n1335 ^ n632 ;
  assign n10806 = ( n512 & n1553 ) | ( n512 & n4697 ) | ( n1553 & n4697 ) ;
  assign n10807 = ( n5129 & n6168 ) | ( n5129 & n10806 ) | ( n6168 & n10806 ) ;
  assign n10804 = n8815 ^ n3246 ^ 1'b0 ;
  assign n10805 = ~n4416 & n10804 ;
  assign n10808 = n10807 ^ n10805 ^ n6673 ;
  assign n10809 = n6170 ^ n2071 ^ 1'b0 ;
  assign n10810 = n10809 ^ n9249 ^ 1'b0 ;
  assign n10811 = ( n2483 & n4793 ) | ( n2483 & n9061 ) | ( n4793 & n9061 ) ;
  assign n10812 = n10811 ^ n8412 ^ n6598 ;
  assign n10813 = ( ~n1764 & n2662 ) | ( ~n1764 & n10812 ) | ( n2662 & n10812 ) ;
  assign n10814 = ( ~n512 & n2596 ) | ( ~n512 & n8580 ) | ( n2596 & n8580 ) ;
  assign n10815 = n7729 ^ n5431 ^ n449 ;
  assign n10817 = ( ~n1690 & n2311 ) | ( ~n1690 & n4533 ) | ( n2311 & n4533 ) ;
  assign n10818 = n10817 ^ n7180 ^ n169 ;
  assign n10816 = n9510 ^ n7481 ^ n1086 ;
  assign n10819 = n10818 ^ n10816 ^ n2458 ;
  assign n10820 = ( n2149 & ~n10815 ) | ( n2149 & n10819 ) | ( ~n10815 & n10819 ) ;
  assign n10821 = ( ~n7543 & n10814 ) | ( ~n7543 & n10820 ) | ( n10814 & n10820 ) ;
  assign n10822 = n10821 ^ n6227 ^ n3682 ;
  assign n10823 = n3885 | n4546 ;
  assign n10824 = ( n1230 & n10516 ) | ( n1230 & ~n10823 ) | ( n10516 & ~n10823 ) ;
  assign n10825 = n10824 ^ n5014 ^ n3152 ;
  assign n10826 = n10825 ^ n10247 ^ n7815 ;
  assign n10827 = ~n10822 & n10826 ;
  assign n10828 = n7963 ^ n2171 ^ n2015 ;
  assign n10829 = n10630 & ~n10828 ;
  assign n10830 = n10600 ^ n2773 ^ 1'b0 ;
  assign n10831 = ~n10829 & n10830 ;
  assign n10832 = ( ~n5197 & n9076 ) | ( ~n5197 & n10831 ) | ( n9076 & n10831 ) ;
  assign n10833 = ( n856 & n6733 ) | ( n856 & n7136 ) | ( n6733 & n7136 ) ;
  assign n10834 = ( n8290 & n8877 ) | ( n8290 & n10833 ) | ( n8877 & n10833 ) ;
  assign n10835 = n10834 ^ n9933 ^ n2173 ;
  assign n10836 = n2874 ^ n1016 ^ n816 ;
  assign n10837 = n10836 ^ n10487 ^ n2082 ;
  assign n10845 = ( n1324 & n1375 ) | ( n1324 & n2274 ) | ( n1375 & n2274 ) ;
  assign n10840 = ~n2175 & n4566 ;
  assign n10841 = n5997 & n10840 ;
  assign n10838 = n311 & n3257 ;
  assign n10839 = n10838 ^ n5235 ^ 1'b0 ;
  assign n10842 = n10841 ^ n10839 ^ n5476 ;
  assign n10843 = ( n3616 & n6597 ) | ( n3616 & ~n10842 ) | ( n6597 & ~n10842 ) ;
  assign n10844 = n10843 ^ n4075 ^ n253 ;
  assign n10846 = n10845 ^ n10844 ^ n4467 ;
  assign n10847 = n6466 ^ n1275 ^ 1'b0 ;
  assign n10848 = ~n4943 & n10847 ;
  assign n10849 = ( n3135 & n8315 ) | ( n3135 & ~n9977 ) | ( n8315 & ~n9977 ) ;
  assign n10850 = ( n5072 & n10848 ) | ( n5072 & ~n10849 ) | ( n10848 & ~n10849 ) ;
  assign n10851 = ( n3973 & n8317 ) | ( n3973 & ~n9861 ) | ( n8317 & ~n9861 ) ;
  assign n10852 = n5562 ^ n398 ^ 1'b0 ;
  assign n10853 = n10852 ^ n5188 ^ n4400 ;
  assign n10854 = ( ~n171 & n3211 ) | ( ~n171 & n4830 ) | ( n3211 & n4830 ) ;
  assign n10855 = n10395 ^ n6556 ^ n3816 ;
  assign n10856 = ~n6609 & n10855 ;
  assign n10857 = ~n4979 & n10856 ;
  assign n10858 = n10854 & ~n10857 ;
  assign n10859 = n9101 ^ n4028 ^ n1768 ;
  assign n10860 = n10859 ^ n5548 ^ n4259 ;
  assign n10861 = n10860 ^ n5270 ^ n1309 ;
  assign n10862 = n3898 | n10861 ;
  assign n10863 = n3707 ^ n1128 ^ 1'b0 ;
  assign n10864 = ( ~n1715 & n2943 ) | ( ~n1715 & n10863 ) | ( n2943 & n10863 ) ;
  assign n10865 = ( ~n1355 & n3617 ) | ( ~n1355 & n6719 ) | ( n3617 & n6719 ) ;
  assign n10866 = ( ~n4399 & n9673 ) | ( ~n4399 & n10865 ) | ( n9673 & n10865 ) ;
  assign n10867 = n10235 ^ n8878 ^ n3905 ;
  assign n10868 = n6213 ^ n5703 ^ n376 ;
  assign n10869 = ( ~n4891 & n10867 ) | ( ~n4891 & n10868 ) | ( n10867 & n10868 ) ;
  assign n10872 = n1546 & n2465 ;
  assign n10873 = n10872 ^ n2476 ^ 1'b0 ;
  assign n10874 = n10873 ^ n6136 ^ n5830 ;
  assign n10875 = ( n2970 & ~n4180 ) | ( n2970 & n10874 ) | ( ~n4180 & n10874 ) ;
  assign n10870 = ( n5677 & n6536 ) | ( n5677 & ~n8877 ) | ( n6536 & ~n8877 ) ;
  assign n10871 = ( n5544 & n9089 ) | ( n5544 & n10870 ) | ( n9089 & n10870 ) ;
  assign n10876 = n10875 ^ n10871 ^ n339 ;
  assign n10884 = n4863 ^ n227 ^ 1'b0 ;
  assign n10877 = n5930 ^ n4880 ^ n188 ;
  assign n10878 = ( n946 & n7063 ) | ( n946 & n10877 ) | ( n7063 & n10877 ) ;
  assign n10879 = n8757 ^ n3376 ^ n1258 ;
  assign n10880 = n4175 ^ n3381 ^ 1'b0 ;
  assign n10881 = ( n2855 & n4230 ) | ( n2855 & ~n10880 ) | ( n4230 & ~n10880 ) ;
  assign n10882 = ( n5731 & n10718 ) | ( n5731 & n10881 ) | ( n10718 & n10881 ) ;
  assign n10883 = ( ~n10878 & n10879 ) | ( ~n10878 & n10882 ) | ( n10879 & n10882 ) ;
  assign n10885 = n10884 ^ n10883 ^ n1707 ;
  assign n10886 = n2965 ^ n2607 ^ n666 ;
  assign n10887 = n10886 ^ n3103 ^ n1946 ;
  assign n10888 = n10887 ^ n6837 ^ 1'b0 ;
  assign n10889 = ~n3764 & n10888 ;
  assign n10890 = ( n3241 & ~n3742 ) | ( n3241 & n10889 ) | ( ~n3742 & n10889 ) ;
  assign n10891 = ~n2763 & n10890 ;
  assign n10892 = n10891 ^ n2008 ^ 1'b0 ;
  assign n10893 = n4983 & n6436 ;
  assign n10894 = n10893 ^ n9555 ^ n5274 ;
  assign n10895 = n10894 ^ n852 ^ 1'b0 ;
  assign n10896 = ( n9487 & n10474 ) | ( n9487 & ~n10895 ) | ( n10474 & ~n10895 ) ;
  assign n10897 = ( n297 & n1037 ) | ( n297 & n7862 ) | ( n1037 & n7862 ) ;
  assign n10898 = ( n8165 & n10896 ) | ( n8165 & n10897 ) | ( n10896 & n10897 ) ;
  assign n10899 = ( n898 & ~n9346 ) | ( n898 & n9587 ) | ( ~n9346 & n9587 ) ;
  assign n10900 = ~n1277 & n2875 ;
  assign n10901 = n10900 ^ n2609 ^ 1'b0 ;
  assign n10902 = ( n683 & ~n5857 ) | ( n683 & n10901 ) | ( ~n5857 & n10901 ) ;
  assign n10903 = n10902 ^ n2540 ^ n757 ;
  assign n10905 = n3359 ^ n1590 ^ n734 ;
  assign n10904 = ( n3319 & ~n5908 ) | ( n3319 & n7966 ) | ( ~n5908 & n7966 ) ;
  assign n10906 = n10905 ^ n10904 ^ n9424 ;
  assign n10907 = ( n2343 & n10903 ) | ( n2343 & ~n10906 ) | ( n10903 & ~n10906 ) ;
  assign n10908 = ( ~n7810 & n8407 ) | ( ~n7810 & n8947 ) | ( n8407 & n8947 ) ;
  assign n10909 = n1254 & n10908 ;
  assign n10910 = ~n3621 & n10909 ;
  assign n10911 = ~n6228 & n9588 ;
  assign n10912 = n10910 & n10911 ;
  assign n10913 = n10912 ^ n4088 ^ n2773 ;
  assign n10914 = ( n2396 & n5168 ) | ( n2396 & ~n10913 ) | ( n5168 & ~n10913 ) ;
  assign n10915 = n2381 ^ n710 ^ n200 ;
  assign n10919 = ( n3351 & n6976 ) | ( n3351 & ~n9759 ) | ( n6976 & ~n9759 ) ;
  assign n10916 = ( n1812 & n2129 ) | ( n1812 & ~n9462 ) | ( n2129 & ~n9462 ) ;
  assign n10917 = ~n9046 & n10916 ;
  assign n10918 = n2379 & n10917 ;
  assign n10920 = n10919 ^ n10918 ^ x117 ;
  assign n10921 = n6068 & n7184 ;
  assign n10922 = n10921 ^ n9877 ^ n3060 ;
  assign n10929 = n890 | n7592 ;
  assign n10930 = ( ~n3939 & n6434 ) | ( ~n3939 & n10929 ) | ( n6434 & n10929 ) ;
  assign n10924 = n8696 ^ n2074 ^ x64 ;
  assign n10925 = n10924 ^ n4557 ^ n3939 ;
  assign n10923 = ( n2520 & ~n7401 ) | ( n2520 & n9118 ) | ( ~n7401 & n9118 ) ;
  assign n10926 = n10925 ^ n10923 ^ n2058 ;
  assign n10927 = ( n2120 & ~n6611 ) | ( n2120 & n8848 ) | ( ~n6611 & n8848 ) ;
  assign n10928 = ( n3329 & ~n10926 ) | ( n3329 & n10927 ) | ( ~n10926 & n10927 ) ;
  assign n10931 = n10930 ^ n10928 ^ n3578 ;
  assign n10932 = n10931 ^ n10132 ^ n9948 ;
  assign n10933 = ( ~n4174 & n10922 ) | ( ~n4174 & n10932 ) | ( n10922 & n10932 ) ;
  assign n10934 = ( n2288 & ~n4583 ) | ( n2288 & n8166 ) | ( ~n4583 & n8166 ) ;
  assign n10935 = ~n228 & n10934 ;
  assign n10940 = n5702 ^ n4087 ^ n2678 ;
  assign n10936 = ( n810 & n5512 ) | ( n810 & n6457 ) | ( n5512 & n6457 ) ;
  assign n10937 = n8903 ^ n5733 ^ n4532 ;
  assign n10938 = n10936 | n10937 ;
  assign n10939 = n10938 ^ n5444 ^ 1'b0 ;
  assign n10941 = n10940 ^ n10939 ^ n8323 ;
  assign n10944 = n10720 ^ n8232 ^ n2077 ;
  assign n10942 = n6534 ^ n1285 ^ n812 ;
  assign n10943 = ~n10572 & n10942 ;
  assign n10945 = n10944 ^ n10943 ^ n6947 ;
  assign n10946 = n4939 ^ n2757 ^ n870 ;
  assign n10947 = ( n405 & n1470 ) | ( n405 & ~n10946 ) | ( n1470 & ~n10946 ) ;
  assign n10948 = ~n803 & n10947 ;
  assign n10949 = n10945 & n10948 ;
  assign n10959 = n4914 ^ n2709 ^ n719 ;
  assign n10960 = n6559 ^ n2853 ^ 1'b0 ;
  assign n10961 = n703 & n10960 ;
  assign n10962 = ( ~n4730 & n10959 ) | ( ~n4730 & n10961 ) | ( n10959 & n10961 ) ;
  assign n10951 = ( ~n2094 & n5259 ) | ( ~n2094 & n5414 ) | ( n5259 & n5414 ) ;
  assign n10955 = n7851 ^ n1103 ^ 1'b0 ;
  assign n10952 = ( n974 & n3796 ) | ( n974 & n10877 ) | ( n3796 & n10877 ) ;
  assign n10953 = n6028 & ~n7074 ;
  assign n10954 = n10952 & n10953 ;
  assign n10956 = n10955 ^ n10954 ^ n5971 ;
  assign n10957 = ( n937 & n10951 ) | ( n937 & ~n10956 ) | ( n10951 & ~n10956 ) ;
  assign n10950 = n5894 ^ n5006 ^ n1840 ;
  assign n10958 = n10957 ^ n10950 ^ n487 ;
  assign n10963 = n10962 ^ n10958 ^ n1555 ;
  assign n10964 = ( n3551 & n4528 ) | ( n3551 & n10619 ) | ( n4528 & n10619 ) ;
  assign n10965 = n10964 ^ n9494 ^ n3415 ;
  assign n10966 = n5919 ^ n4479 ^ 1'b0 ;
  assign n10967 = n5515 & n10966 ;
  assign n10968 = n3373 & ~n3635 ;
  assign n10969 = n10968 ^ n5742 ^ n4422 ;
  assign n10970 = n5817 & ~n7196 ;
  assign n10971 = ( n3773 & ~n4390 ) | ( n3773 & n10970 ) | ( ~n4390 & n10970 ) ;
  assign n10972 = ( n9573 & n10969 ) | ( n9573 & n10971 ) | ( n10969 & n10971 ) ;
  assign n10973 = n189 & ~n3614 ;
  assign n10974 = n3908 | n7494 ;
  assign n10975 = n9995 & ~n10974 ;
  assign n10976 = n10975 ^ n8451 ^ n8344 ;
  assign n10977 = n6987 ^ n2868 ^ 1'b0 ;
  assign n10978 = n2488 & n10977 ;
  assign n10979 = n2381 | n7533 ;
  assign n10980 = n10979 ^ n10061 ^ 1'b0 ;
  assign n10981 = n8770 ^ n2516 ^ n1913 ;
  assign n10982 = ( n2928 & ~n3454 ) | ( n2928 & n10981 ) | ( ~n3454 & n10981 ) ;
  assign n10983 = ~n10449 & n10982 ;
  assign n10984 = n10983 ^ n6281 ^ 1'b0 ;
  assign n10985 = ~n1357 & n2207 ;
  assign n10986 = ~n10984 & n10985 ;
  assign n10987 = ( n3210 & ~n4368 ) | ( n3210 & n5009 ) | ( ~n4368 & n5009 ) ;
  assign n10988 = n4452 ^ n3434 ^ 1'b0 ;
  assign n10989 = n10988 ^ n10956 ^ n3984 ;
  assign n10990 = n2935 ^ n1727 ^ n1558 ;
  assign n10991 = n10990 ^ n8579 ^ n8352 ;
  assign n10993 = ( n2205 & ~n3083 ) | ( n2205 & n7971 ) | ( ~n3083 & n7971 ) ;
  assign n10992 = ( n157 & n4243 ) | ( n157 & n10576 ) | ( n4243 & n10576 ) ;
  assign n10994 = n10993 ^ n10992 ^ n6568 ;
  assign n10995 = n10991 & n10994 ;
  assign n10996 = n10995 ^ n9341 ^ 1'b0 ;
  assign n10997 = n551 & ~n9995 ;
  assign n10998 = ~n10996 & n10997 ;
  assign n10999 = n7388 ^ n1731 ^ n888 ;
  assign n11000 = ( ~n938 & n9090 ) | ( ~n938 & n10999 ) | ( n9090 & n10999 ) ;
  assign n11001 = ( ~n1048 & n3432 ) | ( ~n1048 & n11000 ) | ( n3432 & n11000 ) ;
  assign n11003 = n3822 ^ n2447 ^ 1'b0 ;
  assign n11004 = ( ~n474 & n653 ) | ( ~n474 & n11003 ) | ( n653 & n11003 ) ;
  assign n11005 = n11004 ^ n10750 ^ n5105 ;
  assign n11002 = n630 & n9360 ;
  assign n11006 = n11005 ^ n11002 ^ 1'b0 ;
  assign n11007 = n6705 ^ n1465 ^ n1157 ;
  assign n11008 = ( n1336 & n2296 ) | ( n1336 & ~n11007 ) | ( n2296 & ~n11007 ) ;
  assign n11009 = ( n2516 & n8902 ) | ( n2516 & ~n11008 ) | ( n8902 & ~n11008 ) ;
  assign n11010 = n10814 ^ n3627 ^ n1031 ;
  assign n11011 = n3086 ^ n2602 ^ n1429 ;
  assign n11012 = ( n896 & n2888 ) | ( n896 & ~n3777 ) | ( n2888 & ~n3777 ) ;
  assign n11013 = n11012 ^ n9975 ^ n4562 ;
  assign n11018 = ( ~n5865 & n6271 ) | ( ~n5865 & n9709 ) | ( n6271 & n9709 ) ;
  assign n11015 = n9140 ^ n6311 ^ n178 ;
  assign n11014 = ( n2435 & n2763 ) | ( n2435 & n4617 ) | ( n2763 & n4617 ) ;
  assign n11016 = n11015 ^ n11014 ^ n3429 ;
  assign n11017 = n4533 & n11016 ;
  assign n11019 = n11018 ^ n11017 ^ n4043 ;
  assign n11020 = n11019 ^ n2484 ^ n2396 ;
  assign n11021 = ( n874 & n5161 ) | ( n874 & n10174 ) | ( n5161 & n10174 ) ;
  assign n11022 = n9177 ^ n2936 ^ n754 ;
  assign n11023 = ~n4377 & n4683 ;
  assign n11024 = ~n4351 & n11023 ;
  assign n11025 = ( n7059 & n10481 ) | ( n7059 & n11024 ) | ( n10481 & n11024 ) ;
  assign n11026 = ( n2216 & n3363 ) | ( n2216 & n6201 ) | ( n3363 & n6201 ) ;
  assign n11027 = ( n2928 & ~n7359 ) | ( n2928 & n11026 ) | ( ~n7359 & n11026 ) ;
  assign n11028 = n11027 ^ n8252 ^ n4224 ;
  assign n11029 = n5477 ^ n1751 ^ n1333 ;
  assign n11030 = n980 & n10778 ;
  assign n11031 = n11029 & ~n11030 ;
  assign n11032 = n11031 ^ n580 ^ 1'b0 ;
  assign n11033 = ~n387 & n5541 ;
  assign n11034 = ~n11032 & n11033 ;
  assign n11035 = ( n1468 & ~n2011 ) | ( n1468 & n4505 ) | ( ~n2011 & n4505 ) ;
  assign n11036 = n9482 ^ n5233 ^ n1738 ;
  assign n11037 = n1838 & n5024 ;
  assign n11038 = n11037 ^ n6504 ^ n2447 ;
  assign n11039 = n5678 & ~n6114 ;
  assign n11040 = n4574 | n11039 ;
  assign n11041 = n689 | n11040 ;
  assign n11042 = ( n4002 & n11038 ) | ( n4002 & ~n11041 ) | ( n11038 & ~n11041 ) ;
  assign n11043 = ( n10797 & n11036 ) | ( n10797 & n11042 ) | ( n11036 & n11042 ) ;
  assign n11044 = n11043 ^ n9165 ^ 1'b0 ;
  assign n11045 = n11035 & ~n11044 ;
  assign n11054 = n11038 ^ n3429 ^ x34 ;
  assign n11055 = n4804 & n11054 ;
  assign n11052 = ( ~n2630 & n2998 ) | ( ~n2630 & n4387 ) | ( n2998 & n4387 ) ;
  assign n11048 = ( n2447 & n6220 ) | ( n2447 & n6322 ) | ( n6220 & n6322 ) ;
  assign n11049 = ( n6114 & n10595 ) | ( n6114 & ~n11048 ) | ( n10595 & ~n11048 ) ;
  assign n11050 = n9275 & ~n11049 ;
  assign n11047 = n3601 & n6425 ;
  assign n11046 = n9256 ^ n8933 ^ n4790 ;
  assign n11051 = n11050 ^ n11047 ^ n11046 ;
  assign n11053 = n11052 ^ n11051 ^ n5957 ;
  assign n11056 = n11055 ^ n11053 ^ n4161 ;
  assign n11057 = n10305 ^ n8201 ^ n5495 ;
  assign n11058 = ( n583 & n773 ) | ( n583 & n5262 ) | ( n773 & n5262 ) ;
  assign n11059 = ~n3294 & n11058 ;
  assign n11060 = ~n11057 & n11059 ;
  assign n11061 = ( n4767 & n6981 ) | ( n4767 & n11060 ) | ( n6981 & n11060 ) ;
  assign n11062 = n6862 ^ n1940 ^ n722 ;
  assign n11066 = ( n1269 & n3302 ) | ( n1269 & ~n10051 ) | ( n3302 & ~n10051 ) ;
  assign n11067 = ( n5322 & ~n8232 ) | ( n5322 & n11066 ) | ( ~n8232 & n11066 ) ;
  assign n11063 = ( n1144 & n6726 ) | ( n1144 & n6928 ) | ( n6726 & n6928 ) ;
  assign n11064 = n11063 ^ n3873 ^ n2989 ;
  assign n11065 = ( n1704 & n5259 ) | ( n1704 & ~n11064 ) | ( n5259 & ~n11064 ) ;
  assign n11068 = n11067 ^ n11065 ^ n10426 ;
  assign n11069 = ( ~n4285 & n11062 ) | ( ~n4285 & n11068 ) | ( n11062 & n11068 ) ;
  assign n11071 = ( ~n781 & n2638 ) | ( ~n781 & n3086 ) | ( n2638 & n3086 ) ;
  assign n11070 = n6454 & ~n9184 ;
  assign n11072 = n11071 ^ n11070 ^ 1'b0 ;
  assign n11073 = n11072 ^ n1895 ^ n733 ;
  assign n11074 = ~n4408 & n11073 ;
  assign n11075 = ~n11069 & n11074 ;
  assign n11076 = n1834 & ~n3098 ;
  assign n11077 = ( n183 & ~n5147 ) | ( n183 & n11076 ) | ( ~n5147 & n11076 ) ;
  assign n11078 = x82 & ~n11077 ;
  assign n11079 = n2567 & n11078 ;
  assign n11080 = ( ~n826 & n3611 ) | ( ~n826 & n11079 ) | ( n3611 & n11079 ) ;
  assign n11084 = n5607 ^ n632 ^ 1'b0 ;
  assign n11085 = n1633 | n11084 ;
  assign n11081 = ( n3523 & ~n6320 ) | ( n3523 & n8095 ) | ( ~n6320 & n8095 ) ;
  assign n11082 = n11081 ^ n4704 ^ 1'b0 ;
  assign n11083 = ( ~n2438 & n8942 ) | ( ~n2438 & n11082 ) | ( n8942 & n11082 ) ;
  assign n11086 = n11085 ^ n11083 ^ n2007 ;
  assign n11087 = ( ~n914 & n1352 ) | ( ~n914 & n2185 ) | ( n1352 & n2185 ) ;
  assign n11088 = n11087 ^ n6751 ^ n1303 ;
  assign n11089 = ( n9446 & n9530 ) | ( n9446 & ~n11088 ) | ( n9530 & ~n11088 ) ;
  assign n11090 = n2723 & n3286 ;
  assign n11091 = n11090 ^ x34 ^ 1'b0 ;
  assign n11092 = n7895 ^ n5906 ^ 1'b0 ;
  assign n11093 = ~n11091 & n11092 ;
  assign n11094 = n7534 & n11093 ;
  assign n11095 = n6372 & n11094 ;
  assign n11096 = ( ~n2167 & n2755 ) | ( ~n2167 & n3304 ) | ( n2755 & n3304 ) ;
  assign n11097 = n8725 ^ n1955 ^ 1'b0 ;
  assign n11098 = ( n7015 & ~n11096 ) | ( n7015 & n11097 ) | ( ~n11096 & n11097 ) ;
  assign n11100 = n825 & ~n4830 ;
  assign n11101 = n5335 & n11100 ;
  assign n11102 = n11101 ^ n6042 ^ 1'b0 ;
  assign n11103 = n4045 | n11102 ;
  assign n11099 = ( n384 & n888 ) | ( n384 & ~n6364 ) | ( n888 & ~n6364 ) ;
  assign n11104 = n11103 ^ n11099 ^ n10742 ;
  assign n11105 = n11104 ^ n2551 ^ n2133 ;
  assign n11110 = ~n2139 & n3084 ;
  assign n11111 = n11110 ^ n8639 ^ 1'b0 ;
  assign n11106 = ( n3222 & n5795 ) | ( n3222 & n6607 ) | ( n5795 & n6607 ) ;
  assign n11107 = n11106 ^ n6751 ^ 1'b0 ;
  assign n11108 = n6476 ^ n4454 ^ n1479 ;
  assign n11109 = ( n1522 & n11107 ) | ( n1522 & ~n11108 ) | ( n11107 & ~n11108 ) ;
  assign n11112 = n11111 ^ n11109 ^ n4318 ;
  assign n11113 = n2545 ^ n382 ^ 1'b0 ;
  assign n11114 = ~n435 & n2878 ;
  assign n11115 = n3218 & n11114 ;
  assign n11116 = n8650 ^ n6041 ^ n2547 ;
  assign n11117 = ( n1362 & ~n11115 ) | ( n1362 & n11116 ) | ( ~n11115 & n11116 ) ;
  assign n11118 = ( n2716 & n7546 ) | ( n2716 & n11117 ) | ( n7546 & n11117 ) ;
  assign n11119 = n11118 ^ n9069 ^ n4591 ;
  assign n11120 = ( n1337 & ~n8591 ) | ( n1337 & n11119 ) | ( ~n8591 & n11119 ) ;
  assign n11121 = n7988 ^ n4241 ^ n2436 ;
  assign n11122 = n11121 ^ n2314 ^ n793 ;
  assign n11123 = ( ~n7094 & n8580 ) | ( ~n7094 & n11122 ) | ( n8580 & n11122 ) ;
  assign n11124 = n11123 ^ n4461 ^ n4116 ;
  assign n11125 = n11124 ^ n10710 ^ n755 ;
  assign n11126 = n5365 ^ x86 ^ 1'b0 ;
  assign n11127 = ( n8639 & n8772 ) | ( n8639 & ~n11126 ) | ( n8772 & ~n11126 ) ;
  assign n11128 = n5514 ^ n635 ^ 1'b0 ;
  assign n11129 = ( ~n477 & n4213 ) | ( ~n477 & n11128 ) | ( n4213 & n11128 ) ;
  assign n11130 = n11129 ^ n6616 ^ n3679 ;
  assign n11131 = ( n6816 & n7927 ) | ( n6816 & n11130 ) | ( n7927 & n11130 ) ;
  assign n11132 = ( n584 & ~n3528 ) | ( n584 & n5349 ) | ( ~n3528 & n5349 ) ;
  assign n11133 = n11132 ^ n4166 ^ n372 ;
  assign n11140 = ( n345 & n850 ) | ( n345 & n1055 ) | ( n850 & n1055 ) ;
  assign n11139 = n9226 ^ n2109 ^ n1792 ;
  assign n11137 = ~n947 & n2171 ;
  assign n11138 = n2152 & n11137 ;
  assign n11141 = n11140 ^ n11139 ^ n11138 ;
  assign n11134 = n2179 & n2481 ;
  assign n11135 = n2048 & n11134 ;
  assign n11136 = n4756 & ~n11135 ;
  assign n11142 = n11141 ^ n11136 ^ 1'b0 ;
  assign n11155 = n3107 ^ n1619 ^ n1517 ;
  assign n11154 = n3376 ^ n685 ^ 1'b0 ;
  assign n11143 = n1139 ^ n864 ^ n245 ;
  assign n11144 = ( n5895 & ~n6623 ) | ( n5895 & n11143 ) | ( ~n6623 & n11143 ) ;
  assign n11145 = ~n3501 & n3639 ;
  assign n11146 = ~n2816 & n11145 ;
  assign n11147 = ( ~n791 & n11144 ) | ( ~n791 & n11146 ) | ( n11144 & n11146 ) ;
  assign n11148 = n1728 ^ n310 ^ x122 ;
  assign n11149 = n11148 ^ n3009 ^ n2806 ;
  assign n11150 = n2568 ^ n226 ^ 1'b0 ;
  assign n11151 = n11149 & n11150 ;
  assign n11152 = n11147 & n11151 ;
  assign n11153 = n11152 ^ n9312 ^ 1'b0 ;
  assign n11156 = n11155 ^ n11154 ^ n11153 ;
  assign n11157 = n11156 ^ n9280 ^ n5985 ;
  assign n11158 = n11144 ^ n3815 ^ 1'b0 ;
  assign n11159 = n3631 & ~n11158 ;
  assign n11160 = ( n3240 & n11157 ) | ( n3240 & n11159 ) | ( n11157 & n11159 ) ;
  assign n11161 = ( n2516 & n3154 ) | ( n2516 & ~n4083 ) | ( n3154 & ~n4083 ) ;
  assign n11162 = n11161 ^ n757 ^ n586 ;
  assign n11163 = ( n6295 & n10918 ) | ( n6295 & n11162 ) | ( n10918 & n11162 ) ;
  assign n11170 = ( n2106 & n3466 ) | ( n2106 & n4152 ) | ( n3466 & n4152 ) ;
  assign n11164 = n9402 ^ n7961 ^ n3084 ;
  assign n11165 = ( x81 & n9817 ) | ( x81 & ~n11164 ) | ( n9817 & ~n11164 ) ;
  assign n11166 = ( ~n1345 & n3104 ) | ( ~n1345 & n4053 ) | ( n3104 & n4053 ) ;
  assign n11167 = n11166 ^ n10887 ^ n7952 ;
  assign n11168 = ( ~n1319 & n11165 ) | ( ~n1319 & n11167 ) | ( n11165 & n11167 ) ;
  assign n11169 = n9282 | n11168 ;
  assign n11171 = n11170 ^ n11169 ^ 1'b0 ;
  assign n11172 = n6843 ^ n4430 ^ n1774 ;
  assign n11173 = n1657 ^ n847 ^ 1'b0 ;
  assign n11174 = ( n383 & n6184 ) | ( n383 & n11173 ) | ( n6184 & n11173 ) ;
  assign n11175 = n11174 ^ n8996 ^ n5903 ;
  assign n11176 = ( n5504 & n7131 ) | ( n5504 & ~n11175 ) | ( n7131 & ~n11175 ) ;
  assign n11177 = ( n1847 & n2327 ) | ( n1847 & ~n2466 ) | ( n2327 & ~n2466 ) ;
  assign n11178 = n11177 ^ n8747 ^ 1'b0 ;
  assign n11179 = n11178 ^ n1039 ^ 1'b0 ;
  assign n11180 = n4978 & n11179 ;
  assign n11181 = n11180 ^ n10179 ^ n5133 ;
  assign n11182 = ( n3379 & ~n3414 ) | ( n3379 & n5717 ) | ( ~n3414 & n5717 ) ;
  assign n11183 = ( ~n1819 & n3709 ) | ( ~n1819 & n11182 ) | ( n3709 & n11182 ) ;
  assign n11184 = n3685 & ~n3925 ;
  assign n11185 = n9235 ^ n5434 ^ x31 ;
  assign n11186 = n11185 ^ n526 ^ 1'b0 ;
  assign n11189 = ( n1400 & ~n1874 ) | ( n1400 & n10689 ) | ( ~n1874 & n10689 ) ;
  assign n11187 = n7304 ^ n1609 ^ n783 ;
  assign n11188 = n11187 ^ n10734 ^ n1188 ;
  assign n11190 = n11189 ^ n11188 ^ n9559 ;
  assign n11194 = ( n4566 & ~n5682 ) | ( n4566 & n8585 ) | ( ~n5682 & n8585 ) ;
  assign n11195 = ( n8740 & n8803 ) | ( n8740 & n11194 ) | ( n8803 & n11194 ) ;
  assign n11191 = ( n5669 & n8956 ) | ( n5669 & ~n10129 ) | ( n8956 & ~n10129 ) ;
  assign n11192 = n11191 ^ n10384 ^ n5358 ;
  assign n11193 = ( n3954 & n5793 ) | ( n3954 & ~n11192 ) | ( n5793 & ~n11192 ) ;
  assign n11196 = n11195 ^ n11193 ^ n6602 ;
  assign n11197 = n5471 | n6302 ;
  assign n11198 = n7374 ^ n5879 ^ 1'b0 ;
  assign n11199 = ~n2121 & n11198 ;
  assign n11200 = n7563 ^ n4790 ^ n739 ;
  assign n11201 = ( n4517 & n11199 ) | ( n4517 & n11200 ) | ( n11199 & n11200 ) ;
  assign n11202 = n649 & ~n9915 ;
  assign n11203 = ( n10947 & ~n11201 ) | ( n10947 & n11202 ) | ( ~n11201 & n11202 ) ;
  assign n11205 = n7786 ^ n3280 ^ n638 ;
  assign n11204 = ( n2891 & n3707 ) | ( n2891 & ~n5610 ) | ( n3707 & ~n5610 ) ;
  assign n11206 = n11205 ^ n11204 ^ n3715 ;
  assign n11207 = ( ~n2156 & n2936 ) | ( ~n2156 & n11206 ) | ( n2936 & n11206 ) ;
  assign n11208 = n7009 ^ n3620 ^ n2640 ;
  assign n11209 = n11208 ^ n9573 ^ n3392 ;
  assign n11210 = ( n307 & n5150 ) | ( n307 & ~n11209 ) | ( n5150 & ~n11209 ) ;
  assign n11211 = n6545 ^ n2127 ^ n1719 ;
  assign n11212 = ( n4136 & n7829 ) | ( n4136 & n11211 ) | ( n7829 & n11211 ) ;
  assign n11213 = n7506 & n8607 ;
  assign n11214 = ~n6916 & n11213 ;
  assign n11215 = n8788 ^ n2424 ^ n1437 ;
  assign n11216 = ( n2744 & n5850 ) | ( n2744 & n7242 ) | ( n5850 & n7242 ) ;
  assign n11217 = ( n213 & ~n963 ) | ( n213 & n11216 ) | ( ~n963 & n11216 ) ;
  assign n11218 = n11217 ^ n556 ^ 1'b0 ;
  assign n11219 = n11215 & n11218 ;
  assign n11220 = n10359 & n11219 ;
  assign n11221 = n7012 & ~n8718 ;
  assign n11222 = n11221 ^ n400 ^ 1'b0 ;
  assign n11223 = n5931 ^ n3746 ^ n2987 ;
  assign n11224 = n5026 ^ n2179 ^ n2003 ;
  assign n11225 = n11224 ^ n165 ^ 1'b0 ;
  assign n11226 = ( n534 & ~n1324 ) | ( n534 & n4610 ) | ( ~n1324 & n4610 ) ;
  assign n11227 = ( n1603 & n3593 ) | ( n1603 & n11226 ) | ( n3593 & n11226 ) ;
  assign n11228 = n2380 & n3037 ;
  assign n11229 = ~n11227 & n11228 ;
  assign n11230 = ( n11223 & n11225 ) | ( n11223 & ~n11229 ) | ( n11225 & ~n11229 ) ;
  assign n11231 = n11222 & ~n11230 ;
  assign n11232 = ~n7746 & n11231 ;
  assign n11233 = ( ~n907 & n4546 ) | ( ~n907 & n5562 ) | ( n4546 & n5562 ) ;
  assign n11234 = n11233 ^ n10124 ^ n3879 ;
  assign n11235 = ( n707 & n2879 ) | ( n707 & n5674 ) | ( n2879 & n5674 ) ;
  assign n11236 = n686 | n1179 ;
  assign n11237 = n2496 | n11236 ;
  assign n11238 = ( n2044 & n11235 ) | ( n2044 & n11237 ) | ( n11235 & n11237 ) ;
  assign n11239 = ( n8340 & n11234 ) | ( n8340 & n11238 ) | ( n11234 & n11238 ) ;
  assign n11240 = ( n767 & n9661 ) | ( n767 & ~n10291 ) | ( n9661 & ~n10291 ) ;
  assign n11241 = n7185 ^ n1474 ^ n358 ;
  assign n11242 = n11241 ^ n7686 ^ n7000 ;
  assign n11243 = n11242 ^ n11076 ^ n6257 ;
  assign n11244 = n3615 ^ n3000 ^ n968 ;
  assign n11245 = ( n2042 & ~n4539 ) | ( n2042 & n11244 ) | ( ~n4539 & n11244 ) ;
  assign n11246 = ( n310 & n10906 ) | ( n310 & n11245 ) | ( n10906 & n11245 ) ;
  assign n11248 = ~n323 & n2493 ;
  assign n11249 = ~n5132 & n11248 ;
  assign n11250 = ( n3407 & n6057 ) | ( n3407 & n11249 ) | ( n6057 & n11249 ) ;
  assign n11247 = ( ~n541 & n2878 ) | ( ~n541 & n9562 ) | ( n2878 & n9562 ) ;
  assign n11251 = n11250 ^ n11247 ^ n5208 ;
  assign n11252 = n5119 ^ n3707 ^ n1619 ;
  assign n11253 = n11252 ^ n4266 ^ n289 ;
  assign n11254 = ( n4085 & n6688 ) | ( n4085 & n11253 ) | ( n6688 & n11253 ) ;
  assign n11258 = ( n646 & n5418 ) | ( n646 & n7660 ) | ( n5418 & n7660 ) ;
  assign n11259 = ( n4358 & n8305 ) | ( n4358 & ~n11258 ) | ( n8305 & ~n11258 ) ;
  assign n11255 = ( n199 & n4175 ) | ( n199 & ~n5463 ) | ( n4175 & ~n5463 ) ;
  assign n11256 = n11255 ^ n6668 ^ 1'b0 ;
  assign n11257 = n11256 ^ n7766 ^ n1992 ;
  assign n11260 = n11259 ^ n11257 ^ n8968 ;
  assign n11261 = ( n9617 & n11254 ) | ( n9617 & ~n11260 ) | ( n11254 & ~n11260 ) ;
  assign n11262 = n7786 ^ n3817 ^ n2900 ;
  assign n11263 = n11262 ^ n8127 ^ n7389 ;
  assign n11264 = n3830 ^ n800 ^ 1'b0 ;
  assign n11265 = ( n7026 & n9247 ) | ( n7026 & ~n11264 ) | ( n9247 & ~n11264 ) ;
  assign n11269 = n9178 ^ n2956 ^ n853 ;
  assign n11270 = n11269 ^ n7309 ^ n7265 ;
  assign n11271 = ( n7571 & n10591 ) | ( n7571 & n11270 ) | ( n10591 & n11270 ) ;
  assign n11266 = n3537 & n5837 ;
  assign n11267 = ~n10207 & n11266 ;
  assign n11268 = ( n417 & n8858 ) | ( n417 & ~n11267 ) | ( n8858 & ~n11267 ) ;
  assign n11272 = n11271 ^ n11268 ^ n3957 ;
  assign n11273 = n11272 ^ n6130 ^ 1'b0 ;
  assign n11274 = n8831 ^ n1821 ^ n212 ;
  assign n11275 = ( n907 & n7609 ) | ( n907 & ~n11274 ) | ( n7609 & ~n11274 ) ;
  assign n11276 = n8253 ^ n4533 ^ n595 ;
  assign n11279 = ( x107 & ~n2267 ) | ( x107 & n6796 ) | ( ~n2267 & n6796 ) ;
  assign n11280 = n8998 ^ n7210 ^ n224 ;
  assign n11281 = n11279 & ~n11280 ;
  assign n11277 = n7365 ^ n1634 ^ n1176 ;
  assign n11278 = n11277 ^ n7930 ^ n7180 ;
  assign n11282 = n11281 ^ n11278 ^ 1'b0 ;
  assign n11283 = n1379 ^ n997 ^ n514 ;
  assign n11284 = ( n279 & n5562 ) | ( n279 & ~n5795 ) | ( n5562 & ~n5795 ) ;
  assign n11285 = n8612 ^ n4466 ^ n4413 ;
  assign n11286 = ( n2027 & n8387 ) | ( n2027 & ~n11285 ) | ( n8387 & ~n11285 ) ;
  assign n11287 = n4348 & ~n5683 ;
  assign n11288 = ( n11284 & ~n11286 ) | ( n11284 & n11287 ) | ( ~n11286 & n11287 ) ;
  assign n11292 = x102 | n8664 ;
  assign n11293 = n11292 ^ n6409 ^ n2336 ;
  assign n11289 = n9949 ^ n5716 ^ 1'b0 ;
  assign n11290 = ~n3888 & n11289 ;
  assign n11291 = n11290 ^ n8405 ^ n7577 ;
  assign n11294 = n11293 ^ n11291 ^ n6230 ;
  assign n11295 = ( n1169 & n6823 ) | ( n1169 & n10981 ) | ( n6823 & n10981 ) ;
  assign n11297 = n1589 ^ n1429 ^ n1267 ;
  assign n11298 = ( n1140 & n1441 ) | ( n1140 & n11297 ) | ( n1441 & n11297 ) ;
  assign n11299 = n11298 ^ n4071 ^ n3054 ;
  assign n11296 = ( n440 & ~n1098 ) | ( n440 & n10465 ) | ( ~n1098 & n10465 ) ;
  assign n11300 = n11299 ^ n11296 ^ n1465 ;
  assign n11301 = n5137 | n11300 ;
  assign n11302 = n11301 ^ n5779 ^ 1'b0 ;
  assign n11303 = ( n2505 & n4397 ) | ( n2505 & n5085 ) | ( n4397 & n5085 ) ;
  assign n11304 = n3391 ^ n2304 ^ n1884 ;
  assign n11305 = n11304 ^ n6118 ^ n491 ;
  assign n11306 = ( n2085 & n8089 ) | ( n2085 & n11305 ) | ( n8089 & n11305 ) ;
  assign n11307 = ( ~n3197 & n4794 ) | ( ~n3197 & n11306 ) | ( n4794 & n11306 ) ;
  assign n11308 = ( n3679 & n4267 ) | ( n3679 & ~n5844 ) | ( n4267 & ~n5844 ) ;
  assign n11309 = ( n2250 & ~n9054 ) | ( n2250 & n11308 ) | ( ~n9054 & n11308 ) ;
  assign n11310 = ( n7580 & ~n7883 ) | ( n7580 & n11309 ) | ( ~n7883 & n11309 ) ;
  assign n11311 = ( n1361 & n3679 ) | ( n1361 & n11310 ) | ( n3679 & n11310 ) ;
  assign n11312 = n782 & ~n11311 ;
  assign n11313 = n10206 ^ n8742 ^ n8205 ;
  assign n11314 = n11313 ^ n3909 ^ n3263 ;
  assign n11319 = ( n1083 & n4113 ) | ( n1083 & ~n10726 ) | ( n4113 & ~n10726 ) ;
  assign n11317 = n6155 ^ n2805 ^ n873 ;
  assign n11318 = n11317 ^ n8447 ^ n263 ;
  assign n11315 = n5965 ^ n2831 ^ x47 ;
  assign n11316 = n5282 | n11315 ;
  assign n11320 = n11319 ^ n11318 ^ n11316 ;
  assign n11321 = n4766 ^ n975 ^ n167 ;
  assign n11322 = n1026 & ~n11321 ;
  assign n11323 = ~n11320 & n11322 ;
  assign n11324 = n7930 & ~n11323 ;
  assign n11325 = n11324 ^ n687 ^ 1'b0 ;
  assign n11326 = ( n11312 & n11314 ) | ( n11312 & ~n11325 ) | ( n11314 & ~n11325 ) ;
  assign n11327 = ( n1123 & n7330 ) | ( n1123 & n8510 ) | ( n7330 & n8510 ) ;
  assign n11328 = ( n5104 & n5414 ) | ( n5104 & n11327 ) | ( n5414 & n11327 ) ;
  assign n11329 = ( n1499 & ~n1528 ) | ( n1499 & n2750 ) | ( ~n1528 & n2750 ) ;
  assign n11330 = n3480 & n11329 ;
  assign n11331 = n11330 ^ n4711 ^ 1'b0 ;
  assign n11333 = n3048 ^ n537 ^ n328 ;
  assign n11332 = ( n4293 & n4378 ) | ( n4293 & ~n7015 ) | ( n4378 & ~n7015 ) ;
  assign n11334 = n11333 ^ n11332 ^ n10069 ;
  assign n11335 = ( n1973 & n4029 ) | ( n1973 & ~n5479 ) | ( n4029 & ~n5479 ) ;
  assign n11336 = ( ~n4038 & n10307 ) | ( ~n4038 & n11335 ) | ( n10307 & n11335 ) ;
  assign n11337 = n3824 ^ n1732 ^ n524 ;
  assign n11338 = ( ~n2048 & n7122 ) | ( ~n2048 & n8901 ) | ( n7122 & n8901 ) ;
  assign n11339 = ( n717 & ~n8053 ) | ( n717 & n11338 ) | ( ~n8053 & n11338 ) ;
  assign n11340 = ( n11336 & n11337 ) | ( n11336 & ~n11339 ) | ( n11337 & ~n11339 ) ;
  assign n11341 = n8669 ^ n8053 ^ n6897 ;
  assign n11342 = ( ~n2448 & n3778 ) | ( ~n2448 & n3779 ) | ( n3778 & n3779 ) ;
  assign n11343 = n2077 ^ n1682 ^ n349 ;
  assign n11344 = n11343 ^ n5826 ^ x96 ;
  assign n11348 = n3969 ^ n1330 ^ n1323 ;
  assign n11349 = ( n534 & n3905 ) | ( n534 & ~n4321 ) | ( n3905 & ~n4321 ) ;
  assign n11350 = ( n1939 & n11348 ) | ( n1939 & n11349 ) | ( n11348 & n11349 ) ;
  assign n11345 = n350 & n4010 ;
  assign n11346 = ~n6206 & n11345 ;
  assign n11347 = n11346 ^ n2505 ^ n988 ;
  assign n11351 = n11350 ^ n11347 ^ n3413 ;
  assign n11352 = ( n1408 & n3417 ) | ( n1408 & n6339 ) | ( n3417 & n6339 ) ;
  assign n11353 = n11352 ^ n7847 ^ n336 ;
  assign n11354 = ( n11344 & n11351 ) | ( n11344 & n11353 ) | ( n11351 & n11353 ) ;
  assign n11355 = n8987 ^ n6586 ^ n6098 ;
  assign n11356 = n11355 ^ n3267 ^ n2248 ;
  assign n11357 = n11356 ^ n3987 ^ n2845 ;
  assign n11358 = n11357 ^ n10243 ^ n5662 ;
  assign n11359 = n9520 ^ n6551 ^ n4680 ;
  assign n11360 = ( ~n3185 & n7256 ) | ( ~n3185 & n9124 ) | ( n7256 & n9124 ) ;
  assign n11361 = ( n572 & n7146 ) | ( n572 & ~n11360 ) | ( n7146 & ~n11360 ) ;
  assign n11362 = ( n2802 & n3275 ) | ( n2802 & n3681 ) | ( n3275 & n3681 ) ;
  assign n11363 = ( ~n4188 & n5259 ) | ( ~n4188 & n7048 ) | ( n5259 & n7048 ) ;
  assign n11364 = n11362 | n11363 ;
  assign n11365 = ( ~n9095 & n11361 ) | ( ~n9095 & n11364 ) | ( n11361 & n11364 ) ;
  assign n11366 = n7265 ^ n946 ^ 1'b0 ;
  assign n11367 = n5200 | n11366 ;
  assign n11368 = n8967 ^ n2563 ^ n1941 ;
  assign n11369 = ( ~n6840 & n11367 ) | ( ~n6840 & n11368 ) | ( n11367 & n11368 ) ;
  assign n11370 = n706 | n1517 ;
  assign n11371 = n9319 | n11370 ;
  assign n11372 = n11371 ^ n1961 ^ n171 ;
  assign n11373 = n6467 ^ n2054 ^ 1'b0 ;
  assign n11374 = n11372 & ~n11373 ;
  assign n11375 = ( ~n4528 & n8358 ) | ( ~n4528 & n11374 ) | ( n8358 & n11374 ) ;
  assign n11376 = n11375 ^ n5550 ^ n2176 ;
  assign n11377 = n6154 & n11376 ;
  assign n11378 = n11377 ^ n11122 ^ n10070 ;
  assign n11379 = ( n193 & n8194 ) | ( n193 & n10372 ) | ( n8194 & n10372 ) ;
  assign n11382 = n5480 ^ n2059 ^ 1'b0 ;
  assign n11380 = ( ~x60 & n4232 ) | ( ~x60 & n11264 ) | ( n4232 & n11264 ) ;
  assign n11381 = ( n6344 & n6497 ) | ( n6344 & ~n11380 ) | ( n6497 & ~n11380 ) ;
  assign n11383 = n11382 ^ n11381 ^ n9754 ;
  assign n11384 = ( ~n5950 & n7371 ) | ( ~n5950 & n11383 ) | ( n7371 & n11383 ) ;
  assign n11385 = n5893 ^ n3647 ^ n436 ;
  assign n11386 = ( n2320 & n4750 ) | ( n2320 & ~n11385 ) | ( n4750 & ~n11385 ) ;
  assign n11387 = n11386 ^ n10606 ^ n2039 ;
  assign n11390 = x110 & ~n6853 ;
  assign n11391 = n11390 ^ n3020 ^ 1'b0 ;
  assign n11392 = n11391 ^ n7980 ^ n5905 ;
  assign n11393 = n11392 ^ n6146 ^ n1910 ;
  assign n11388 = n4087 ^ n3901 ^ n567 ;
  assign n11389 = n11388 ^ n3128 ^ n1213 ;
  assign n11394 = n11393 ^ n11389 ^ n5784 ;
  assign n11395 = ( ~n362 & n11387 ) | ( ~n362 & n11394 ) | ( n11387 & n11394 ) ;
  assign n11396 = n11395 ^ n10937 ^ n4931 ;
  assign n11397 = ~n1516 & n10442 ;
  assign n11398 = n9237 ^ n1877 ^ 1'b0 ;
  assign n11399 = x92 & n11398 ;
  assign n11400 = n3413 & n11399 ;
  assign n11401 = n3044 & n11400 ;
  assign n11402 = n11401 ^ n5695 ^ n1639 ;
  assign n11403 = ( n3325 & ~n6378 ) | ( n3325 & n6663 ) | ( ~n6378 & n6663 ) ;
  assign n11404 = ( n142 & ~n10787 ) | ( n142 & n11403 ) | ( ~n10787 & n11403 ) ;
  assign n11405 = ( n6394 & n9357 ) | ( n6394 & n11199 ) | ( n9357 & n11199 ) ;
  assign n11406 = ( n1106 & n3527 ) | ( n1106 & n10745 ) | ( n3527 & n10745 ) ;
  assign n11408 = n7905 ^ n5770 ^ n3502 ;
  assign n11409 = n1263 & n11408 ;
  assign n11407 = ( ~n4871 & n9966 ) | ( ~n4871 & n10538 ) | ( n9966 & n10538 ) ;
  assign n11410 = n11409 ^ n11407 ^ 1'b0 ;
  assign n11413 = n9523 ^ n5887 ^ 1'b0 ;
  assign n11411 = ( x80 & n3924 ) | ( x80 & n7407 ) | ( n3924 & n7407 ) ;
  assign n11412 = n11411 ^ n5200 ^ n3695 ;
  assign n11414 = n11413 ^ n11412 ^ n714 ;
  assign n11419 = n9386 ^ n3722 ^ n2993 ;
  assign n11415 = n6541 ^ n1612 ^ n630 ;
  assign n11416 = ( n414 & n1280 ) | ( n414 & n8987 ) | ( n1280 & n8987 ) ;
  assign n11417 = ( n5945 & n11415 ) | ( n5945 & ~n11416 ) | ( n11415 & ~n11416 ) ;
  assign n11418 = n11417 ^ n10991 ^ n305 ;
  assign n11420 = n11419 ^ n11418 ^ n9598 ;
  assign n11421 = ( n283 & n466 ) | ( n283 & n1211 ) | ( n466 & n1211 ) ;
  assign n11422 = n2970 & n3777 ;
  assign n11423 = ( n11372 & ~n11421 ) | ( n11372 & n11422 ) | ( ~n11421 & n11422 ) ;
  assign n11424 = ~n4009 & n4219 ;
  assign n11425 = ( n3899 & n11423 ) | ( n3899 & n11424 ) | ( n11423 & n11424 ) ;
  assign n11426 = ( n5018 & ~n7694 ) | ( n5018 & n9998 ) | ( ~n7694 & n9998 ) ;
  assign n11427 = n11426 ^ n4758 ^ n333 ;
  assign n11428 = ( n3109 & n3339 ) | ( n3109 & ~n11427 ) | ( n3339 & ~n11427 ) ;
  assign n11429 = n827 | n9001 ;
  assign n11430 = n6116 | n11429 ;
  assign n11431 = ( n1925 & n2701 ) | ( n1925 & ~n10461 ) | ( n2701 & ~n10461 ) ;
  assign n11432 = n11430 | n11431 ;
  assign n11433 = n11144 ^ n1397 ^ x126 ;
  assign n11434 = n6468 & n11433 ;
  assign n11435 = n9901 ^ n4720 ^ n1501 ;
  assign n11436 = ( n3431 & ~n5695 ) | ( n3431 & n11435 ) | ( ~n5695 & n11435 ) ;
  assign n11437 = ( n2152 & ~n9020 ) | ( n2152 & n11436 ) | ( ~n9020 & n11436 ) ;
  assign n11438 = ( n4838 & ~n8915 ) | ( n4838 & n10112 ) | ( ~n8915 & n10112 ) ;
  assign n11448 = ( n1815 & n2122 ) | ( n1815 & n3494 ) | ( n2122 & n3494 ) ;
  assign n11449 = n11448 ^ n2995 ^ 1'b0 ;
  assign n11450 = ~n1859 & n11449 ;
  assign n11451 = ~n4788 & n11450 ;
  assign n11452 = n8008 ^ n7251 ^ n4289 ;
  assign n11453 = n8244 ^ n5039 ^ n3581 ;
  assign n11454 = ( n11451 & ~n11452 ) | ( n11451 & n11453 ) | ( ~n11452 & n11453 ) ;
  assign n11442 = ( n5006 & n7228 ) | ( n5006 & ~n8189 ) | ( n7228 & ~n8189 ) ;
  assign n11444 = n1798 | n2368 ;
  assign n11445 = n1324 & ~n11444 ;
  assign n11443 = n9068 ^ n6777 ^ n5236 ;
  assign n11446 = n11445 ^ n11443 ^ n7139 ;
  assign n11447 = ( n7379 & ~n11442 ) | ( n7379 & n11446 ) | ( ~n11442 & n11446 ) ;
  assign n11440 = n8787 ^ n6417 ^ n3519 ;
  assign n11439 = n8221 ^ n3740 ^ n301 ;
  assign n11441 = n11440 ^ n11439 ^ n6546 ;
  assign n11455 = n11454 ^ n11447 ^ n11441 ;
  assign n11456 = n11455 ^ n9391 ^ n4510 ;
  assign n11459 = ( n4009 & n5843 ) | ( n4009 & n8565 ) | ( n5843 & n8565 ) ;
  assign n11460 = ( n2110 & ~n6804 ) | ( n2110 & n11459 ) | ( ~n6804 & n11459 ) ;
  assign n11461 = n5617 & n11460 ;
  assign n11462 = n7395 & n11461 ;
  assign n11457 = ( n740 & n4287 ) | ( n740 & n6712 ) | ( n4287 & n6712 ) ;
  assign n11458 = n11457 ^ n11123 ^ x118 ;
  assign n11463 = n11462 ^ n11458 ^ n8303 ;
  assign n11464 = x33 & n6097 ;
  assign n11465 = n11464 ^ n2790 ^ 1'b0 ;
  assign n11466 = ( ~n746 & n3060 ) | ( ~n746 & n4897 ) | ( n3060 & n4897 ) ;
  assign n11467 = n5150 | n11466 ;
  assign n11468 = n951 & ~n11467 ;
  assign n11469 = n11468 ^ n8914 ^ 1'b0 ;
  assign n11470 = n889 | n6573 ;
  assign n11471 = n4841 ^ n1732 ^ x8 ;
  assign n11472 = ( n4686 & n7668 ) | ( n4686 & ~n11471 ) | ( n7668 & ~n11471 ) ;
  assign n11473 = ( n1823 & ~n3515 ) | ( n1823 & n6435 ) | ( ~n3515 & n6435 ) ;
  assign n11474 = ( n1975 & ~n11472 ) | ( n1975 & n11473 ) | ( ~n11472 & n11473 ) ;
  assign n11475 = n11474 ^ n9874 ^ n4370 ;
  assign n11476 = ( n10568 & n11470 ) | ( n10568 & n11475 ) | ( n11470 & n11475 ) ;
  assign n11478 = ( ~n347 & n1861 ) | ( ~n347 & n2916 ) | ( n1861 & n2916 ) ;
  assign n11479 = n11478 ^ n9192 ^ n4663 ;
  assign n11480 = ( n1780 & ~n8943 ) | ( n1780 & n11479 ) | ( ~n8943 & n11479 ) ;
  assign n11477 = n6782 & ~n11079 ;
  assign n11481 = n11480 ^ n11477 ^ 1'b0 ;
  assign n11482 = ( n4273 & n9532 ) | ( n4273 & n11481 ) | ( n9532 & n11481 ) ;
  assign n11485 = n2154 ^ n617 ^ 1'b0 ;
  assign n11486 = n3744 | n11485 ;
  assign n11484 = ( n2581 & n4106 ) | ( n2581 & n9915 ) | ( n4106 & n9915 ) ;
  assign n11483 = ( ~n2902 & n7442 ) | ( ~n2902 & n9978 ) | ( n7442 & n9978 ) ;
  assign n11487 = n11486 ^ n11484 ^ n11483 ;
  assign n11488 = ( x19 & ~n5406 ) | ( x19 & n10371 ) | ( ~n5406 & n10371 ) ;
  assign n11489 = n11488 ^ n8557 ^ n5826 ;
  assign n11490 = n11489 ^ n10624 ^ n443 ;
  assign n11491 = ( ~x92 & n671 ) | ( ~x92 & n6648 ) | ( n671 & n6648 ) ;
  assign n11492 = n4213 & ~n11491 ;
  assign n11493 = n5256 & n11492 ;
  assign n11494 = n2901 ^ n2116 ^ n445 ;
  assign n11495 = ( n4841 & n9556 ) | ( n4841 & ~n11494 ) | ( n9556 & ~n11494 ) ;
  assign n11496 = n11495 ^ n8470 ^ n5243 ;
  assign n11497 = ( n4816 & n11493 ) | ( n4816 & ~n11496 ) | ( n11493 & ~n11496 ) ;
  assign n11498 = ~n1119 & n10040 ;
  assign n11499 = ( n3293 & ~n5485 ) | ( n3293 & n11498 ) | ( ~n5485 & n11498 ) ;
  assign n11500 = n8688 ^ n2913 ^ n2486 ;
  assign n11501 = n3224 ^ n2806 ^ n643 ;
  assign n11502 = ( ~n517 & n1155 ) | ( ~n517 & n1785 ) | ( n1155 & n1785 ) ;
  assign n11503 = ( n2467 & n11501 ) | ( n2467 & n11502 ) | ( n11501 & n11502 ) ;
  assign n11504 = n2273 | n11503 ;
  assign n11505 = n11500 | n11504 ;
  assign n11508 = n2623 ^ n2329 ^ 1'b0 ;
  assign n11509 = n3233 & n11508 ;
  assign n11506 = ( ~n3526 & n4978 ) | ( ~n3526 & n9780 ) | ( n4978 & n9780 ) ;
  assign n11507 = n11506 ^ n1671 ^ n1245 ;
  assign n11510 = n11509 ^ n11507 ^ n248 ;
  assign n11511 = n7481 ^ n1421 ^ n923 ;
  assign n11512 = ( ~n1964 & n7876 ) | ( ~n1964 & n11511 ) | ( n7876 & n11511 ) ;
  assign n11513 = ( n627 & n1705 ) | ( n627 & n8490 ) | ( n1705 & n8490 ) ;
  assign n11514 = n6316 ^ n6300 ^ n5505 ;
  assign n11515 = n11514 ^ n5655 ^ n3175 ;
  assign n11516 = ( n5894 & n11513 ) | ( n5894 & n11515 ) | ( n11513 & n11515 ) ;
  assign n11517 = n9362 ^ n7599 ^ n952 ;
  assign n11518 = n9479 ^ n5150 ^ n2607 ;
  assign n11519 = n11518 ^ n6625 ^ n2641 ;
  assign n11520 = ( ~n3323 & n3449 ) | ( ~n3323 & n8285 ) | ( n3449 & n8285 ) ;
  assign n11521 = n11520 ^ n2444 ^ n1289 ;
  assign n11522 = ( ~n3245 & n4693 ) | ( ~n3245 & n11521 ) | ( n4693 & n11521 ) ;
  assign n11523 = ( ~n568 & n11519 ) | ( ~n568 & n11522 ) | ( n11519 & n11522 ) ;
  assign n11524 = n9077 & ~n11523 ;
  assign n11525 = n1217 ^ n1089 ^ 1'b0 ;
  assign n11526 = n4426 ^ n1311 ^ n1103 ;
  assign n11527 = n4518 ^ n2709 ^ n2178 ;
  assign n11528 = ( n330 & n11526 ) | ( n330 & ~n11527 ) | ( n11526 & ~n11527 ) ;
  assign n11529 = n5713 ^ n4225 ^ 1'b0 ;
  assign n11530 = n11529 ^ n9802 ^ n6115 ;
  assign n11531 = n5891 & n7199 ;
  assign n11532 = ( n3232 & n10020 ) | ( n3232 & ~n11531 ) | ( n10020 & ~n11531 ) ;
  assign n11533 = ( n4014 & n4884 ) | ( n4014 & n7573 ) | ( n4884 & n7573 ) ;
  assign n11535 = n3582 | n4463 ;
  assign n11534 = n3167 & ~n6784 ;
  assign n11536 = n11535 ^ n11534 ^ 1'b0 ;
  assign n11537 = n11536 ^ n8103 ^ n355 ;
  assign n11538 = ( n2729 & n4451 ) | ( n2729 & n11537 ) | ( n4451 & n11537 ) ;
  assign n11539 = ( n2404 & n11533 ) | ( n2404 & n11538 ) | ( n11533 & n11538 ) ;
  assign n11540 = n5376 ^ n3052 ^ n884 ;
  assign n11541 = ( n3774 & n7726 ) | ( n3774 & n9061 ) | ( n7726 & n9061 ) ;
  assign n11542 = ( n1957 & ~n2837 ) | ( n1957 & n10623 ) | ( ~n2837 & n10623 ) ;
  assign n11543 = n11541 | n11542 ;
  assign n11544 = n11540 | n11543 ;
  assign n11545 = ( n2193 & n3120 ) | ( n2193 & ~n10942 ) | ( n3120 & ~n10942 ) ;
  assign n11546 = ( ~n8341 & n9780 ) | ( ~n8341 & n11545 ) | ( n9780 & n11545 ) ;
  assign n11547 = n3724 ^ n1932 ^ 1'b0 ;
  assign n11548 = n4334 & n11547 ;
  assign n11549 = n11548 ^ n1743 ^ n144 ;
  assign n11550 = n9470 ^ n933 ^ 1'b0 ;
  assign n11551 = n788 & n3013 ;
  assign n11552 = n5741 & n11551 ;
  assign n11553 = n11552 ^ n9399 ^ n9258 ;
  assign n11554 = n11553 ^ n10297 ^ n1591 ;
  assign n11555 = n10944 ^ n4587 ^ n1751 ;
  assign n11556 = n11555 ^ n10682 ^ n929 ;
  assign n11557 = n11556 ^ n8653 ^ n8521 ;
  assign n11568 = n2013 & ~n2598 ;
  assign n11569 = ~n8980 & n11568 ;
  assign n11570 = n5884 ^ n3494 ^ 1'b0 ;
  assign n11571 = ( ~n2656 & n3240 ) | ( ~n2656 & n3677 ) | ( n3240 & n3677 ) ;
  assign n11572 = ( ~n4127 & n11570 ) | ( ~n4127 & n11571 ) | ( n11570 & n11571 ) ;
  assign n11573 = ( n4184 & n4413 ) | ( n4184 & n11572 ) | ( n4413 & n11572 ) ;
  assign n11574 = ( n6307 & n11569 ) | ( n6307 & n11573 ) | ( n11569 & n11573 ) ;
  assign n11567 = ( n830 & ~n6306 ) | ( n830 & n8643 ) | ( ~n6306 & n8643 ) ;
  assign n11563 = ( n917 & n4014 ) | ( n917 & ~n8024 ) | ( n4014 & ~n8024 ) ;
  assign n11558 = n2386 & n4760 ;
  assign n11559 = n5705 ^ n5426 ^ n2683 ;
  assign n11560 = ( n7076 & n7449 ) | ( n7076 & ~n7587 ) | ( n7449 & ~n7587 ) ;
  assign n11561 = ~n11559 & n11560 ;
  assign n11562 = n11558 & n11561 ;
  assign n11564 = n11563 ^ n11562 ^ n2687 ;
  assign n11565 = n5793 ^ n3463 ^ n1483 ;
  assign n11566 = ( ~n10584 & n11564 ) | ( ~n10584 & n11565 ) | ( n11564 & n11565 ) ;
  assign n11575 = n11574 ^ n11567 ^ n11566 ;
  assign n11576 = n3674 ^ n2710 ^ n1335 ;
  assign n11583 = ( n2203 & n2942 ) | ( n2203 & n8682 ) | ( n2942 & n8682 ) ;
  assign n11582 = ~n3387 & n5093 ;
  assign n11584 = n11583 ^ n11582 ^ 1'b0 ;
  assign n11585 = ( n7342 & n9395 ) | ( n7342 & ~n11584 ) | ( n9395 & ~n11584 ) ;
  assign n11580 = ( n3740 & n5517 ) | ( n3740 & ~n7449 ) | ( n5517 & ~n7449 ) ;
  assign n11581 = ( n1013 & n6911 ) | ( n1013 & ~n11580 ) | ( n6911 & ~n11580 ) ;
  assign n11577 = n11317 ^ n8496 ^ 1'b0 ;
  assign n11578 = n5610 & ~n11577 ;
  assign n11579 = ( n5069 & n10716 ) | ( n5069 & n11578 ) | ( n10716 & n11578 ) ;
  assign n11586 = n11585 ^ n11581 ^ n11579 ;
  assign n11587 = ( n5278 & ~n11576 ) | ( n5278 & n11586 ) | ( ~n11576 & n11586 ) ;
  assign n11588 = n7057 ^ n3086 ^ 1'b0 ;
  assign n11589 = ~n2483 & n11588 ;
  assign n11590 = n7465 & ~n11299 ;
  assign n11591 = n2757 & ~n4195 ;
  assign n11592 = n6487 & n11591 ;
  assign n11593 = ( n7905 & ~n11590 ) | ( n7905 & n11592 ) | ( ~n11590 & n11592 ) ;
  assign n11594 = n264 & ~n9547 ;
  assign n11595 = n11594 ^ n10360 ^ n6686 ;
  assign n11596 = n11595 ^ n3528 ^ n3351 ;
  assign n11597 = n1154 & ~n8679 ;
  assign n11598 = n3813 & n11597 ;
  assign n11599 = ( n339 & n3352 ) | ( n339 & ~n11598 ) | ( n3352 & ~n11598 ) ;
  assign n11600 = n11599 ^ n8071 ^ n5278 ;
  assign n11603 = n2468 ^ n2211 ^ 1'b0 ;
  assign n11604 = ~n4464 & n11603 ;
  assign n11601 = n10139 ^ n6743 ^ 1'b0 ;
  assign n11602 = n2322 & n11601 ;
  assign n11605 = n11604 ^ n11602 ^ 1'b0 ;
  assign n11606 = n11605 ^ n6379 ^ n795 ;
  assign n11610 = ( ~n1193 & n4404 ) | ( ~n1193 & n9805 ) | ( n4404 & n9805 ) ;
  assign n11611 = n11610 ^ n1825 ^ n982 ;
  assign n11607 = n1061 | n8912 ;
  assign n11608 = n10276 | n11607 ;
  assign n11609 = ( n1003 & ~n4660 ) | ( n1003 & n11608 ) | ( ~n4660 & n11608 ) ;
  assign n11612 = n11611 ^ n11609 ^ n1718 ;
  assign n11613 = x82 | n11612 ;
  assign n11617 = ( n1108 & ~n1790 ) | ( n1108 & n5591 ) | ( ~n1790 & n5591 ) ;
  assign n11618 = ( ~n1685 & n7136 ) | ( ~n1685 & n11617 ) | ( n7136 & n11617 ) ;
  assign n11619 = n11618 ^ n169 ^ 1'b0 ;
  assign n11620 = n1218 & n11619 ;
  assign n11621 = n4480 & ~n6822 ;
  assign n11622 = ~n11620 & n11621 ;
  assign n11616 = ( n959 & n5770 ) | ( n959 & n6551 ) | ( n5770 & n6551 ) ;
  assign n11614 = ( n1240 & n2303 ) | ( n1240 & n3847 ) | ( n2303 & n3847 ) ;
  assign n11615 = n11614 ^ n11278 ^ n387 ;
  assign n11623 = n11622 ^ n11616 ^ n11615 ;
  assign n11624 = ( n1403 & ~n3898 ) | ( n1403 & n4076 ) | ( ~n3898 & n4076 ) ;
  assign n11625 = n11624 ^ n11161 ^ 1'b0 ;
  assign n11626 = n2574 & ~n11625 ;
  assign n11627 = n6885 | n11626 ;
  assign n11628 = n2638 ^ n386 ^ 1'b0 ;
  assign n11629 = ( x73 & n881 ) | ( x73 & n11628 ) | ( n881 & n11628 ) ;
  assign n11630 = n1249 & ~n6450 ;
  assign n11631 = n11629 & n11630 ;
  assign n11632 = n11631 ^ n3390 ^ 1'b0 ;
  assign n11633 = n11000 & n11632 ;
  assign n11634 = n5969 ^ n3123 ^ x95 ;
  assign n11635 = ( ~n2402 & n7022 ) | ( ~n2402 & n11634 ) | ( n7022 & n11634 ) ;
  assign n11636 = n5021 ^ n3600 ^ n1494 ;
  assign n11637 = n6276 ^ n4910 ^ n4011 ;
  assign n11638 = n659 & n11637 ;
  assign n11639 = ~n11636 & n11638 ;
  assign n11640 = n11639 ^ n6512 ^ 1'b0 ;
  assign n11641 = ~n1766 & n11640 ;
  assign n11642 = ( n6258 & ~n9042 ) | ( n6258 & n9588 ) | ( ~n9042 & n9588 ) ;
  assign n11643 = ( ~n2946 & n3847 ) | ( ~n2946 & n11642 ) | ( n3847 & n11642 ) ;
  assign n11644 = n3581 ^ n2674 ^ n1483 ;
  assign n11645 = ( n3293 & ~n3771 ) | ( n3293 & n11644 ) | ( ~n3771 & n11644 ) ;
  assign n11646 = n405 | n11645 ;
  assign n11647 = n11643 | n11646 ;
  assign n11652 = ( n2866 & n7480 ) | ( n2866 & ~n9479 ) | ( n7480 & ~n9479 ) ;
  assign n11649 = ( n3363 & n3601 ) | ( n3363 & ~n6282 ) | ( n3601 & ~n6282 ) ;
  assign n11650 = n6409 & ~n11649 ;
  assign n11651 = n11650 ^ n10670 ^ n9365 ;
  assign n11653 = n11652 ^ n11651 ^ n5294 ;
  assign n11648 = ( x75 & n6384 ) | ( x75 & n9718 ) | ( n6384 & n9718 ) ;
  assign n11654 = n11653 ^ n11648 ^ n10066 ;
  assign n11657 = ( n1672 & n2651 ) | ( n1672 & ~n3864 ) | ( n2651 & ~n3864 ) ;
  assign n11658 = n11657 ^ n973 ^ 1'b0 ;
  assign n11659 = n878 & ~n11658 ;
  assign n11655 = ( ~x79 & n2090 ) | ( ~x79 & n4408 ) | ( n2090 & n4408 ) ;
  assign n11656 = n11655 ^ n5042 ^ n4670 ;
  assign n11660 = n11659 ^ n11656 ^ 1'b0 ;
  assign n11661 = n554 & n2327 ;
  assign n11662 = n11661 ^ n10177 ^ n7983 ;
  assign n11663 = ( ~n5640 & n6336 ) | ( ~n5640 & n7579 ) | ( n6336 & n7579 ) ;
  assign n11664 = ( n762 & ~n11258 ) | ( n762 & n11663 ) | ( ~n11258 & n11663 ) ;
  assign n11665 = n10176 ^ n6037 ^ 1'b0 ;
  assign n11666 = ~n7021 & n11665 ;
  assign n11667 = ~n7200 & n11666 ;
  assign n11668 = n11667 ^ n3412 ^ 1'b0 ;
  assign n11669 = n11668 ^ n3212 ^ n915 ;
  assign n11670 = ( n11662 & n11664 ) | ( n11662 & ~n11669 ) | ( n11664 & ~n11669 ) ;
  assign n11671 = n9532 ^ n7486 ^ x30 ;
  assign n11672 = n11671 ^ n2814 ^ n2131 ;
  assign n11673 = n11672 ^ n6616 ^ x109 ;
  assign n11674 = ( n282 & n641 ) | ( n282 & ~n11673 ) | ( n641 & ~n11673 ) ;
  assign n11675 = n11674 ^ n3578 ^ 1'b0 ;
  assign n11676 = n5060 ^ n2387 ^ 1'b0 ;
  assign n11678 = ( ~n2081 & n4376 ) | ( ~n2081 & n4774 ) | ( n4376 & n4774 ) ;
  assign n11679 = n11678 ^ n5993 ^ n5545 ;
  assign n11677 = n6620 ^ n3307 ^ n239 ;
  assign n11680 = n11679 ^ n11677 ^ n5738 ;
  assign n11694 = ( n1000 & ~n2172 ) | ( n1000 & n7531 ) | ( ~n2172 & n7531 ) ;
  assign n11695 = n11694 ^ n4170 ^ n1579 ;
  assign n11693 = n2931 ^ n2659 ^ n1895 ;
  assign n11696 = n11695 ^ n11693 ^ n1544 ;
  assign n11690 = ( n891 & n2670 ) | ( n891 & ~n5088 ) | ( n2670 & ~n5088 ) ;
  assign n11687 = n11274 ^ n2129 ^ n415 ;
  assign n11688 = n11687 ^ n2116 ^ n1734 ;
  assign n11689 = n11688 ^ n2233 ^ 1'b0 ;
  assign n11691 = n11690 ^ n11689 ^ n8275 ;
  assign n11684 = ( ~n254 & n1676 ) | ( ~n254 & n2627 ) | ( n1676 & n2627 ) ;
  assign n11685 = n2360 | n11684 ;
  assign n11686 = ( n5014 & n5172 ) | ( n5014 & n11685 ) | ( n5172 & n11685 ) ;
  assign n11681 = n9820 ^ n6330 ^ n3478 ;
  assign n11682 = n11681 ^ n4566 ^ 1'b0 ;
  assign n11683 = n11682 ^ n507 ^ n178 ;
  assign n11692 = n11691 ^ n11686 ^ n11683 ;
  assign n11697 = n11696 ^ n11692 ^ x81 ;
  assign n11698 = n7988 & ~n8294 ;
  assign n11700 = n7916 ^ n7799 ^ 1'b0 ;
  assign n11699 = n11012 ^ n6809 ^ n5260 ;
  assign n11701 = n11700 ^ n11699 ^ n1577 ;
  assign n11702 = n9091 ^ n3940 ^ n3124 ;
  assign n11704 = ( n356 & n1674 ) | ( n356 & ~n9739 ) | ( n1674 & ~n9739 ) ;
  assign n11703 = ( n803 & n2898 ) | ( n803 & ~n9312 ) | ( n2898 & ~n9312 ) ;
  assign n11705 = n11704 ^ n11703 ^ n9719 ;
  assign n11706 = ( ~n9142 & n11702 ) | ( ~n9142 & n11705 ) | ( n11702 & n11705 ) ;
  assign n11707 = ( n3346 & n6093 ) | ( n3346 & n8622 ) | ( n6093 & n8622 ) ;
  assign n11708 = n3881 ^ n3201 ^ n371 ;
  assign n11709 = n11708 ^ n7192 ^ n2137 ;
  assign n11710 = n11709 ^ n9961 ^ x95 ;
  assign n11711 = n11710 ^ n4315 ^ 1'b0 ;
  assign n11712 = n11707 & n11711 ;
  assign n11713 = ( n6034 & n8573 ) | ( n6034 & ~n11170 ) | ( n8573 & ~n11170 ) ;
  assign n11714 = ( n3244 & n3956 ) | ( n3244 & n9748 ) | ( n3956 & n9748 ) ;
  assign n11715 = ( n440 & n745 ) | ( n440 & n7947 ) | ( n745 & n7947 ) ;
  assign n11716 = ( n1882 & ~n4890 ) | ( n1882 & n11715 ) | ( ~n4890 & n11715 ) ;
  assign n11717 = ( ~n2669 & n11714 ) | ( ~n2669 & n11716 ) | ( n11714 & n11716 ) ;
  assign n11718 = ( n4828 & n9489 ) | ( n4828 & n11717 ) | ( n9489 & n11717 ) ;
  assign n11719 = ( ~n1253 & n6220 ) | ( ~n1253 & n8862 ) | ( n6220 & n8862 ) ;
  assign n11720 = n826 ^ n535 ^ 1'b0 ;
  assign n11721 = ( n6659 & n7504 ) | ( n6659 & ~n8687 ) | ( n7504 & ~n8687 ) ;
  assign n11722 = ( n4153 & n5554 ) | ( n4153 & ~n11721 ) | ( n5554 & ~n11721 ) ;
  assign n11723 = ( n2836 & n11503 ) | ( n2836 & n11722 ) | ( n11503 & n11722 ) ;
  assign n11724 = ( ~n914 & n5466 ) | ( ~n914 & n6777 ) | ( n5466 & n6777 ) ;
  assign n11725 = ( n3068 & n7183 ) | ( n3068 & ~n11724 ) | ( n7183 & ~n11724 ) ;
  assign n11726 = n3120 ^ n1838 ^ n1682 ;
  assign n11727 = n11725 & ~n11726 ;
  assign n11728 = n11727 ^ n1038 ^ 1'b0 ;
  assign n11729 = ( ~n11720 & n11723 ) | ( ~n11720 & n11728 ) | ( n11723 & n11728 ) ;
  assign n11730 = n5092 ^ n3721 ^ 1'b0 ;
  assign n11731 = n11730 ^ n3771 ^ 1'b0 ;
  assign n11732 = n11731 ^ n10275 ^ n4009 ;
  assign n11735 = ( ~n2148 & n3264 ) | ( ~n2148 & n6541 ) | ( n3264 & n6541 ) ;
  assign n11736 = n10780 & n11735 ;
  assign n11733 = ( n1674 & n1686 ) | ( n1674 & n7652 ) | ( n1686 & n7652 ) ;
  assign n11734 = n11733 ^ n9814 ^ n3596 ;
  assign n11737 = n11736 ^ n11734 ^ n5191 ;
  assign n11739 = n5197 ^ n3387 ^ n2929 ;
  assign n11740 = ( n5740 & n5845 ) | ( n5740 & n11739 ) | ( n5845 & n11739 ) ;
  assign n11738 = ~n6532 & n7302 ;
  assign n11741 = n11740 ^ n11738 ^ n5515 ;
  assign n11742 = ( n1562 & n11737 ) | ( n1562 & n11741 ) | ( n11737 & n11741 ) ;
  assign n11743 = n5538 & ~n11313 ;
  assign n11744 = n11743 ^ n5217 ^ 1'b0 ;
  assign n11745 = n11744 ^ n9229 ^ n9094 ;
  assign n11746 = n9330 ^ n5747 ^ n2136 ;
  assign n11747 = ( n7769 & n7930 ) | ( n7769 & n11746 ) | ( n7930 & n11746 ) ;
  assign n11748 = n1947 | n6485 ;
  assign n11749 = n1140 | n11748 ;
  assign n11750 = ( n5434 & n8180 ) | ( n5434 & n11749 ) | ( n8180 & n11749 ) ;
  assign n11751 = ( n2076 & n5201 ) | ( n2076 & ~n11750 ) | ( n5201 & ~n11750 ) ;
  assign n11752 = n11337 ^ n3442 ^ n2795 ;
  assign n11753 = n11752 ^ n7349 ^ n4805 ;
  assign n11754 = ( ~n2429 & n4235 ) | ( ~n2429 & n11693 ) | ( n4235 & n11693 ) ;
  assign n11755 = n11754 ^ n10529 ^ n3692 ;
  assign n11756 = n9535 ^ n3078 ^ 1'b0 ;
  assign n11757 = n3078 | n11756 ;
  assign n11758 = n7274 ^ n4204 ^ n2267 ;
  assign n11759 = n4514 ^ n3613 ^ 1'b0 ;
  assign n11760 = n4962 & n11759 ;
  assign n11761 = ( n1407 & n2703 ) | ( n1407 & n7639 ) | ( n2703 & n7639 ) ;
  assign n11762 = ( n10418 & n11760 ) | ( n10418 & ~n11761 ) | ( n11760 & ~n11761 ) ;
  assign n11763 = ( n3322 & ~n8645 ) | ( n3322 & n11762 ) | ( ~n8645 & n11762 ) ;
  assign n11764 = ( n3372 & n8483 ) | ( n3372 & ~n11763 ) | ( n8483 & ~n11763 ) ;
  assign n11765 = ( n7832 & n11758 ) | ( n7832 & ~n11764 ) | ( n11758 & ~n11764 ) ;
  assign n11766 = n11765 ^ n7599 ^ 1'b0 ;
  assign n11767 = n2097 & n11766 ;
  assign n11776 = n9029 ^ n401 ^ 1'b0 ;
  assign n11777 = ( n7372 & n7932 ) | ( n7372 & ~n11776 ) | ( n7932 & ~n11776 ) ;
  assign n11768 = n11313 ^ n10578 ^ n5673 ;
  assign n11772 = n8505 ^ n5884 ^ n5756 ;
  assign n11769 = n9519 ^ n1749 ^ 1'b0 ;
  assign n11770 = n6004 & ~n6807 ;
  assign n11771 = ~n11769 & n11770 ;
  assign n11773 = n11772 ^ n11771 ^ 1'b0 ;
  assign n11774 = ( ~n9814 & n11768 ) | ( ~n9814 & n11773 ) | ( n11768 & n11773 ) ;
  assign n11775 = ( ~n8298 & n8461 ) | ( ~n8298 & n11774 ) | ( n8461 & n11774 ) ;
  assign n11778 = n11777 ^ n11775 ^ n3581 ;
  assign n11779 = n6863 & n11381 ;
  assign n11780 = n706 & n11779 ;
  assign n11781 = n6023 ^ n1920 ^ 1'b0 ;
  assign n11782 = ~n2152 & n11781 ;
  assign n11783 = ( n1337 & ~n3545 ) | ( n1337 & n6403 ) | ( ~n3545 & n6403 ) ;
  assign n11784 = n4148 | n11783 ;
  assign n11785 = n11784 ^ n210 ^ 1'b0 ;
  assign n11786 = ( n3612 & n11555 ) | ( n3612 & n11785 ) | ( n11555 & n11785 ) ;
  assign n11787 = n11786 ^ n11639 ^ 1'b0 ;
  assign n11788 = n11782 & ~n11787 ;
  assign n11789 = ( n2552 & ~n6425 ) | ( n2552 & n10618 ) | ( ~n6425 & n10618 ) ;
  assign n11790 = ( ~n6991 & n10393 ) | ( ~n6991 & n11789 ) | ( n10393 & n11789 ) ;
  assign n11791 = ~n6640 & n11790 ;
  assign n11792 = n9124 ^ n3074 ^ 1'b0 ;
  assign n11793 = ( n8935 & n9896 ) | ( n8935 & n11792 ) | ( n9896 & n11792 ) ;
  assign n11794 = n10175 ^ n9517 ^ n1672 ;
  assign n11795 = ( n1393 & n7966 ) | ( n1393 & ~n11794 ) | ( n7966 & ~n11794 ) ;
  assign n11796 = n9616 ^ n5295 ^ 1'b0 ;
  assign n11797 = n2864 ^ n929 ^ 1'b0 ;
  assign n11798 = ( ~x13 & n1079 ) | ( ~x13 & n10908 ) | ( n1079 & n10908 ) ;
  assign n11799 = ( n4374 & n11797 ) | ( n4374 & ~n11798 ) | ( n11797 & ~n11798 ) ;
  assign n11800 = ( n1866 & n3214 ) | ( n1866 & n11799 ) | ( n3214 & n11799 ) ;
  assign n11801 = n11800 ^ n9025 ^ n2942 ;
  assign n11802 = n917 & ~n2579 ;
  assign n11803 = n7040 & n11802 ;
  assign n11807 = ( n729 & n2932 ) | ( n729 & n6429 ) | ( n2932 & n6429 ) ;
  assign n11804 = n4038 ^ n2188 ^ n554 ;
  assign n11805 = ( n1328 & ~n2824 ) | ( n1328 & n4536 ) | ( ~n2824 & n4536 ) ;
  assign n11806 = ( ~n7670 & n11804 ) | ( ~n7670 & n11805 ) | ( n11804 & n11805 ) ;
  assign n11808 = n11807 ^ n11806 ^ n3866 ;
  assign n11809 = n11116 ^ n4750 ^ n2417 ;
  assign n11810 = ( x40 & ~n3721 ) | ( x40 & n5858 ) | ( ~n3721 & n5858 ) ;
  assign n11811 = n6211 & n11810 ;
  assign n11812 = n10163 & n11811 ;
  assign n11813 = ( n8297 & n11809 ) | ( n8297 & n11812 ) | ( n11809 & n11812 ) ;
  assign n11814 = ( n2413 & ~n8300 ) | ( n2413 & n11097 ) | ( ~n8300 & n11097 ) ;
  assign n11815 = ~n6689 & n11814 ;
  assign n11816 = n11815 ^ n337 ^ 1'b0 ;
  assign n11817 = n10170 ^ n8437 ^ 1'b0 ;
  assign n11818 = ( n5695 & n7207 ) | ( n5695 & ~n7855 ) | ( n7207 & ~n7855 ) ;
  assign n11819 = ( n1112 & ~n5734 ) | ( n1112 & n7240 ) | ( ~n5734 & n7240 ) ;
  assign n11820 = n10649 ^ n5715 ^ 1'b0 ;
  assign n11821 = ( ~n3288 & n8947 ) | ( ~n3288 & n11820 ) | ( n8947 & n11820 ) ;
  assign n11822 = ~n3754 & n7234 ;
  assign n11823 = n7525 & n11822 ;
  assign n11824 = n11193 ^ n9914 ^ n4622 ;
  assign n11825 = ( ~n446 & n1862 ) | ( ~n446 & n2712 ) | ( n1862 & n2712 ) ;
  assign n11826 = ( n962 & n2557 ) | ( n962 & n11825 ) | ( n2557 & n11825 ) ;
  assign n11827 = n11826 ^ n6405 ^ n4847 ;
  assign n11828 = ( n3500 & n4025 ) | ( n3500 & n9474 ) | ( n4025 & n9474 ) ;
  assign n11829 = ( n1299 & n1615 ) | ( n1299 & ~n11828 ) | ( n1615 & ~n11828 ) ;
  assign n11830 = n2717 & n7303 ;
  assign n11831 = ( n11012 & n11829 ) | ( n11012 & ~n11830 ) | ( n11829 & ~n11830 ) ;
  assign n11832 = n11831 ^ n371 ^ 1'b0 ;
  assign n11833 = n8933 & n11832 ;
  assign n11842 = n2456 ^ n2219 ^ n1388 ;
  assign n11843 = n5094 & n11842 ;
  assign n11834 = ~n1003 & n1167 ;
  assign n11835 = n7536 & n11834 ;
  assign n11836 = x29 & ~n3041 ;
  assign n11837 = n11836 ^ n5658 ^ 1'b0 ;
  assign n11838 = ( ~n10545 & n11835 ) | ( ~n10545 & n11837 ) | ( n11835 & n11837 ) ;
  assign n11839 = ( ~x41 & n7480 ) | ( ~x41 & n11838 ) | ( n7480 & n11838 ) ;
  assign n11840 = n11839 ^ n11637 ^ n8228 ;
  assign n11841 = ( n2347 & n11250 ) | ( n2347 & n11840 ) | ( n11250 & n11840 ) ;
  assign n11844 = n11843 ^ n11841 ^ n9760 ;
  assign n11845 = ( n3431 & n3687 ) | ( n3431 & ~n11844 ) | ( n3687 & ~n11844 ) ;
  assign n11846 = n5765 & ~n7912 ;
  assign n11847 = n8191 ^ n592 ^ 1'b0 ;
  assign n11848 = n11847 ^ n7008 ^ n1220 ;
  assign n11849 = n5228 ^ n5189 ^ n3377 ;
  assign n11850 = n11849 ^ n10277 ^ n2286 ;
  assign n11851 = n1197 & ~n11850 ;
  assign n11852 = n11851 ^ n2378 ^ 1'b0 ;
  assign n11860 = n10823 ^ n3717 ^ n3090 ;
  assign n11861 = n11860 ^ n11385 ^ n2002 ;
  assign n11857 = n5209 ^ x71 ^ 1'b0 ;
  assign n11858 = n11857 ^ n2408 ^ n1053 ;
  assign n11859 = n11858 ^ n3891 ^ n980 ;
  assign n11853 = n1109 | n5475 ;
  assign n11854 = n11853 ^ n6524 ^ n1260 ;
  assign n11855 = n11854 ^ n8219 ^ 1'b0 ;
  assign n11856 = ~n4624 & n11855 ;
  assign n11862 = n11861 ^ n11859 ^ n11856 ;
  assign n11863 = ( n3654 & n11852 ) | ( n3654 & n11862 ) | ( n11852 & n11862 ) ;
  assign n11864 = n3791 ^ n2813 ^ 1'b0 ;
  assign n11865 = n5216 | n7365 ;
  assign n11866 = n11864 & ~n11865 ;
  assign n11870 = ~n1583 & n3611 ;
  assign n11867 = n2170 | n2511 ;
  assign n11868 = n791 & ~n11867 ;
  assign n11869 = n9585 | n11868 ;
  assign n11871 = n11870 ^ n11869 ^ n11107 ;
  assign n11872 = ( n9132 & ~n11866 ) | ( n9132 & n11871 ) | ( ~n11866 & n11871 ) ;
  assign n11874 = ( n530 & n4521 ) | ( n530 & ~n7518 ) | ( n4521 & ~n7518 ) ;
  assign n11873 = ( n3995 & ~n8456 ) | ( n3995 & n10685 ) | ( ~n8456 & n10685 ) ;
  assign n11875 = n11874 ^ n11873 ^ 1'b0 ;
  assign n11876 = n10622 & n11875 ;
  assign n11877 = n9095 ^ n4996 ^ n3357 ;
  assign n11878 = n659 & n959 ;
  assign n11879 = n2714 ^ n1964 ^ x123 ;
  assign n11880 = n3491 ^ n2785 ^ n582 ;
  assign n11881 = n11880 ^ n6606 ^ n5569 ;
  assign n11882 = ( n2962 & ~n11879 ) | ( n2962 & n11881 ) | ( ~n11879 & n11881 ) ;
  assign n11883 = ( n6965 & n11878 ) | ( n6965 & n11882 ) | ( n11878 & n11882 ) ;
  assign n11884 = n11810 ^ n4875 ^ n4282 ;
  assign n11885 = ( n1077 & ~n1323 ) | ( n1077 & n6837 ) | ( ~n1323 & n6837 ) ;
  assign n11886 = n2256 | n7442 ;
  assign n11887 = n11885 | n11886 ;
  assign n11888 = n11138 ^ n10003 ^ n4433 ;
  assign n11889 = ( n4914 & n11346 ) | ( n4914 & n11888 ) | ( n11346 & n11888 ) ;
  assign n11890 = n4054 ^ n1850 ^ n1320 ;
  assign n11891 = n2206 & n6255 ;
  assign n11892 = n11298 ^ n1346 ^ 1'b0 ;
  assign n11893 = ~n11891 & n11892 ;
  assign n11894 = n11893 ^ n4392 ^ n4087 ;
  assign n11895 = ( n7734 & n11890 ) | ( n7734 & n11894 ) | ( n11890 & n11894 ) ;
  assign n11896 = n8725 ^ n7990 ^ n2373 ;
  assign n11897 = ( n6127 & n11895 ) | ( n6127 & ~n11896 ) | ( n11895 & ~n11896 ) ;
  assign n11898 = n11897 ^ n9816 ^ 1'b0 ;
  assign n11899 = ~n11889 & n11898 ;
  assign n11900 = ( n6622 & n11887 ) | ( n6622 & ~n11899 ) | ( n11887 & ~n11899 ) ;
  assign n11901 = ( n1871 & ~n7785 ) | ( n1871 & n9484 ) | ( ~n7785 & n9484 ) ;
  assign n11902 = n11901 ^ n1768 ^ 1'b0 ;
  assign n11903 = n11902 ^ n7981 ^ n1415 ;
  assign n11904 = n11062 ^ n7577 ^ n1729 ;
  assign n11911 = n10263 ^ n5378 ^ n1270 ;
  assign n11912 = ( n3237 & ~n5064 ) | ( n3237 & n11911 ) | ( ~n5064 & n11911 ) ;
  assign n11913 = ( n1139 & ~n2101 ) | ( n1139 & n11912 ) | ( ~n2101 & n11912 ) ;
  assign n11914 = ( n2504 & n9080 ) | ( n2504 & ~n11913 ) | ( n9080 & ~n11913 ) ;
  assign n11905 = ~n1462 & n5902 ;
  assign n11906 = ~n3554 & n11905 ;
  assign n11907 = n11847 ^ n7978 ^ n6111 ;
  assign n11908 = ( n10356 & n10402 ) | ( n10356 & ~n11907 ) | ( n10402 & ~n11907 ) ;
  assign n11909 = ( ~n1686 & n6479 ) | ( ~n1686 & n11908 ) | ( n6479 & n11908 ) ;
  assign n11910 = ( ~n8857 & n11906 ) | ( ~n8857 & n11909 ) | ( n11906 & n11909 ) ;
  assign n11915 = n11914 ^ n11910 ^ n469 ;
  assign n11916 = ~n3593 & n8365 ;
  assign n11917 = n11916 ^ n6492 ^ n3468 ;
  assign n11918 = n5113 & n6631 ;
  assign n11919 = ~n4780 & n11918 ;
  assign n11920 = n11917 | n11919 ;
  assign n11921 = ( n605 & ~n7595 ) | ( n605 & n10199 ) | ( ~n7595 & n10199 ) ;
  assign n11922 = ( n6610 & n6928 ) | ( n6610 & ~n8606 ) | ( n6928 & ~n8606 ) ;
  assign n11923 = ( n2369 & ~n5644 ) | ( n2369 & n7858 ) | ( ~n5644 & n7858 ) ;
  assign n11925 = n6034 ^ n1712 ^ n191 ;
  assign n11924 = ( ~n1803 & n9545 ) | ( ~n1803 & n10955 ) | ( n9545 & n10955 ) ;
  assign n11926 = n11925 ^ n11924 ^ n2209 ;
  assign n11927 = n11926 ^ n4897 ^ n2010 ;
  assign n11928 = ( n1128 & n9364 ) | ( n1128 & ~n11927 ) | ( n9364 & ~n11927 ) ;
  assign n11929 = ( n7749 & n11923 ) | ( n7749 & n11928 ) | ( n11923 & n11928 ) ;
  assign n11930 = n10263 ^ n4540 ^ 1'b0 ;
  assign n11931 = n6876 ^ n3686 ^ 1'b0 ;
  assign n11932 = ( ~n5234 & n11930 ) | ( ~n5234 & n11931 ) | ( n11930 & n11931 ) ;
  assign n11933 = ( n4916 & n9145 ) | ( n4916 & ~n9650 ) | ( n9145 & ~n9650 ) ;
  assign n11934 = n11933 ^ n11718 ^ n1776 ;
  assign n11935 = n2185 & n6794 ;
  assign n11936 = n5536 & n11935 ;
  assign n11937 = n542 | n11936 ;
  assign n11938 = n11937 ^ n2969 ^ 1'b0 ;
  assign n11939 = n9517 ^ n8100 ^ n1452 ;
  assign n11940 = ~n7027 & n11939 ;
  assign n11941 = n9315 & n11940 ;
  assign n11942 = ( ~n3564 & n5050 ) | ( ~n3564 & n11941 ) | ( n5050 & n11941 ) ;
  assign n11943 = n5198 & n11942 ;
  assign n11944 = n1520 & n7785 ;
  assign n11945 = n11944 ^ n3559 ^ 1'b0 ;
  assign n11946 = ( n2838 & n4621 ) | ( n2838 & n11945 ) | ( n4621 & n11945 ) ;
  assign n11947 = n11685 ^ n1442 ^ n535 ;
  assign n11948 = ( ~n676 & n2861 ) | ( ~n676 & n6056 ) | ( n2861 & n6056 ) ;
  assign n11949 = n7651 | n11948 ;
  assign n11953 = n2262 | n6765 ;
  assign n11950 = ( n263 & n1919 ) | ( n263 & ~n2010 ) | ( n1919 & ~n2010 ) ;
  assign n11951 = n5725 ^ n4631 ^ n2967 ;
  assign n11952 = n11950 & n11951 ;
  assign n11954 = n11953 ^ n11952 ^ n4089 ;
  assign n11955 = ( ~n1299 & n2596 ) | ( ~n1299 & n4757 ) | ( n2596 & n4757 ) ;
  assign n11956 = ~n1633 & n11955 ;
  assign n11957 = n11956 ^ n10131 ^ n6862 ;
  assign n11958 = n3060 ^ n2248 ^ n1754 ;
  assign n11959 = ( n352 & ~n5669 ) | ( n352 & n11958 ) | ( ~n5669 & n11958 ) ;
  assign n11960 = n700 & ~n11959 ;
  assign n11961 = ( n1870 & n2923 ) | ( n1870 & n3526 ) | ( n2923 & n3526 ) ;
  assign n11962 = ( n4160 & ~n7647 ) | ( n4160 & n11961 ) | ( ~n7647 & n11961 ) ;
  assign n11966 = n276 ^ n139 ^ 1'b0 ;
  assign n11967 = n399 & ~n11966 ;
  assign n11965 = ~n2466 & n4096 ;
  assign n11963 = n8150 ^ n2560 ^ n1726 ;
  assign n11964 = ( n2386 & ~n4451 ) | ( n2386 & n11963 ) | ( ~n4451 & n11963 ) ;
  assign n11968 = n11967 ^ n11965 ^ n11964 ;
  assign n11969 = ( n985 & n1183 ) | ( n985 & ~n1720 ) | ( n1183 & ~n1720 ) ;
  assign n11970 = ( n3739 & ~n4582 ) | ( n3739 & n11024 ) | ( ~n4582 & n11024 ) ;
  assign n11971 = n11970 ^ n1460 ^ 1'b0 ;
  assign n11972 = ( n3023 & n11969 ) | ( n3023 & ~n11971 ) | ( n11969 & ~n11971 ) ;
  assign n11973 = n6725 ^ n3642 ^ n565 ;
  assign n11975 = n9219 ^ n9182 ^ n1284 ;
  assign n11976 = n11975 ^ n1591 ^ n1523 ;
  assign n11974 = n6768 ^ n4359 ^ n3928 ;
  assign n11977 = n11976 ^ n11974 ^ n11555 ;
  assign n11978 = ( n847 & ~n4068 ) | ( n847 & n4189 ) | ( ~n4068 & n4189 ) ;
  assign n11979 = ( n1426 & n4059 ) | ( n1426 & n10886 ) | ( n4059 & n10886 ) ;
  assign n11980 = ~n2958 & n6962 ;
  assign n11981 = n7447 & n11980 ;
  assign n11984 = ( n903 & n8584 ) | ( n903 & n8718 ) | ( n8584 & n8718 ) ;
  assign n11985 = n11984 ^ n997 ^ 1'b0 ;
  assign n11986 = ( ~n6092 & n6475 ) | ( ~n6092 & n11985 ) | ( n6475 & n11985 ) ;
  assign n11982 = n7678 ^ n4426 ^ n1907 ;
  assign n11983 = n11982 ^ n4129 ^ n1026 ;
  assign n11987 = n11986 ^ n11983 ^ 1'b0 ;
  assign n11988 = ( ~n11979 & n11981 ) | ( ~n11979 & n11987 ) | ( n11981 & n11987 ) ;
  assign n11989 = n6044 ^ n1036 ^ n566 ;
  assign n11990 = ( n4862 & n9780 ) | ( n4862 & ~n10783 ) | ( n9780 & ~n10783 ) ;
  assign n11991 = n452 | n6698 ;
  assign n11992 = n3862 | n11991 ;
  assign n11993 = ( ~n4039 & n11990 ) | ( ~n4039 & n11992 ) | ( n11990 & n11992 ) ;
  assign n11994 = n9730 ^ n3014 ^ n1978 ;
  assign n11995 = n11473 ^ n5270 ^ n3131 ;
  assign n11996 = n4604 ^ n2931 ^ n2761 ;
  assign n11997 = n11996 ^ n11772 ^ n10828 ;
  assign n12003 = ~n7301 & n11147 ;
  assign n12000 = ( n1147 & n1545 ) | ( n1147 & ~n1618 ) | ( n1545 & ~n1618 ) ;
  assign n12001 = ( n5603 & n7335 ) | ( n5603 & n12000 ) | ( n7335 & n12000 ) ;
  assign n12002 = n12001 ^ n3619 ^ n3599 ;
  assign n11998 = n3181 ^ n1523 ^ n345 ;
  assign n11999 = n11998 ^ n7796 ^ n5827 ;
  assign n12004 = n12003 ^ n12002 ^ n11999 ;
  assign n12005 = n10008 ^ n8567 ^ 1'b0 ;
  assign n12006 = n7515 & n12005 ;
  assign n12007 = n12006 ^ n5969 ^ n270 ;
  assign n12008 = ( ~n314 & n1898 ) | ( ~n314 & n12007 ) | ( n1898 & n12007 ) ;
  assign n12009 = n12008 ^ n10668 ^ n3949 ;
  assign n12010 = n1336 | n6903 ;
  assign n12011 = n2378 & n7713 ;
  assign n12012 = n2709 & ~n4243 ;
  assign n12013 = n12012 ^ n3570 ^ 1'b0 ;
  assign n12014 = n2186 | n12013 ;
  assign n12015 = n12014 ^ n4820 ^ n3455 ;
  assign n12016 = ( n496 & n8153 ) | ( n496 & ~n12015 ) | ( n8153 & ~n12015 ) ;
  assign n12017 = n5828 ^ n4776 ^ n4485 ;
  assign n12018 = ( n2359 & n4761 ) | ( n2359 & ~n12017 ) | ( n4761 & ~n12017 ) ;
  assign n12019 = n12018 ^ n10536 ^ n5186 ;
  assign n12020 = ( ~n1901 & n10168 ) | ( ~n1901 & n12019 ) | ( n10168 & n12019 ) ;
  assign n12021 = n10012 | n12020 ;
  assign n12022 = ( ~n12011 & n12016 ) | ( ~n12011 & n12021 ) | ( n12016 & n12021 ) ;
  assign n12023 = n11418 ^ n10959 ^ 1'b0 ;
  assign n12027 = ( ~n780 & n1002 ) | ( ~n780 & n4045 ) | ( n1002 & n4045 ) ;
  assign n12026 = n7544 ^ n6327 ^ x47 ;
  assign n12024 = n3180 ^ n1072 ^ 1'b0 ;
  assign n12025 = ~n3618 & n12024 ;
  assign n12028 = n12027 ^ n12026 ^ n12025 ;
  assign n12029 = n2705 & n3731 ;
  assign n12030 = ( n282 & n2374 ) | ( n282 & ~n8653 ) | ( n2374 & ~n8653 ) ;
  assign n12031 = n12030 ^ n4503 ^ 1'b0 ;
  assign n12032 = n12029 | n12031 ;
  assign n12033 = n12032 ^ n9056 ^ n1397 ;
  assign n12034 = ( n8118 & n9730 ) | ( n8118 & ~n12033 ) | ( n9730 & ~n12033 ) ;
  assign n12037 = n4649 ^ n4602 ^ n403 ;
  assign n12036 = n11526 ^ n5694 ^ n3724 ;
  assign n12035 = x106 & ~n8168 ;
  assign n12038 = n12037 ^ n12036 ^ n12035 ;
  assign n12039 = ( ~n6572 & n10704 ) | ( ~n6572 & n12038 ) | ( n10704 & n12038 ) ;
  assign n12040 = n1587 | n12039 ;
  assign n12051 = ( n1373 & ~n2392 ) | ( n1373 & n10197 ) | ( ~n2392 & n10197 ) ;
  assign n12052 = ( n918 & n3939 ) | ( n918 & n12051 ) | ( n3939 & n12051 ) ;
  assign n12053 = n12052 ^ n10114 ^ 1'b0 ;
  assign n12054 = n571 | n12053 ;
  assign n12055 = ( n3614 & ~n7655 ) | ( n3614 & n12054 ) | ( ~n7655 & n12054 ) ;
  assign n12045 = n7117 ^ n6900 ^ n3442 ;
  assign n12046 = n12045 ^ n8541 ^ n3985 ;
  assign n12047 = n4910 ^ n2133 ^ x99 ;
  assign n12048 = ( n2927 & ~n11552 ) | ( n2927 & n12047 ) | ( ~n11552 & n12047 ) ;
  assign n12049 = ( n479 & n8156 ) | ( n479 & n12048 ) | ( n8156 & n12048 ) ;
  assign n12050 = ( n5262 & n12046 ) | ( n5262 & ~n12049 ) | ( n12046 & ~n12049 ) ;
  assign n12041 = n4582 ^ n3530 ^ n393 ;
  assign n12042 = n6384 ^ n6032 ^ n5853 ;
  assign n12043 = ( n1477 & n2929 ) | ( n1477 & n12042 ) | ( n2929 & n12042 ) ;
  assign n12044 = n12041 & ~n12043 ;
  assign n12056 = n12055 ^ n12050 ^ n12044 ;
  assign n12057 = ~n1198 & n1897 ;
  assign n12059 = ( x65 & n4422 ) | ( x65 & n7033 ) | ( n4422 & n7033 ) ;
  assign n12058 = ~n2733 & n6768 ;
  assign n12060 = n12059 ^ n12058 ^ 1'b0 ;
  assign n12061 = n12057 & ~n12060 ;
  assign n12062 = n12061 ^ n912 ^ n508 ;
  assign n12063 = n8212 ^ n2706 ^ n2246 ;
  assign n12064 = n12063 ^ n3712 ^ n634 ;
  assign n12065 = ( x16 & ~n2220 ) | ( x16 & n10008 ) | ( ~n2220 & n10008 ) ;
  assign n12066 = ( n1432 & n1985 ) | ( n1432 & n3794 ) | ( n1985 & n3794 ) ;
  assign n12067 = ( ~n4210 & n6317 ) | ( ~n4210 & n12066 ) | ( n6317 & n12066 ) ;
  assign n12068 = ( n2219 & ~n12065 ) | ( n2219 & n12067 ) | ( ~n12065 & n12067 ) ;
  assign n12069 = n12068 ^ n664 ^ 1'b0 ;
  assign n12070 = ( ~n3403 & n5149 ) | ( ~n3403 & n6537 ) | ( n5149 & n6537 ) ;
  assign n12071 = ( n3929 & ~n5396 ) | ( n3929 & n12070 ) | ( ~n5396 & n12070 ) ;
  assign n12072 = ( ~n2650 & n4301 ) | ( ~n2650 & n12071 ) | ( n4301 & n12071 ) ;
  assign n12073 = ( ~n732 & n3795 ) | ( ~n732 & n12072 ) | ( n3795 & n12072 ) ;
  assign n12074 = n12073 ^ n3916 ^ 1'b0 ;
  assign n12075 = n9046 ^ n4518 ^ n442 ;
  assign n12076 = ( n5833 & ~n9548 ) | ( n5833 & n12075 ) | ( ~n9548 & n12075 ) ;
  assign n12077 = ( n748 & n1008 ) | ( n748 & n8460 ) | ( n1008 & n8460 ) ;
  assign n12078 = ( n4338 & n5656 ) | ( n4338 & ~n12077 ) | ( n5656 & ~n12077 ) ;
  assign n12079 = n12078 ^ n325 ^ 1'b0 ;
  assign n12080 = n12076 | n12079 ;
  assign n12083 = n390 | n11739 ;
  assign n12084 = n1255 & ~n12083 ;
  assign n12081 = ( n1410 & ~n3030 ) | ( n1410 & n3104 ) | ( ~n3030 & n3104 ) ;
  assign n12082 = n9024 & ~n12081 ;
  assign n12085 = n12084 ^ n12082 ^ n2491 ;
  assign n12086 = ~n11941 & n12085 ;
  assign n12091 = ( ~n2041 & n3107 ) | ( ~n2041 & n7032 ) | ( n3107 & n7032 ) ;
  assign n12092 = ( ~n818 & n2844 ) | ( ~n818 & n12091 ) | ( n2844 & n12091 ) ;
  assign n12087 = ( n373 & n1339 ) | ( n373 & n4660 ) | ( n1339 & n4660 ) ;
  assign n12088 = n12087 ^ n5432 ^ n1550 ;
  assign n12089 = ( n4622 & n5216 ) | ( n4622 & ~n12088 ) | ( n5216 & ~n12088 ) ;
  assign n12090 = n5466 & ~n12089 ;
  assign n12093 = n12092 ^ n12090 ^ 1'b0 ;
  assign n12094 = ( n2897 & n3670 ) | ( n2897 & n12093 ) | ( n3670 & n12093 ) ;
  assign n12095 = ( n1361 & ~n2254 ) | ( n1361 & n3986 ) | ( ~n2254 & n3986 ) ;
  assign n12096 = ( n5227 & ~n11500 ) | ( n5227 & n12095 ) | ( ~n11500 & n12095 ) ;
  assign n12097 = n12094 | n12096 ;
  assign n12098 = n12097 ^ n9064 ^ n2127 ;
  assign n12099 = n1701 ^ n1592 ^ 1'b0 ;
  assign n12100 = n6044 | n12099 ;
  assign n12101 = ( n5974 & ~n6738 ) | ( n5974 & n12100 ) | ( ~n6738 & n12100 ) ;
  assign n12103 = n5655 ^ n5304 ^ 1'b0 ;
  assign n12104 = n9143 | n12103 ;
  assign n12102 = ~n3756 & n4888 ;
  assign n12105 = n12104 ^ n12102 ^ n3533 ;
  assign n12107 = ( n3250 & ~n4257 ) | ( n3250 & n9474 ) | ( ~n4257 & n9474 ) ;
  assign n12106 = n8035 ^ n5860 ^ n1176 ;
  assign n12108 = n12107 ^ n12106 ^ n8225 ;
  assign n12115 = n5437 ^ n1520 ^ 1'b0 ;
  assign n12113 = ( n2029 & n4010 ) | ( n2029 & n6767 ) | ( n4010 & n6767 ) ;
  assign n12114 = n12113 ^ n7071 ^ n706 ;
  assign n12109 = ( n359 & n3105 ) | ( n359 & n4794 ) | ( n3105 & n4794 ) ;
  assign n12110 = ( x103 & ~n574 ) | ( x103 & n3516 ) | ( ~n574 & n3516 ) ;
  assign n12111 = n604 & ~n12110 ;
  assign n12112 = n12109 & n12111 ;
  assign n12116 = n12115 ^ n12114 ^ n12112 ;
  assign n12117 = ( n9049 & ~n10964 ) | ( n9049 & n12116 ) | ( ~n10964 & n12116 ) ;
  assign n12118 = ( n4144 & ~n6606 ) | ( n4144 & n10321 ) | ( ~n6606 & n10321 ) ;
  assign n12124 = n9399 ^ n8302 ^ n2775 ;
  assign n12125 = ( n5227 & ~n10674 ) | ( n5227 & n12124 ) | ( ~n10674 & n12124 ) ;
  assign n12119 = ( n233 & ~n2908 ) | ( n233 & n3741 ) | ( ~n2908 & n3741 ) ;
  assign n12120 = ( ~n719 & n5060 ) | ( ~n719 & n12119 ) | ( n5060 & n12119 ) ;
  assign n12121 = ( n818 & n2814 ) | ( n818 & n3327 ) | ( n2814 & n3327 ) ;
  assign n12122 = n12120 & ~n12121 ;
  assign n12123 = ~n2351 & n12122 ;
  assign n12126 = n12125 ^ n12123 ^ n3137 ;
  assign n12127 = ( n2317 & n5898 ) | ( n2317 & n12126 ) | ( n5898 & n12126 ) ;
  assign n12129 = n11014 ^ n10591 ^ n933 ;
  assign n12128 = ( n252 & n5569 ) | ( n252 & n8520 ) | ( n5569 & n8520 ) ;
  assign n12130 = n12129 ^ n12128 ^ n7152 ;
  assign n12131 = n12130 ^ n3365 ^ n2391 ;
  assign n12141 = n10680 ^ n8028 ^ 1'b0 ;
  assign n12136 = n11628 ^ n8064 ^ n4039 ;
  assign n12137 = n2245 & ~n12136 ;
  assign n12138 = n12137 ^ n10729 ^ 1'b0 ;
  assign n12139 = ~n801 & n12138 ;
  assign n12140 = n12139 ^ n11790 ^ n6158 ;
  assign n12132 = ( ~n293 & n3090 ) | ( ~n293 & n4128 ) | ( n3090 & n4128 ) ;
  assign n12133 = n12132 ^ n11270 ^ n3956 ;
  assign n12134 = ( n2875 & n4050 ) | ( n2875 & ~n12133 ) | ( n4050 & ~n12133 ) ;
  assign n12135 = n12134 ^ n5763 ^ n3525 ;
  assign n12142 = n12141 ^ n12140 ^ n12135 ;
  assign n12143 = n12142 ^ n11961 ^ n4929 ;
  assign n12144 = ( n6111 & n10934 ) | ( n6111 & n12143 ) | ( n10934 & n12143 ) ;
  assign n12150 = ( n205 & n10197 ) | ( n205 & n11540 ) | ( n10197 & n11540 ) ;
  assign n12149 = n8205 ^ n3689 ^ n656 ;
  assign n12147 = ( n3557 & n5647 ) | ( n3557 & ~n10472 ) | ( n5647 & ~n10472 ) ;
  assign n12145 = n7550 ^ n4042 ^ n736 ;
  assign n12146 = ( n1635 & n7502 ) | ( n1635 & ~n12145 ) | ( n7502 & ~n12145 ) ;
  assign n12148 = n12147 ^ n12146 ^ n8462 ;
  assign n12151 = n12150 ^ n12149 ^ n12148 ;
  assign n12152 = n7569 ^ n4822 ^ 1'b0 ;
  assign n12153 = ( n3696 & n6986 ) | ( n3696 & ~n12152 ) | ( n6986 & ~n12152 ) ;
  assign n12161 = ( n2763 & n6413 ) | ( n2763 & n6598 ) | ( n6413 & n6598 ) ;
  assign n12156 = ( n186 & ~n3867 ) | ( n186 & n5942 ) | ( ~n3867 & n5942 ) ;
  assign n12157 = n12156 ^ n10744 ^ n4456 ;
  assign n12158 = ( n6516 & n8022 ) | ( n6516 & ~n12157 ) | ( n8022 & ~n12157 ) ;
  assign n12154 = ( n5516 & n6627 ) | ( n5516 & ~n8435 ) | ( n6627 & ~n8435 ) ;
  assign n12155 = ( n3196 & n4030 ) | ( n3196 & n12154 ) | ( n4030 & n12154 ) ;
  assign n12159 = n12158 ^ n12155 ^ 1'b0 ;
  assign n12160 = n6758 | n12159 ;
  assign n12162 = n12161 ^ n12160 ^ n3085 ;
  assign n12163 = ( n2280 & ~n2435 ) | ( n2280 & n10505 ) | ( ~n2435 & n10505 ) ;
  assign n12164 = n173 & ~n3308 ;
  assign n12165 = n3066 & n12164 ;
  assign n12166 = n12165 ^ n5666 ^ 1'b0 ;
  assign n12167 = ( ~n7009 & n12163 ) | ( ~n7009 & n12166 ) | ( n12163 & n12166 ) ;
  assign n12168 = n11026 ^ n4581 ^ 1'b0 ;
  assign n12169 = n12168 ^ n11064 ^ 1'b0 ;
  assign n12170 = n3012 & ~n12169 ;
  assign n12171 = n4956 ^ n3993 ^ n3189 ;
  assign n12172 = ( x94 & n3189 ) | ( x94 & ~n5767 ) | ( n3189 & ~n5767 ) ;
  assign n12173 = n12172 ^ n7469 ^ n2657 ;
  assign n12174 = ( n11454 & n12171 ) | ( n11454 & ~n12173 ) | ( n12171 & ~n12173 ) ;
  assign n12175 = n9529 ^ n4438 ^ n4168 ;
  assign n12177 = n6490 ^ n6391 ^ n858 ;
  assign n12176 = n10492 ^ n8298 ^ n1230 ;
  assign n12178 = n12177 ^ n12176 ^ n301 ;
  assign n12179 = n12178 ^ n6047 ^ n5672 ;
  assign n12180 = n503 & ~n6397 ;
  assign n12181 = ~n411 & n12180 ;
  assign n12182 = n7553 & ~n10669 ;
  assign n12183 = ~n2873 & n6105 ;
  assign n12184 = n12183 ^ n8323 ^ 1'b0 ;
  assign n12185 = n4358 & ~n12184 ;
  assign n12186 = n12182 & n12185 ;
  assign n12187 = n10688 ^ n8764 ^ n5379 ;
  assign n12188 = x4 & ~n2026 ;
  assign n12191 = n6598 ^ n4638 ^ 1'b0 ;
  assign n12189 = ( n1572 & n3931 ) | ( n1572 & n5613 ) | ( n3931 & n5613 ) ;
  assign n12190 = ( n1939 & n6604 ) | ( n1939 & ~n12189 ) | ( n6604 & ~n12189 ) ;
  assign n12192 = n12191 ^ n12190 ^ n195 ;
  assign n12193 = ( n7311 & n12188 ) | ( n7311 & n12192 ) | ( n12188 & n12192 ) ;
  assign n12194 = n11004 & ~n12193 ;
  assign n12195 = n12194 ^ n5901 ^ 1'b0 ;
  assign n12196 = ( n7676 & n11206 ) | ( n7676 & ~n12195 ) | ( n11206 & ~n12195 ) ;
  assign n12197 = n6630 ^ n1517 ^ n375 ;
  assign n12198 = n12197 ^ n2712 ^ 1'b0 ;
  assign n12199 = ~n5966 & n12198 ;
  assign n12200 = ( n3435 & ~n6624 ) | ( n3435 & n12199 ) | ( ~n6624 & n12199 ) ;
  assign n12201 = n10373 ^ n9247 ^ 1'b0 ;
  assign n12202 = n7877 ^ n6685 ^ 1'b0 ;
  assign n12203 = n12202 ^ n10670 ^ n4871 ;
  assign n12206 = n2787 ^ n1179 ^ n1165 ;
  assign n12204 = n1744 & ~n3560 ;
  assign n12205 = n12204 ^ n2843 ^ 1'b0 ;
  assign n12207 = n12206 ^ n12205 ^ 1'b0 ;
  assign n12208 = ~n12203 & n12207 ;
  assign n12209 = n1988 ^ n605 ^ 1'b0 ;
  assign n12210 = n9456 ^ n4496 ^ 1'b0 ;
  assign n12211 = n3190 ^ n1743 ^ n340 ;
  assign n12212 = n7768 & n12211 ;
  assign n12213 = ( ~n1390 & n3067 ) | ( ~n1390 & n8804 ) | ( n3067 & n8804 ) ;
  assign n12214 = n7094 & n12213 ;
  assign n12215 = n1562 & n12214 ;
  assign n12216 = n3679 ^ n3674 ^ n3459 ;
  assign n12217 = n12216 ^ n6596 ^ n6286 ;
  assign n12218 = ( n7652 & n8884 ) | ( n7652 & ~n10353 ) | ( n8884 & ~n10353 ) ;
  assign n12219 = n12218 ^ n6958 ^ 1'b0 ;
  assign n12220 = n4196 ^ n1793 ^ n1623 ;
  assign n12221 = ( n1144 & n10800 ) | ( n1144 & n12220 ) | ( n10800 & n12220 ) ;
  assign n12222 = ~n2116 & n7185 ;
  assign n12223 = n12222 ^ n10472 ^ 1'b0 ;
  assign n12232 = ( ~n2000 & n2347 ) | ( ~n2000 & n3082 ) | ( n2347 & n3082 ) ;
  assign n12225 = n7229 ^ n1486 ^ n433 ;
  assign n12226 = n4682 ^ n4344 ^ n337 ;
  assign n12227 = ~n10347 & n12226 ;
  assign n12228 = ~n6282 & n12227 ;
  assign n12229 = ( n12166 & n12225 ) | ( n12166 & ~n12228 ) | ( n12225 & ~n12228 ) ;
  assign n12230 = n12229 ^ n7118 ^ 1'b0 ;
  assign n12231 = n1062 | n12230 ;
  assign n12224 = n6458 ^ n757 ^ n404 ;
  assign n12233 = n12232 ^ n12231 ^ n12224 ;
  assign n12236 = n8446 ^ n5589 ^ n4801 ;
  assign n12234 = ( ~n974 & n3623 ) | ( ~n974 & n8770 ) | ( n3623 & n8770 ) ;
  assign n12235 = n12234 ^ n12148 ^ n4801 ;
  assign n12237 = n12236 ^ n12235 ^ n10446 ;
  assign n12238 = ( n393 & n3970 ) | ( n393 & ~n7990 ) | ( n3970 & ~n7990 ) ;
  assign n12239 = ( n691 & n9486 ) | ( n691 & n12238 ) | ( n9486 & n12238 ) ;
  assign n12240 = n4761 ^ n4417 ^ n146 ;
  assign n12241 = n4184 ^ n2696 ^ n2065 ;
  assign n12242 = n11066 ^ n5294 ^ n4712 ;
  assign n12243 = ( ~n381 & n7176 ) | ( ~n381 & n7756 ) | ( n7176 & n7756 ) ;
  assign n12244 = ( ~n12241 & n12242 ) | ( ~n12241 & n12243 ) | ( n12242 & n12243 ) ;
  assign n12245 = ~n12240 & n12244 ;
  assign n12246 = n9731 ^ n9119 ^ n2732 ;
  assign n12247 = n12246 ^ n9927 ^ n5156 ;
  assign n12248 = ( n2137 & n8881 ) | ( n2137 & ~n12247 ) | ( n8881 & ~n12247 ) ;
  assign n12249 = n8777 ^ n3352 ^ n1876 ;
  assign n12250 = n10429 ^ n7879 ^ n1721 ;
  assign n12252 = ( ~n1207 & n4380 ) | ( ~n1207 & n6575 ) | ( n4380 & n6575 ) ;
  assign n12253 = ( ~n3117 & n6168 ) | ( ~n3117 & n12252 ) | ( n6168 & n12252 ) ;
  assign n12251 = n10073 ^ n9378 ^ n9008 ;
  assign n12254 = n12253 ^ n12251 ^ n10025 ;
  assign n12258 = n8101 ^ n6821 ^ n2748 ;
  assign n12259 = n4046 | n4369 ;
  assign n12260 = n10452 | n12259 ;
  assign n12261 = ( ~n11139 & n12258 ) | ( ~n11139 & n12260 ) | ( n12258 & n12260 ) ;
  assign n12255 = ( ~x24 & n272 ) | ( ~x24 & n3181 ) | ( n272 & n3181 ) ;
  assign n12256 = ( n1474 & n7148 ) | ( n1474 & n12255 ) | ( n7148 & n12255 ) ;
  assign n12257 = ( n646 & n9151 ) | ( n646 & n12256 ) | ( n9151 & n12256 ) ;
  assign n12262 = n12261 ^ n12257 ^ n1895 ;
  assign n12263 = n12262 ^ n8387 ^ n4301 ;
  assign n12264 = ( ~n1289 & n1842 ) | ( ~n1289 & n10131 ) | ( n1842 & n10131 ) ;
  assign n12265 = n6027 ^ n5860 ^ n1182 ;
  assign n12266 = n11467 | n12265 ;
  assign n12267 = n12264 & ~n12266 ;
  assign n12268 = n5868 | n7826 ;
  assign n12269 = n12267 & ~n12268 ;
  assign n12278 = n490 & ~n3397 ;
  assign n12279 = n12278 ^ n721 ^ 1'b0 ;
  assign n12280 = n12279 ^ n4787 ^ n1642 ;
  assign n12277 = n3964 ^ n3417 ^ 1'b0 ;
  assign n12281 = n12280 ^ n12277 ^ n6648 ;
  assign n12274 = n150 & n4557 ;
  assign n12275 = n2570 & n12274 ;
  assign n12276 = ( ~n1239 & n8205 ) | ( ~n1239 & n12275 ) | ( n8205 & n12275 ) ;
  assign n12270 = n5323 ^ n1825 ^ n1057 ;
  assign n12271 = n10413 & n12270 ;
  assign n12272 = n12271 ^ n2642 ^ 1'b0 ;
  assign n12273 = n12272 ^ n2563 ^ 1'b0 ;
  assign n12282 = n12281 ^ n12276 ^ n12273 ;
  assign n12283 = ( ~n7926 & n12269 ) | ( ~n7926 & n12282 ) | ( n12269 & n12282 ) ;
  assign n12284 = ( n677 & n1865 ) | ( n677 & ~n5703 ) | ( n1865 & ~n5703 ) ;
  assign n12285 = ( n789 & n1855 ) | ( n789 & n12284 ) | ( n1855 & n12284 ) ;
  assign n12286 = x15 & n3831 ;
  assign n12287 = ~n6142 & n12286 ;
  assign n12288 = n12287 ^ n10745 ^ 1'b0 ;
  assign n12289 = ( n5026 & n7769 ) | ( n5026 & ~n8521 ) | ( n7769 & ~n8521 ) ;
  assign n12290 = n6965 ^ n3117 ^ n448 ;
  assign n12291 = n9239 & ~n10945 ;
  assign n12292 = n12291 ^ n11234 ^ 1'b0 ;
  assign n12293 = ( ~n10595 & n12290 ) | ( ~n10595 & n12292 ) | ( n12290 & n12292 ) ;
  assign n12294 = n6395 ^ n1817 ^ n1494 ;
  assign n12295 = ( n1818 & ~n6118 ) | ( n1818 & n11233 ) | ( ~n6118 & n11233 ) ;
  assign n12296 = ( n8389 & n9705 ) | ( n8389 & ~n12295 ) | ( n9705 & ~n12295 ) ;
  assign n12297 = ( ~n1516 & n12294 ) | ( ~n1516 & n12296 ) | ( n12294 & n12296 ) ;
  assign n12298 = n9522 ^ n9279 ^ n4446 ;
  assign n12299 = ~n5771 & n6358 ;
  assign n12300 = n12299 ^ n10393 ^ 1'b0 ;
  assign n12301 = n3407 ^ n1003 ^ x64 ;
  assign n12302 = n12301 ^ n3581 ^ n2564 ;
  assign n12303 = ( n6099 & n11752 ) | ( n6099 & ~n12302 ) | ( n11752 & ~n12302 ) ;
  assign n12305 = ( n528 & n3469 ) | ( n528 & n5293 ) | ( n3469 & n5293 ) ;
  assign n12304 = n9719 ^ n8770 ^ n2207 ;
  assign n12306 = n12305 ^ n12304 ^ n1154 ;
  assign n12307 = n11480 ^ n4459 ^ n2186 ;
  assign n12308 = n10222 ^ n7412 ^ n2411 ;
  assign n12309 = n12308 ^ n6497 ^ n1468 ;
  assign n12310 = ( n1814 & n6252 ) | ( n1814 & ~n12309 ) | ( n6252 & ~n12309 ) ;
  assign n12317 = n5225 ^ n2991 ^ x90 ;
  assign n12314 = n4940 ^ n2446 ^ x90 ;
  assign n12315 = n12314 ^ n12182 ^ n2837 ;
  assign n12316 = n6884 & ~n12315 ;
  assign n12312 = ( ~n980 & n6253 ) | ( ~n980 & n7707 ) | ( n6253 & n7707 ) ;
  assign n12311 = n4805 ^ n2397 ^ n1085 ;
  assign n12313 = n12312 ^ n12311 ^ n9337 ;
  assign n12318 = n12317 ^ n12316 ^ n12313 ;
  assign n12319 = ( n5064 & n5137 ) | ( n5064 & n6024 ) | ( n5137 & n6024 ) ;
  assign n12320 = n6543 & n11601 ;
  assign n12321 = n1315 & n12320 ;
  assign n12322 = n10749 | n12321 ;
  assign n12323 = n12322 ^ n11356 ^ 1'b0 ;
  assign n12324 = ( n8463 & n12319 ) | ( n8463 & n12323 ) | ( n12319 & n12323 ) ;
  assign n12329 = ( n1431 & n3484 ) | ( n1431 & n12106 ) | ( n3484 & n12106 ) ;
  assign n12326 = n7077 ^ n6182 ^ n3478 ;
  assign n12327 = n12326 ^ n6698 ^ n130 ;
  assign n12325 = ~n2301 & n6452 ;
  assign n12328 = n12327 ^ n12325 ^ 1'b0 ;
  assign n12330 = n12329 ^ n12328 ^ n6480 ;
  assign n12331 = n2357 ^ n2330 ^ n1378 ;
  assign n12332 = n12331 ^ n6972 ^ n3640 ;
  assign n12333 = ( ~n4445 & n6790 ) | ( ~n4445 & n8300 ) | ( n6790 & n8300 ) ;
  assign n12334 = n4446 ^ n469 ^ 1'b0 ;
  assign n12338 = ( n812 & ~n9165 ) | ( n812 & n11572 ) | ( ~n9165 & n11572 ) ;
  assign n12336 = n11155 ^ n5262 ^ n2770 ;
  assign n12335 = n2916 & n9903 ;
  assign n12337 = n12336 ^ n12335 ^ 1'b0 ;
  assign n12339 = n12338 ^ n12337 ^ n8823 ;
  assign n12340 = n7536 ^ n2297 ^ n363 ;
  assign n12341 = n12340 ^ n6169 ^ n2335 ;
  assign n12344 = n5888 ^ n5562 ^ n4249 ;
  assign n12343 = ( ~n371 & n947 ) | ( ~n371 & n4165 ) | ( n947 & n4165 ) ;
  assign n12342 = n7266 ^ n5625 ^ n2935 ;
  assign n12345 = n12344 ^ n12343 ^ n12342 ;
  assign n12346 = n3362 ^ n1084 ^ n560 ;
  assign n12347 = ( n3587 & n4484 ) | ( n3587 & n5852 ) | ( n4484 & n5852 ) ;
  assign n12354 = ( n309 & n860 ) | ( n309 & ~n1982 ) | ( n860 & ~n1982 ) ;
  assign n12355 = ( n1429 & ~n3474 ) | ( n1429 & n12354 ) | ( ~n3474 & n12354 ) ;
  assign n12353 = ( n1223 & n5566 ) | ( n1223 & n8647 ) | ( n5566 & n8647 ) ;
  assign n12356 = n12355 ^ n12353 ^ 1'b0 ;
  assign n12348 = ( n3300 & ~n3953 ) | ( n3300 & n6055 ) | ( ~n3953 & n6055 ) ;
  assign n12349 = n193 & n12348 ;
  assign n12350 = n12349 ^ n6422 ^ 1'b0 ;
  assign n12351 = n12178 ^ n7983 ^ n5998 ;
  assign n12352 = n12350 & ~n12351 ;
  assign n12357 = n12356 ^ n12352 ^ 1'b0 ;
  assign n12358 = n582 & n859 ;
  assign n12359 = ( n1623 & ~n10508 ) | ( n1623 & n12358 ) | ( ~n10508 & n12358 ) ;
  assign n12360 = ~n437 & n12359 ;
  assign n12361 = n6970 ^ n6288 ^ n4668 ;
  assign n12362 = ~n5194 & n9900 ;
  assign n12363 = n12362 ^ n7923 ^ 1'b0 ;
  assign n12364 = n12363 ^ n9842 ^ n5036 ;
  assign n12365 = ( n4660 & n8083 ) | ( n4660 & ~n8194 ) | ( n8083 & ~n8194 ) ;
  assign n12366 = ( n312 & n3597 ) | ( n312 & n12365 ) | ( n3597 & n12365 ) ;
  assign n12369 = n8638 ^ n5063 ^ n454 ;
  assign n12367 = ( ~n963 & n2410 ) | ( ~n963 & n2997 ) | ( n2410 & n2997 ) ;
  assign n12368 = ( ~n1441 & n1893 ) | ( ~n1441 & n12367 ) | ( n1893 & n12367 ) ;
  assign n12370 = n12369 ^ n12368 ^ n8028 ;
  assign n12371 = ( n3691 & ~n8087 ) | ( n3691 & n12370 ) | ( ~n8087 & n12370 ) ;
  assign n12372 = n12371 ^ n8520 ^ n5023 ;
  assign n12376 = n5879 ^ n1856 ^ n513 ;
  assign n12377 = n12376 ^ n2064 ^ 1'b0 ;
  assign n12378 = n10546 ^ n8570 ^ 1'b0 ;
  assign n12379 = ~n12377 & n12378 ;
  assign n12374 = n6370 ^ n6077 ^ n5305 ;
  assign n12375 = n9811 & ~n12374 ;
  assign n12373 = ( ~n3373 & n6804 ) | ( ~n3373 & n7539 ) | ( n6804 & n7539 ) ;
  assign n12380 = n12379 ^ n12375 ^ n12373 ;
  assign n12381 = n3992 ^ n3154 ^ n302 ;
  assign n12382 = n12381 ^ n3459 ^ n1122 ;
  assign n12383 = n12382 ^ n3264 ^ 1'b0 ;
  assign n12386 = ( x94 & n1388 ) | ( x94 & ~n2612 ) | ( n1388 & ~n2612 ) ;
  assign n12387 = n12386 ^ n3211 ^ n2653 ;
  assign n12388 = ~n1578 & n12387 ;
  assign n12384 = n2591 ^ n1209 ^ 1'b0 ;
  assign n12385 = n1450 & n12384 ;
  assign n12389 = n12388 ^ n12385 ^ n6296 ;
  assign n12390 = n12289 & ~n12389 ;
  assign n12391 = ( n995 & n7408 ) | ( n995 & ~n12311 ) | ( n7408 & ~n12311 ) ;
  assign n12392 = n12391 ^ n12039 ^ n8490 ;
  assign n12393 = ( n3620 & n3630 ) | ( n3620 & ~n4275 ) | ( n3630 & ~n4275 ) ;
  assign n12394 = n2406 | n6840 ;
  assign n12395 = n12393 & ~n12394 ;
  assign n12396 = n790 & ~n3002 ;
  assign n12397 = n7930 ^ n5016 ^ n1292 ;
  assign n12398 = ( ~n12395 & n12396 ) | ( ~n12395 & n12397 ) | ( n12396 & n12397 ) ;
  assign n12399 = n8075 ^ n5828 ^ n1813 ;
  assign n12400 = ( n2039 & ~n8287 ) | ( n2039 & n8802 ) | ( ~n8287 & n8802 ) ;
  assign n12401 = ( n960 & ~n4448 ) | ( n960 & n12400 ) | ( ~n4448 & n12400 ) ;
  assign n12402 = ( ~n2657 & n3999 ) | ( ~n2657 & n12401 ) | ( n3999 & n12401 ) ;
  assign n12403 = n5793 ^ n1099 ^ 1'b0 ;
  assign n12404 = ( ~n9359 & n12402 ) | ( ~n9359 & n12403 ) | ( n12402 & n12403 ) ;
  assign n12406 = n6282 ^ n5368 ^ n4370 ;
  assign n12407 = n12406 ^ n6426 ^ n3435 ;
  assign n12405 = ( ~n542 & n1277 ) | ( ~n542 & n9035 ) | ( n1277 & n9035 ) ;
  assign n12408 = n12407 ^ n12405 ^ n8043 ;
  assign n12412 = n9633 ^ n5052 ^ n761 ;
  assign n12413 = n12412 ^ n8482 ^ n3389 ;
  assign n12409 = n5085 ^ n3123 ^ n1055 ;
  assign n12410 = n4091 | n6812 ;
  assign n12411 = n12409 | n12410 ;
  assign n12414 = n12413 ^ n12411 ^ n578 ;
  assign n12415 = n10924 ^ n8729 ^ 1'b0 ;
  assign n12416 = ( n2256 & n9374 ) | ( n2256 & n10224 ) | ( n9374 & n10224 ) ;
  assign n12417 = ( ~n6496 & n9426 ) | ( ~n6496 & n12416 ) | ( n9426 & n12416 ) ;
  assign n12418 = n12417 ^ n9478 ^ n7108 ;
  assign n12419 = n12418 ^ n7340 ^ n2373 ;
  assign n12420 = ( n12414 & ~n12415 ) | ( n12414 & n12419 ) | ( ~n12415 & n12419 ) ;
  assign n12423 = n4347 ^ n1341 ^ n288 ;
  assign n12421 = n1890 ^ x122 ^ 1'b0 ;
  assign n12422 = n12421 ^ n8828 ^ n1316 ;
  assign n12424 = n12423 ^ n12422 ^ n8847 ;
  assign n12441 = ( ~n1855 & n2488 ) | ( ~n1855 & n4052 ) | ( n2488 & n4052 ) ;
  assign n12442 = ( n1977 & n6748 ) | ( n1977 & ~n12441 ) | ( n6748 & ~n12441 ) ;
  assign n12443 = ( n1725 & n5646 ) | ( n1725 & n12442 ) | ( n5646 & n12442 ) ;
  assign n12436 = n1767 ^ n1212 ^ n1128 ;
  assign n12437 = ( ~n2069 & n8686 ) | ( ~n2069 & n12436 ) | ( n8686 & n12436 ) ;
  assign n12438 = ~n1790 & n12437 ;
  assign n12439 = n12438 ^ n7944 ^ 1'b0 ;
  assign n12431 = n1520 | n1983 ;
  assign n12432 = n12431 ^ n558 ^ 1'b0 ;
  assign n12433 = ( n2028 & ~n5384 ) | ( n2028 & n8199 ) | ( ~n5384 & n8199 ) ;
  assign n12434 = n12433 ^ n6901 ^ 1'b0 ;
  assign n12435 = n12432 | n12434 ;
  assign n12426 = n11391 ^ n3934 ^ n2486 ;
  assign n12427 = ~n3459 & n8863 ;
  assign n12428 = n4359 & n12427 ;
  assign n12429 = ( ~n3060 & n12426 ) | ( ~n3060 & n12428 ) | ( n12426 & n12428 ) ;
  assign n12425 = n4702 ^ n2241 ^ n1817 ;
  assign n12430 = n12429 ^ n12425 ^ n5458 ;
  assign n12440 = n12439 ^ n12435 ^ n12430 ;
  assign n12444 = n12443 ^ n12440 ^ n3484 ;
  assign n12445 = ( n6439 & n8982 ) | ( n6439 & ~n10545 ) | ( n8982 & ~n10545 ) ;
  assign n12446 = ( n2476 & ~n9397 ) | ( n2476 & n10393 ) | ( ~n9397 & n10393 ) ;
  assign n12447 = ( n388 & ~n864 ) | ( n388 & n920 ) | ( ~n864 & n920 ) ;
  assign n12448 = n12447 ^ n5761 ^ n1220 ;
  assign n12449 = ~n1897 & n12448 ;
  assign n12450 = n12449 ^ n2218 ^ n1645 ;
  assign n12451 = ( n619 & ~n1423 ) | ( n619 & n4285 ) | ( ~n1423 & n4285 ) ;
  assign n12452 = ( n6982 & n9945 ) | ( n6982 & n11332 ) | ( n9945 & n11332 ) ;
  assign n12453 = n12451 & ~n12452 ;
  assign n12454 = n12453 ^ n5251 ^ 1'b0 ;
  assign n12455 = ( ~n6109 & n6502 ) | ( ~n6109 & n10467 ) | ( n6502 & n10467 ) ;
  assign n12456 = ( n1581 & n11255 ) | ( n1581 & n12455 ) | ( n11255 & n12455 ) ;
  assign n12457 = n2978 ^ n2397 ^ n1485 ;
  assign n12458 = n12457 ^ n8223 ^ n1885 ;
  assign n12460 = n2067 ^ n624 ^ n481 ;
  assign n12461 = n2898 | n12460 ;
  assign n12462 = n2491 | n12461 ;
  assign n12459 = ( n701 & n4492 ) | ( n701 & ~n7818 ) | ( n4492 & ~n7818 ) ;
  assign n12463 = n12462 ^ n12459 ^ n2305 ;
  assign n12464 = n12463 ^ n9726 ^ n8253 ;
  assign n12465 = n1528 | n3156 ;
  assign n12466 = n7652 | n12465 ;
  assign n12467 = ( x61 & ~n1377 ) | ( x61 & n1749 ) | ( ~n1377 & n1749 ) ;
  assign n12468 = n12467 ^ n3665 ^ 1'b0 ;
  assign n12469 = n12468 ^ n10281 ^ n542 ;
  assign n12470 = ( ~n9893 & n12466 ) | ( ~n9893 & n12469 ) | ( n12466 & n12469 ) ;
  assign n12471 = ~n401 & n514 ;
  assign n12472 = n12471 ^ n1722 ^ 1'b0 ;
  assign n12473 = n6941 | n10314 ;
  assign n12474 = n3560 & ~n12473 ;
  assign n12475 = ( n5021 & n5450 ) | ( n5021 & ~n12474 ) | ( n5450 & ~n12474 ) ;
  assign n12476 = ( n4922 & ~n12472 ) | ( n4922 & n12475 ) | ( ~n12472 & n12475 ) ;
  assign n12477 = n12476 ^ n1085 ^ 1'b0 ;
  assign n12478 = n7888 ^ n5122 ^ n3746 ;
  assign n12479 = n12478 ^ n7802 ^ n6265 ;
  assign n12480 = ( n362 & ~n2353 ) | ( n362 & n4042 ) | ( ~n2353 & n4042 ) ;
  assign n12481 = ( n597 & n10826 ) | ( n597 & n12480 ) | ( n10826 & n12480 ) ;
  assign n12482 = ( n7467 & ~n10093 ) | ( n7467 & n12481 ) | ( ~n10093 & n12481 ) ;
  assign n12483 = ( n5083 & n12479 ) | ( n5083 & n12482 ) | ( n12479 & n12482 ) ;
  assign n12487 = ( n1349 & n7104 ) | ( n1349 & n7504 ) | ( n7104 & n7504 ) ;
  assign n12485 = ( n4002 & ~n4521 ) | ( n4002 & n5381 ) | ( ~n4521 & n5381 ) ;
  assign n12484 = n1911 & ~n5538 ;
  assign n12486 = n12485 ^ n12484 ^ 1'b0 ;
  assign n12488 = n12487 ^ n12486 ^ n3356 ;
  assign n12489 = ( ~n5810 & n12184 ) | ( ~n5810 & n12488 ) | ( n12184 & n12488 ) ;
  assign n12490 = n1501 & ~n8783 ;
  assign n12497 = n9858 ^ n9587 ^ n3638 ;
  assign n12498 = n12497 ^ n4897 ^ n3920 ;
  assign n12491 = ( n704 & n4158 ) | ( n704 & ~n4864 ) | ( n4158 & ~n4864 ) ;
  assign n12492 = n198 & n4392 ;
  assign n12493 = n12492 ^ n5895 ^ 1'b0 ;
  assign n12494 = ( n8473 & ~n8576 ) | ( n8473 & n12493 ) | ( ~n8576 & n12493 ) ;
  assign n12495 = ( n8359 & n12491 ) | ( n8359 & n12494 ) | ( n12491 & n12494 ) ;
  assign n12496 = ~n3416 & n12495 ;
  assign n12499 = n12498 ^ n12496 ^ 1'b0 ;
  assign n12500 = ( n4730 & ~n10811 ) | ( n4730 & n11388 ) | ( ~n10811 & n11388 ) ;
  assign n12501 = ( n2397 & n3248 ) | ( n2397 & ~n3893 ) | ( n3248 & ~n3893 ) ;
  assign n12506 = ( ~n2151 & n2965 ) | ( ~n2151 & n3183 ) | ( n2965 & n3183 ) ;
  assign n12503 = n3611 ^ n698 ^ 1'b0 ;
  assign n12504 = ~n2918 & n12503 ;
  assign n12502 = ( n8243 & n9567 ) | ( n8243 & n9628 ) | ( n9567 & n9628 ) ;
  assign n12505 = n12504 ^ n12502 ^ n8651 ;
  assign n12507 = n12506 ^ n12505 ^ n7251 ;
  assign n12508 = ( n7544 & n8928 ) | ( n7544 & ~n12507 ) | ( n8928 & ~n12507 ) ;
  assign n12510 = n5728 ^ n2224 ^ 1'b0 ;
  assign n12511 = ~n7859 & n12510 ;
  assign n12509 = n2356 & n8691 ;
  assign n12512 = n12511 ^ n12509 ^ 1'b0 ;
  assign n12513 = n12512 ^ n2656 ^ n1658 ;
  assign n12514 = n3494 & n7823 ;
  assign n12515 = n12514 ^ n7758 ^ 1'b0 ;
  assign n12516 = n5190 | n9837 ;
  assign n12517 = n12516 ^ n733 ^ 1'b0 ;
  assign n12518 = n12517 ^ n3359 ^ 1'b0 ;
  assign n12519 = ( n4960 & n12515 ) | ( n4960 & ~n12518 ) | ( n12515 & ~n12518 ) ;
  assign n12520 = ( ~n12321 & n12513 ) | ( ~n12321 & n12519 ) | ( n12513 & n12519 ) ;
  assign n12521 = n8946 ^ x114 ^ 1'b0 ;
  assign n12522 = n12520 & n12521 ;
  assign n12523 = ( ~n3876 & n6627 ) | ( ~n3876 & n12460 ) | ( n6627 & n12460 ) ;
  assign n12524 = n12523 ^ n6040 ^ n3868 ;
  assign n12525 = n12524 ^ n4130 ^ n3642 ;
  assign n12526 = n1626 | n4310 ;
  assign n12527 = n12526 ^ n8747 ^ 1'b0 ;
  assign n12528 = n8159 & ~n12527 ;
  assign n12529 = n12528 ^ n3784 ^ n1125 ;
  assign n12530 = n5259 ^ n175 ^ 1'b0 ;
  assign n12531 = ( n12525 & ~n12529 ) | ( n12525 & n12530 ) | ( ~n12529 & n12530 ) ;
  assign n12532 = ( n3160 & n5771 ) | ( n3160 & n12531 ) | ( n5771 & n12531 ) ;
  assign n12533 = n10905 ^ n6798 ^ n4581 ;
  assign n12534 = n12533 ^ n953 ^ n333 ;
  assign n12535 = ( n1249 & ~n2487 ) | ( n1249 & n12534 ) | ( ~n2487 & n12534 ) ;
  assign n12536 = n12535 ^ n6943 ^ 1'b0 ;
  assign n12537 = n10981 & ~n12536 ;
  assign n12538 = ( n868 & ~n7833 ) | ( n868 & n12537 ) | ( ~n7833 & n12537 ) ;
  assign n12539 = n4463 ^ n2640 ^ n1668 ;
  assign n12540 = ( n11961 & ~n12158 ) | ( n11961 & n12539 ) | ( ~n12158 & n12539 ) ;
  assign n12541 = ( n1087 & n5688 ) | ( n1087 & ~n7476 ) | ( n5688 & ~n7476 ) ;
  assign n12542 = n7456 ^ n3379 ^ 1'b0 ;
  assign n12543 = n12541 & n12542 ;
  assign n12544 = n1208 & ~n2640 ;
  assign n12545 = n12544 ^ n12232 ^ 1'b0 ;
  assign n12546 = n5959 ^ n1738 ^ n1414 ;
  assign n12547 = n12546 ^ n8927 ^ n4424 ;
  assign n12548 = n7709 ^ n6088 ^ 1'b0 ;
  assign n12549 = ( n1978 & ~n8603 ) | ( n1978 & n12548 ) | ( ~n8603 & n12548 ) ;
  assign n12550 = ( ~n1412 & n7477 ) | ( ~n1412 & n12046 ) | ( n7477 & n12046 ) ;
  assign n12551 = ( n5479 & n7851 ) | ( n5479 & n11881 ) | ( n7851 & n11881 ) ;
  assign n12552 = ( ~n1714 & n1771 ) | ( ~n1714 & n3175 ) | ( n1771 & n3175 ) ;
  assign n12553 = n12552 ^ n3784 ^ n1834 ;
  assign n12554 = ( ~n2094 & n5567 ) | ( ~n2094 & n12553 ) | ( n5567 & n12553 ) ;
  assign n12555 = n4374 & n6217 ;
  assign n12556 = ( n7440 & n11652 ) | ( n7440 & n12555 ) | ( n11652 & n12555 ) ;
  assign n12557 = n12556 ^ n8320 ^ 1'b0 ;
  assign n12558 = n9870 & n12557 ;
  assign n12559 = ( n1350 & n10386 ) | ( n1350 & n12558 ) | ( n10386 & n12558 ) ;
  assign n12563 = n161 | n2885 ;
  assign n12564 = n8770 | n12563 ;
  assign n12560 = n7689 & ~n10655 ;
  assign n12561 = n480 & n12560 ;
  assign n12562 = n12561 ^ n5865 ^ n2236 ;
  assign n12565 = n12564 ^ n12562 ^ n2942 ;
  assign n12566 = n12565 ^ n6455 ^ n1424 ;
  assign n12567 = n12566 ^ n6494 ^ n5749 ;
  assign n12568 = ( n9478 & n12455 ) | ( n9478 & n12567 ) | ( n12455 & n12567 ) ;
  assign n12569 = n12001 ^ n11317 ^ 1'b0 ;
  assign n12570 = n5357 ^ n4074 ^ n881 ;
  assign n12571 = ( n5113 & ~n8457 ) | ( n5113 & n12570 ) | ( ~n8457 & n12570 ) ;
  assign n12572 = ( ~n5949 & n9128 ) | ( ~n5949 & n10817 ) | ( n9128 & n10817 ) ;
  assign n12573 = n12572 ^ n4342 ^ n3237 ;
  assign n12576 = n5793 ^ n144 ^ 1'b0 ;
  assign n12574 = n7818 ^ n7407 ^ n416 ;
  assign n12575 = n11604 & ~n12574 ;
  assign n12577 = n12576 ^ n12575 ^ 1'b0 ;
  assign n12578 = n6952 ^ n5454 ^ n4465 ;
  assign n12579 = ( n5541 & ~n11151 ) | ( n5541 & n12578 ) | ( ~n11151 & n12578 ) ;
  assign n12582 = ( n2147 & n3303 ) | ( n2147 & ~n8662 ) | ( n3303 & ~n8662 ) ;
  assign n12581 = n9976 ^ n3094 ^ n759 ;
  assign n12580 = ( ~n6253 & n9137 ) | ( ~n6253 & n9208 ) | ( n9137 & n9208 ) ;
  assign n12583 = n12582 ^ n12581 ^ n12580 ;
  assign n12584 = ( n664 & n5405 ) | ( n664 & ~n6627 ) | ( n5405 & ~n6627 ) ;
  assign n12585 = ( n4485 & ~n6221 ) | ( n4485 & n12584 ) | ( ~n6221 & n12584 ) ;
  assign n12586 = n6891 ^ n6407 ^ 1'b0 ;
  assign n12587 = ( n2879 & n5591 ) | ( n2879 & ~n9618 ) | ( n5591 & ~n9618 ) ;
  assign n12588 = n6217 & n12587 ;
  assign n12589 = ( n6982 & n12586 ) | ( n6982 & n12588 ) | ( n12586 & n12588 ) ;
  assign n12595 = n3656 ^ n3224 ^ 1'b0 ;
  assign n12590 = ( n3660 & ~n6139 ) | ( n3660 & n12125 ) | ( ~n6139 & n12125 ) ;
  assign n12591 = n12590 ^ n4118 ^ n1080 ;
  assign n12592 = ( n2278 & ~n8625 ) | ( n2278 & n12591 ) | ( ~n8625 & n12591 ) ;
  assign n12593 = ~n9833 & n12592 ;
  assign n12594 = n12593 ^ n5703 ^ 1'b0 ;
  assign n12596 = n12595 ^ n12594 ^ n1619 ;
  assign n12598 = n4232 | n5615 ;
  assign n12599 = n12598 ^ n7841 ^ 1'b0 ;
  assign n12600 = ~n5613 & n12599 ;
  assign n12597 = ( ~n5102 & n10001 ) | ( ~n5102 & n11885 ) | ( n10001 & n11885 ) ;
  assign n12601 = n12600 ^ n12597 ^ n4887 ;
  assign n12602 = n5748 & n11527 ;
  assign n12603 = n1393 & n3011 ;
  assign n12604 = ~n1203 & n12603 ;
  assign n12605 = n10044 ^ n6217 ^ n1808 ;
  assign n12606 = n1568 | n2270 ;
  assign n12607 = n12605 & ~n12606 ;
  assign n12608 = ( n6001 & n12604 ) | ( n6001 & n12607 ) | ( n12604 & n12607 ) ;
  assign n12609 = n12608 ^ n10844 ^ n1016 ;
  assign n12610 = n6163 ^ n4543 ^ n228 ;
  assign n12611 = n12610 ^ n9563 ^ n4720 ;
  assign n12618 = n5470 ^ n143 ^ x53 ;
  assign n12619 = n12618 ^ n5620 ^ n1911 ;
  assign n12620 = ~n1135 & n12619 ;
  assign n12621 = n3120 & n12620 ;
  assign n12613 = n1877 | n5913 ;
  assign n12614 = n5146 | n12613 ;
  assign n12615 = n12614 ^ n6926 ^ n5870 ;
  assign n12616 = ( n3088 & n7200 ) | ( n3088 & n12615 ) | ( n7200 & n12615 ) ;
  assign n12612 = ( n2553 & n5062 ) | ( n2553 & n8874 ) | ( n5062 & n8874 ) ;
  assign n12617 = n12616 ^ n12612 ^ 1'b0 ;
  assign n12622 = n12621 ^ n12617 ^ n11284 ;
  assign n12623 = ( n1867 & n8651 ) | ( n1867 & n11143 ) | ( n8651 & n11143 ) ;
  assign n12624 = ( n2358 & n5961 ) | ( n2358 & n12368 ) | ( n5961 & n12368 ) ;
  assign n12625 = n12624 ^ n11543 ^ n5737 ;
  assign n12626 = n12625 ^ n5375 ^ n2794 ;
  assign n12627 = n4269 | n12626 ;
  assign n12628 = n6426 ^ n1674 ^ 1'b0 ;
  assign n12629 = ~n12627 & n12628 ;
  assign n12638 = n7570 ^ n3119 ^ n2357 ;
  assign n12636 = n11435 ^ n9396 ^ n5695 ;
  assign n12637 = n12636 ^ n4354 ^ n2336 ;
  assign n12639 = n12638 ^ n12637 ^ n6292 ;
  assign n12640 = n12639 ^ n10547 ^ n6173 ;
  assign n12630 = n6917 ^ n5258 ^ n2186 ;
  assign n12631 = ( n1520 & ~n5861 ) | ( n1520 & n9948 ) | ( ~n5861 & n9948 ) ;
  assign n12632 = n3016 & ~n3859 ;
  assign n12633 = n12632 ^ n8317 ^ 1'b0 ;
  assign n12634 = ( ~n1912 & n12631 ) | ( ~n1912 & n12633 ) | ( n12631 & n12633 ) ;
  assign n12635 = n12630 | n12634 ;
  assign n12641 = n12640 ^ n12635 ^ 1'b0 ;
  assign n12645 = ( ~n3874 & n9327 ) | ( ~n3874 & n9964 ) | ( n9327 & n9964 ) ;
  assign n12642 = ( ~x36 & n1992 ) | ( ~x36 & n5309 ) | ( n1992 & n5309 ) ;
  assign n12643 = n12642 ^ n10447 ^ n2400 ;
  assign n12644 = ~n3655 & n12643 ;
  assign n12646 = n12645 ^ n12644 ^ n11584 ;
  assign n12647 = n1887 | n3764 ;
  assign n12648 = n5869 | n12647 ;
  assign n12649 = ( n727 & n6533 ) | ( n727 & n12648 ) | ( n6533 & n12648 ) ;
  assign n12650 = n9456 ^ n4408 ^ n524 ;
  assign n12651 = n4030 & n9073 ;
  assign n12652 = n12651 ^ n8397 ^ 1'b0 ;
  assign n12653 = n12652 ^ n8795 ^ 1'b0 ;
  assign n12654 = n3406 & n12653 ;
  assign n12657 = ~n1006 & n2144 ;
  assign n12655 = ( n3071 & n4054 ) | ( n3071 & n12460 ) | ( n4054 & n12460 ) ;
  assign n12656 = n12655 ^ n6255 ^ n3911 ;
  assign n12658 = n12657 ^ n12656 ^ n6788 ;
  assign n12659 = n12658 ^ n7709 ^ n1774 ;
  assign n12660 = n4844 ^ n2932 ^ n1657 ;
  assign n12661 = n4144 ^ n1064 ^ n797 ;
  assign n12662 = ( n9454 & n12660 ) | ( n9454 & ~n12661 ) | ( n12660 & ~n12661 ) ;
  assign n12663 = n12662 ^ n9871 ^ n3776 ;
  assign n12664 = ~n2378 & n12663 ;
  assign n12665 = ( ~n2875 & n6876 ) | ( ~n2875 & n11473 ) | ( n6876 & n11473 ) ;
  assign n12666 = ( ~n5245 & n6422 ) | ( ~n5245 & n9386 ) | ( n6422 & n9386 ) ;
  assign n12667 = n2937 ^ n2154 ^ 1'b0 ;
  assign n12668 = n12667 ^ n8384 ^ n1273 ;
  assign n12669 = n12668 ^ n1413 ^ 1'b0 ;
  assign n12670 = n7404 & n12669 ;
  assign n12671 = n12670 ^ n1610 ^ 1'b0 ;
  assign n12672 = ( n5557 & ~n12666 ) | ( n5557 & n12671 ) | ( ~n12666 & n12671 ) ;
  assign n12673 = ( n3681 & ~n12665 ) | ( n3681 & n12672 ) | ( ~n12665 & n12672 ) ;
  assign n12674 = ( ~n1175 & n3937 ) | ( ~n1175 & n6209 ) | ( n3937 & n6209 ) ;
  assign n12675 = n12674 ^ n11895 ^ n366 ;
  assign n12676 = n2454 ^ n328 ^ 1'b0 ;
  assign n12677 = n5000 & n9552 ;
  assign n12678 = ( n5009 & n12676 ) | ( n5009 & ~n12677 ) | ( n12676 & ~n12677 ) ;
  assign n12679 = n5853 ^ n474 ^ 1'b0 ;
  assign n12680 = x29 & n12679 ;
  assign n12681 = n12680 ^ n5383 ^ 1'b0 ;
  assign n12683 = n11509 ^ n5831 ^ n2100 ;
  assign n12682 = n7197 ^ n2970 ^ n1027 ;
  assign n12684 = n12683 ^ n12682 ^ n11866 ;
  assign n12685 = ( ~x91 & n5341 ) | ( ~x91 & n7419 ) | ( n5341 & n7419 ) ;
  assign n12686 = n12685 ^ n8829 ^ 1'b0 ;
  assign n12687 = n4285 & ~n12686 ;
  assign n12688 = ( n3598 & n10070 ) | ( n3598 & n12687 ) | ( n10070 & n12687 ) ;
  assign n12689 = n12688 ^ n11538 ^ n3647 ;
  assign n12690 = n5076 ^ n2490 ^ 1'b0 ;
  assign n12691 = n12504 ^ n3963 ^ n2801 ;
  assign n12692 = ~n5121 & n6633 ;
  assign n12693 = n12691 & n12692 ;
  assign n12694 = n8307 ^ n8004 ^ n1354 ;
  assign n12695 = n5719 ^ n1922 ^ n1874 ;
  assign n12696 = n12695 ^ n2977 ^ n2116 ;
  assign n12697 = ( n1281 & n2698 ) | ( n1281 & n12696 ) | ( n2698 & n12696 ) ;
  assign n12698 = ( n5551 & n9593 ) | ( n5551 & n12697 ) | ( n9593 & n12697 ) ;
  assign n12699 = n9897 ^ n8118 ^ n7123 ;
  assign n12700 = n1776 & n8827 ;
  assign n12701 = n12700 ^ n11529 ^ n2734 ;
  assign n12702 = ( n702 & n3891 ) | ( n702 & n5514 ) | ( n3891 & n5514 ) ;
  assign n12703 = n12702 ^ n7783 ^ n6243 ;
  assign n12704 = ( n2390 & ~n12701 ) | ( n2390 & n12703 ) | ( ~n12701 & n12703 ) ;
  assign n12705 = ~n2872 & n12704 ;
  assign n12706 = n8782 ^ n4344 ^ x88 ;
  assign n12707 = ~n12633 & n12706 ;
  assign n12708 = ~n1151 & n4504 ;
  assign n12709 = n12708 ^ n8542 ^ n6763 ;
  assign n12710 = ( x79 & n4014 ) | ( x79 & n12709 ) | ( n4014 & n12709 ) ;
  assign n12711 = n9813 ^ n3811 ^ 1'b0 ;
  assign n12712 = ~n280 & n12711 ;
  assign n12713 = ~n12710 & n12712 ;
  assign n12714 = ( ~n4639 & n12707 ) | ( ~n4639 & n12713 ) | ( n12707 & n12713 ) ;
  assign n12715 = ( n4044 & ~n4569 ) | ( n4044 & n7228 ) | ( ~n4569 & n7228 ) ;
  assign n12716 = n12715 ^ n8601 ^ n1846 ;
  assign n12717 = n11707 & n12502 ;
  assign n12718 = n12716 & n12717 ;
  assign n12719 = n5146 ^ n3992 ^ 1'b0 ;
  assign n12720 = n12719 ^ n8791 ^ n3380 ;
  assign n12721 = ( n1173 & n4683 ) | ( n1173 & ~n12720 ) | ( n4683 & ~n12720 ) ;
  assign n12722 = n10482 ^ n9483 ^ n7434 ;
  assign n12723 = ( n551 & n2343 ) | ( n551 & n12722 ) | ( n2343 & n12722 ) ;
  assign n12724 = n12655 ^ n11891 ^ n9050 ;
  assign n12725 = n3898 ^ n2503 ^ n1280 ;
  assign n12726 = n12725 ^ n2066 ^ n751 ;
  assign n12727 = n12726 ^ n5716 ^ n4760 ;
  assign n12728 = n12727 ^ n5763 ^ n5507 ;
  assign n12732 = n2235 | n4825 ;
  assign n12733 = n12732 ^ n778 ^ 1'b0 ;
  assign n12734 = ( n1929 & n2165 ) | ( n1929 & ~n7657 ) | ( n2165 & ~n7657 ) ;
  assign n12735 = ( ~n9520 & n12733 ) | ( ~n9520 & n12734 ) | ( n12733 & n12734 ) ;
  assign n12729 = ( n2768 & ~n5594 ) | ( n2768 & n6570 ) | ( ~n5594 & n6570 ) ;
  assign n12730 = ~n12203 & n12729 ;
  assign n12731 = ( ~n1074 & n11498 ) | ( ~n1074 & n12730 ) | ( n11498 & n12730 ) ;
  assign n12736 = n12735 ^ n12731 ^ n4974 ;
  assign n12738 = n12052 ^ n7249 ^ n4028 ;
  assign n12739 = ~n1908 & n3419 ;
  assign n12740 = n12739 ^ n8525 ^ 1'b0 ;
  assign n12741 = ( ~n6571 & n12738 ) | ( ~n6571 & n12740 ) | ( n12738 & n12740 ) ;
  assign n12737 = n8764 | n11250 ;
  assign n12742 = n12741 ^ n12737 ^ 1'b0 ;
  assign n12750 = n6666 ^ n1255 ^ 1'b0 ;
  assign n12751 = n2835 & n12750 ;
  assign n12748 = ~n3529 & n9458 ;
  assign n12749 = n12748 ^ n12685 ^ 1'b0 ;
  assign n12743 = n10785 ^ n5007 ^ 1'b0 ;
  assign n12744 = ( n1406 & n2437 ) | ( n1406 & n6665 ) | ( n2437 & n6665 ) ;
  assign n12745 = ( ~n2836 & n8796 ) | ( ~n2836 & n12744 ) | ( n8796 & n12744 ) ;
  assign n12746 = n645 | n12745 ;
  assign n12747 = n12743 | n12746 ;
  assign n12752 = n12751 ^ n12749 ^ n12747 ;
  assign n12753 = ~n2171 & n3121 ;
  assign n12754 = ( n3138 & n4692 ) | ( n3138 & n9893 ) | ( n4692 & n9893 ) ;
  assign n12759 = n7505 ^ n6116 ^ n1543 ;
  assign n12760 = ( n620 & ~n9905 ) | ( n620 & n12759 ) | ( ~n9905 & n12759 ) ;
  assign n12761 = n12760 ^ n5655 ^ n5091 ;
  assign n12755 = ( n359 & n2891 ) | ( n359 & n8406 ) | ( n2891 & n8406 ) ;
  assign n12756 = n3938 & n12755 ;
  assign n12757 = ~n7512 & n12756 ;
  assign n12758 = n12757 ^ n4065 ^ n812 ;
  assign n12762 = n12761 ^ n12758 ^ n7301 ;
  assign n12763 = n2406 | n10712 ;
  assign n12764 = ( ~n785 & n8092 ) | ( ~n785 & n12763 ) | ( n8092 & n12763 ) ;
  assign n12765 = ( ~n2522 & n4575 ) | ( ~n2522 & n12764 ) | ( n4575 & n12764 ) ;
  assign n12766 = ( n288 & n5646 ) | ( n288 & ~n10105 ) | ( n5646 & ~n10105 ) ;
  assign n12767 = ~n5567 & n12766 ;
  assign n12768 = n12767 ^ n836 ^ 1'b0 ;
  assign n12769 = ( n555 & n3758 ) | ( n555 & n7229 ) | ( n3758 & n7229 ) ;
  assign n12770 = n12769 ^ n7564 ^ n4940 ;
  assign n12771 = n12770 ^ n7848 ^ n1884 ;
  assign n12772 = ( ~n2395 & n4090 ) | ( ~n2395 & n5065 ) | ( n4090 & n5065 ) ;
  assign n12773 = ( n1347 & n4906 ) | ( n1347 & ~n6941 ) | ( n4906 & ~n6941 ) ;
  assign n12774 = n12773 ^ n11736 ^ 1'b0 ;
  assign n12775 = ( n9080 & n12772 ) | ( n9080 & ~n12774 ) | ( n12772 & ~n12774 ) ;
  assign n12776 = n8510 ^ n2466 ^ n988 ;
  assign n12777 = ( n2424 & n2821 ) | ( n2424 & ~n12776 ) | ( n2821 & ~n12776 ) ;
  assign n12778 = ( n1257 & n5361 ) | ( n1257 & n11192 ) | ( n5361 & n11192 ) ;
  assign n12779 = ( n196 & ~n1863 ) | ( n196 & n2451 ) | ( ~n1863 & n2451 ) ;
  assign n12780 = n12779 ^ n2450 ^ 1'b0 ;
  assign n12781 = n1703 ^ n1623 ^ n240 ;
  assign n12782 = n12781 ^ n6906 ^ 1'b0 ;
  assign n12783 = n12780 & n12782 ;
  assign n12784 = ~n8080 & n10302 ;
  assign n12785 = n12784 ^ n7704 ^ 1'b0 ;
  assign n12786 = n8814 | n12785 ;
  assign n12787 = n12786 ^ n12699 ^ 1'b0 ;
  assign n12788 = n2048 | n8489 ;
  assign n12789 = n5039 | n12788 ;
  assign n12790 = ( n5874 & ~n5900 ) | ( n5874 & n12789 ) | ( ~n5900 & n12789 ) ;
  assign n12791 = ( n9294 & n11389 ) | ( n9294 & ~n12790 ) | ( n11389 & ~n12790 ) ;
  assign n12792 = n1201 & ~n5332 ;
  assign n12793 = ( n457 & n1491 ) | ( n457 & ~n12792 ) | ( n1491 & ~n12792 ) ;
  assign n12794 = ( n671 & n2167 ) | ( n671 & n12793 ) | ( n2167 & n12793 ) ;
  assign n12795 = ( n568 & n788 ) | ( n568 & n2256 ) | ( n788 & n2256 ) ;
  assign n12796 = n12795 ^ n1432 ^ 1'b0 ;
  assign n12797 = ( ~n2753 & n6306 ) | ( ~n2753 & n7600 ) | ( n6306 & n7600 ) ;
  assign n12798 = ( n8447 & ~n10228 ) | ( n8447 & n12797 ) | ( ~n10228 & n12797 ) ;
  assign n12804 = ( ~n1978 & n7813 ) | ( ~n1978 & n12336 ) | ( n7813 & n12336 ) ;
  assign n12805 = n12804 ^ n5634 ^ n4259 ;
  assign n12801 = n5493 ^ n5338 ^ 1'b0 ;
  assign n12802 = n6284 & ~n12801 ;
  assign n12799 = n9622 ^ n1538 ^ 1'b0 ;
  assign n12800 = ( ~n1206 & n3783 ) | ( ~n1206 & n12799 ) | ( n3783 & n12799 ) ;
  assign n12803 = n12802 ^ n12800 ^ n8205 ;
  assign n12806 = n12805 ^ n12803 ^ n8155 ;
  assign n12807 = n2075 ^ n1314 ^ x83 ;
  assign n12808 = n9211 & ~n12807 ;
  assign n12809 = n12808 ^ n9517 ^ n3147 ;
  assign n12810 = ( ~n806 & n1946 ) | ( ~n806 & n12809 ) | ( n1946 & n12809 ) ;
  assign n12811 = ( ~n1482 & n6839 ) | ( ~n1482 & n11349 ) | ( n6839 & n11349 ) ;
  assign n12812 = ~n6406 & n12811 ;
  assign n12813 = n12812 ^ n10795 ^ n8487 ;
  assign n12814 = n5407 ^ n1779 ^ n203 ;
  assign n12815 = n12814 ^ n9658 ^ n8073 ;
  assign n12816 = n12815 ^ n8987 ^ n222 ;
  assign n12817 = ( n2728 & n4117 ) | ( n2728 & ~n12816 ) | ( n4117 & ~n12816 ) ;
  assign n12823 = n10075 ^ n9748 ^ n6960 ;
  assign n12818 = ( ~n3286 & n3463 ) | ( ~n3286 & n8363 ) | ( n3463 & n8363 ) ;
  assign n12819 = n12818 ^ n297 ^ 1'b0 ;
  assign n12820 = ~n2785 & n12819 ;
  assign n12821 = n12820 ^ n4801 ^ n3716 ;
  assign n12822 = ( ~n10469 & n10699 ) | ( ~n10469 & n12821 ) | ( n10699 & n12821 ) ;
  assign n12824 = n12823 ^ n12822 ^ n9321 ;
  assign n12825 = n2090 ^ n1503 ^ n272 ;
  assign n12826 = n12825 ^ n12703 ^ n2218 ;
  assign n12827 = n8059 ^ n3068 ^ n1422 ;
  assign n12828 = n12827 ^ n9794 ^ n4979 ;
  assign n12829 = n12828 ^ n10792 ^ n3530 ;
  assign n12830 = n411 & ~n3352 ;
  assign n12831 = n10969 ^ n7667 ^ n3843 ;
  assign n12834 = n4984 ^ n4688 ^ n373 ;
  assign n12833 = ( ~x61 & n3977 ) | ( ~x61 & n7196 ) | ( n3977 & n7196 ) ;
  assign n12835 = n12834 ^ n12833 ^ n2638 ;
  assign n12832 = n3414 ^ n2511 ^ n656 ;
  assign n12836 = n12835 ^ n12832 ^ n2869 ;
  assign n12837 = n12836 ^ n740 ^ 1'b0 ;
  assign n12838 = ( n12830 & ~n12831 ) | ( n12830 & n12837 ) | ( ~n12831 & n12837 ) ;
  assign n12839 = n8518 ^ n5515 ^ n2802 ;
  assign n12840 = n5074 ^ n2134 ^ n914 ;
  assign n12841 = ~n12839 & n12840 ;
  assign n12842 = ( n3484 & n5146 ) | ( n3484 & n12841 ) | ( n5146 & n12841 ) ;
  assign n12843 = n5282 ^ n3916 ^ 1'b0 ;
  assign n12844 = n10442 & ~n12843 ;
  assign n12845 = n2465 & n12844 ;
  assign n12846 = n6598 ^ n4817 ^ 1'b0 ;
  assign n12847 = ( n1499 & n10423 ) | ( n1499 & ~n12529 ) | ( n10423 & ~n12529 ) ;
  assign n12848 = n5662 | n12847 ;
  assign n12849 = n12848 ^ n3759 ^ 1'b0 ;
  assign n12852 = ( n4733 & n5800 ) | ( n4733 & ~n7301 ) | ( n5800 & ~n7301 ) ;
  assign n12853 = n12852 ^ n7813 ^ n4465 ;
  assign n12850 = ( n430 & ~n1985 ) | ( n430 & n4426 ) | ( ~n1985 & n4426 ) ;
  assign n12851 = n12850 ^ n11244 ^ n10038 ;
  assign n12854 = n12853 ^ n12851 ^ n7642 ;
  assign n12855 = n1721 & ~n2268 ;
  assign n12856 = n722 | n4097 ;
  assign n12857 = ( ~n2729 & n4072 ) | ( ~n2729 & n6114 ) | ( n4072 & n6114 ) ;
  assign n12858 = ( n12855 & n12856 ) | ( n12855 & ~n12857 ) | ( n12856 & ~n12857 ) ;
  assign n12860 = ( n2368 & n2371 ) | ( n2368 & ~n6217 ) | ( n2371 & ~n6217 ) ;
  assign n12859 = n12075 ^ n10955 ^ n5629 ;
  assign n12861 = n12860 ^ n12859 ^ n5132 ;
  assign n12862 = ( n5189 & ~n12858 ) | ( n5189 & n12861 ) | ( ~n12858 & n12861 ) ;
  assign n12863 = n4925 & n9847 ;
  assign n12864 = ( x36 & n9257 ) | ( x36 & n10109 ) | ( n9257 & n10109 ) ;
  assign n12865 = n12864 ^ n3615 ^ x61 ;
  assign n12866 = n1606 & n2457 ;
  assign n12867 = n12866 ^ n1395 ^ 1'b0 ;
  assign n12868 = ( n848 & ~n5147 ) | ( n848 & n12867 ) | ( ~n5147 & n12867 ) ;
  assign n12869 = n12865 | n12868 ;
  assign n12870 = n12863 & ~n12869 ;
  assign n12871 = ( n5458 & n5828 ) | ( n5458 & n9128 ) | ( n5828 & n9128 ) ;
  assign n12873 = n6224 ^ n4449 ^ n3361 ;
  assign n12872 = ( n2701 & n9484 ) | ( n2701 & ~n11155 ) | ( n9484 & ~n11155 ) ;
  assign n12874 = n12873 ^ n12872 ^ n1255 ;
  assign n12876 = ~n7649 & n11304 ;
  assign n12875 = n7158 & n7448 ;
  assign n12877 = n12876 ^ n12875 ^ 1'b0 ;
  assign n12878 = n11459 ^ n7042 ^ n2658 ;
  assign n12879 = n12878 ^ n11761 ^ n3891 ;
  assign n12880 = ( n2773 & n3487 ) | ( n2773 & ~n7201 ) | ( n3487 & ~n7201 ) ;
  assign n12881 = n8884 ^ n2425 ^ 1'b0 ;
  assign n12882 = n12881 ^ n8455 ^ 1'b0 ;
  assign n12883 = n5149 & ~n11481 ;
  assign n12884 = ~n2600 & n12883 ;
  assign n12885 = ( n772 & ~n868 ) | ( n772 & n3623 ) | ( ~n868 & n3623 ) ;
  assign n12886 = n12885 ^ n3740 ^ n1406 ;
  assign n12887 = n12457 ^ n3745 ^ 1'b0 ;
  assign n12889 = n11916 ^ n889 ^ n656 ;
  assign n12890 = ( n3289 & n4025 ) | ( n3289 & n12889 ) | ( n4025 & n12889 ) ;
  assign n12888 = n12165 ^ n11313 ^ n1494 ;
  assign n12891 = n12890 ^ n12888 ^ n5850 ;
  assign n12892 = ( n12886 & n12887 ) | ( n12886 & ~n12891 ) | ( n12887 & ~n12891 ) ;
  assign n12893 = ~n3501 & n6570 ;
  assign n12894 = ( n11218 & n11870 ) | ( n11218 & n12893 ) | ( n11870 & n12893 ) ;
  assign n12895 = n5821 | n10742 ;
  assign n12896 = ( ~n6460 & n10480 ) | ( ~n6460 & n12895 ) | ( n10480 & n12895 ) ;
  assign n12897 = n7072 ^ n5796 ^ n2585 ;
  assign n12899 = ( ~n2348 & n6253 ) | ( ~n2348 & n6863 ) | ( n6253 & n6863 ) ;
  assign n12900 = n12899 ^ n7687 ^ n1587 ;
  assign n12898 = ( n5727 & n8422 ) | ( n5727 & n12403 ) | ( n8422 & n12403 ) ;
  assign n12901 = n12900 ^ n12898 ^ n5140 ;
  assign n12902 = n12901 ^ n8297 ^ n1925 ;
  assign n12905 = ( n296 & n1790 ) | ( n296 & ~n10278 ) | ( n1790 & ~n10278 ) ;
  assign n12903 = n12388 ^ n2150 ^ n1395 ;
  assign n12904 = ( n4863 & n8462 ) | ( n4863 & ~n12903 ) | ( n8462 & ~n12903 ) ;
  assign n12906 = n12905 ^ n12904 ^ n2541 ;
  assign n12907 = ( n755 & n1940 ) | ( n755 & n2306 ) | ( n1940 & n2306 ) ;
  assign n12908 = n6174 ^ n1709 ^ 1'b0 ;
  assign n12909 = ~n5024 & n6869 ;
  assign n12910 = ( n12907 & ~n12908 ) | ( n12907 & n12909 ) | ( ~n12908 & n12909 ) ;
  assign n12911 = ( n11063 & n12906 ) | ( n11063 & ~n12910 ) | ( n12906 & ~n12910 ) ;
  assign n12912 = ( ~n1447 & n2028 ) | ( ~n1447 & n5183 ) | ( n2028 & n5183 ) ;
  assign n12913 = n4456 & n5886 ;
  assign n12914 = ( ~n8782 & n12912 ) | ( ~n8782 & n12913 ) | ( n12912 & n12913 ) ;
  assign n12917 = ( n2245 & ~n4297 ) | ( n2245 & n8149 ) | ( ~n4297 & n8149 ) ;
  assign n12915 = n11052 ^ n3409 ^ n2576 ;
  assign n12916 = n9670 & ~n12915 ;
  assign n12918 = n12917 ^ n12916 ^ 1'b0 ;
  assign n12919 = n12811 ^ n7418 ^ 1'b0 ;
  assign n12920 = ( n2463 & ~n9114 ) | ( n2463 & n12272 ) | ( ~n9114 & n12272 ) ;
  assign n12921 = n6044 ^ n1180 ^ n628 ;
  assign n12922 = n12921 ^ n7107 ^ 1'b0 ;
  assign n12923 = ~n11979 & n12922 ;
  assign n12924 = ( n7308 & n7513 ) | ( n7308 & n12923 ) | ( n7513 & n12923 ) ;
  assign n12925 = ( n11964 & n12920 ) | ( n11964 & n12924 ) | ( n12920 & n12924 ) ;
  assign n12926 = n12925 ^ n4512 ^ n4066 ;
  assign n12927 = n12926 ^ n12626 ^ n5364 ;
  assign n12928 = n10442 ^ n574 ^ n326 ;
  assign n12929 = n2301 | n12928 ;
  assign n12930 = n8308 | n11233 ;
  assign n12931 = n12930 ^ n6822 ^ 1'b0 ;
  assign n12932 = n10124 ^ n7629 ^ n1059 ;
  assign n12933 = n12932 ^ n6372 ^ n3235 ;
  assign n12934 = n9530 ^ n8509 ^ n4189 ;
  assign n12935 = n6152 & ~n10785 ;
  assign n12936 = ( n3796 & n6686 ) | ( n3796 & n12935 ) | ( n6686 & n12935 ) ;
  assign n12937 = n7101 ^ n2974 ^ n1524 ;
  assign n12941 = n10578 ^ n6352 ^ n3129 ;
  assign n12942 = ( n8122 & n8990 ) | ( n8122 & n12941 ) | ( n8990 & n12941 ) ;
  assign n12938 = n635 ^ x42 ^ 1'b0 ;
  assign n12939 = n12938 ^ n3892 ^ n2341 ;
  assign n12940 = ( n2465 & ~n10506 ) | ( n2465 & n12939 ) | ( ~n10506 & n12939 ) ;
  assign n12943 = n12942 ^ n12940 ^ n2925 ;
  assign n12944 = n136 & ~n1657 ;
  assign n12945 = n3274 & n12944 ;
  assign n12947 = n3390 ^ x32 ^ 1'b0 ;
  assign n12948 = n12947 ^ n6698 ^ 1'b0 ;
  assign n12949 = n12041 | n12948 ;
  assign n12946 = ( n3069 & ~n4771 ) | ( n3069 & n9860 ) | ( ~n4771 & n9860 ) ;
  assign n12950 = n12949 ^ n12946 ^ 1'b0 ;
  assign n12951 = n11595 ^ n9130 ^ n426 ;
  assign n12952 = ( n12945 & n12950 ) | ( n12945 & n12951 ) | ( n12950 & n12951 ) ;
  assign n12953 = n12952 ^ n3478 ^ n2136 ;
  assign n12958 = n9534 ^ n7149 ^ n2996 ;
  assign n12959 = n12958 ^ n2099 ^ 1'b0 ;
  assign n12954 = ( n550 & ~n717 ) | ( n550 & n9749 ) | ( ~n717 & n9749 ) ;
  assign n12955 = ( ~n3165 & n5245 ) | ( ~n3165 & n7532 ) | ( n5245 & n7532 ) ;
  assign n12956 = n12955 ^ n5479 ^ n732 ;
  assign n12957 = ( n3688 & ~n12954 ) | ( n3688 & n12956 ) | ( ~n12954 & n12956 ) ;
  assign n12960 = n12959 ^ n12957 ^ n3968 ;
  assign n12963 = n8747 ^ x87 ^ 1'b0 ;
  assign n12964 = n12963 ^ n9245 ^ 1'b0 ;
  assign n12965 = n414 | n12964 ;
  assign n12961 = n7200 ^ n5672 ^ 1'b0 ;
  assign n12962 = n12961 ^ n2541 ^ n824 ;
  assign n12966 = n12965 ^ n12962 ^ n1848 ;
  assign n12967 = n12085 ^ n7335 ^ n2905 ;
  assign n12968 = ( n5275 & n12966 ) | ( n5275 & ~n12967 ) | ( n12966 & ~n12967 ) ;
  assign n12969 = ( n444 & n4076 ) | ( n444 & n5062 ) | ( n4076 & n5062 ) ;
  assign n12970 = n10759 ^ n2181 ^ n266 ;
  assign n12971 = ( n2005 & ~n12969 ) | ( n2005 & n12970 ) | ( ~n12969 & n12970 ) ;
  assign n12972 = ~n12968 & n12971 ;
  assign n12973 = ~n255 & n12972 ;
  assign n12979 = ( ~n7692 & n10570 ) | ( ~n7692 & n11371 ) | ( n10570 & n11371 ) ;
  assign n12976 = n12665 ^ n11839 ^ n7050 ;
  assign n12974 = n12700 ^ n10016 ^ n6378 ;
  assign n12975 = ( n2427 & n3089 ) | ( n2427 & ~n12974 ) | ( n3089 & ~n12974 ) ;
  assign n12977 = n12976 ^ n12975 ^ 1'b0 ;
  assign n12978 = ~n3254 & n12977 ;
  assign n12980 = n12979 ^ n12978 ^ n3565 ;
  assign n12985 = ( n1363 & ~n5463 ) | ( n1363 & n6422 ) | ( ~n5463 & n6422 ) ;
  assign n12981 = ( n2107 & ~n2650 ) | ( n2107 & n3551 ) | ( ~n2650 & n3551 ) ;
  assign n12982 = n10373 ^ n5837 ^ n595 ;
  assign n12983 = n4252 | n4444 ;
  assign n12984 = ( ~n12981 & n12982 ) | ( ~n12981 & n12983 ) | ( n12982 & n12983 ) ;
  assign n12986 = n12985 ^ n12984 ^ 1'b0 ;
  assign n12987 = n8007 | n12986 ;
  assign n12988 = n8915 ^ n3307 ^ n2985 ;
  assign n12989 = n7254 & ~n12988 ;
  assign n12990 = n12989 ^ n2213 ^ 1'b0 ;
  assign n12991 = ( n1633 & n5284 ) | ( n1633 & ~n10652 ) | ( n5284 & ~n10652 ) ;
  assign n12992 = n7460 ^ n7203 ^ n6384 ;
  assign n12993 = n1130 | n7898 ;
  assign n12994 = n12993 ^ n4049 ^ 1'b0 ;
  assign n12995 = n12994 ^ n3463 ^ x89 ;
  assign n12996 = ( n12991 & n12992 ) | ( n12991 & n12995 ) | ( n12992 & n12995 ) ;
  assign n12997 = ( ~n1205 & n4057 ) | ( ~n1205 & n10880 ) | ( n4057 & n10880 ) ;
  assign n12998 = n12958 ^ n4168 ^ n4053 ;
  assign n12999 = n12998 ^ n12216 ^ n4949 ;
  assign n13004 = ( n1089 & n1369 ) | ( n1089 & ~n6458 ) | ( n1369 & ~n6458 ) ;
  assign n13001 = n6242 ^ n2768 ^ 1'b0 ;
  assign n13002 = ~n6760 & n13001 ;
  assign n13000 = n7589 & ~n7974 ;
  assign n13003 = n13002 ^ n13000 ^ 1'b0 ;
  assign n13005 = n13004 ^ n13003 ^ n7171 ;
  assign n13006 = ( n5017 & n9451 ) | ( n5017 & ~n12476 ) | ( n9451 & ~n12476 ) ;
  assign n13007 = n13006 ^ n843 ^ 1'b0 ;
  assign n13008 = ~n5547 & n13007 ;
  assign n13009 = ( ~n5338 & n5869 ) | ( ~n5338 & n7377 ) | ( n5869 & n7377 ) ;
  assign n13010 = ( n422 & n5507 ) | ( n422 & n7106 ) | ( n5507 & n7106 ) ;
  assign n13011 = ( n3746 & n11257 ) | ( n3746 & n13010 ) | ( n11257 & n13010 ) ;
  assign n13012 = ~n13009 & n13011 ;
  assign n13013 = n13012 ^ n4962 ^ 1'b0 ;
  assign n13016 = n10052 ^ n8563 ^ 1'b0 ;
  assign n13017 = n1155 & ~n13016 ;
  assign n13015 = ~n1131 & n3819 ;
  assign n13018 = n13017 ^ n13015 ^ n4220 ;
  assign n13014 = n1110 & n5335 ;
  assign n13019 = n13018 ^ n13014 ^ n227 ;
  assign n13020 = n12356 ^ n11466 ^ n8209 ;
  assign n13022 = ~n1580 & n11450 ;
  assign n13023 = ~n11644 & n13022 ;
  assign n13021 = ( n5094 & n8405 ) | ( n5094 & ~n8457 ) | ( n8405 & ~n8457 ) ;
  assign n13024 = n13023 ^ n13021 ^ n9334 ;
  assign n13025 = ( n7237 & n9212 ) | ( n7237 & ~n11433 ) | ( n9212 & ~n11433 ) ;
  assign n13026 = n13025 ^ n8900 ^ n6272 ;
  assign n13027 = ( n4588 & n4698 ) | ( n4588 & ~n13026 ) | ( n4698 & ~n13026 ) ;
  assign n13028 = ( n4857 & n6336 ) | ( n4857 & ~n8472 ) | ( n6336 & ~n8472 ) ;
  assign n13029 = n13028 ^ n12070 ^ n5088 ;
  assign n13030 = ~n12224 & n12548 ;
  assign n13031 = ( ~n2741 & n13029 ) | ( ~n2741 & n13030 ) | ( n13029 & n13030 ) ;
  assign n13032 = ( n2619 & n7569 ) | ( n2619 & n8308 ) | ( n7569 & n8308 ) ;
  assign n13033 = ( n440 & n5547 ) | ( n440 & n12046 ) | ( n5547 & n12046 ) ;
  assign n13036 = ( n5015 & ~n6330 ) | ( n5015 & n6417 ) | ( ~n6330 & n6417 ) ;
  assign n13037 = ( n2607 & n3460 ) | ( n2607 & ~n13036 ) | ( n3460 & ~n13036 ) ;
  assign n13034 = n6837 & n8022 ;
  assign n13035 = n7270 & n13034 ;
  assign n13038 = n13037 ^ n13035 ^ n2551 ;
  assign n13039 = n13038 ^ n6152 ^ 1'b0 ;
  assign n13040 = n11064 & ~n13039 ;
  assign n13041 = n2035 | n4485 ;
  assign n13042 = n8185 ^ n7944 ^ n5180 ;
  assign n13043 = n3178 | n13042 ;
  assign n13047 = ( ~n11417 & n11507 ) | ( ~n11417 & n12534 ) | ( n11507 & n12534 ) ;
  assign n13048 = n13047 ^ n8458 ^ n3060 ;
  assign n13044 = n744 & n4848 ;
  assign n13045 = n13044 ^ n2627 ^ 1'b0 ;
  assign n13046 = n3795 & n13045 ;
  assign n13049 = n13048 ^ n13046 ^ n6427 ;
  assign n13050 = n1203 & n4541 ;
  assign n13051 = n9300 ^ n7161 ^ n1813 ;
  assign n13052 = n5196 & ~n13051 ;
  assign n13053 = n13052 ^ n11919 ^ n5779 ;
  assign n13054 = n10411 ^ n9909 ^ 1'b0 ;
  assign n13055 = n8256 | n13054 ;
  assign n13056 = n10893 ^ n10328 ^ n9414 ;
  assign n13057 = n5922 & n13056 ;
  assign n13058 = n13057 ^ n4634 ^ 1'b0 ;
  assign n13059 = n9642 ^ n7438 ^ 1'b0 ;
  assign n13060 = n13059 ^ n4066 ^ 1'b0 ;
  assign n13061 = ( n13055 & n13058 ) | ( n13055 & ~n13060 ) | ( n13058 & ~n13060 ) ;
  assign n13062 = ( n5791 & n8942 ) | ( n5791 & n10541 ) | ( n8942 & n10541 ) ;
  assign n13063 = ( ~n4865 & n8259 ) | ( ~n4865 & n9723 ) | ( n8259 & n9723 ) ;
  assign n13065 = ( ~n1427 & n4392 ) | ( ~n1427 & n12472 ) | ( n4392 & n12472 ) ;
  assign n13064 = ( ~n523 & n1103 ) | ( ~n523 & n4665 ) | ( n1103 & n4665 ) ;
  assign n13066 = n13065 ^ n13064 ^ n5919 ;
  assign n13067 = ( n4887 & ~n5700 ) | ( n4887 & n6172 ) | ( ~n5700 & n6172 ) ;
  assign n13068 = ( n293 & n10131 ) | ( n293 & ~n10215 ) | ( n10131 & ~n10215 ) ;
  assign n13072 = n7479 | n8947 ;
  assign n13073 = n13072 ^ n7541 ^ 1'b0 ;
  assign n13074 = ( n4781 & ~n6270 ) | ( n4781 & n13073 ) | ( ~n6270 & n13073 ) ;
  assign n13069 = n3220 ^ n1594 ^ n912 ;
  assign n13070 = ( n1152 & ~n5405 ) | ( n1152 & n13069 ) | ( ~n5405 & n13069 ) ;
  assign n13071 = ~n7808 & n13070 ;
  assign n13075 = n13074 ^ n13071 ^ n4984 ;
  assign n13076 = ( n5684 & n7076 ) | ( n5684 & ~n13075 ) | ( n7076 & ~n13075 ) ;
  assign n13077 = ( n7001 & n10386 ) | ( n7001 & ~n10685 ) | ( n10386 & ~n10685 ) ;
  assign n13078 = n13077 ^ n11542 ^ n1492 ;
  assign n13079 = ( n2917 & ~n5087 ) | ( n2917 & n7668 ) | ( ~n5087 & n7668 ) ;
  assign n13080 = ( n7387 & n8624 ) | ( n7387 & n13079 ) | ( n8624 & n13079 ) ;
  assign n13081 = n10809 ^ n4695 ^ n3141 ;
  assign n13082 = n11422 ^ x91 ^ 1'b0 ;
  assign n13083 = ( n4793 & n13081 ) | ( n4793 & n13082 ) | ( n13081 & n13082 ) ;
  assign n13084 = ( ~n13078 & n13080 ) | ( ~n13078 & n13083 ) | ( n13080 & n13083 ) ;
  assign n13085 = ( n326 & n2216 ) | ( n326 & n12984 ) | ( n2216 & n12984 ) ;
  assign n13086 = ( n164 & n535 ) | ( n164 & n12478 ) | ( n535 & n12478 ) ;
  assign n13087 = n13086 ^ n10299 ^ n735 ;
  assign n13088 = n13087 ^ n10879 ^ n3925 ;
  assign n13089 = n11433 ^ n9080 ^ n5659 ;
  assign n13090 = ( ~n7841 & n10089 ) | ( ~n7841 & n13089 ) | ( n10089 & n13089 ) ;
  assign n13092 = n12000 ^ n11650 ^ n1556 ;
  assign n13091 = ( n1119 & n1710 ) | ( n1119 & n3630 ) | ( n1710 & n3630 ) ;
  assign n13093 = n13092 ^ n13091 ^ 1'b0 ;
  assign n13094 = ( n4517 & n13090 ) | ( n4517 & n13093 ) | ( n13090 & n13093 ) ;
  assign n13095 = n2652 & n5611 ;
  assign n13096 = n13095 ^ n2500 ^ 1'b0 ;
  assign n13097 = ( n1565 & ~n13094 ) | ( n1565 & n13096 ) | ( ~n13094 & n13096 ) ;
  assign n13098 = n13097 ^ n12592 ^ n11269 ;
  assign n13099 = n5942 ^ n2623 ^ n2265 ;
  assign n13100 = n13099 ^ n12287 ^ n1160 ;
  assign n13101 = ( n6515 & n12003 ) | ( n6515 & n12975 ) | ( n12003 & n12975 ) ;
  assign n13102 = n8911 ^ n2015 ^ n529 ;
  assign n13115 = n8006 ^ n6752 ^ n3102 ;
  assign n13116 = n8875 ^ n4797 ^ n4646 ;
  assign n13117 = ( ~n1911 & n13115 ) | ( ~n1911 & n13116 ) | ( n13115 & n13116 ) ;
  assign n13109 = n7443 ^ n4877 ^ n173 ;
  assign n13111 = n5026 ^ n1427 ^ n373 ;
  assign n13110 = ( n2794 & ~n6169 ) | ( n2794 & n9172 ) | ( ~n6169 & n9172 ) ;
  assign n13112 = n13111 ^ n13110 ^ n4618 ;
  assign n13113 = n13109 & n13112 ;
  assign n13103 = n2498 ^ n544 ^ n368 ;
  assign n13104 = ( n521 & ~n11270 ) | ( n521 & n13103 ) | ( ~n11270 & n13103 ) ;
  assign n13105 = ( ~n2997 & n8355 ) | ( ~n2997 & n13104 ) | ( n8355 & n13104 ) ;
  assign n13106 = n9228 ^ n3889 ^ n1373 ;
  assign n13107 = n13106 ^ n11052 ^ n7824 ;
  assign n13108 = ( ~n9079 & n13105 ) | ( ~n9079 & n13107 ) | ( n13105 & n13107 ) ;
  assign n13114 = n13113 ^ n13108 ^ x95 ;
  assign n13118 = n13117 ^ n13114 ^ n11572 ;
  assign n13119 = n294 & ~n8838 ;
  assign n13120 = ~n1459 & n4145 ;
  assign n13121 = n13120 ^ n1921 ^ 1'b0 ;
  assign n13122 = n6253 & ~n13121 ;
  assign n13123 = n13122 ^ n6722 ^ n2436 ;
  assign n13124 = ( ~n1085 & n1990 ) | ( ~n1085 & n2630 ) | ( n1990 & n2630 ) ;
  assign n13125 = n13124 ^ n2458 ^ n2078 ;
  assign n13126 = ( n1742 & n3620 ) | ( n1742 & ~n13125 ) | ( n3620 & ~n13125 ) ;
  assign n13127 = n13126 ^ n5316 ^ n627 ;
  assign n13128 = ~n2393 & n9854 ;
  assign n13129 = ( n8212 & n10107 ) | ( n8212 & n13128 ) | ( n10107 & n13128 ) ;
  assign n13130 = ( n2340 & ~n2460 ) | ( n2340 & n7706 ) | ( ~n2460 & n7706 ) ;
  assign n13131 = n13130 ^ n10686 ^ 1'b0 ;
  assign n13132 = n5829 & n13131 ;
  assign n13137 = n8809 ^ n3629 ^ 1'b0 ;
  assign n13133 = n4486 ^ n2290 ^ n997 ;
  assign n13134 = n9107 ^ n5959 ^ n4149 ;
  assign n13135 = n13134 ^ n1310 ^ n954 ;
  assign n13136 = ~n13133 & n13135 ;
  assign n13138 = n13137 ^ n13136 ^ n1844 ;
  assign n13139 = n9356 ^ n7207 ^ n790 ;
  assign n13145 = n6665 ^ n4221 ^ n2216 ;
  assign n13140 = n3604 & n12047 ;
  assign n13141 = n12277 ^ n8924 ^ n685 ;
  assign n13142 = ( n232 & ~n13140 ) | ( n232 & n13141 ) | ( ~n13140 & n13141 ) ;
  assign n13143 = n13142 ^ n3329 ^ n393 ;
  assign n13144 = ( ~n6832 & n11375 ) | ( ~n6832 & n13143 ) | ( n11375 & n13143 ) ;
  assign n13146 = n13145 ^ n13144 ^ n345 ;
  assign n13147 = ( ~n4577 & n13139 ) | ( ~n4577 & n13146 ) | ( n13139 & n13146 ) ;
  assign n13148 = n12774 ^ n12607 ^ n7807 ;
  assign n13149 = n9212 ^ n6685 ^ n2589 ;
  assign n13150 = n13149 ^ n4648 ^ n477 ;
  assign n13151 = ~n3386 & n6777 ;
  assign n13152 = ~n5848 & n7006 ;
  assign n13153 = n13152 ^ n3602 ^ 1'b0 ;
  assign n13154 = n13153 ^ n7345 ^ n535 ;
  assign n13155 = n2913 | n5488 ;
  assign n13156 = n6221 & ~n13155 ;
  assign n13162 = ( n953 & n5194 ) | ( n953 & n12429 ) | ( n5194 & n12429 ) ;
  assign n13161 = n11422 ^ n906 ^ 1'b0 ;
  assign n13163 = n13162 ^ n13161 ^ n6192 ;
  assign n13164 = ( n3214 & ~n6393 ) | ( n3214 & n13163 ) | ( ~n6393 & n13163 ) ;
  assign n13157 = ( ~n837 & n5085 ) | ( ~n837 & n6406 ) | ( n5085 & n6406 ) ;
  assign n13158 = n8550 & ~n13157 ;
  assign n13159 = ~n5078 & n13158 ;
  assign n13160 = n13159 ^ n9904 ^ n1547 ;
  assign n13165 = n13164 ^ n13160 ^ 1'b0 ;
  assign n13166 = n9913 ^ n2452 ^ n139 ;
  assign n13167 = ( n4827 & n5159 ) | ( n4827 & ~n9590 ) | ( n5159 & ~n9590 ) ;
  assign n13168 = n6546 & ~n13167 ;
  assign n13174 = n2354 ^ n2241 ^ x28 ;
  assign n13175 = n13174 ^ n1985 ^ n550 ;
  assign n13170 = n4197 & ~n10066 ;
  assign n13171 = ( n3604 & n4235 ) | ( n3604 & ~n6055 ) | ( n4235 & ~n6055 ) ;
  assign n13172 = ~n1434 & n13171 ;
  assign n13173 = ~n13170 & n13172 ;
  assign n13169 = ( n5083 & n10207 ) | ( n5083 & ~n11614 ) | ( n10207 & ~n11614 ) ;
  assign n13176 = n13175 ^ n13173 ^ n13169 ;
  assign n13178 = ( n1999 & n7278 ) | ( n1999 & ~n10021 ) | ( n7278 & ~n10021 ) ;
  assign n13177 = n10218 ^ n6846 ^ n1897 ;
  assign n13179 = n13178 ^ n13177 ^ n4550 ;
  assign n13180 = n6920 ^ n3408 ^ n1844 ;
  assign n13181 = n13180 ^ n11321 ^ n5248 ;
  assign n13187 = n8191 ^ n6783 ^ n2019 ;
  assign n13185 = ( n5398 & n5562 ) | ( n5398 & n7600 ) | ( n5562 & n7600 ) ;
  assign n13186 = n13185 ^ n12388 ^ n4527 ;
  assign n13182 = ( n2604 & n3616 ) | ( n2604 & ~n5476 ) | ( n3616 & ~n5476 ) ;
  assign n13183 = n13182 ^ n4469 ^ 1'b0 ;
  assign n13184 = ~n3039 & n13183 ;
  assign n13188 = n13187 ^ n13186 ^ n13184 ;
  assign n13189 = n10878 ^ n5018 ^ n632 ;
  assign n13190 = n13189 ^ n12451 ^ n5027 ;
  assign n13191 = ( n367 & n5704 ) | ( n367 & ~n7622 ) | ( n5704 & ~n7622 ) ;
  assign n13192 = ( n952 & ~n8476 ) | ( n952 & n9959 ) | ( ~n8476 & n9959 ) ;
  assign n13193 = n13192 ^ n6059 ^ n2462 ;
  assign n13194 = ( n932 & n1301 ) | ( n932 & ~n8458 ) | ( n1301 & ~n8458 ) ;
  assign n13195 = n6608 ^ n981 ^ 1'b0 ;
  assign n13196 = n13195 ^ n11939 ^ 1'b0 ;
  assign n13197 = ( n13193 & n13194 ) | ( n13193 & ~n13196 ) | ( n13194 & ~n13196 ) ;
  assign n13198 = n11349 ^ n5491 ^ n1653 ;
  assign n13199 = ( n3631 & n3791 ) | ( n3631 & n8247 ) | ( n3791 & n8247 ) ;
  assign n13200 = n13199 ^ n9127 ^ n482 ;
  assign n13201 = n13200 ^ n5501 ^ 1'b0 ;
  assign n13202 = n13198 & ~n13201 ;
  assign n13203 = ( n1621 & n3583 ) | ( n1621 & n13202 ) | ( n3583 & n13202 ) ;
  assign n13204 = n13203 ^ n9753 ^ n7074 ;
  assign n13209 = ( n255 & ~n563 ) | ( n255 & n9237 ) | ( ~n563 & n9237 ) ;
  assign n13206 = n4513 ^ n657 ^ n575 ;
  assign n13205 = n6138 ^ n5916 ^ n474 ;
  assign n13207 = n13206 ^ n13205 ^ n729 ;
  assign n13208 = n13207 ^ n7590 ^ n705 ;
  assign n13210 = n13209 ^ n13208 ^ n12922 ;
  assign n13211 = ( n1130 & ~n3718 ) | ( n1130 & n9142 ) | ( ~n3718 & n9142 ) ;
  assign n13214 = ( n1208 & ~n5508 ) | ( n1208 & n8407 ) | ( ~n5508 & n8407 ) ;
  assign n13215 = ( ~n3868 & n4064 ) | ( ~n3868 & n13214 ) | ( n4064 & n13214 ) ;
  assign n13216 = ( ~n2679 & n12437 ) | ( ~n2679 & n13215 ) | ( n12437 & n13215 ) ;
  assign n13212 = ( n2016 & n4852 ) | ( n2016 & n6787 ) | ( n4852 & n6787 ) ;
  assign n13213 = n9359 | n13212 ;
  assign n13217 = n13216 ^ n13213 ^ 1'b0 ;
  assign n13218 = n5443 ^ n1180 ^ 1'b0 ;
  assign n13219 = ~n3504 & n11749 ;
  assign n13220 = n13219 ^ n4574 ^ 1'b0 ;
  assign n13221 = ( ~n4331 & n10131 ) | ( ~n4331 & n13220 ) | ( n10131 & n13220 ) ;
  assign n13222 = ( n3734 & n4561 ) | ( n3734 & ~n5095 ) | ( n4561 & ~n5095 ) ;
  assign n13223 = n13222 ^ n12767 ^ n4982 ;
  assign n13224 = n10190 ^ n7933 ^ n2178 ;
  assign n13225 = ( n6133 & ~n13223 ) | ( n6133 & n13224 ) | ( ~n13223 & n13224 ) ;
  assign n13226 = ( n855 & n1522 ) | ( n855 & ~n2908 ) | ( n1522 & ~n2908 ) ;
  assign n13227 = ( ~n2091 & n8505 ) | ( ~n2091 & n11139 ) | ( n8505 & n11139 ) ;
  assign n13228 = ( n10349 & n13226 ) | ( n10349 & ~n13227 ) | ( n13226 & ~n13227 ) ;
  assign n13229 = ( n1207 & ~n7645 ) | ( n1207 & n13228 ) | ( ~n7645 & n13228 ) ;
  assign n13230 = ( n1632 & ~n5727 ) | ( n1632 & n12733 ) | ( ~n5727 & n12733 ) ;
  assign n13231 = n5865 ^ n3643 ^ n914 ;
  assign n13232 = ~n9806 & n13231 ;
  assign n13233 = ( n939 & n7429 ) | ( n939 & n9361 ) | ( n7429 & n9361 ) ;
  assign n13234 = n13233 ^ n2988 ^ n1655 ;
  assign n13235 = n6554 & ~n12683 ;
  assign n13236 = ( n3972 & n10550 ) | ( n3972 & n13235 ) | ( n10550 & n13235 ) ;
  assign n13237 = n3412 & n9595 ;
  assign n13238 = ~n5673 & n13237 ;
  assign n13239 = n12319 ^ n6484 ^ n5747 ;
  assign n13240 = ( n4480 & n4633 ) | ( n4480 & n13239 ) | ( n4633 & n13239 ) ;
  assign n13241 = ( ~n10599 & n13238 ) | ( ~n10599 & n13240 ) | ( n13238 & n13240 ) ;
  assign n13245 = n9784 ^ n1310 ^ n1230 ;
  assign n13246 = ( n2501 & n6893 ) | ( n2501 & ~n13245 ) | ( n6893 & ~n13245 ) ;
  assign n13242 = n9235 ^ n9171 ^ n4723 ;
  assign n13243 = n13242 ^ n10257 ^ n4207 ;
  assign n13244 = ( ~n3406 & n11277 ) | ( ~n3406 & n13243 ) | ( n11277 & n13243 ) ;
  assign n13247 = n13246 ^ n13244 ^ 1'b0 ;
  assign n13248 = n11816 & ~n13247 ;
  assign n13255 = n2744 ^ n2297 ^ n309 ;
  assign n13256 = ( ~n2574 & n2614 ) | ( ~n2574 & n13255 ) | ( n2614 & n13255 ) ;
  assign n13253 = n10044 ^ n2229 ^ x18 ;
  assign n13254 = n13253 ^ n11797 ^ n4512 ;
  assign n13249 = n7640 ^ n5535 ^ n1993 ;
  assign n13250 = ( ~n3123 & n8446 ) | ( ~n3123 & n13249 ) | ( n8446 & n13249 ) ;
  assign n13251 = n13250 ^ n9967 ^ n992 ;
  assign n13252 = n13251 ^ n10189 ^ 1'b0 ;
  assign n13257 = n13256 ^ n13254 ^ n13252 ;
  assign n13258 = n3301 ^ n2629 ^ n1359 ;
  assign n13259 = n7364 ^ n6119 ^ n599 ;
  assign n13260 = n608 & n13259 ;
  assign n13261 = ( n711 & ~n2009 ) | ( n711 & n2243 ) | ( ~n2009 & n2243 ) ;
  assign n13262 = n13261 ^ n10228 ^ n5564 ;
  assign n13267 = ( n3522 & ~n3570 ) | ( n3522 & n4759 ) | ( ~n3570 & n4759 ) ;
  assign n13266 = ( n174 & ~n3588 ) | ( n174 & n13140 ) | ( ~n3588 & n13140 ) ;
  assign n13264 = ( n493 & n3874 ) | ( n493 & n8677 ) | ( n3874 & n8677 ) ;
  assign n13263 = ( x82 & n7692 ) | ( x82 & n12685 ) | ( n7692 & n12685 ) ;
  assign n13265 = n13264 ^ n13263 ^ n743 ;
  assign n13268 = n13267 ^ n13266 ^ n13265 ;
  assign n13269 = ( n8408 & n13094 ) | ( n8408 & ~n13268 ) | ( n13094 & ~n13268 ) ;
  assign n13270 = n4518 ^ n2243 ^ 1'b0 ;
  assign n13271 = n761 & n13270 ;
  assign n13272 = ~n1511 & n4140 ;
  assign n13273 = ( n4325 & n5606 ) | ( n4325 & n13272 ) | ( n5606 & n13272 ) ;
  assign n13274 = ( ~n6446 & n12412 ) | ( ~n6446 & n13273 ) | ( n12412 & n13273 ) ;
  assign n13275 = ( ~n5622 & n13271 ) | ( ~n5622 & n13274 ) | ( n13271 & n13274 ) ;
  assign n13276 = n2262 ^ n1836 ^ 1'b0 ;
  assign n13277 = n874 & n13276 ;
  assign n13278 = n13277 ^ n12479 ^ n4278 ;
  assign n13279 = n11661 ^ n10314 ^ n2493 ;
  assign n13280 = ( n13275 & n13278 ) | ( n13275 & n13279 ) | ( n13278 & n13279 ) ;
  assign n13281 = n8279 ^ n3574 ^ n1056 ;
  assign n13282 = ( n557 & ~n10344 ) | ( n557 & n10444 ) | ( ~n10344 & n10444 ) ;
  assign n13283 = n8344 ^ n3553 ^ n145 ;
  assign n13284 = ( ~n11882 & n13282 ) | ( ~n11882 & n13283 ) | ( n13282 & n13283 ) ;
  assign n13285 = n13284 ^ n7572 ^ 1'b0 ;
  assign n13286 = n9200 & ~n13285 ;
  assign n13287 = ( n12020 & n13281 ) | ( n12020 & n13286 ) | ( n13281 & n13286 ) ;
  assign n13288 = n13287 ^ n13227 ^ n6631 ;
  assign n13290 = n5093 ^ n1297 ^ n1157 ;
  assign n13291 = n13290 ^ n6347 ^ 1'b0 ;
  assign n13292 = n8147 & n13291 ;
  assign n13289 = n4408 ^ n4134 ^ 1'b0 ;
  assign n13293 = n13292 ^ n13289 ^ n5052 ;
  assign n13294 = ( n237 & ~n437 ) | ( n237 & n4178 ) | ( ~n437 & n4178 ) ;
  assign n13295 = n8007 & ~n13294 ;
  assign n13296 = n6523 ^ n5033 ^ n4132 ;
  assign n13297 = ( n1472 & n2636 ) | ( n1472 & n3079 ) | ( n2636 & n3079 ) ;
  assign n13298 = ( n10124 & ~n10401 ) | ( n10124 & n13297 ) | ( ~n10401 & n13297 ) ;
  assign n13299 = ( n3101 & n3204 ) | ( n3101 & n13298 ) | ( n3204 & n13298 ) ;
  assign n13300 = n12343 & ~n13299 ;
  assign n13301 = ~n12966 & n13300 ;
  assign n13302 = ( n7916 & n13296 ) | ( n7916 & n13301 ) | ( n13296 & n13301 ) ;
  assign n13303 = n7648 ^ n2902 ^ n2573 ;
  assign n13304 = n3795 ^ n1711 ^ n1640 ;
  assign n13305 = n13304 ^ n806 ^ n342 ;
  assign n13306 = n3708 | n13305 ;
  assign n13307 = n13306 ^ n3374 ^ 1'b0 ;
  assign n13308 = n12387 ^ n3665 ^ n2692 ;
  assign n13309 = ( n5771 & n9034 ) | ( n5771 & n12451 ) | ( n9034 & n12451 ) ;
  assign n13310 = n13309 ^ n759 ^ 1'b0 ;
  assign n13311 = n13308 | n13310 ;
  assign n13312 = ( n13303 & ~n13307 ) | ( n13303 & n13311 ) | ( ~n13307 & n13311 ) ;
  assign n13319 = ( n6126 & n8750 ) | ( n6126 & ~n9052 ) | ( n8750 & ~n9052 ) ;
  assign n13317 = ( n585 & n7411 ) | ( n585 & n7841 ) | ( n7411 & n7841 ) ;
  assign n13318 = n13317 ^ n7587 ^ n2162 ;
  assign n13313 = n5843 & n12409 ;
  assign n13314 = n13313 ^ n6565 ^ 1'b0 ;
  assign n13315 = n8096 ^ n2570 ^ n2351 ;
  assign n13316 = ( n726 & n13314 ) | ( n726 & ~n13315 ) | ( n13314 & ~n13315 ) ;
  assign n13320 = n13319 ^ n13318 ^ n13316 ;
  assign n13321 = n13320 ^ n4285 ^ n4226 ;
  assign n13322 = ( ~n987 & n3102 ) | ( ~n987 & n3397 ) | ( n3102 & n3397 ) ;
  assign n13324 = n1298 ^ n969 ^ 1'b0 ;
  assign n13325 = n13324 ^ n5637 ^ n715 ;
  assign n13323 = n4589 ^ n2117 ^ n1131 ;
  assign n13326 = n13325 ^ n13323 ^ n2833 ;
  assign n13327 = ( n6480 & n10652 ) | ( n6480 & ~n13326 ) | ( n10652 & ~n13326 ) ;
  assign n13328 = ( ~n6105 & n6299 ) | ( ~n6105 & n13327 ) | ( n6299 & n13327 ) ;
  assign n13329 = n3237 & ~n6706 ;
  assign n13330 = n13329 ^ n9614 ^ n6228 ;
  assign n13335 = ( ~n1083 & n3421 ) | ( ~n1083 & n8827 ) | ( n3421 & n8827 ) ;
  assign n13331 = ( n6243 & ~n8495 ) | ( n6243 & n9325 ) | ( ~n8495 & n9325 ) ;
  assign n13332 = n13331 ^ n6715 ^ n391 ;
  assign n13333 = n1847 & n7700 ;
  assign n13334 = n13332 & n13333 ;
  assign n13336 = n13335 ^ n13334 ^ n1313 ;
  assign n13337 = ( n3289 & n3552 ) | ( n3289 & ~n6760 ) | ( n3552 & ~n6760 ) ;
  assign n13338 = ( n8470 & ~n8828 ) | ( n8470 & n13337 ) | ( ~n8828 & n13337 ) ;
  assign n13339 = ( ~n5373 & n7071 ) | ( ~n5373 & n8222 ) | ( n7071 & n8222 ) ;
  assign n13340 = ( ~n5632 & n9819 ) | ( ~n5632 & n13339 ) | ( n9819 & n13339 ) ;
  assign n13341 = n12581 ^ n5785 ^ n649 ;
  assign n13342 = ~n3665 & n13341 ;
  assign n13343 = ( ~n2524 & n13340 ) | ( ~n2524 & n13342 ) | ( n13340 & n13342 ) ;
  assign n13344 = n11666 ^ n4663 ^ n3237 ;
  assign n13345 = ( ~n1327 & n3202 ) | ( ~n1327 & n4958 ) | ( n3202 & n4958 ) ;
  assign n13346 = ( n1295 & n7368 ) | ( n1295 & n13345 ) | ( n7368 & n13345 ) ;
  assign n13347 = ( n7514 & ~n10353 ) | ( n7514 & n13346 ) | ( ~n10353 & n13346 ) ;
  assign n13348 = n12872 ^ n11480 ^ n10842 ;
  assign n13349 = n13348 ^ n2674 ^ n2189 ;
  assign n13355 = n11608 ^ n2775 ^ n1934 ;
  assign n13356 = ( n1547 & ~n8134 ) | ( n1547 & n13355 ) | ( ~n8134 & n13355 ) ;
  assign n13351 = ~n1105 & n2890 ;
  assign n13352 = ~n9569 & n13351 ;
  assign n13353 = n13352 ^ n1796 ^ 1'b0 ;
  assign n13354 = n13353 ^ n9962 ^ n6600 ;
  assign n13350 = n12363 ^ n4537 ^ n3640 ;
  assign n13357 = n13356 ^ n13354 ^ n13350 ;
  assign n13358 = ~n6397 & n13357 ;
  assign n13359 = ~n5111 & n13358 ;
  assign n13366 = n2897 & n7695 ;
  assign n13367 = ~n1721 & n13366 ;
  assign n13368 = n13367 ^ n6188 ^ n5337 ;
  assign n13363 = n4540 ^ n4128 ^ n1277 ;
  assign n13364 = ( ~n9603 & n10893 ) | ( ~n9603 & n13363 ) | ( n10893 & n13363 ) ;
  assign n13361 = ~n1813 & n3793 ;
  assign n13362 = n4188 & n13361 ;
  assign n13360 = ( n387 & n1026 ) | ( n387 & ~n11439 ) | ( n1026 & ~n11439 ) ;
  assign n13365 = n13364 ^ n13362 ^ n13360 ;
  assign n13369 = n13368 ^ n13365 ^ n9012 ;
  assign n13370 = ( n588 & ~n2032 ) | ( n588 & n4707 ) | ( ~n2032 & n4707 ) ;
  assign n13371 = n13370 ^ n3916 ^ 1'b0 ;
  assign n13372 = ~n13369 & n13371 ;
  assign n13373 = ( n575 & ~n6192 ) | ( n575 & n9333 ) | ( ~n6192 & n9333 ) ;
  assign n13374 = ( n6171 & n7342 ) | ( n6171 & ~n7375 ) | ( n7342 & ~n7375 ) ;
  assign n13375 = ~n4832 & n13374 ;
  assign n13376 = n3261 ^ n3105 ^ n781 ;
  assign n13382 = ( n3055 & n5974 ) | ( n3055 & n11161 ) | ( n5974 & n11161 ) ;
  assign n13383 = ( n881 & n10216 ) | ( n881 & n13382 ) | ( n10216 & n13382 ) ;
  assign n13384 = ( n3637 & n4860 ) | ( n3637 & ~n13383 ) | ( n4860 & ~n13383 ) ;
  assign n13377 = ( n2153 & n4189 ) | ( n2153 & ~n8518 ) | ( n4189 & ~n8518 ) ;
  assign n13378 = ( n1004 & ~n5260 ) | ( n1004 & n13377 ) | ( ~n5260 & n13377 ) ;
  assign n13379 = ( ~n990 & n2377 ) | ( ~n990 & n13378 ) | ( n2377 & n13378 ) ;
  assign n13380 = n4171 & ~n13379 ;
  assign n13381 = ~x86 & n13380 ;
  assign n13385 = n13384 ^ n13381 ^ 1'b0 ;
  assign n13386 = ~n13376 & n13385 ;
  assign n13387 = n2513 ^ n1441 ^ n1114 ;
  assign n13388 = n13387 ^ n11738 ^ n4269 ;
  assign n13396 = n11769 ^ n3702 ^ n1261 ;
  assign n13397 = ( n3257 & ~n10718 ) | ( n3257 & n13396 ) | ( ~n10718 & n13396 ) ;
  assign n13394 = n3989 ^ n1014 ^ n700 ;
  assign n13389 = ( n1016 & n3982 ) | ( n1016 & ~n10179 ) | ( n3982 & ~n10179 ) ;
  assign n13390 = n13389 ^ n3704 ^ n2498 ;
  assign n13391 = ( ~n3392 & n12912 ) | ( ~n3392 & n13390 ) | ( n12912 & n13390 ) ;
  assign n13392 = n13391 ^ n3438 ^ 1'b0 ;
  assign n13393 = ( x5 & ~n3709 ) | ( x5 & n13392 ) | ( ~n3709 & n13392 ) ;
  assign n13395 = n13394 ^ n13393 ^ n9876 ;
  assign n13398 = n13397 ^ n13395 ^ n3537 ;
  assign n13399 = n5497 & n13398 ;
  assign n13402 = n2331 & n5494 ;
  assign n13403 = ~n13325 & n13402 ;
  assign n13404 = ( n3485 & n3824 ) | ( n3485 & n13403 ) | ( n3824 & n13403 ) ;
  assign n13400 = n10852 ^ n929 ^ 1'b0 ;
  assign n13401 = n13400 ^ n11975 ^ n3395 ;
  assign n13405 = n13404 ^ n13401 ^ n12252 ;
  assign n13406 = n9130 ^ n2237 ^ n258 ;
  assign n13407 = n4790 | n13406 ;
  assign n13408 = n12171 | n13407 ;
  assign n13411 = ~n9324 & n9881 ;
  assign n13412 = ( n829 & n1390 ) | ( n829 & n13411 ) | ( n1390 & n13411 ) ;
  assign n13409 = n8754 ^ n4245 ^ 1'b0 ;
  assign n13410 = n2698 & ~n13409 ;
  assign n13413 = n13412 ^ n13410 ^ n5249 ;
  assign n13414 = n5693 ^ n5257 ^ n2525 ;
  assign n13415 = ( n3647 & ~n4958 ) | ( n3647 & n6217 ) | ( ~n4958 & n6217 ) ;
  assign n13416 = n4028 ^ n3957 ^ n687 ;
  assign n13417 = ( n4463 & n5865 ) | ( n4463 & n8221 ) | ( n5865 & n8221 ) ;
  assign n13418 = ( n13415 & ~n13416 ) | ( n13415 & n13417 ) | ( ~n13416 & n13417 ) ;
  assign n13419 = ( ~n155 & n13414 ) | ( ~n155 & n13418 ) | ( n13414 & n13418 ) ;
  assign n13420 = ( n480 & n1032 ) | ( n480 & n1585 ) | ( n1032 & n1585 ) ;
  assign n13421 = n12638 ^ n10975 ^ 1'b0 ;
  assign n13422 = n13420 & ~n13421 ;
  assign n13423 = n9212 ^ n4049 ^ n2243 ;
  assign n13424 = n10566 ^ n8584 ^ n6932 ;
  assign n13425 = n7976 | n13424 ;
  assign n13426 = n2451 & ~n13425 ;
  assign n13427 = ( n11507 & n13423 ) | ( n11507 & ~n13426 ) | ( n13423 & ~n13426 ) ;
  assign n13428 = n11864 ^ n7389 ^ n3317 ;
  assign n13429 = ~n4896 & n13428 ;
  assign n13430 = n13429 ^ n8659 ^ 1'b0 ;
  assign n13431 = n10581 ^ n3873 ^ n1814 ;
  assign n13432 = ( ~n2471 & n2981 ) | ( ~n2471 & n3811 ) | ( n2981 & n3811 ) ;
  assign n13433 = n13432 ^ n4245 ^ n4055 ;
  assign n13434 = ( x103 & n13431 ) | ( x103 & n13433 ) | ( n13431 & n13433 ) ;
  assign n13435 = n11381 ^ n9522 ^ n6459 ;
  assign n13436 = n2178 | n13435 ;
  assign n13437 = n11066 ^ n7130 ^ 1'b0 ;
  assign n13438 = ( ~n7859 & n8080 ) | ( ~n7859 & n13437 ) | ( n8080 & n13437 ) ;
  assign n13439 = ( n5174 & ~n7341 ) | ( n5174 & n8713 ) | ( ~n7341 & n8713 ) ;
  assign n13440 = ( n9352 & n11721 ) | ( n9352 & n13439 ) | ( n11721 & n13439 ) ;
  assign n13441 = n12493 | n13440 ;
  assign n13442 = ( ~n740 & n13438 ) | ( ~n740 & n13441 ) | ( n13438 & n13441 ) ;
  assign n13446 = n4483 | n10841 ;
  assign n13447 = n5850 | n13446 ;
  assign n13443 = n3104 ^ n1951 ^ n793 ;
  assign n13444 = ( ~n2094 & n2636 ) | ( ~n2094 & n13443 ) | ( n2636 & n13443 ) ;
  assign n13445 = ~n6919 & n13444 ;
  assign n13448 = n13447 ^ n13445 ^ n13195 ;
  assign n13449 = n12281 ^ n9084 ^ n2435 ;
  assign n13450 = n4844 ^ n2658 ^ n949 ;
  assign n13451 = ( n259 & n941 ) | ( n259 & ~n13450 ) | ( n941 & ~n13450 ) ;
  assign n13452 = n8379 ^ n2308 ^ n301 ;
  assign n13453 = ( n9346 & ~n13451 ) | ( n9346 & n13452 ) | ( ~n13451 & n13452 ) ;
  assign n13459 = n5544 ^ n5039 ^ n1845 ;
  assign n13460 = n13459 ^ n13308 ^ 1'b0 ;
  assign n13456 = n9465 ^ n7208 ^ n4082 ;
  assign n13454 = n5486 ^ n2937 ^ n160 ;
  assign n13455 = n13454 ^ n10103 ^ n8620 ;
  assign n13457 = n13456 ^ n13455 ^ n3602 ;
  assign n13458 = ( ~n3297 & n9972 ) | ( ~n3297 & n13457 ) | ( n9972 & n13457 ) ;
  assign n13461 = n13460 ^ n13458 ^ n1110 ;
  assign n13462 = n13461 ^ n10033 ^ n5217 ;
  assign n13463 = ( n1680 & n9909 ) | ( n1680 & ~n12065 ) | ( n9909 & ~n12065 ) ;
  assign n13464 = n252 | n3593 ;
  assign n13465 = n6379 | n13464 ;
  assign n13466 = n13465 ^ n9208 ^ 1'b0 ;
  assign n13467 = n13466 ^ n10189 ^ n7600 ;
  assign n13468 = ( ~n4011 & n5608 ) | ( ~n4011 & n9966 ) | ( n5608 & n9966 ) ;
  assign n13469 = ( n229 & n7015 ) | ( n229 & n13468 ) | ( n7015 & n13468 ) ;
  assign n13470 = ( n238 & n4546 ) | ( n238 & ~n10143 ) | ( n4546 & ~n10143 ) ;
  assign n13471 = n12633 ^ n3998 ^ n741 ;
  assign n13472 = ( n2288 & n9372 ) | ( n2288 & ~n13471 ) | ( n9372 & ~n13471 ) ;
  assign n13473 = ( n4423 & ~n4766 ) | ( n4423 & n12666 ) | ( ~n4766 & n12666 ) ;
  assign n13474 = ( ~x127 & n2295 ) | ( ~x127 & n13473 ) | ( n2295 & n13473 ) ;
  assign n13475 = n13474 ^ n7544 ^ n3280 ;
  assign n13476 = n9733 & ~n13475 ;
  assign n13477 = ~n13472 & n13476 ;
  assign n13489 = n10772 ^ n222 ^ 1'b0 ;
  assign n13485 = n3366 ^ n2622 ^ 1'b0 ;
  assign n13486 = n2410 & n13485 ;
  assign n13480 = ( ~n206 & n3451 ) | ( ~n206 & n5442 ) | ( n3451 & n5442 ) ;
  assign n13481 = n13480 ^ n7407 ^ n6504 ;
  assign n13482 = n13481 ^ n3446 ^ n519 ;
  assign n13479 = n8147 ^ n3912 ^ 1'b0 ;
  assign n13478 = ~n8926 & n11450 ;
  assign n13483 = n13482 ^ n13479 ^ n13478 ;
  assign n13484 = n6619 & ~n13483 ;
  assign n13487 = n13486 ^ n13484 ^ n6211 ;
  assign n13488 = ( n8530 & n9020 ) | ( n8530 & ~n13487 ) | ( n9020 & ~n13487 ) ;
  assign n13490 = n13489 ^ n13488 ^ n8197 ;
  assign n13491 = ( n500 & n2686 ) | ( n500 & n4656 ) | ( n2686 & n4656 ) ;
  assign n13492 = ( n1745 & n3081 ) | ( n1745 & ~n13491 ) | ( n3081 & ~n13491 ) ;
  assign n13493 = ( n1769 & n5362 ) | ( n1769 & ~n13492 ) | ( n5362 & ~n13492 ) ;
  assign n13494 = n13493 ^ n6233 ^ n4085 ;
  assign n13495 = n11693 ^ n10380 ^ n8635 ;
  assign n13496 = ( n903 & n1234 ) | ( n903 & ~n5834 ) | ( n1234 & ~n5834 ) ;
  assign n13497 = n13496 ^ n1943 ^ n699 ;
  assign n13498 = ( n2708 & n5164 ) | ( n2708 & n13497 ) | ( n5164 & n13497 ) ;
  assign n13499 = n8775 ^ n6630 ^ n2906 ;
  assign n13500 = n13499 ^ n10797 ^ 1'b0 ;
  assign n13501 = ( n2142 & ~n3115 ) | ( n2142 & n9280 ) | ( ~n3115 & n9280 ) ;
  assign n13502 = n7511 ^ n6606 ^ n1128 ;
  assign n13503 = n13502 ^ n4342 ^ n3716 ;
  assign n13504 = n7564 ^ n6285 ^ n5113 ;
  assign n13505 = n13504 ^ n9760 ^ n7876 ;
  assign n13506 = ( n8951 & ~n9436 ) | ( n8951 & n13505 ) | ( ~n9436 & n13505 ) ;
  assign n13507 = x90 | n3236 ;
  assign n13508 = n13507 ^ n12108 ^ n6366 ;
  assign n13509 = ( n3877 & n11316 ) | ( n3877 & ~n13240 ) | ( n11316 & ~n13240 ) ;
  assign n13510 = ( ~n654 & n3451 ) | ( ~n654 & n13509 ) | ( n3451 & n13509 ) ;
  assign n13511 = ( n3557 & ~n7118 ) | ( n3557 & n13277 ) | ( ~n7118 & n13277 ) ;
  assign n13512 = ( ~n2967 & n6473 ) | ( ~n2967 & n13511 ) | ( n6473 & n13511 ) ;
  assign n13513 = n5180 & n13512 ;
  assign n13514 = n12556 & n13513 ;
  assign n13515 = n13514 ^ n5381 ^ n2683 ;
  assign n13516 = n12011 ^ n10344 ^ n8579 ;
  assign n13517 = ( n867 & ~n2449 ) | ( n867 & n4043 ) | ( ~n2449 & n4043 ) ;
  assign n13518 = n13517 ^ n1719 ^ 1'b0 ;
  assign n13519 = ( ~n7226 & n8220 ) | ( ~n7226 & n13518 ) | ( n8220 & n13518 ) ;
  assign n13520 = n2697 ^ n1414 ^ n246 ;
  assign n13521 = n13520 ^ n7233 ^ n3112 ;
  assign n13522 = n8035 ^ n2757 ^ x113 ;
  assign n13523 = ( n5112 & n6952 ) | ( n5112 & n13522 ) | ( n6952 & n13522 ) ;
  assign n13524 = ( n7461 & n8877 ) | ( n7461 & ~n13523 ) | ( n8877 & ~n13523 ) ;
  assign n13529 = n6821 ^ n1897 ^ n1013 ;
  assign n13526 = ( n4486 & n8740 ) | ( n4486 & ~n10728 ) | ( n8740 & ~n10728 ) ;
  assign n13527 = n13526 ^ n2075 ^ 1'b0 ;
  assign n13525 = n11690 ^ n6536 ^ n5444 ;
  assign n13528 = n13527 ^ n13525 ^ n6986 ;
  assign n13530 = n13529 ^ n13528 ^ n9020 ;
  assign n13531 = n10842 ^ n7792 ^ n1352 ;
  assign n13532 = ( n10561 & ~n10734 ) | ( n10561 & n13531 ) | ( ~n10734 & n13531 ) ;
  assign n13533 = n13532 ^ n6689 ^ n4029 ;
  assign n13534 = n4358 ^ n650 ^ 1'b0 ;
  assign n13535 = ~n3232 & n13534 ;
  assign n13536 = n5087 & n13535 ;
  assign n13537 = n7458 & ~n13536 ;
  assign n13538 = ( n1020 & n4355 ) | ( n1020 & n13537 ) | ( n4355 & n13537 ) ;
  assign n13539 = n627 & n11331 ;
  assign n13540 = n13539 ^ n1166 ^ 1'b0 ;
  assign n13541 = n9237 ^ n7544 ^ n1081 ;
  assign n13545 = x80 & n6624 ;
  assign n13546 = n366 & n13545 ;
  assign n13547 = n2395 & n13546 ;
  assign n13542 = ( n3889 & n6837 ) | ( n3889 & n10447 ) | ( n6837 & n10447 ) ;
  assign n13543 = ( n5468 & ~n7324 ) | ( n5468 & n13542 ) | ( ~n7324 & n13542 ) ;
  assign n13544 = n13543 ^ n10833 ^ n3386 ;
  assign n13548 = n13547 ^ n13544 ^ n1888 ;
  assign n13549 = n13541 & n13548 ;
  assign n13550 = n13549 ^ n11527 ^ 1'b0 ;
  assign n13552 = n7403 ^ n4537 ^ n988 ;
  assign n13551 = ( n3444 & n6253 ) | ( n3444 & ~n7860 ) | ( n6253 & ~n7860 ) ;
  assign n13553 = n13552 ^ n13551 ^ n11859 ;
  assign n13554 = n10216 ^ n5618 ^ n1803 ;
  assign n13555 = n13554 ^ n11881 ^ 1'b0 ;
  assign n13556 = ( n8875 & ~n13553 ) | ( n8875 & n13555 ) | ( ~n13553 & n13555 ) ;
  assign n13557 = n13556 ^ n13357 ^ 1'b0 ;
  assign n13560 = ( n2440 & ~n2821 ) | ( n2440 & n6523 ) | ( ~n2821 & n6523 ) ;
  assign n13561 = n2090 ^ n1492 ^ n688 ;
  assign n13562 = ( n1649 & ~n1659 ) | ( n1649 & n2820 ) | ( ~n1659 & n2820 ) ;
  assign n13563 = ( n833 & n13561 ) | ( n833 & n13562 ) | ( n13561 & n13562 ) ;
  assign n13564 = ( n2931 & n13560 ) | ( n2931 & n13563 ) | ( n13560 & n13563 ) ;
  assign n13558 = n1783 & ~n9758 ;
  assign n13559 = n13558 ^ n12195 ^ 1'b0 ;
  assign n13565 = n13564 ^ n13559 ^ 1'b0 ;
  assign n13566 = n6828 ^ n3720 ^ 1'b0 ;
  assign n13567 = n4697 & ~n7255 ;
  assign n13568 = ~n13566 & n13567 ;
  assign n13569 = n13568 ^ n12548 ^ 1'b0 ;
  assign n13570 = n13112 & n13569 ;
  assign n13571 = n8317 ^ n1529 ^ n1201 ;
  assign n13572 = ( n6958 & n8571 ) | ( n6958 & n13571 ) | ( n8571 & n13571 ) ;
  assign n13574 = ( n4563 & n10222 ) | ( n4563 & n13261 ) | ( n10222 & n13261 ) ;
  assign n13573 = ( n1994 & n6006 ) | ( n1994 & n7455 ) | ( n6006 & n7455 ) ;
  assign n13575 = n13574 ^ n13573 ^ 1'b0 ;
  assign n13576 = ~n8881 & n13575 ;
  assign n13577 = n7948 ^ n1591 ^ 1'b0 ;
  assign n13578 = ( n2568 & n11128 ) | ( n2568 & n11511 ) | ( n11128 & n11511 ) ;
  assign n13579 = ( ~n1839 & n2223 ) | ( ~n1839 & n5966 ) | ( n2223 & n5966 ) ;
  assign n13580 = ~n1813 & n5040 ;
  assign n13581 = n13579 & n13580 ;
  assign n13582 = n13581 ^ n8795 ^ n7310 ;
  assign n13583 = ( ~n2416 & n13133 ) | ( ~n2416 & n13582 ) | ( n13133 & n13582 ) ;
  assign n13584 = n13583 ^ n11217 ^ n5364 ;
  assign n13585 = n13584 ^ n4875 ^ n1057 ;
  assign n13586 = n13585 ^ n6296 ^ n3615 ;
  assign n13587 = ( n13577 & n13578 ) | ( n13577 & ~n13586 ) | ( n13578 & ~n13586 ) ;
  assign n13588 = ( n634 & ~n9748 ) | ( n634 & n13587 ) | ( ~n9748 & n13587 ) ;
  assign n13589 = ( ~n5065 & n5538 ) | ( ~n5065 & n13058 ) | ( n5538 & n13058 ) ;
  assign n13590 = n6221 ^ n2888 ^ n1668 ;
  assign n13591 = ( ~n2916 & n5848 ) | ( ~n2916 & n5911 ) | ( n5848 & n5911 ) ;
  assign n13592 = n13591 ^ n8000 ^ n2155 ;
  assign n13593 = n13592 ^ n1562 ^ 1'b0 ;
  assign n13594 = n13590 & ~n13593 ;
  assign n13595 = n2473 | n2882 ;
  assign n13596 = n13595 ^ n459 ^ 1'b0 ;
  assign n13597 = n13596 ^ n3113 ^ n1602 ;
  assign n13598 = n8566 ^ n6202 ^ n437 ;
  assign n13599 = ( ~n9343 & n13597 ) | ( ~n9343 & n13598 ) | ( n13597 & n13598 ) ;
  assign n13600 = ( ~n463 & n720 ) | ( ~n463 & n9480 ) | ( n720 & n9480 ) ;
  assign n13604 = n7661 ^ n5132 ^ n2615 ;
  assign n13602 = n4755 ^ n1804 ^ n1292 ;
  assign n13601 = ( n426 & ~n1059 ) | ( n426 & n6255 ) | ( ~n1059 & n6255 ) ;
  assign n13603 = n13602 ^ n13601 ^ n10152 ;
  assign n13605 = n13604 ^ n13603 ^ n4929 ;
  assign n13606 = ( n3633 & n10021 ) | ( n3633 & ~n13605 ) | ( n10021 & ~n13605 ) ;
  assign n13607 = ( n8365 & ~n13600 ) | ( n8365 & n13606 ) | ( ~n13600 & n13606 ) ;
  assign n13609 = ( ~n1963 & n2596 ) | ( ~n1963 & n3676 ) | ( n2596 & n3676 ) ;
  assign n13608 = n1390 | n11555 ;
  assign n13610 = n13609 ^ n13608 ^ 1'b0 ;
  assign n13611 = ( ~n3963 & n13607 ) | ( ~n3963 & n13610 ) | ( n13607 & n13610 ) ;
  assign n13612 = n8392 & n13346 ;
  assign n13613 = n8502 & n13612 ;
  assign n13614 = n13613 ^ n9495 ^ n2394 ;
  assign n13615 = n6346 | n9288 ;
  assign n13626 = n6770 ^ n4020 ^ n1015 ;
  assign n13627 = ( n7665 & ~n11714 ) | ( n7665 & n13626 ) | ( ~n11714 & n13626 ) ;
  assign n13624 = n3658 ^ n1281 ^ 1'b0 ;
  assign n13623 = ( ~n1934 & n2998 ) | ( ~n1934 & n9513 ) | ( n2998 & n9513 ) ;
  assign n13622 = n13273 ^ n8872 ^ n5182 ;
  assign n13625 = n13624 ^ n13623 ^ n13622 ;
  assign n13616 = ( n1587 & n3162 ) | ( n1587 & ~n3365 ) | ( n3162 & ~n3365 ) ;
  assign n13617 = n13616 ^ n3249 ^ n3004 ;
  assign n13618 = n13617 ^ n2605 ^ n287 ;
  assign n13619 = n2984 ^ n1158 ^ n240 ;
  assign n13620 = ( ~n3919 & n12036 ) | ( ~n3919 & n13619 ) | ( n12036 & n13619 ) ;
  assign n13621 = ( ~n10553 & n13618 ) | ( ~n10553 & n13620 ) | ( n13618 & n13620 ) ;
  assign n13628 = n13627 ^ n13625 ^ n13621 ;
  assign n13635 = n10623 ^ n3898 ^ n2543 ;
  assign n13630 = n3478 ^ n572 ^ n438 ;
  assign n13631 = ( n6065 & n10277 ) | ( n6065 & ~n13630 ) | ( n10277 & ~n13630 ) ;
  assign n13629 = n4328 ^ n1015 ^ n769 ;
  assign n13632 = n13631 ^ n13629 ^ n11579 ;
  assign n13633 = ( n8672 & n13292 ) | ( n8672 & n13632 ) | ( n13292 & n13632 ) ;
  assign n13634 = ( n4730 & ~n13091 ) | ( n4730 & n13633 ) | ( ~n13091 & n13633 ) ;
  assign n13636 = n13635 ^ n13634 ^ n4056 ;
  assign n13637 = ( n13615 & ~n13628 ) | ( n13615 & n13636 ) | ( ~n13628 & n13636 ) ;
  assign n13638 = ( ~n2259 & n8682 ) | ( ~n2259 & n10321 ) | ( n8682 & n10321 ) ;
  assign n13639 = n3543 ^ n3086 ^ n2724 ;
  assign n13640 = ~n431 & n13639 ;
  assign n13641 = n13638 & n13640 ;
  assign n13642 = ( n2562 & ~n6233 ) | ( n2562 & n8317 ) | ( ~n6233 & n8317 ) ;
  assign n13643 = n6265 ^ n4929 ^ n2449 ;
  assign n13644 = n13643 ^ n11457 ^ n8607 ;
  assign n13645 = n13644 ^ n10027 ^ n3908 ;
  assign n13646 = ( n2557 & n11789 ) | ( n2557 & ~n13145 ) | ( n11789 & ~n13145 ) ;
  assign n13647 = ( n13642 & n13645 ) | ( n13642 & n13646 ) | ( n13645 & n13646 ) ;
  assign n13648 = n8118 ^ n7331 ^ 1'b0 ;
  assign n13649 = n10268 ^ n6364 ^ n3169 ;
  assign n13650 = n12430 ^ n6645 ^ x79 ;
  assign n13651 = ( n11474 & n13649 ) | ( n11474 & n13650 ) | ( n13649 & n13650 ) ;
  assign n13653 = n2157 ^ n2013 ^ n491 ;
  assign n13652 = ( n2314 & n6702 ) | ( n2314 & n13133 ) | ( n6702 & n13133 ) ;
  assign n13654 = n13653 ^ n13652 ^ n2699 ;
  assign n13655 = ( n255 & ~n7731 ) | ( n255 & n12839 ) | ( ~n7731 & n12839 ) ;
  assign n13656 = ( n2051 & n9523 ) | ( n2051 & ~n13655 ) | ( n9523 & ~n13655 ) ;
  assign n13657 = ( n3698 & n5142 ) | ( n3698 & ~n13596 ) | ( n5142 & ~n13596 ) ;
  assign n13658 = n13657 ^ n7875 ^ n5274 ;
  assign n13659 = n4144 ^ n1777 ^ 1'b0 ;
  assign n13660 = n13658 | n13659 ;
  assign n13661 = ( n13654 & n13656 ) | ( n13654 & ~n13660 ) | ( n13656 & ~n13660 ) ;
  assign n13662 = ( n423 & n945 ) | ( n423 & ~n12967 ) | ( n945 & ~n12967 ) ;
  assign n13663 = n13662 ^ n9049 ^ n8086 ;
  assign n13664 = ~n4006 & n13663 ;
  assign n13666 = ( ~n3710 & n5290 ) | ( ~n3710 & n8550 ) | ( n5290 & n8550 ) ;
  assign n13667 = n13666 ^ n4598 ^ n1690 ;
  assign n13665 = ( n1723 & n5398 ) | ( n1723 & n10735 ) | ( n5398 & n10735 ) ;
  assign n13668 = n13667 ^ n13665 ^ n4367 ;
  assign n13669 = n3801 ^ n3227 ^ 1'b0 ;
  assign n13670 = ~n13668 & n13669 ;
  assign n13671 = n8405 ^ n3139 ^ n1586 ;
  assign n13672 = n13671 ^ n5245 ^ 1'b0 ;
  assign n13673 = n3466 | n12634 ;
  assign n13674 = n13673 ^ n9173 ^ 1'b0 ;
  assign n13675 = ( n168 & n929 ) | ( n168 & n13674 ) | ( n929 & n13674 ) ;
  assign n13683 = ( n2943 & n6871 ) | ( n2943 & n11478 ) | ( n6871 & n11478 ) ;
  assign n13681 = n12120 ^ n2716 ^ n956 ;
  assign n13682 = n13681 ^ n8365 ^ n4598 ;
  assign n13679 = ( n4955 & ~n10065 ) | ( n4955 & n11471 ) | ( ~n10065 & n11471 ) ;
  assign n13677 = n1044 | n5153 ;
  assign n13676 = n4256 ^ n1288 ^ 1'b0 ;
  assign n13678 = n13677 ^ n13676 ^ n11132 ;
  assign n13680 = n13679 ^ n13678 ^ n6253 ;
  assign n13684 = n13683 ^ n13682 ^ n13680 ;
  assign n13685 = n13684 ^ n9776 ^ n8153 ;
  assign n13686 = n10716 ^ n5775 ^ n468 ;
  assign n13687 = n4470 ^ n1642 ^ 1'b0 ;
  assign n13688 = n1812 & n13687 ;
  assign n13689 = ( n1866 & ~n13686 ) | ( n1866 & n13688 ) | ( ~n13686 & n13688 ) ;
  assign n13691 = n5780 ^ n3160 ^ n1727 ;
  assign n13692 = ( n2055 & n2914 ) | ( n2055 & n13691 ) | ( n2914 & n13691 ) ;
  assign n13693 = n13692 ^ n3629 ^ 1'b0 ;
  assign n13694 = n681 | n13693 ;
  assign n13695 = n13694 ^ n4230 ^ n1300 ;
  assign n13690 = ( n4130 & n9201 ) | ( n4130 & ~n10884 ) | ( n9201 & ~n10884 ) ;
  assign n13696 = n13695 ^ n13690 ^ n8208 ;
  assign n13697 = ( n12922 & n13689 ) | ( n12922 & ~n13696 ) | ( n13689 & ~n13696 ) ;
  assign n13698 = ( n9696 & n13685 ) | ( n9696 & n13697 ) | ( n13685 & n13697 ) ;
  assign n13699 = ( n13672 & n13675 ) | ( n13672 & ~n13698 ) | ( n13675 & ~n13698 ) ;
  assign n13700 = n9816 ^ n5376 ^ n1114 ;
  assign n13701 = n13700 ^ n10268 ^ n534 ;
  assign n13702 = ( n3369 & n8241 ) | ( n3369 & n13701 ) | ( n8241 & n13701 ) ;
  assign n13703 = ( n194 & ~n200 ) | ( n194 & n9416 ) | ( ~n200 & n9416 ) ;
  assign n13704 = n13703 ^ n12779 ^ n7583 ;
  assign n13705 = ( n11220 & n13702 ) | ( n11220 & n13704 ) | ( n13702 & n13704 ) ;
  assign n13708 = ( n1679 & ~n2969 ) | ( n1679 & n5164 ) | ( ~n2969 & n5164 ) ;
  assign n13706 = n304 & n3178 ;
  assign n13707 = n13706 ^ n7633 ^ 1'b0 ;
  assign n13709 = n13708 ^ n13707 ^ n11175 ;
  assign n13710 = n3582 ^ n1654 ^ 1'b0 ;
  assign n13711 = n13710 ^ n13643 ^ n5875 ;
  assign n13712 = n8240 ^ n7410 ^ 1'b0 ;
  assign n13713 = n716 ^ n343 ^ x72 ;
  assign n13714 = ( n218 & n11291 ) | ( n218 & ~n13713 ) | ( n11291 & ~n13713 ) ;
  assign n13716 = ( ~n3333 & n4319 ) | ( ~n3333 & n7629 ) | ( n4319 & n7629 ) ;
  assign n13715 = ( n7088 & n8506 ) | ( n7088 & ~n8747 ) | ( n8506 & ~n8747 ) ;
  assign n13717 = n13716 ^ n13715 ^ n2279 ;
  assign n13718 = n12986 ^ n9391 ^ 1'b0 ;
  assign n13719 = n9520 | n13718 ;
  assign n13720 = ( n7333 & n7858 ) | ( n7333 & n8168 ) | ( n7858 & n8168 ) ;
  assign n13721 = n8223 ^ n5131 ^ 1'b0 ;
  assign n13722 = n13720 & ~n13721 ;
  assign n13723 = n13722 ^ n2118 ^ n1179 ;
  assign n13724 = ( ~n2037 & n3645 ) | ( ~n2037 & n5195 ) | ( n3645 & n5195 ) ;
  assign n13725 = ( n5161 & n10783 ) | ( n5161 & n13724 ) | ( n10783 & n13724 ) ;
  assign n13726 = ( ~n4063 & n4939 ) | ( ~n4063 & n13725 ) | ( n4939 & n13725 ) ;
  assign n13727 = ( n1603 & n10623 ) | ( n1603 & n11230 ) | ( n10623 & n11230 ) ;
  assign n13728 = n13727 ^ n13311 ^ n6622 ;
  assign n13729 = n9785 ^ n7346 ^ 1'b0 ;
  assign n13730 = n13729 ^ n11925 ^ 1'b0 ;
  assign n13731 = ( n4094 & n8241 ) | ( n4094 & ~n13730 ) | ( n8241 & ~n13730 ) ;
  assign n13732 = n13731 ^ n13249 ^ n3667 ;
  assign n13733 = n11580 ^ n9612 ^ n2617 ;
  assign n13734 = n11817 ^ n11489 ^ 1'b0 ;
  assign n13735 = ~n13733 & n13734 ;
  assign n13737 = ( x91 & n1162 ) | ( x91 & n2314 ) | ( n1162 & n2314 ) ;
  assign n13736 = n9224 ^ n6364 ^ n4291 ;
  assign n13738 = n13737 ^ n13736 ^ n6352 ;
  assign n13739 = n10334 ^ n6959 ^ n4799 ;
  assign n13740 = ( n2876 & n12385 ) | ( n2876 & ~n13739 ) | ( n12385 & ~n13739 ) ;
  assign n13743 = n6125 ^ n2211 ^ 1'b0 ;
  assign n13741 = n4222 ^ n2301 ^ n806 ;
  assign n13742 = ( ~n2520 & n9135 ) | ( ~n2520 & n13741 ) | ( n9135 & n13741 ) ;
  assign n13744 = n13743 ^ n13742 ^ n2103 ;
  assign n13748 = n9622 ^ n9153 ^ n7305 ;
  assign n13745 = n6275 & n10060 ;
  assign n13746 = n13745 ^ n12747 ^ n1970 ;
  assign n13747 = n10258 & n13746 ;
  assign n13749 = n13748 ^ n13747 ^ 1'b0 ;
  assign n13750 = ( ~n5241 & n7333 ) | ( ~n5241 & n12132 ) | ( n7333 & n12132 ) ;
  assign n13755 = n8687 ^ n943 ^ 1'b0 ;
  assign n13756 = n2180 | n13755 ;
  assign n13751 = ( ~n455 & n2431 ) | ( ~n455 & n5059 ) | ( n2431 & n5059 ) ;
  assign n13752 = n1616 ^ n448 ^ 1'b0 ;
  assign n13753 = n5278 & n13752 ;
  assign n13754 = ( n8327 & n13751 ) | ( n8327 & ~n13753 ) | ( n13751 & ~n13753 ) ;
  assign n13757 = n13756 ^ n13754 ^ n10994 ;
  assign n13758 = n13757 ^ n10131 ^ n3377 ;
  assign n13760 = n10601 ^ n5903 ^ n519 ;
  assign n13761 = n1477 | n13760 ;
  assign n13762 = n13761 ^ n10120 ^ 1'b0 ;
  assign n13759 = n6205 & ~n7194 ;
  assign n13763 = n13762 ^ n13759 ^ n1782 ;
  assign n13764 = n13763 ^ n7833 ^ n887 ;
  assign n13765 = n4739 ^ n1574 ^ n1404 ;
  assign n13766 = n3400 ^ n2041 ^ 1'b0 ;
  assign n13767 = n3406 & ~n13766 ;
  assign n13768 = ( n10408 & ~n13765 ) | ( n10408 & n13767 ) | ( ~n13765 & n13767 ) ;
  assign n13769 = n8139 ^ n6608 ^ n1885 ;
  assign n13770 = n11604 ^ n7597 ^ n410 ;
  assign n13771 = n7639 & n13770 ;
  assign n13772 = n13771 ^ n13481 ^ 1'b0 ;
  assign n13773 = ( ~n2771 & n11858 ) | ( ~n2771 & n12611 ) | ( n11858 & n12611 ) ;
  assign n13774 = n7411 ^ n2689 ^ n2565 ;
  assign n13775 = ( ~n612 & n1812 ) | ( ~n612 & n3046 ) | ( n1812 & n3046 ) ;
  assign n13776 = ( n5974 & n12401 ) | ( n5974 & n13775 ) | ( n12401 & n13775 ) ;
  assign n13777 = ( n3211 & ~n9886 ) | ( n3211 & n13776 ) | ( ~n9886 & n13776 ) ;
  assign n13778 = ( n11472 & n13774 ) | ( n11472 & ~n13777 ) | ( n13774 & ~n13777 ) ;
  assign n13779 = ( ~n1975 & n2718 ) | ( ~n1975 & n5304 ) | ( n2718 & n5304 ) ;
  assign n13780 = n13779 ^ n6543 ^ 1'b0 ;
  assign n13781 = n13780 ^ n4343 ^ n190 ;
  assign n13782 = ( n7979 & ~n8073 ) | ( n7979 & n11467 ) | ( ~n8073 & n11467 ) ;
  assign n13783 = ( n5659 & n6458 ) | ( n5659 & ~n8920 ) | ( n6458 & ~n8920 ) ;
  assign n13784 = n13783 ^ n6587 ^ n969 ;
  assign n13785 = n13784 ^ n12133 ^ 1'b0 ;
  assign n13786 = ~n4269 & n13785 ;
  assign n13787 = n5166 | n6230 ;
  assign n13788 = n9445 ^ n459 ^ 1'b0 ;
  assign n13789 = n11332 ^ n4093 ^ n3186 ;
  assign n13790 = n9149 ^ n6492 ^ n4196 ;
  assign n13791 = n12097 ^ n8090 ^ n2922 ;
  assign n13792 = ~n3968 & n8142 ;
  assign n13793 = n8207 ^ n3041 ^ 1'b0 ;
  assign n13794 = ~n13792 & n13793 ;
  assign n13795 = n2232 & ~n2473 ;
  assign n13796 = ~n13794 & n13795 ;
  assign n13797 = n11226 ^ n6964 ^ n2027 ;
  assign n13798 = n7801 ^ n4807 ^ n2063 ;
  assign n13799 = n13798 ^ n3709 ^ n2092 ;
  assign n13801 = ( n528 & ~n1697 ) | ( n528 & n2535 ) | ( ~n1697 & n2535 ) ;
  assign n13800 = n11689 ^ n6461 ^ n3597 ;
  assign n13802 = n13801 ^ n13800 ^ n5741 ;
  assign n13803 = ( n1183 & ~n2213 ) | ( n1183 & n5999 ) | ( ~n2213 & n5999 ) ;
  assign n13804 = n10852 ^ n2549 ^ n812 ;
  assign n13805 = n4775 ^ n3808 ^ n3750 ;
  assign n13806 = n13805 ^ n11274 ^ 1'b0 ;
  assign n13807 = ~n4575 & n13806 ;
  assign n13808 = n13807 ^ n10783 ^ 1'b0 ;
  assign n13809 = ~n319 & n13808 ;
  assign n13810 = ~n13804 & n13809 ;
  assign n13811 = n13803 | n13810 ;
  assign n13812 = n13802 & ~n13811 ;
  assign n13813 = ( n3988 & ~n8229 ) | ( n3988 & n9350 ) | ( ~n8229 & n9350 ) ;
  assign n13814 = ( ~n4008 & n5986 ) | ( ~n4008 & n12491 ) | ( n5986 & n12491 ) ;
  assign n13815 = ( n2099 & ~n8617 ) | ( n2099 & n13814 ) | ( ~n8617 & n13814 ) ;
  assign n13816 = ~n3198 & n10736 ;
  assign n13817 = n13816 ^ n9966 ^ n9480 ;
  assign n13818 = ( ~n499 & n6253 ) | ( ~n499 & n9657 ) | ( n6253 & n9657 ) ;
  assign n13819 = ( n1868 & n2138 ) | ( n1868 & n5682 ) | ( n2138 & n5682 ) ;
  assign n13821 = n987 & ~n2339 ;
  assign n13820 = n7479 & n13492 ;
  assign n13822 = n13821 ^ n13820 ^ n7758 ;
  assign n13823 = n13415 ^ n7724 ^ n3968 ;
  assign n13824 = n3739 ^ n2753 ^ 1'b0 ;
  assign n13825 = n2117 & ~n13824 ;
  assign n13826 = ( n12992 & n13038 ) | ( n12992 & ~n13825 ) | ( n13038 & ~n13825 ) ;
  assign n13827 = ( ~n1114 & n2065 ) | ( ~n1114 & n2637 ) | ( n2065 & n2637 ) ;
  assign n13828 = n13827 ^ n3150 ^ 1'b0 ;
  assign n13829 = n2544 | n13828 ;
  assign n13830 = ( n271 & ~n1002 ) | ( n271 & n9811 ) | ( ~n1002 & n9811 ) ;
  assign n13831 = n13830 ^ n7033 ^ 1'b0 ;
  assign n13832 = n8629 | n13831 ;
  assign n13835 = n6606 | n8953 ;
  assign n13836 = n4359 & ~n13835 ;
  assign n13833 = x74 & n5023 ;
  assign n13834 = n13833 ^ n8422 ^ 1'b0 ;
  assign n13837 = n13836 ^ n13834 ^ n4181 ;
  assign n13838 = ( ~n9861 & n13832 ) | ( ~n9861 & n13837 ) | ( n13832 & n13837 ) ;
  assign n13839 = n2861 ^ n589 ^ 1'b0 ;
  assign n13840 = ~n7536 & n13839 ;
  assign n13841 = ~n1730 & n2625 ;
  assign n13842 = ~n4282 & n13841 ;
  assign n13843 = ( n603 & n10670 ) | ( n603 & n13842 ) | ( n10670 & n13842 ) ;
  assign n13844 = n8591 ^ n1280 ^ n289 ;
  assign n13845 = ( ~n7880 & n12422 ) | ( ~n7880 & n13844 ) | ( n12422 & n13844 ) ;
  assign n13846 = ( n6455 & n6750 ) | ( n6455 & ~n13845 ) | ( n6750 & ~n13845 ) ;
  assign n13847 = n13846 ^ n8076 ^ n1515 ;
  assign n13848 = n13847 ^ n4575 ^ 1'b0 ;
  assign n13849 = ~n13843 & n13848 ;
  assign n13850 = ( n4924 & n13840 ) | ( n4924 & n13849 ) | ( n13840 & n13849 ) ;
  assign n13851 = ( n6383 & n6754 ) | ( n6383 & n8578 ) | ( n6754 & n8578 ) ;
  assign n13852 = n6130 ^ n4541 ^ n2450 ;
  assign n13853 = n13852 ^ n2701 ^ 1'b0 ;
  assign n13854 = n13851 | n13853 ;
  assign n13855 = ( n4629 & n5808 ) | ( n4629 & n6205 ) | ( n5808 & n6205 ) ;
  assign n13856 = ( x125 & n6366 ) | ( x125 & n7925 ) | ( n6366 & n7925 ) ;
  assign n13857 = ~n13855 & n13856 ;
  assign n13858 = n13857 ^ n13547 ^ 1'b0 ;
  assign n13859 = n13858 ^ n11368 ^ x108 ;
  assign n13860 = n3616 ^ n2558 ^ 1'b0 ;
  assign n13861 = n12872 ^ n12795 ^ n1359 ;
  assign n13862 = ( n4967 & n13860 ) | ( n4967 & n13861 ) | ( n13860 & n13861 ) ;
  assign n13863 = ( n3066 & ~n7708 ) | ( n3066 & n9228 ) | ( ~n7708 & n9228 ) ;
  assign n13864 = n13863 ^ n7410 ^ 1'b0 ;
  assign n13865 = n7345 | n13864 ;
  assign n13866 = n9897 ^ n4271 ^ 1'b0 ;
  assign n13867 = ( n4195 & n9808 ) | ( n4195 & n13866 ) | ( n9808 & n13866 ) ;
  assign n13868 = n7628 ^ n5932 ^ n5368 ;
  assign n13872 = ( n2206 & n2447 ) | ( n2206 & ~n3014 ) | ( n2447 & ~n3014 ) ;
  assign n13869 = n7345 ^ n4088 ^ 1'b0 ;
  assign n13870 = n2686 | n13869 ;
  assign n13871 = n13870 ^ n4425 ^ n197 ;
  assign n13873 = n13872 ^ n13871 ^ n10359 ;
  assign n13874 = ( n5047 & n8407 ) | ( n5047 & n13873 ) | ( n8407 & n13873 ) ;
  assign n13875 = n10351 ^ n7855 ^ n3814 ;
  assign n13876 = n8514 ^ n4201 ^ n4099 ;
  assign n13877 = n5626 & ~n6978 ;
  assign n13878 = n13876 & n13877 ;
  assign n13879 = ( n4154 & ~n4647 ) | ( n4154 & n13878 ) | ( ~n4647 & n13878 ) ;
  assign n13880 = n11720 ^ n5161 ^ n3628 ;
  assign n13881 = ( n1042 & n2618 ) | ( n1042 & n10204 ) | ( n2618 & n10204 ) ;
  assign n13882 = n13881 ^ n6525 ^ n3352 ;
  assign n13883 = ( n767 & n1395 ) | ( n767 & ~n9995 ) | ( n1395 & ~n9995 ) ;
  assign n13884 = n13883 ^ n2567 ^ 1'b0 ;
  assign n13885 = n8036 & ~n13884 ;
  assign n13886 = n13882 | n13885 ;
  assign n13887 = ( ~n9997 & n13880 ) | ( ~n9997 & n13886 ) | ( n13880 & n13886 ) ;
  assign n13888 = ( n13875 & ~n13879 ) | ( n13875 & n13887 ) | ( ~n13879 & n13887 ) ;
  assign n13889 = n12974 ^ n7068 ^ n2017 ;
  assign n13890 = n2981 & ~n7862 ;
  assign n13891 = n13890 ^ n10992 ^ 1'b0 ;
  assign n13892 = n13891 ^ n13163 ^ n5377 ;
  assign n13894 = x22 & n8211 ;
  assign n13895 = n13894 ^ n3259 ^ 1'b0 ;
  assign n13893 = ( ~n7257 & n8163 ) | ( ~n7257 & n10093 ) | ( n8163 & n10093 ) ;
  assign n13896 = n13895 ^ n13893 ^ n12277 ;
  assign n13897 = n9268 ^ n7046 ^ n3102 ;
  assign n13899 = n2598 | n5504 ;
  assign n13900 = n3316 | n13899 ;
  assign n13898 = ~n1114 & n4626 ;
  assign n13901 = n13900 ^ n13898 ^ 1'b0 ;
  assign n13902 = ( n2507 & ~n10044 ) | ( n2507 & n13901 ) | ( ~n10044 & n13901 ) ;
  assign n13918 = n6354 ^ n5645 ^ n3199 ;
  assign n13914 = n874 ^ n684 ^ 1'b0 ;
  assign n13915 = n2604 | n13914 ;
  assign n13913 = ( ~n403 & n1422 ) | ( ~n403 & n5630 ) | ( n1422 & n5630 ) ;
  assign n13916 = n13915 ^ n13913 ^ n13692 ;
  assign n13917 = ( n5970 & ~n13677 ) | ( n5970 & n13916 ) | ( ~n13677 & n13916 ) ;
  assign n13919 = n13918 ^ n13917 ^ n832 ;
  assign n13920 = n13919 ^ n11555 ^ n3010 ;
  assign n13907 = ( ~n907 & n1155 ) | ( ~n907 & n2695 ) | ( n1155 & n2695 ) ;
  assign n13908 = ( n288 & ~n1620 ) | ( n288 & n1902 ) | ( ~n1620 & n1902 ) ;
  assign n13909 = ( n3207 & n4822 ) | ( n3207 & ~n13908 ) | ( n4822 & ~n13908 ) ;
  assign n13910 = ~n13907 & n13909 ;
  assign n13903 = ~n5290 & n11837 ;
  assign n13904 = n13903 ^ n5341 ^ 1'b0 ;
  assign n13905 = ( n2304 & n10431 ) | ( n2304 & n13904 ) | ( n10431 & n13904 ) ;
  assign n13906 = ( n4461 & ~n12963 ) | ( n4461 & n13905 ) | ( ~n12963 & n13905 ) ;
  assign n13911 = n13910 ^ n13906 ^ 1'b0 ;
  assign n13912 = n13644 & ~n13911 ;
  assign n13921 = n13920 ^ n13912 ^ 1'b0 ;
  assign n13922 = ( n881 & n13902 ) | ( n881 & n13921 ) | ( n13902 & n13921 ) ;
  assign n13923 = ( ~n961 & n2952 ) | ( ~n961 & n6493 ) | ( n2952 & n6493 ) ;
  assign n13924 = ( ~n2115 & n12125 ) | ( ~n2115 & n13923 ) | ( n12125 & n13923 ) ;
  assign n13925 = n10306 ^ n3571 ^ x108 ;
  assign n13926 = n13925 ^ n7477 ^ n4583 ;
  assign n13927 = ( n423 & ~n1083 ) | ( n423 & n1506 ) | ( ~n1083 & n1506 ) ;
  assign n13928 = ( n8886 & n12913 ) | ( n8886 & ~n13927 ) | ( n12913 & ~n13927 ) ;
  assign n13929 = n6072 | n13928 ;
  assign n13930 = n4183 | n13929 ;
  assign n13931 = ( n199 & ~n1853 ) | ( n199 & n13930 ) | ( ~n1853 & n13930 ) ;
  assign n13932 = n11521 ^ n5880 ^ 1'b0 ;
  assign n13933 = ( n1669 & n4370 ) | ( n1669 & ~n13932 ) | ( n4370 & ~n13932 ) ;
  assign n13934 = ( n5718 & ~n10356 ) | ( n5718 & n10616 ) | ( ~n10356 & n10616 ) ;
  assign n13935 = n9115 ^ n5597 ^ n4218 ;
  assign n13936 = n2758 ^ n941 ^ 1'b0 ;
  assign n13937 = n13936 ^ n3342 ^ n1538 ;
  assign n13938 = ( n9379 & n13935 ) | ( n9379 & n13937 ) | ( n13935 & n13937 ) ;
  assign n13939 = x85 & n175 ;
  assign n13940 = ~n3596 & n13939 ;
  assign n13941 = n13940 ^ n9315 ^ n5020 ;
  assign n13942 = ( n1369 & ~n5981 ) | ( n1369 & n13941 ) | ( ~n5981 & n13941 ) ;
  assign n13943 = ( n1440 & n3065 ) | ( n1440 & n5194 ) | ( n3065 & n5194 ) ;
  assign n13944 = n13943 ^ n10918 ^ n4843 ;
  assign n13945 = n3167 & ~n9365 ;
  assign n13946 = n8932 ^ n2704 ^ 1'b0 ;
  assign n13947 = n13946 ^ n12226 ^ n2086 ;
  assign n13948 = n13947 ^ n5781 ^ n2121 ;
  assign n13949 = n12840 ^ n6310 ^ n381 ;
  assign n13950 = ( n12511 & n13642 ) | ( n12511 & n13949 ) | ( n13642 & n13949 ) ;
  assign n13951 = n3535 ^ n2314 ^ 1'b0 ;
  assign n13952 = ( n8696 & n10080 ) | ( n8696 & ~n13951 ) | ( n10080 & ~n13951 ) ;
  assign n13953 = ( n2538 & ~n5510 ) | ( n2538 & n10264 ) | ( ~n5510 & n10264 ) ;
  assign n13954 = ( ~n3815 & n9504 ) | ( ~n3815 & n13953 ) | ( n9504 & n13953 ) ;
  assign n13955 = ( ~n11858 & n13649 ) | ( ~n11858 & n13954 ) | ( n13649 & n13954 ) ;
  assign n13956 = n3188 & n3558 ;
  assign n13957 = ~n3868 & n13956 ;
  assign n13958 = n9013 ^ n2563 ^ n175 ;
  assign n13959 = n13958 ^ n10616 ^ 1'b0 ;
  assign n13960 = n13959 ^ n13055 ^ 1'b0 ;
  assign n13961 = n2245 & n13960 ;
  assign n13962 = n6059 ^ n5309 ^ n2047 ;
  assign n13965 = ( n3711 & n3851 ) | ( n3711 & n4874 ) | ( n3851 & n4874 ) ;
  assign n13966 = ( n1365 & ~n4024 ) | ( n1365 & n13965 ) | ( ~n4024 & n13965 ) ;
  assign n13963 = n3499 ^ n1443 ^ 1'b0 ;
  assign n13964 = n1097 & n13963 ;
  assign n13967 = n13966 ^ n13964 ^ n13943 ;
  assign n13968 = ( n2304 & n2849 ) | ( n2304 & n13967 ) | ( n2849 & n13967 ) ;
  assign n13969 = n13290 ^ n7625 ^ n428 ;
  assign n13970 = n13969 ^ n9657 ^ n3976 ;
  assign n13971 = n10363 ^ n9265 ^ n2364 ;
  assign n13972 = n13971 ^ n7602 ^ n7162 ;
  assign n13973 = ( n4189 & ~n4978 ) | ( n4189 & n12604 ) | ( ~n4978 & n12604 ) ;
  assign n13974 = ( n1175 & ~n3786 ) | ( n1175 & n5121 ) | ( ~n3786 & n5121 ) ;
  assign n13975 = ( ~n1207 & n4827 ) | ( ~n1207 & n13974 ) | ( n4827 & n13974 ) ;
  assign n13976 = ( n964 & n1012 ) | ( n964 & n4435 ) | ( n1012 & n4435 ) ;
  assign n13977 = n11789 | n13976 ;
  assign n13978 = n8616 | n13977 ;
  assign n13979 = n13978 ^ n6811 ^ n2002 ;
  assign n13980 = ( n7944 & ~n13975 ) | ( n7944 & n13979 ) | ( ~n13975 & n13979 ) ;
  assign n13981 = n2534 & ~n3788 ;
  assign n13982 = n7516 ^ n1982 ^ 1'b0 ;
  assign n13983 = n7026 & n13982 ;
  assign n13984 = n13981 & n13983 ;
  assign n13986 = n4307 ^ n4121 ^ n2528 ;
  assign n13985 = n6310 ^ n5860 ^ n3264 ;
  assign n13987 = n13986 ^ n13985 ^ n2048 ;
  assign n13988 = n10505 ^ n9964 ^ n370 ;
  assign n13989 = n12505 ^ n5486 ^ n331 ;
  assign n13994 = ( n5158 & ~n6787 ) | ( n5158 & n9205 ) | ( ~n6787 & n9205 ) ;
  assign n13990 = ( n2045 & n4992 ) | ( n2045 & ~n5039 ) | ( n4992 & ~n5039 ) ;
  assign n13991 = n4217 | n13990 ;
  assign n13992 = n8515 & ~n13991 ;
  assign n13993 = n13992 ^ n9170 ^ n321 ;
  assign n13995 = n13994 ^ n13993 ^ n5259 ;
  assign n13996 = n7739 ^ n5638 ^ 1'b0 ;
  assign n13997 = ~n3314 & n8438 ;
  assign n13998 = n9857 ^ n5519 ^ n1295 ;
  assign n13999 = n13998 ^ n11879 ^ n5365 ;
  assign n14000 = ( n6625 & n12799 ) | ( n6625 & ~n13999 ) | ( n12799 & ~n13999 ) ;
  assign n14001 = ( n5139 & ~n8165 ) | ( n5139 & n14000 ) | ( ~n8165 & n14000 ) ;
  assign n14002 = n8224 ^ n838 ^ 1'b0 ;
  assign n14003 = n14002 ^ n1358 ^ 1'b0 ;
  assign n14004 = n14001 | n14003 ;
  assign n14005 = ( n13996 & ~n13997 ) | ( n13996 & n14004 ) | ( ~n13997 & n14004 ) ;
  assign n14006 = n8395 ^ n1736 ^ 1'b0 ;
  assign n14007 = ( n2149 & n7952 ) | ( n2149 & ~n14006 ) | ( n7952 & ~n14006 ) ;
  assign n14008 = ( n131 & ~n4034 ) | ( n131 & n4707 ) | ( ~n4034 & n4707 ) ;
  assign n14009 = ( ~n1072 & n9294 ) | ( ~n1072 & n14008 ) | ( n9294 & n14008 ) ;
  assign n14010 = n14009 ^ n1600 ^ 1'b0 ;
  assign n14011 = ( n3963 & n13901 ) | ( n3963 & n14010 ) | ( n13901 & n14010 ) ;
  assign n14012 = n14011 ^ n10700 ^ 1'b0 ;
  assign n14013 = n14007 & ~n14012 ;
  assign n14014 = ( n1201 & n4945 ) | ( n1201 & ~n14013 ) | ( n4945 & ~n14013 ) ;
  assign n14015 = n11253 ^ n5308 ^ n2701 ;
  assign n14016 = ( n5439 & ~n11837 ) | ( n5439 & n14015 ) | ( ~n11837 & n14015 ) ;
  assign n14017 = n5036 ^ n3878 ^ n3697 ;
  assign n14018 = n14017 ^ n6961 ^ n254 ;
  assign n14019 = n13821 ^ n12815 ^ n2229 ;
  assign n14020 = n14019 ^ n10481 ^ n4247 ;
  assign n14021 = n11620 & n12436 ;
  assign n14022 = n4393 & n14021 ;
  assign n14023 = ( n6471 & ~n13339 ) | ( n6471 & n14022 ) | ( ~n13339 & n14022 ) ;
  assign n14034 = n172 | n2322 ;
  assign n14035 = n524 | n14034 ;
  assign n14029 = ( n2554 & ~n2662 ) | ( n2554 & n13454 ) | ( ~n2662 & n13454 ) ;
  assign n14030 = ( x96 & ~n1122 ) | ( x96 & n3560 ) | ( ~n1122 & n3560 ) ;
  assign n14031 = n14030 ^ n10968 ^ n1223 ;
  assign n14032 = n14031 ^ n12708 ^ n5077 ;
  assign n14033 = ( n11237 & ~n14029 ) | ( n11237 & n14032 ) | ( ~n14029 & n14032 ) ;
  assign n14024 = n10134 ^ n2884 ^ 1'b0 ;
  assign n14025 = n261 & ~n14024 ;
  assign n14026 = n14025 ^ n7787 ^ n5514 ;
  assign n14027 = n10189 ^ n648 ^ 1'b0 ;
  assign n14028 = ( n5452 & ~n14026 ) | ( n5452 & n14027 ) | ( ~n14026 & n14027 ) ;
  assign n14036 = n14035 ^ n14033 ^ n14028 ;
  assign n14037 = ( n9292 & n12730 ) | ( n9292 & n12978 ) | ( n12730 & n12978 ) ;
  assign n14038 = n6428 ^ n5379 ^ x42 ;
  assign n14039 = n14038 ^ n3199 ^ n295 ;
  assign n14040 = n8613 ^ n7756 ^ n508 ;
  assign n14041 = ( n630 & ~n14039 ) | ( n630 & n14040 ) | ( ~n14039 & n14040 ) ;
  assign n14042 = ( ~n2568 & n10264 ) | ( ~n2568 & n14041 ) | ( n10264 & n14041 ) ;
  assign n14043 = ( n7012 & ~n10500 ) | ( n7012 & n14042 ) | ( ~n10500 & n14042 ) ;
  assign n14044 = n4195 | n12553 ;
  assign n14045 = n5722 ^ n555 ^ 1'b0 ;
  assign n14046 = n5008 ^ n2641 ^ 1'b0 ;
  assign n14047 = ( n10712 & ~n14045 ) | ( n10712 & n14046 ) | ( ~n14045 & n14046 ) ;
  assign n14048 = n719 | n14047 ;
  assign n14049 = ( n1199 & ~n6697 ) | ( n1199 & n14048 ) | ( ~n6697 & n14048 ) ;
  assign n14050 = n7793 & n14049 ;
  assign n14052 = n6590 ^ n4727 ^ n2531 ;
  assign n14053 = n14052 ^ n13655 ^ n1386 ;
  assign n14051 = ( ~n1247 & n4133 ) | ( ~n1247 & n14030 ) | ( n4133 & n14030 ) ;
  assign n14054 = n14053 ^ n14051 ^ n9797 ;
  assign n14055 = n12463 ^ n12094 ^ n2002 ;
  assign n14056 = ( n13177 & ~n14054 ) | ( n13177 & n14055 ) | ( ~n14054 & n14055 ) ;
  assign n14057 = n10402 ^ n3243 ^ n1068 ;
  assign n14058 = n10989 ^ n1443 ^ 1'b0 ;
  assign n14059 = n14058 ^ n14032 ^ n11445 ;
  assign n14060 = n6119 ^ n2109 ^ 1'b0 ;
  assign n14061 = n3277 & ~n14060 ;
  assign n14062 = n14061 ^ n5829 ^ n1645 ;
  assign n14063 = ( ~n169 & n2162 ) | ( ~n169 & n7079 ) | ( n2162 & n7079 ) ;
  assign n14064 = ( ~x122 & n14062 ) | ( ~x122 & n14063 ) | ( n14062 & n14063 ) ;
  assign n14065 = n5830 ^ n4107 ^ n1819 ;
  assign n14066 = n8848 ^ n7893 ^ n5486 ;
  assign n14067 = ( n12011 & n14065 ) | ( n12011 & n14066 ) | ( n14065 & n14066 ) ;
  assign n14068 = n11409 ^ n10466 ^ n4901 ;
  assign n14069 = ( n2670 & ~n5508 ) | ( n2670 & n11331 ) | ( ~n5508 & n11331 ) ;
  assign n14070 = ( n13163 & n14068 ) | ( n13163 & n14069 ) | ( n14068 & n14069 ) ;
  assign n14072 = n6587 ^ n6466 ^ n3969 ;
  assign n14071 = n1633 | n3977 ;
  assign n14073 = n14072 ^ n14071 ^ n14068 ;
  assign n14074 = ( ~n1729 & n7541 ) | ( ~n1729 & n14073 ) | ( n7541 & n14073 ) ;
  assign n14075 = n3369 ^ n736 ^ 1'b0 ;
  assign n14076 = n7302 ^ n373 ^ 1'b0 ;
  assign n14077 = ( n1279 & n14075 ) | ( n1279 & n14076 ) | ( n14075 & n14076 ) ;
  assign n14078 = ( n3648 & n9414 ) | ( n3648 & ~n14077 ) | ( n9414 & ~n14077 ) ;
  assign n14079 = ( n7827 & n10411 ) | ( n7827 & n14078 ) | ( n10411 & n14078 ) ;
  assign n14080 = n692 & n4910 ;
  assign n14081 = n3114 ^ n2879 ^ 1'b0 ;
  assign n14084 = ~n5738 & n12134 ;
  assign n14085 = ~n12134 & n14084 ;
  assign n14082 = ( ~n960 & n1036 ) | ( ~n960 & n3293 ) | ( n1036 & n3293 ) ;
  assign n14083 = ( n7895 & n9587 ) | ( n7895 & n14082 ) | ( n9587 & n14082 ) ;
  assign n14086 = n14085 ^ n14083 ^ n13283 ;
  assign n14087 = ( n1983 & ~n2048 ) | ( n1983 & n6020 ) | ( ~n2048 & n6020 ) ;
  assign n14088 = ( n1414 & ~n3692 ) | ( n1414 & n6094 ) | ( ~n3692 & n6094 ) ;
  assign n14089 = n14088 ^ n7029 ^ 1'b0 ;
  assign n14090 = n9316 ^ n5425 ^ n2073 ;
  assign n14091 = n11624 & ~n14090 ;
  assign n14092 = ( ~n4152 & n5656 ) | ( ~n4152 & n14091 ) | ( n5656 & n14091 ) ;
  assign n14093 = ( ~n14087 & n14089 ) | ( ~n14087 & n14092 ) | ( n14089 & n14092 ) ;
  assign n14094 = ( n2820 & ~n4436 ) | ( n2820 & n11404 ) | ( ~n4436 & n11404 ) ;
  assign n14095 = n9566 ^ n5187 ^ n4841 ;
  assign n14104 = n197 | n5836 ;
  assign n14103 = ( ~n3369 & n8094 ) | ( ~n3369 & n9858 ) | ( n8094 & n9858 ) ;
  assign n14099 = ~n285 & n342 ;
  assign n14100 = ~n10277 & n14099 ;
  assign n14097 = n12092 ^ n6407 ^ n3307 ;
  assign n14096 = ( n4912 & n5568 ) | ( n4912 & ~n6340 ) | ( n5568 & ~n6340 ) ;
  assign n14098 = n14097 ^ n14096 ^ n3810 ;
  assign n14101 = n14100 ^ n14098 ^ n474 ;
  assign n14102 = n14101 ^ n6249 ^ n3824 ;
  assign n14105 = n14104 ^ n14103 ^ n14102 ;
  assign n14106 = n8768 ^ n3639 ^ n1514 ;
  assign n14107 = n14106 ^ n13266 ^ n2386 ;
  assign n14108 = ( n3667 & n3861 ) | ( n3667 & ~n9914 ) | ( n3861 & ~n9914 ) ;
  assign n14109 = ( x40 & n3208 ) | ( x40 & ~n5050 ) | ( n3208 & ~n5050 ) ;
  assign n14111 = ( n2594 & n4750 ) | ( n2594 & ~n6002 ) | ( n4750 & ~n6002 ) ;
  assign n14110 = n8344 ^ n3320 ^ n2870 ;
  assign n14112 = n14111 ^ n14110 ^ n7833 ;
  assign n14113 = ( n8317 & ~n11264 ) | ( n8317 & n11775 ) | ( ~n11264 & n11775 ) ;
  assign n14114 = ( n3844 & n5424 ) | ( n3844 & ~n11474 ) | ( n5424 & ~n11474 ) ;
  assign n14115 = n7435 ^ n5357 ^ n3499 ;
  assign n14116 = ( n7026 & n11445 ) | ( n7026 & n14115 ) | ( n11445 & n14115 ) ;
  assign n14117 = ( n3289 & ~n8013 ) | ( n3289 & n14116 ) | ( ~n8013 & n14116 ) ;
  assign n14119 = ( n1217 & n2755 ) | ( n1217 & n6640 ) | ( n2755 & n6640 ) ;
  assign n14120 = n4409 | n14119 ;
  assign n14121 = n14120 ^ n6903 ^ 1'b0 ;
  assign n14118 = n6605 ^ n2924 ^ 1'b0 ;
  assign n14122 = n14121 ^ n14118 ^ n6119 ;
  assign n14124 = n167 & ~n10587 ;
  assign n14123 = ( ~n163 & n569 ) | ( ~n163 & n10421 ) | ( n569 & n10421 ) ;
  assign n14125 = n14124 ^ n14123 ^ 1'b0 ;
  assign n14126 = n12531 | n14125 ;
  assign n14127 = ( ~x43 & n14122 ) | ( ~x43 & n14126 ) | ( n14122 & n14126 ) ;
  assign n14128 = ( ~n7606 & n10431 ) | ( ~n7606 & n12147 ) | ( n10431 & n12147 ) ;
  assign n14130 = n10720 ^ n3670 ^ n475 ;
  assign n14129 = n5070 ^ n4624 ^ n3519 ;
  assign n14131 = n14130 ^ n14129 ^ n12428 ;
  assign n14132 = n3272 ^ n3128 ^ n728 ;
  assign n14133 = n3319 ^ n1477 ^ n1355 ;
  assign n14134 = ( ~n5122 & n14132 ) | ( ~n5122 & n14133 ) | ( n14132 & n14133 ) ;
  assign n14135 = ( n5209 & n14131 ) | ( n5209 & n14134 ) | ( n14131 & n14134 ) ;
  assign n14136 = ( n3510 & ~n3813 ) | ( n3510 & n8240 ) | ( ~n3813 & n8240 ) ;
  assign n14137 = n14136 ^ n12301 ^ n3897 ;
  assign n14138 = ( n3557 & n8877 ) | ( n3557 & ~n10077 ) | ( n8877 & ~n10077 ) ;
  assign n14139 = ( ~n683 & n14137 ) | ( ~n683 & n14138 ) | ( n14137 & n14138 ) ;
  assign n14144 = n9140 ^ n2389 ^ n209 ;
  assign n14140 = n977 & ~n1679 ;
  assign n14141 = ~n4940 & n14140 ;
  assign n14142 = n14141 ^ n5121 ^ n442 ;
  assign n14143 = n14142 ^ n8602 ^ n4839 ;
  assign n14145 = n14144 ^ n14143 ^ n9739 ;
  assign n14146 = n14145 ^ n13959 ^ n12025 ;
  assign n14147 = n5013 ^ n4123 ^ 1'b0 ;
  assign n14148 = ( n5483 & n10355 ) | ( n5483 & ~n13739 ) | ( n10355 & ~n13739 ) ;
  assign n14165 = n5566 & n7785 ;
  assign n14166 = n14165 ^ n3057 ^ 1'b0 ;
  assign n14162 = n8677 ^ n7438 ^ 1'b0 ;
  assign n14158 = n8651 ^ n4876 ^ n3407 ;
  assign n14159 = n8019 ^ n3497 ^ n1867 ;
  assign n14160 = ( n12965 & n14158 ) | ( n12965 & ~n14159 ) | ( n14158 & ~n14159 ) ;
  assign n14157 = n2179 ^ n962 ^ n864 ;
  assign n14161 = n14160 ^ n14157 ^ n5807 ;
  assign n14151 = ( ~n3566 & n3660 ) | ( ~n3566 & n6164 ) | ( n3660 & n6164 ) ;
  assign n14152 = ~n8228 & n12893 ;
  assign n14153 = ~n5197 & n14152 ;
  assign n14154 = ( n2388 & n4721 ) | ( n2388 & ~n14153 ) | ( n4721 & ~n14153 ) ;
  assign n14155 = ( n8480 & ~n14151 ) | ( n8480 & n14154 ) | ( ~n14151 & n14154 ) ;
  assign n14156 = n14155 ^ n13579 ^ n6193 ;
  assign n14163 = n14162 ^ n14161 ^ n14156 ;
  assign n14149 = n6804 & n10178 ;
  assign n14150 = n2804 | n14149 ;
  assign n14164 = n14163 ^ n14150 ^ 1'b0 ;
  assign n14167 = n14166 ^ n14164 ^ n3693 ;
  assign n14168 = ( n790 & ~n10244 ) | ( n790 & n14167 ) | ( ~n10244 & n14167 ) ;
  assign n14169 = n14168 ^ n4266 ^ n4231 ;
  assign n14170 = n11035 ^ n8366 ^ n5009 ;
  assign n14171 = n3322 ^ n1757 ^ 1'b0 ;
  assign n14172 = ( n8567 & n10937 ) | ( n8567 & ~n13554 ) | ( n10937 & ~n13554 ) ;
  assign n14173 = n13028 ^ n9080 ^ 1'b0 ;
  assign n14174 = n6893 ^ n6093 ^ n3163 ;
  assign n14175 = ( n586 & n4798 ) | ( n586 & ~n7416 ) | ( n4798 & ~n7416 ) ;
  assign n14176 = ( n10129 & n14174 ) | ( n10129 & n14175 ) | ( n14174 & n14175 ) ;
  assign n14177 = n3693 & n8996 ;
  assign n14178 = n14177 ^ n3926 ^ 1'b0 ;
  assign n14179 = n14178 ^ n4401 ^ n1437 ;
  assign n14180 = n9819 ^ n8420 ^ n3137 ;
  assign n14181 = n7654 ^ n5389 ^ n1049 ;
  assign n14187 = n1174 ^ n783 ^ n440 ;
  assign n14183 = ( n1125 & n1500 ) | ( n1125 & ~n10725 ) | ( n1500 & ~n10725 ) ;
  assign n14184 = ( n4511 & n12630 ) | ( n4511 & n14183 ) | ( n12630 & n14183 ) ;
  assign n14182 = n6144 & n7405 ;
  assign n14185 = n14184 ^ n14182 ^ 1'b0 ;
  assign n14186 = ( ~n6050 & n9740 ) | ( ~n6050 & n14185 ) | ( n9740 & n14185 ) ;
  assign n14188 = n14187 ^ n14186 ^ n4398 ;
  assign n14189 = n14071 ^ n8664 ^ n5875 ;
  assign n14190 = ( n563 & n2224 ) | ( n563 & ~n10749 ) | ( n2224 & ~n10749 ) ;
  assign n14191 = ( n2489 & n13195 ) | ( n2489 & n14190 ) | ( n13195 & n14190 ) ;
  assign n14193 = ( n1918 & ~n2475 ) | ( n1918 & n5901 ) | ( ~n2475 & n5901 ) ;
  assign n14194 = n14193 ^ n3631 ^ n1080 ;
  assign n14192 = ( ~n1985 & n5923 ) | ( ~n1985 & n10088 ) | ( n5923 & n10088 ) ;
  assign n14195 = n14194 ^ n14192 ^ n1994 ;
  assign n14196 = n14191 & ~n14195 ;
  assign n14197 = n5351 & n14196 ;
  assign n14198 = n8936 ^ n1572 ^ 1'b0 ;
  assign n14199 = n14198 ^ n6037 ^ n4414 ;
  assign n14200 = n13996 ^ n8913 ^ n3905 ;
  assign n14201 = ( n4243 & n12561 ) | ( n4243 & n14200 ) | ( n12561 & n14200 ) ;
  assign n14202 = ( n3517 & n6753 ) | ( n3517 & n14201 ) | ( n6753 & n14201 ) ;
  assign n14203 = ( n2825 & ~n4121 ) | ( n2825 & n7048 ) | ( ~n4121 & n7048 ) ;
  assign n14204 = ( ~x68 & n3580 ) | ( ~x68 & n4349 ) | ( n3580 & n4349 ) ;
  assign n14208 = n11537 ^ n8978 ^ 1'b0 ;
  assign n14206 = ( n2623 & ~n4063 ) | ( n2623 & n6107 ) | ( ~n4063 & n6107 ) ;
  assign n14205 = ( n1685 & ~n3653 ) | ( n1685 & n7382 ) | ( ~n3653 & n7382 ) ;
  assign n14207 = n14206 ^ n14205 ^ n9476 ;
  assign n14209 = n14208 ^ n14207 ^ n5931 ;
  assign n14210 = n14204 & n14209 ;
  assign n14211 = ( n2255 & n14203 ) | ( n2255 & ~n14210 ) | ( n14203 & ~n14210 ) ;
  assign n14212 = n5224 ^ n1927 ^ n547 ;
  assign n14213 = n14212 ^ n10124 ^ n5605 ;
  assign n14214 = n14213 ^ n6663 ^ n2917 ;
  assign n14215 = n10066 ^ n9087 ^ n2127 ;
  assign n14216 = n7072 ^ n4357 ^ n1708 ;
  assign n14217 = ( n9341 & n10003 ) | ( n9341 & n14216 ) | ( n10003 & n14216 ) ;
  assign n14218 = ( n8984 & n14215 ) | ( n8984 & ~n14217 ) | ( n14215 & ~n14217 ) ;
  assign n14219 = n11925 ^ n10924 ^ n1865 ;
  assign n14220 = n427 & ~n14219 ;
  assign n14221 = ~n7140 & n14220 ;
  assign n14222 = ( n6430 & n8496 ) | ( n6430 & ~n11576 ) | ( n8496 & ~n11576 ) ;
  assign n14223 = n3683 & n4051 ;
  assign n14224 = n14222 & n14223 ;
  assign n14225 = ( n2712 & ~n11663 ) | ( n2712 & n14224 ) | ( ~n11663 & n14224 ) ;
  assign n14226 = ( n2703 & n8134 ) | ( n2703 & ~n11501 ) | ( n8134 & ~n11501 ) ;
  assign n14227 = ( n2334 & ~n3297 ) | ( n2334 & n14226 ) | ( ~n3297 & n14226 ) ;
  assign n14228 = n11641 & ~n14227 ;
  assign n14229 = n14228 ^ n5087 ^ 1'b0 ;
  assign n14230 = ( n3570 & n14225 ) | ( n3570 & ~n14229 ) | ( n14225 & ~n14229 ) ;
  assign n14238 = n12029 ^ n2108 ^ n1974 ;
  assign n14231 = ( n428 & ~n11242 ) | ( n428 & n12904 ) | ( ~n11242 & n12904 ) ;
  assign n14232 = ( x17 & n2329 ) | ( x17 & ~n12739 ) | ( n2329 & ~n12739 ) ;
  assign n14233 = n14232 ^ n5087 ^ n4864 ;
  assign n14234 = n1659 & ~n2683 ;
  assign n14235 = n14234 ^ n4956 ^ 1'b0 ;
  assign n14236 = ( n13532 & n14233 ) | ( n13532 & ~n14235 ) | ( n14233 & ~n14235 ) ;
  assign n14237 = ( ~n13863 & n14231 ) | ( ~n13863 & n14236 ) | ( n14231 & n14236 ) ;
  assign n14239 = n14238 ^ n14237 ^ n5761 ;
  assign n14240 = n3704 ^ n3183 ^ n130 ;
  assign n14241 = n14240 ^ n5820 ^ n3525 ;
  assign n14242 = n14241 ^ n10561 ^ n5627 ;
  assign n14243 = n13394 ^ n1411 ^ n406 ;
  assign n14244 = ( ~n7157 & n10276 ) | ( ~n7157 & n14243 ) | ( n10276 & n14243 ) ;
  assign n14245 = n10794 ^ n9354 ^ 1'b0 ;
  assign n14247 = ~n1615 & n2306 ;
  assign n14248 = ~n7136 & n14247 ;
  assign n14246 = ~n4190 & n9951 ;
  assign n14249 = n14248 ^ n14246 ^ n9552 ;
  assign n14250 = n14249 ^ n3695 ^ 1'b0 ;
  assign n14251 = x14 & ~n14250 ;
  assign n14252 = n1894 & n12154 ;
  assign n14253 = n14252 ^ n310 ^ 1'b0 ;
  assign n14254 = ( n1151 & n13683 ) | ( n1151 & n14253 ) | ( n13683 & n14253 ) ;
  assign n14255 = ~n1568 & n4159 ;
  assign n14256 = ~n8754 & n14255 ;
  assign n14257 = ( n697 & ~n10686 ) | ( n697 & n14256 ) | ( ~n10686 & n14256 ) ;
  assign n14259 = n10863 ^ n6727 ^ n2262 ;
  assign n14258 = n10278 ^ n3084 ^ n2353 ;
  assign n14260 = n14259 ^ n14258 ^ n905 ;
  assign n14261 = ~n5649 & n14078 ;
  assign n14262 = n14261 ^ n1964 ^ 1'b0 ;
  assign n14263 = n10848 ^ n5121 ^ 1'b0 ;
  assign n14264 = n7539 & ~n14263 ;
  assign n14265 = n1004 & n14264 ;
  assign n14266 = ( ~n5823 & n6837 ) | ( ~n5823 & n10413 ) | ( n6837 & n10413 ) ;
  assign n14267 = n14266 ^ n6351 ^ n1151 ;
  assign n14268 = ( x121 & ~n9688 ) | ( x121 & n14267 ) | ( ~n9688 & n14267 ) ;
  assign n14270 = ( n5143 & n5844 ) | ( n5143 & ~n11690 ) | ( n5844 & ~n11690 ) ;
  assign n14269 = ( n2946 & n9513 ) | ( n2946 & n14143 ) | ( n9513 & n14143 ) ;
  assign n14271 = n14270 ^ n14269 ^ n9512 ;
  assign n14272 = n3300 & ~n6407 ;
  assign n14273 = ( ~n6307 & n7818 ) | ( ~n6307 & n14272 ) | ( n7818 & n14272 ) ;
  assign n14274 = ~n6440 & n10071 ;
  assign n14275 = n11694 ^ n4123 ^ n1853 ;
  assign n14276 = ( ~n4776 & n13825 ) | ( ~n4776 & n14275 ) | ( n13825 & n14275 ) ;
  assign n14277 = ( n14273 & n14274 ) | ( n14273 & n14276 ) | ( n14274 & n14276 ) ;
  assign n14278 = ( ~n4816 & n7930 ) | ( ~n4816 & n13927 ) | ( n7930 & n13927 ) ;
  assign n14279 = ( n1359 & ~n4116 ) | ( n1359 & n14278 ) | ( ~n4116 & n14278 ) ;
  assign n14280 = n10861 ^ n129 ^ 1'b0 ;
  assign n14281 = n14280 ^ n333 ^ x17 ;
  assign n14284 = n9385 ^ n8184 ^ n735 ;
  assign n14286 = n5285 ^ n3136 ^ n3067 ;
  assign n14287 = ( ~n2838 & n6935 ) | ( ~n2838 & n14286 ) | ( n6935 & n14286 ) ;
  assign n14288 = ( n3383 & n7209 ) | ( n3383 & ~n14287 ) | ( n7209 & ~n14287 ) ;
  assign n14285 = ( ~n1979 & n3254 ) | ( ~n1979 & n12696 ) | ( n3254 & n12696 ) ;
  assign n14289 = n14288 ^ n14285 ^ n3325 ;
  assign n14290 = n8407 ^ n997 ^ x55 ;
  assign n14291 = n14290 ^ n10873 ^ 1'b0 ;
  assign n14292 = ~n9334 & n14291 ;
  assign n14293 = ( n12700 & ~n14289 ) | ( n12700 & n14292 ) | ( ~n14289 & n14292 ) ;
  assign n14294 = ~n14284 & n14293 ;
  assign n14295 = n14294 ^ n13840 ^ 1'b0 ;
  assign n14282 = n3807 ^ n1165 ^ 1'b0 ;
  assign n14283 = ~n6213 & n14282 ;
  assign n14296 = n14295 ^ n14283 ^ n5933 ;
  assign n14298 = n2412 ^ n1510 ^ 1'b0 ;
  assign n14299 = n1302 | n14298 ;
  assign n14297 = n6372 ^ n3978 ^ n2812 ;
  assign n14300 = n14299 ^ n14297 ^ n8073 ;
  assign n14304 = ( ~n1421 & n4319 ) | ( ~n1421 & n7442 ) | ( n4319 & n7442 ) ;
  assign n14301 = ( ~n1928 & n7281 ) | ( ~n1928 & n11893 ) | ( n7281 & n11893 ) ;
  assign n14302 = n14301 ^ n2973 ^ x69 ;
  assign n14303 = n14302 ^ n10278 ^ n7170 ;
  assign n14305 = n14304 ^ n14303 ^ n5381 ;
  assign n14306 = ( n4688 & ~n6761 ) | ( n4688 & n9371 ) | ( ~n6761 & n9371 ) ;
  assign n14309 = ( n3865 & ~n6330 ) | ( n3865 & n13655 ) | ( ~n6330 & n13655 ) ;
  assign n14307 = ~n2453 & n6752 ;
  assign n14308 = ( n1110 & n13604 ) | ( n1110 & n14307 ) | ( n13604 & n14307 ) ;
  assign n14310 = n14309 ^ n14308 ^ n1680 ;
  assign n14314 = n9775 ^ n2705 ^ n454 ;
  assign n14311 = n2492 ^ n2330 ^ 1'b0 ;
  assign n14312 = n10224 | n14311 ;
  assign n14313 = ( n8382 & ~n9370 ) | ( n8382 & n14312 ) | ( ~n9370 & n14312 ) ;
  assign n14315 = n14314 ^ n14313 ^ n4279 ;
  assign n14316 = ( n14306 & n14310 ) | ( n14306 & ~n14315 ) | ( n14310 & ~n14315 ) ;
  assign n14317 = ( n1946 & ~n6818 ) | ( n1946 & n12942 ) | ( ~n6818 & n12942 ) ;
  assign n14318 = n8566 ^ n5551 ^ n4149 ;
  assign n14319 = n10586 ^ n9136 ^ n1585 ;
  assign n14320 = n14319 ^ n8330 ^ n3437 ;
  assign n14321 = n14320 ^ n6274 ^ 1'b0 ;
  assign n14322 = ~n14318 & n14321 ;
  assign n14323 = n3170 ^ n2786 ^ n474 ;
  assign n14324 = n14323 ^ n12893 ^ n6076 ;
  assign n14325 = n10470 & n14324 ;
  assign n14326 = ( ~n1289 & n3215 ) | ( ~n1289 & n3320 ) | ( n3215 & n3320 ) ;
  assign n14327 = ~n508 & n14326 ;
  assign n14328 = n14327 ^ n6020 ^ 1'b0 ;
  assign n14329 = n10117 ^ n9784 ^ n1615 ;
  assign n14330 = ( n2068 & n13069 ) | ( n2068 & ~n14329 ) | ( n13069 & ~n14329 ) ;
  assign n14331 = ( n2850 & n3318 ) | ( n2850 & ~n3654 ) | ( n3318 & ~n3654 ) ;
  assign n14332 = n14331 ^ n2054 ^ 1'b0 ;
  assign n14333 = ( ~n1525 & n4181 ) | ( ~n1525 & n7514 ) | ( n4181 & n7514 ) ;
  assign n14334 = n14333 ^ n11014 ^ n4362 ;
  assign n14335 = ( n2248 & ~n7137 ) | ( n2248 & n14334 ) | ( ~n7137 & n14334 ) ;
  assign n14336 = ( ~n6224 & n7401 ) | ( ~n6224 & n14335 ) | ( n7401 & n14335 ) ;
  assign n14339 = n6998 ^ n3667 ^ 1'b0 ;
  assign n14337 = n3498 ^ n1171 ^ n708 ;
  assign n14338 = n2004 & n14337 ;
  assign n14340 = n14339 ^ n14338 ^ n3072 ;
  assign n14341 = n14340 ^ n7817 ^ n889 ;
  assign n14342 = ( n1255 & n3997 ) | ( n1255 & n10029 ) | ( n3997 & n10029 ) ;
  assign n14343 = ( ~n4457 & n13324 ) | ( ~n4457 & n14342 ) | ( n13324 & n14342 ) ;
  assign n14344 = n5125 ^ n5047 ^ x27 ;
  assign n14345 = ( n1352 & n10245 ) | ( n1352 & n14344 ) | ( n10245 & n14344 ) ;
  assign n14346 = n140 & n11155 ;
  assign n14347 = ~n3741 & n14346 ;
  assign n14350 = ( ~n3437 & n6623 ) | ( ~n3437 & n8711 ) | ( n6623 & n8711 ) ;
  assign n14349 = n4210 ^ n2320 ^ n1523 ;
  assign n14348 = n12433 ^ n4844 ^ n962 ;
  assign n14351 = n14350 ^ n14349 ^ n14348 ;
  assign n14352 = ( n1591 & ~n14347 ) | ( n1591 & n14351 ) | ( ~n14347 & n14351 ) ;
  assign n14353 = n10943 | n13353 ;
  assign n14354 = n2683 & ~n14353 ;
  assign n14355 = n3673 ^ n1580 ^ 1'b0 ;
  assign n14356 = n1077 | n14355 ;
  assign n14357 = ( x70 & n549 ) | ( x70 & ~n1379 ) | ( n549 & ~n1379 ) ;
  assign n14358 = ( ~n7799 & n13151 ) | ( ~n7799 & n14357 ) | ( n13151 & n14357 ) ;
  assign n14359 = n14356 | n14358 ;
  assign n14360 = n14359 ^ n13378 ^ 1'b0 ;
  assign n14361 = n11319 ^ n8189 ^ n2330 ;
  assign n14362 = ( ~n3995 & n4830 ) | ( ~n3995 & n14361 ) | ( n4830 & n14361 ) ;
  assign n14363 = ( ~n567 & n8284 ) | ( ~n567 & n14362 ) | ( n8284 & n14362 ) ;
  assign n14364 = n10408 ^ n2714 ^ n495 ;
  assign n14365 = ( ~n8990 & n14363 ) | ( ~n8990 & n14364 ) | ( n14363 & n14364 ) ;
  assign n14366 = n1995 | n9650 ;
  assign n14367 = ( n3256 & n13836 ) | ( n3256 & ~n14366 ) | ( n13836 & ~n14366 ) ;
  assign n14368 = n14367 ^ n7322 ^ n2858 ;
  assign n14369 = ( n848 & ~n9184 ) | ( n848 & n14368 ) | ( ~n9184 & n14368 ) ;
  assign n14370 = ( n747 & n14365 ) | ( n747 & ~n14369 ) | ( n14365 & ~n14369 ) ;
  assign n14371 = n9780 ^ n6857 ^ n3875 ;
  assign n14372 = ( ~n6283 & n12184 ) | ( ~n6283 & n14371 ) | ( n12184 & n14371 ) ;
  assign n14373 = ( n1634 & ~n9520 ) | ( n1634 & n13700 ) | ( ~n9520 & n13700 ) ;
  assign n14374 = n6568 ^ n6468 ^ n577 ;
  assign n14375 = n14374 ^ n7923 ^ n2480 ;
  assign n14376 = n2407 & n9395 ;
  assign n14377 = n14376 ^ n5872 ^ 1'b0 ;
  assign n14378 = ( n1406 & n2877 ) | ( n1406 & ~n4304 ) | ( n2877 & ~n4304 ) ;
  assign n14380 = n9178 ^ n6947 ^ n5578 ;
  assign n14379 = ( n1616 & ~n3980 ) | ( n1616 & n4196 ) | ( ~n3980 & n4196 ) ;
  assign n14381 = n14380 ^ n14379 ^ n8447 ;
  assign n14382 = ( n14377 & n14378 ) | ( n14377 & n14381 ) | ( n14378 & n14381 ) ;
  assign n14383 = ( n1749 & n5084 ) | ( n1749 & n5259 ) | ( n5084 & n5259 ) ;
  assign n14384 = ( n5847 & n6752 ) | ( n5847 & n6772 ) | ( n6752 & n6772 ) ;
  assign n14385 = n14384 ^ n7412 ^ 1'b0 ;
  assign n14386 = ( ~n8582 & n14383 ) | ( ~n8582 & n14385 ) | ( n14383 & n14385 ) ;
  assign n14387 = n3723 & ~n3986 ;
  assign n14388 = n14387 ^ n4679 ^ 1'b0 ;
  assign n14389 = ( n3615 & n9211 ) | ( n3615 & n14388 ) | ( n9211 & n14388 ) ;
  assign n14390 = n14389 ^ n7609 ^ x117 ;
  assign n14391 = n14205 ^ n9602 ^ n1175 ;
  assign n14392 = n14391 ^ n254 ^ 1'b0 ;
  assign n14393 = n13663 | n14392 ;
  assign n14394 = n14390 | n14393 ;
  assign n14395 = ( n5613 & n8848 ) | ( n5613 & ~n9723 ) | ( n8848 & ~n9723 ) ;
  assign n14399 = n7766 ^ n7001 ^ n421 ;
  assign n14400 = ( n5026 & n13657 ) | ( n5026 & ~n14399 ) | ( n13657 & ~n14399 ) ;
  assign n14396 = ( n1666 & n2166 ) | ( n1666 & ~n8783 ) | ( n2166 & ~n8783 ) ;
  assign n14397 = n14396 ^ n10234 ^ n3453 ;
  assign n14398 = n14397 ^ n7265 ^ n5237 ;
  assign n14401 = n14400 ^ n14398 ^ n7921 ;
  assign n14402 = ( ~n11683 & n14395 ) | ( ~n11683 & n14401 ) | ( n14395 & n14401 ) ;
  assign n14406 = n8850 ^ n8642 ^ n3736 ;
  assign n14404 = n7356 ^ n5890 ^ n3889 ;
  assign n14405 = n14404 ^ n14338 ^ n8865 ;
  assign n14403 = n12082 ^ n4761 ^ n2671 ;
  assign n14407 = n14406 ^ n14405 ^ n14403 ;
  assign n14408 = ( n8476 & ~n9802 ) | ( n8476 & n14407 ) | ( ~n9802 & n14407 ) ;
  assign n14410 = n10991 ^ n7944 ^ 1'b0 ;
  assign n14409 = n4234 & ~n7118 ;
  assign n14411 = n14410 ^ n14409 ^ 1'b0 ;
  assign n14412 = n7818 ^ n5235 ^ n3970 ;
  assign n14413 = n7362 ^ n5416 ^ n1353 ;
  assign n14414 = n14412 | n14413 ;
  assign n14415 = ( n445 & n14166 ) | ( n445 & n14414 ) | ( n14166 & n14414 ) ;
  assign n14418 = ( n271 & n2771 ) | ( n271 & n7818 ) | ( n2771 & n7818 ) ;
  assign n14416 = n8803 ^ n1860 ^ n460 ;
  assign n14417 = ( n6236 & ~n8138 ) | ( n6236 & n14416 ) | ( ~n8138 & n14416 ) ;
  assign n14419 = n14418 ^ n14417 ^ n1203 ;
  assign n14420 = n14419 ^ n12112 ^ n636 ;
  assign n14421 = n5454 ^ n2569 ^ n2371 ;
  assign n14422 = ( n4210 & n7284 ) | ( n4210 & n14421 ) | ( n7284 & n14421 ) ;
  assign n14423 = ( ~n2492 & n3567 ) | ( ~n2492 & n14422 ) | ( n3567 & n14422 ) ;
  assign n14424 = n2664 ^ n1169 ^ n705 ;
  assign n14425 = ( n2107 & n2928 ) | ( n2107 & n14424 ) | ( n2928 & n14424 ) ;
  assign n14426 = ( n5124 & ~n6555 ) | ( n5124 & n7079 ) | ( ~n6555 & n7079 ) ;
  assign n14427 = n14426 ^ n14224 ^ n3240 ;
  assign n14428 = n9866 ^ n565 ^ 1'b0 ;
  assign n14429 = n2088 & ~n14428 ;
  assign n14436 = n12302 ^ n6173 ^ n6040 ;
  assign n14433 = n7822 ^ n1055 ^ 1'b0 ;
  assign n14431 = ( n7751 & n11830 ) | ( n7751 & ~n13261 ) | ( n11830 & ~n13261 ) ;
  assign n14430 = n2758 | n5139 ;
  assign n14432 = n14431 ^ n14430 ^ 1'b0 ;
  assign n14434 = n14433 ^ n14432 ^ n11004 ;
  assign n14435 = n14434 ^ n12505 ^ n9226 ;
  assign n14437 = n14436 ^ n14435 ^ n6688 ;
  assign n14438 = ( n1737 & n4657 ) | ( n1737 & ~n9725 ) | ( n4657 & ~n9725 ) ;
  assign n14439 = n10193 ^ n6435 ^ n2150 ;
  assign n14440 = ( n5412 & n7172 ) | ( n5412 & ~n11442 ) | ( n7172 & ~n11442 ) ;
  assign n14441 = n14099 ^ n1461 ^ 1'b0 ;
  assign n14442 = ~n14440 & n14441 ;
  assign n14443 = n14442 ^ n9352 ^ n1532 ;
  assign n14444 = n14443 ^ n11071 ^ 1'b0 ;
  assign n14445 = n14439 | n14444 ;
  assign n14446 = ( ~n1543 & n4256 ) | ( ~n1543 & n9143 ) | ( n4256 & n9143 ) ;
  assign n14447 = ( n7121 & ~n14270 ) | ( n7121 & n14446 ) | ( ~n14270 & n14446 ) ;
  assign n14448 = ( n2889 & ~n3617 ) | ( n2889 & n4034 ) | ( ~n3617 & n4034 ) ;
  assign n14449 = ( n315 & n1303 ) | ( n315 & ~n9001 ) | ( n1303 & ~n9001 ) ;
  assign n14450 = ( ~n3201 & n14448 ) | ( ~n3201 & n14449 ) | ( n14448 & n14449 ) ;
  assign n14451 = n14450 ^ n10919 ^ n541 ;
  assign n14452 = ( n2763 & ~n3072 ) | ( n2763 & n10697 ) | ( ~n3072 & n10697 ) ;
  assign n14453 = n5050 & n9872 ;
  assign n14454 = ~n14452 & n14453 ;
  assign n14455 = n2457 ^ n1967 ^ n1765 ;
  assign n14456 = ( n1349 & n8686 ) | ( n1349 & ~n12429 ) | ( n8686 & ~n12429 ) ;
  assign n14457 = ( n8172 & ~n9753 ) | ( n8172 & n14456 ) | ( ~n9753 & n14456 ) ;
  assign n14458 = ( n3104 & n9877 ) | ( n3104 & n14457 ) | ( n9877 & n14457 ) ;
  assign n14459 = ( x68 & n14455 ) | ( x68 & ~n14458 ) | ( n14455 & ~n14458 ) ;
  assign n14460 = n8196 ^ n3873 ^ 1'b0 ;
  assign n14461 = ( n3227 & n9786 ) | ( n3227 & n14460 ) | ( n9786 & n14460 ) ;
  assign n14462 = ( n2410 & n2604 ) | ( n2410 & ~n11121 ) | ( n2604 & ~n11121 ) ;
  assign n14463 = n14462 ^ n10681 ^ x118 ;
  assign n14464 = ( ~n2466 & n3134 ) | ( ~n2466 & n4282 ) | ( n3134 & n4282 ) ;
  assign n14465 = n14464 ^ n9805 ^ 1'b0 ;
  assign n14468 = n4725 & n9321 ;
  assign n14466 = n7198 & ~n7796 ;
  assign n14467 = ~n11790 & n14466 ;
  assign n14469 = n14468 ^ n14467 ^ n3415 ;
  assign n14470 = n3709 ^ n3631 ^ n1339 ;
  assign n14471 = ( n4096 & ~n14469 ) | ( n4096 & n14470 ) | ( ~n14469 & n14470 ) ;
  assign n14472 = n1747 ^ n537 ^ n331 ;
  assign n14473 = n6111 ^ n5222 ^ 1'b0 ;
  assign n14475 = n3888 ^ n3035 ^ n2501 ;
  assign n14474 = ~n5667 & n11116 ;
  assign n14476 = n14475 ^ n14474 ^ 1'b0 ;
  assign n14477 = n14476 ^ n5431 ^ 1'b0 ;
  assign n14478 = ( n14472 & n14473 ) | ( n14472 & n14477 ) | ( n14473 & n14477 ) ;
  assign n14479 = n14478 ^ n12437 ^ n2798 ;
  assign n14480 = ( n995 & n3275 ) | ( n995 & ~n3864 ) | ( n3275 & ~n3864 ) ;
  assign n14481 = n14480 ^ n3857 ^ n1738 ;
  assign n14482 = ( ~n1121 & n1671 ) | ( ~n1121 & n7498 ) | ( n1671 & n7498 ) ;
  assign n14483 = n6635 & n14482 ;
  assign n14484 = n9607 ^ n7449 ^ n4466 ;
  assign n14485 = ( ~n1044 & n11416 ) | ( ~n1044 & n14484 ) | ( n11416 & n14484 ) ;
  assign n14486 = ( ~n3325 & n5696 ) | ( ~n3325 & n8687 ) | ( n5696 & n8687 ) ;
  assign n14487 = n14486 ^ n7077 ^ n3378 ;
  assign n14488 = n7346 ^ n1520 ^ n344 ;
  assign n14489 = n7511 ^ n6042 ^ n633 ;
  assign n14490 = ( n4018 & ~n4040 ) | ( n4018 & n14489 ) | ( ~n4040 & n14489 ) ;
  assign n14491 = n8958 ^ n4916 ^ n4078 ;
  assign n14492 = n2894 ^ n1257 ^ 1'b0 ;
  assign n14493 = n350 & n14492 ;
  assign n14494 = ( n161 & n14491 ) | ( n161 & n14493 ) | ( n14491 & n14493 ) ;
  assign n14495 = ( n14488 & n14490 ) | ( n14488 & n14494 ) | ( n14490 & n14494 ) ;
  assign n14496 = ( n4344 & n5802 ) | ( n4344 & n9883 ) | ( n5802 & n9883 ) ;
  assign n14497 = ( n9321 & ~n10870 ) | ( n9321 & n12365 ) | ( ~n10870 & n12365 ) ;
  assign n14498 = ~n10836 & n13783 ;
  assign n14499 = n14498 ^ n7369 ^ 1'b0 ;
  assign n14500 = n14499 ^ n13625 ^ n12395 ;
  assign n14501 = n13660 ^ n4044 ^ n1321 ;
  assign n14502 = n8212 ^ n6406 ^ n5051 ;
  assign n14503 = ( ~n2238 & n4846 ) | ( ~n2238 & n14502 ) | ( n4846 & n14502 ) ;
  assign n14504 = ~n5922 & n14503 ;
  assign n14505 = n14145 ^ n8011 ^ n5160 ;
  assign n14506 = ( n4937 & n8526 ) | ( n4937 & n10461 ) | ( n8526 & n10461 ) ;
  assign n14507 = n14505 | n14506 ;
  assign n14508 = n14507 ^ n8745 ^ 1'b0 ;
  assign n14509 = n13432 ^ n8410 ^ n5515 ;
  assign n14510 = n14509 ^ n10400 ^ n7216 ;
  assign n14511 = n3507 ^ n1379 ^ 1'b0 ;
  assign n14512 = ~n7028 & n14511 ;
  assign n14513 = ( n4104 & n7440 ) | ( n4104 & n14512 ) | ( n7440 & n14512 ) ;
  assign n14514 = ( n3969 & n8691 ) | ( n3969 & n14513 ) | ( n8691 & n14513 ) ;
  assign n14515 = n14514 ^ n9821 ^ n8475 ;
  assign n14516 = n12425 ^ n10083 ^ n1193 ;
  assign n14517 = n14516 ^ n6103 ^ n996 ;
  assign n14522 = ( n2913 & n3431 ) | ( n2913 & ~n5702 ) | ( n3431 & ~n5702 ) ;
  assign n14523 = ( ~n4555 & n6160 ) | ( ~n4555 & n14522 ) | ( n6160 & n14522 ) ;
  assign n14518 = n1421 | n12133 ;
  assign n14519 = n8540 | n14518 ;
  assign n14520 = n7515 & ~n10782 ;
  assign n14521 = ~n14519 & n14520 ;
  assign n14524 = n14523 ^ n14521 ^ n10843 ;
  assign n14526 = ( ~n2032 & n6036 ) | ( ~n2032 & n10921 ) | ( n6036 & n10921 ) ;
  assign n14527 = n14526 ^ n3338 ^ n495 ;
  assign n14525 = n3591 | n6139 ;
  assign n14528 = n14527 ^ n14525 ^ 1'b0 ;
  assign n14529 = ~n1698 & n14528 ;
  assign n14530 = ~n5634 & n10057 ;
  assign n14531 = n14530 ^ n9022 ^ 1'b0 ;
  assign n14532 = ( n568 & n4604 ) | ( n568 & ~n14531 ) | ( n4604 & ~n14531 ) ;
  assign n14533 = ( n2321 & ~n4191 ) | ( n2321 & n13958 ) | ( ~n4191 & n13958 ) ;
  assign n14534 = ( ~n6853 & n11235 ) | ( ~n6853 & n14533 ) | ( n11235 & n14533 ) ;
  assign n14535 = ( n14142 & ~n14532 ) | ( n14142 & n14534 ) | ( ~n14532 & n14534 ) ;
  assign n14536 = n14535 ^ n13208 ^ n2180 ;
  assign n14537 = n3855 | n10897 ;
  assign n14538 = n9444 & ~n14537 ;
  assign n14539 = n8445 ^ n3143 ^ n2633 ;
  assign n14540 = ( x17 & ~n1618 ) | ( x17 & n14539 ) | ( ~n1618 & n14539 ) ;
  assign n14541 = ( n4916 & n7761 ) | ( n4916 & n13337 ) | ( n7761 & n13337 ) ;
  assign n14546 = n11529 ^ n8902 ^ n8026 ;
  assign n14547 = ( n2194 & n11735 ) | ( n2194 & ~n14546 ) | ( n11735 & ~n14546 ) ;
  assign n14542 = ( n1974 & n2604 ) | ( n1974 & ~n12605 ) | ( n2604 & ~n12605 ) ;
  assign n14543 = n14542 ^ n13655 ^ n5128 ;
  assign n14544 = n14543 ^ n2338 ^ n1343 ;
  assign n14545 = ( n3907 & ~n8565 ) | ( n3907 & n14544 ) | ( ~n8565 & n14544 ) ;
  assign n14548 = n14547 ^ n14545 ^ n8492 ;
  assign n14550 = ( n4204 & n7858 ) | ( n4204 & n13677 ) | ( n7858 & n13677 ) ;
  assign n14549 = ( ~n2787 & n5878 ) | ( ~n2787 & n7766 ) | ( n5878 & n7766 ) ;
  assign n14551 = n14550 ^ n14549 ^ 1'b0 ;
  assign n14552 = n5378 ^ n2337 ^ x106 ;
  assign n14553 = n14552 ^ n7173 ^ n2665 ;
  assign n14554 = ( n4385 & ~n8538 ) | ( n4385 & n14553 ) | ( ~n8538 & n14553 ) ;
  assign n14555 = n14554 ^ n12449 ^ n5808 ;
  assign n14556 = n14253 ^ n13741 ^ n732 ;
  assign n14557 = ( n719 & n8978 ) | ( n719 & n11861 ) | ( n8978 & n11861 ) ;
  assign n14558 = n8206 ^ n7029 ^ n5441 ;
  assign n14559 = ~n5313 & n14558 ;
  assign n14560 = n14559 ^ n6125 ^ n1152 ;
  assign n14561 = ( ~n365 & n683 ) | ( ~n365 & n14560 ) | ( n683 & n14560 ) ;
  assign n14562 = n10342 ^ n8307 ^ n1971 ;
  assign n14563 = n14562 ^ n8791 ^ n1939 ;
  assign n14567 = n13733 ^ n3869 ^ n3333 ;
  assign n14564 = ( n319 & ~n3527 ) | ( n319 & n6415 ) | ( ~n3527 & n6415 ) ;
  assign n14565 = ( n3265 & n14153 ) | ( n3265 & ~n14564 ) | ( n14153 & ~n14564 ) ;
  assign n14566 = ( ~n5291 & n7689 ) | ( ~n5291 & n14565 ) | ( n7689 & n14565 ) ;
  assign n14568 = n14567 ^ n14566 ^ n3473 ;
  assign n14569 = n9330 ^ n2473 ^ n1956 ;
  assign n14570 = n7614 ^ n2898 ^ n2573 ;
  assign n14571 = ~n7586 & n14570 ;
  assign n14572 = n14571 ^ n192 ^ 1'b0 ;
  assign n14573 = n14572 ^ n5757 ^ n1199 ;
  assign n14574 = ( ~n732 & n8632 ) | ( ~n732 & n14573 ) | ( n8632 & n14573 ) ;
  assign n14575 = ( n518 & ~n3982 ) | ( n518 & n4836 ) | ( ~n3982 & n4836 ) ;
  assign n14576 = ( ~n1872 & n3239 ) | ( ~n1872 & n9864 ) | ( n3239 & n9864 ) ;
  assign n14577 = ( n13704 & n14575 ) | ( n13704 & n14576 ) | ( n14575 & n14576 ) ;
  assign n14578 = n13805 ^ n2270 ^ 1'b0 ;
  assign n14579 = n14578 ^ n11526 ^ n1858 ;
  assign n14580 = n14579 ^ n4640 ^ n812 ;
  assign n14583 = n6361 & ~n12531 ;
  assign n14581 = n5667 ^ n4007 ^ n2903 ;
  assign n14582 = ( ~n3817 & n7349 ) | ( ~n3817 & n14581 ) | ( n7349 & n14581 ) ;
  assign n14584 = n14583 ^ n14582 ^ n5446 ;
  assign n14585 = ( n3104 & ~n14580 ) | ( n3104 & n14584 ) | ( ~n14580 & n14584 ) ;
  assign n14593 = n13162 ^ n10581 ^ n5444 ;
  assign n14592 = n4977 ^ n3613 ^ n1155 ;
  assign n14594 = n14593 ^ n14592 ^ n9760 ;
  assign n14586 = n10093 ^ n3249 ^ 1'b0 ;
  assign n14587 = n3007 | n14586 ;
  assign n14588 = n14587 ^ n8363 ^ n6642 ;
  assign n14589 = n14588 ^ x54 ^ 1'b0 ;
  assign n14590 = n8290 | n14589 ;
  assign n14591 = ( n3901 & ~n12401 ) | ( n3901 & n14590 ) | ( ~n12401 & n14590 ) ;
  assign n14595 = n14594 ^ n14591 ^ n683 ;
  assign n14596 = n13231 ^ n7066 ^ n4758 ;
  assign n14597 = ( ~n3478 & n4751 ) | ( ~n3478 & n14596 ) | ( n4751 & n14596 ) ;
  assign n14598 = ( n2236 & n10423 ) | ( n2236 & ~n13951 ) | ( n10423 & ~n13951 ) ;
  assign n14600 = ( n1055 & n1326 ) | ( n1055 & n3641 ) | ( n1326 & n3641 ) ;
  assign n14599 = n4779 | n7859 ;
  assign n14601 = n14600 ^ n14599 ^ 1'b0 ;
  assign n14602 = n3069 & n3840 ;
  assign n14603 = n14602 ^ x58 ^ 1'b0 ;
  assign n14604 = ( n4127 & n8268 ) | ( n4127 & n14603 ) | ( n8268 & n14603 ) ;
  assign n14605 = ( n10112 & n10342 ) | ( n10112 & n14604 ) | ( n10342 & n14604 ) ;
  assign n14606 = ( n4429 & ~n7333 ) | ( n4429 & n8370 ) | ( ~n7333 & n8370 ) ;
  assign n14607 = n14606 ^ n10189 ^ n6360 ;
  assign n14608 = n5970 ^ n1012 ^ n469 ;
  assign n14609 = ( n1693 & n2311 ) | ( n1693 & n10189 ) | ( n2311 & n10189 ) ;
  assign n14610 = ( x84 & n14608 ) | ( x84 & ~n14609 ) | ( n14608 & ~n14609 ) ;
  assign n14611 = ( n13334 & ~n14607 ) | ( n13334 & n14610 ) | ( ~n14607 & n14610 ) ;
  assign n14612 = n12984 ^ n8000 ^ n7414 ;
  assign n14613 = ( n4490 & ~n14611 ) | ( n4490 & n14612 ) | ( ~n14611 & n14612 ) ;
  assign n14614 = ( n2514 & n6284 ) | ( n2514 & ~n13305 ) | ( n6284 & ~n13305 ) ;
  assign n14615 = n3178 & ~n3364 ;
  assign n14616 = n14615 ^ n7091 ^ 1'b0 ;
  assign n14617 = n5804 & ~n14616 ;
  assign n14618 = ( ~n2280 & n14614 ) | ( ~n2280 & n14617 ) | ( n14614 & n14617 ) ;
  assign n14619 = n14388 ^ n4136 ^ n2489 ;
  assign n14620 = ~n6759 & n14619 ;
  assign n14621 = n14620 ^ n12763 ^ 1'b0 ;
  assign n14623 = n7577 ^ n4914 ^ n3853 ;
  assign n14624 = n14623 ^ n7531 ^ n3120 ;
  assign n14625 = ( ~n2354 & n9200 ) | ( ~n2354 & n14624 ) | ( n9200 & n14624 ) ;
  assign n14622 = n4513 & ~n5648 ;
  assign n14626 = n14625 ^ n14622 ^ 1'b0 ;
  assign n14630 = n527 | n2928 ;
  assign n14631 = n14630 ^ n679 ^ 1'b0 ;
  assign n14632 = ( ~n12637 & n12991 ) | ( ~n12637 & n14631 ) | ( n12991 & n14631 ) ;
  assign n14633 = n13259 | n14632 ;
  assign n14627 = n8438 ^ n5619 ^ n1326 ;
  assign n14628 = ( n2921 & n6471 ) | ( n2921 & ~n8815 ) | ( n6471 & ~n8815 ) ;
  assign n14629 = ( n7365 & ~n14627 ) | ( n7365 & n14628 ) | ( ~n14627 & n14628 ) ;
  assign n14634 = n14633 ^ n14629 ^ 1'b0 ;
  assign n14635 = n133 & ~n14121 ;
  assign n14636 = n14635 ^ n9818 ^ n4013 ;
  assign n14637 = n9454 ^ n7439 ^ n1882 ;
  assign n14638 = n1640 & ~n6798 ;
  assign n14639 = n4794 ^ n2863 ^ n2324 ;
  assign n14640 = ( n6171 & n14638 ) | ( n6171 & ~n14639 ) | ( n14638 & ~n14639 ) ;
  assign n14641 = ( n1563 & n4892 ) | ( n1563 & ~n14640 ) | ( n4892 & ~n14640 ) ;
  assign n14642 = ( n1543 & ~n2872 ) | ( n1543 & n3986 ) | ( ~n2872 & n3986 ) ;
  assign n14643 = ( n10685 & n14641 ) | ( n10685 & ~n14642 ) | ( n14641 & ~n14642 ) ;
  assign n14644 = ( n1328 & n3509 ) | ( n1328 & n8122 ) | ( n3509 & n8122 ) ;
  assign n14645 = n8075 | n14644 ;
  assign n14646 = n14645 ^ n7665 ^ 1'b0 ;
  assign n14647 = n2554 | n4066 ;
  assign n14648 = ( n2058 & n5972 ) | ( n2058 & ~n12472 ) | ( n5972 & ~n12472 ) ;
  assign n14649 = n14647 & ~n14648 ;
  assign n14650 = n8814 & n14649 ;
  assign n14651 = ( n3022 & n3748 ) | ( n3022 & n8924 ) | ( n3748 & n8924 ) ;
  assign n14652 = ( n3831 & n6069 ) | ( n3831 & ~n14651 ) | ( n6069 & ~n14651 ) ;
  assign n14653 = ( n2868 & n8070 ) | ( n2868 & n14652 ) | ( n8070 & n14652 ) ;
  assign n14654 = n14650 | n14653 ;
  assign n14655 = n14646 & ~n14654 ;
  assign n14656 = ( n3159 & n14643 ) | ( n3159 & ~n14655 ) | ( n14643 & ~n14655 ) ;
  assign n14657 = n11200 ^ n10045 ^ n7535 ;
  assign n14658 = ( ~n14637 & n14656 ) | ( ~n14637 & n14657 ) | ( n14656 & n14657 ) ;
  assign n14660 = ( n1801 & n3504 ) | ( n1801 & ~n5739 ) | ( n3504 & ~n5739 ) ;
  assign n14661 = n14660 ^ n13678 ^ n2852 ;
  assign n14662 = ( n454 & n4439 ) | ( n454 & ~n14661 ) | ( n4439 & ~n14661 ) ;
  assign n14659 = ~n535 & n5886 ;
  assign n14663 = n14662 ^ n14659 ^ 1'b0 ;
  assign n14665 = ( n3101 & n4647 ) | ( n3101 & ~n8134 ) | ( n4647 & ~n8134 ) ;
  assign n14666 = ( n4142 & n10334 ) | ( n4142 & n14665 ) | ( n10334 & n14665 ) ;
  assign n14664 = ( n7456 & n8480 ) | ( n7456 & n10282 ) | ( n8480 & n10282 ) ;
  assign n14667 = n14666 ^ n14664 ^ n691 ;
  assign n14669 = n7472 ^ n4221 ^ n2355 ;
  assign n14668 = n12548 ^ n4948 ^ n4425 ;
  assign n14670 = n14669 ^ n14668 ^ n4554 ;
  assign n14671 = n14670 ^ n11953 ^ n10310 ;
  assign n14674 = n4905 ^ n2896 ^ n913 ;
  assign n14672 = n2232 & n3526 ;
  assign n14673 = ( n10697 & ~n12578 ) | ( n10697 & n14672 ) | ( ~n12578 & n14672 ) ;
  assign n14675 = n14674 ^ n14673 ^ n9733 ;
  assign n14676 = ( n1955 & ~n4993 ) | ( n1955 & n9593 ) | ( ~n4993 & n9593 ) ;
  assign n14677 = ( ~n2596 & n6551 ) | ( ~n2596 & n14676 ) | ( n6551 & n14676 ) ;
  assign n14678 = n14677 ^ n10660 ^ n2107 ;
  assign n14679 = n9348 ^ n6049 ^ n581 ;
  assign n14680 = ~n4899 & n6880 ;
  assign n14681 = ( n6587 & n14141 ) | ( n6587 & n14680 ) | ( n14141 & n14680 ) ;
  assign n14684 = n6743 & n14129 ;
  assign n14682 = n7535 ^ n3581 ^ 1'b0 ;
  assign n14683 = n14682 ^ n10629 ^ 1'b0 ;
  assign n14685 = n14684 ^ n14683 ^ 1'b0 ;
  assign n14686 = ~n12426 & n14685 ;
  assign n14694 = n11439 ^ n7854 ^ 1'b0 ;
  assign n14695 = n2525 & ~n14694 ;
  assign n14696 = ( n882 & n1954 ) | ( n882 & ~n14695 ) | ( n1954 & ~n14695 ) ;
  assign n14697 = n14696 ^ n5414 ^ n1853 ;
  assign n14687 = n9550 ^ n6193 ^ n2428 ;
  assign n14688 = ( n5931 & n8040 ) | ( n5931 & ~n13974 ) | ( n8040 & ~n13974 ) ;
  assign n14689 = n14688 ^ n8393 ^ n278 ;
  assign n14690 = ( n5315 & ~n12524 ) | ( n5315 & n14061 ) | ( ~n12524 & n14061 ) ;
  assign n14691 = n14689 & n14690 ;
  assign n14692 = ~n12006 & n14691 ;
  assign n14693 = n14687 & ~n14692 ;
  assign n14698 = n14697 ^ n14693 ^ 1'b0 ;
  assign n14699 = ~n8341 & n12928 ;
  assign n14700 = n14082 ^ n9590 ^ n589 ;
  assign n14701 = n2392 & n14700 ;
  assign n14703 = n7514 ^ n5654 ^ n4213 ;
  assign n14702 = n1426 | n3042 ;
  assign n14704 = n14703 ^ n14702 ^ 1'b0 ;
  assign n14705 = ( ~n396 & n6883 ) | ( ~n396 & n7164 ) | ( n6883 & n7164 ) ;
  assign n14706 = n14705 ^ n6986 ^ n3311 ;
  assign n14707 = n5349 ^ n1094 ^ n431 ;
  assign n14708 = ( n3998 & n4205 ) | ( n3998 & n6674 ) | ( n4205 & n6674 ) ;
  assign n14709 = n14635 ^ n13976 ^ 1'b0 ;
  assign n14710 = n14708 & n14709 ;
  assign n14711 = ( ~n6795 & n14707 ) | ( ~n6795 & n14710 ) | ( n14707 & n14710 ) ;
  assign n14712 = n14711 ^ n10234 ^ x112 ;
  assign n14713 = n7593 & n8193 ;
  assign n14714 = ( n2459 & n11108 ) | ( n2459 & n14713 ) | ( n11108 & n14713 ) ;
  assign n14716 = n11424 ^ n4134 ^ n4048 ;
  assign n14717 = n14716 ^ n8857 ^ n7695 ;
  assign n14715 = ( ~n1672 & n8787 ) | ( ~n1672 & n12225 ) | ( n8787 & n12225 ) ;
  assign n14718 = n14717 ^ n14715 ^ n5843 ;
  assign n14719 = ( n587 & n14714 ) | ( n587 & ~n14718 ) | ( n14714 & ~n14718 ) ;
  assign n14720 = ( n1337 & n2810 ) | ( n1337 & ~n4212 ) | ( n2810 & ~n4212 ) ;
  assign n14721 = ( n5522 & ~n9618 ) | ( n5522 & n14720 ) | ( ~n9618 & n14720 ) ;
  assign n14722 = n1822 & n2839 ;
  assign n14723 = ~n11733 & n14722 ;
  assign n14724 = ~n3387 & n7438 ;
  assign n14725 = ~n1158 & n14724 ;
  assign n14726 = ( n6330 & n14723 ) | ( n6330 & n14725 ) | ( n14723 & n14725 ) ;
  assign n14727 = n14726 ^ n13491 ^ n12287 ;
  assign n14728 = n14727 ^ n11467 ^ 1'b0 ;
  assign n14729 = n14721 | n14728 ;
  assign n14730 = n8862 ^ n6809 ^ n1286 ;
  assign n14731 = n13304 ^ n4344 ^ 1'b0 ;
  assign n14732 = n4739 & n14731 ;
  assign n14733 = n14732 ^ n10040 ^ n8608 ;
  assign n14734 = ( n556 & n7346 ) | ( n556 & n14733 ) | ( n7346 & n14733 ) ;
  assign n14735 = ( n12581 & n14730 ) | ( n12581 & ~n14734 ) | ( n14730 & ~n14734 ) ;
  assign n14736 = n13548 ^ n687 ^ x88 ;
  assign n14737 = ( n3603 & n11594 ) | ( n3603 & n13411 ) | ( n11594 & n13411 ) ;
  assign n14741 = ( n1294 & ~n12663 ) | ( n1294 & n14078 ) | ( ~n12663 & n14078 ) ;
  assign n14742 = n14741 ^ n14484 ^ n4522 ;
  assign n14738 = n9949 ^ n2902 ^ n279 ;
  assign n14739 = ( n1588 & n10944 ) | ( n1588 & ~n14738 ) | ( n10944 & ~n14738 ) ;
  assign n14740 = n5897 | n14739 ;
  assign n14743 = n14742 ^ n14740 ^ 1'b0 ;
  assign n14744 = n11826 ^ n5164 ^ 1'b0 ;
  assign n14745 = ( n906 & ~n7570 ) | ( n906 & n7606 ) | ( ~n7570 & n7606 ) ;
  assign n14746 = n14745 ^ n7925 ^ n5369 ;
  assign n14747 = n14746 ^ n6513 ^ n5605 ;
  assign n14753 = ( ~n3407 & n3838 ) | ( ~n3407 & n9446 ) | ( n3838 & n9446 ) ;
  assign n14754 = n14753 ^ n10631 ^ n3619 ;
  assign n14750 = n8795 ^ n6838 ^ 1'b0 ;
  assign n14751 = n1110 & ~n14750 ;
  assign n14748 = ( n2166 & n7270 ) | ( n2166 & ~n11961 ) | ( n7270 & ~n11961 ) ;
  assign n14749 = n14748 ^ n2396 ^ 1'b0 ;
  assign n14752 = n14751 ^ n14749 ^ n4331 ;
  assign n14755 = n14754 ^ n14752 ^ n3743 ;
  assign n14756 = ( n4930 & ~n7439 ) | ( n4930 & n14755 ) | ( ~n7439 & n14755 ) ;
  assign n14757 = n5362 ^ n5040 ^ n3564 ;
  assign n14758 = n14757 ^ n12211 ^ n10772 ;
  assign n14760 = ( n1280 & ~n9181 ) | ( n1280 & n14593 ) | ( ~n9181 & n14593 ) ;
  assign n14759 = n7947 & n12157 ;
  assign n14761 = n14760 ^ n14759 ^ n4491 ;
  assign n14762 = ( n1367 & ~n4688 ) | ( n1367 & n14761 ) | ( ~n4688 & n14761 ) ;
  assign n14763 = ( ~n5564 & n13943 ) | ( ~n5564 & n14762 ) | ( n13943 & n14762 ) ;
  assign n14764 = n9512 ^ n3095 ^ n2251 ;
  assign n14765 = ( x14 & n502 ) | ( x14 & n3252 ) | ( n502 & n3252 ) ;
  assign n14766 = ~n14764 & n14765 ;
  assign n14767 = ( n6388 & ~n6681 ) | ( n6388 & n12486 ) | ( ~n6681 & n12486 ) ;
  assign n14768 = n14767 ^ n2503 ^ n192 ;
  assign n14769 = ( n2609 & n3223 ) | ( n2609 & n5168 ) | ( n3223 & n5168 ) ;
  assign n14770 = n14769 ^ n3471 ^ 1'b0 ;
  assign n14771 = n2807 & ~n14770 ;
  assign n14772 = ( ~n6292 & n10090 ) | ( ~n6292 & n10901 ) | ( n10090 & n10901 ) ;
  assign n14773 = n3049 & ~n5064 ;
  assign n14774 = n959 | n14773 ;
  assign n14775 = n14772 | n14774 ;
  assign n14777 = x102 & n297 ;
  assign n14776 = n3261 ^ n2429 ^ n1306 ;
  assign n14778 = n14777 ^ n14776 ^ 1'b0 ;
  assign n14779 = ~n7633 & n11226 ;
  assign n14780 = n14778 & n14779 ;
  assign n14781 = n14780 ^ n10568 ^ n2657 ;
  assign n14782 = ( n4980 & n13526 ) | ( n4980 & n14781 ) | ( n13526 & n14781 ) ;
  assign n14783 = ( n13222 & n14775 ) | ( n13222 & n14782 ) | ( n14775 & n14782 ) ;
  assign n14784 = ( n3466 & n14771 ) | ( n3466 & n14783 ) | ( n14771 & n14783 ) ;
  assign n14786 = ( ~n5385 & n7004 ) | ( ~n5385 & n13566 ) | ( n7004 & n13566 ) ;
  assign n14785 = ( n716 & n1625 ) | ( n716 & ~n1964 ) | ( n1625 & ~n1964 ) ;
  assign n14787 = n14786 ^ n14785 ^ n1181 ;
  assign n14788 = n3416 ^ n2160 ^ x108 ;
  assign n14789 = ( n4594 & n5974 ) | ( n4594 & ~n7184 ) | ( n5974 & ~n7184 ) ;
  assign n14790 = n14789 ^ n14008 ^ n8476 ;
  assign n14791 = ( n2850 & ~n13242 ) | ( n2850 & n14790 ) | ( ~n13242 & n14790 ) ;
  assign n14792 = n14791 ^ n1328 ^ 1'b0 ;
  assign n14793 = ( n8717 & n14788 ) | ( n8717 & ~n14792 ) | ( n14788 & ~n14792 ) ;
  assign n14794 = n3314 & ~n14793 ;
  assign n14799 = n10001 ^ n2913 ^ n879 ;
  assign n14800 = n8074 ^ n6262 ^ 1'b0 ;
  assign n14801 = n14799 | n14800 ;
  assign n14797 = n12955 & ~n13552 ;
  assign n14798 = n14797 ^ n7282 ^ n3462 ;
  assign n14795 = n11628 ^ n11144 ^ n8472 ;
  assign n14796 = ( n1510 & n3544 ) | ( n1510 & ~n14795 ) | ( n3544 & ~n14795 ) ;
  assign n14802 = n14801 ^ n14798 ^ n14796 ;
  assign n14803 = n9552 ^ n9426 ^ n3502 ;
  assign n14804 = n583 & n14803 ;
  assign n14805 = ~n14755 & n14804 ;
  assign n14806 = ( n3236 & n5748 ) | ( n3236 & n9837 ) | ( n5748 & n9837 ) ;
  assign n14807 = ( n5119 & n7552 ) | ( n5119 & n14806 ) | ( n7552 & n14806 ) ;
  assign n14808 = n14807 ^ n1708 ^ n643 ;
  assign n14812 = ( n246 & n8988 ) | ( n246 & n14669 ) | ( n8988 & n14669 ) ;
  assign n14813 = n14812 ^ n2004 ^ x40 ;
  assign n14810 = ( n7793 & n8475 ) | ( n7793 & n8613 ) | ( n8475 & n8613 ) ;
  assign n14811 = n14810 ^ n10265 ^ n10186 ;
  assign n14809 = n2992 | n12636 ;
  assign n14814 = n14813 ^ n14811 ^ n14809 ;
  assign n14815 = ( n1039 & n3010 ) | ( n1039 & n6425 ) | ( n3010 & n6425 ) ;
  assign n14816 = ( n2349 & n13393 ) | ( n2349 & ~n14815 ) | ( n13393 & ~n14815 ) ;
  assign n14817 = n7737 ^ n4614 ^ n581 ;
  assign n14818 = n6189 ^ n3741 ^ n3499 ;
  assign n14819 = ( n730 & ~n1244 ) | ( n730 & n4960 ) | ( ~n1244 & n4960 ) ;
  assign n14820 = ( n1551 & n5128 ) | ( n1551 & n14819 ) | ( n5128 & n14819 ) ;
  assign n14821 = ( n11806 & n14818 ) | ( n11806 & n14820 ) | ( n14818 & n14820 ) ;
  assign n14822 = ( n6964 & n14817 ) | ( n6964 & ~n14821 ) | ( n14817 & ~n14821 ) ;
  assign n14823 = n1796 & ~n14822 ;
  assign n14824 = ~n5039 & n14823 ;
  assign n14826 = n4799 ^ n1632 ^ n1544 ;
  assign n14825 = ~n7021 & n11144 ;
  assign n14827 = n14826 ^ n14825 ^ 1'b0 ;
  assign n14828 = n14827 ^ n398 ^ n207 ;
  assign n14829 = ( ~n465 & n10673 ) | ( ~n465 & n14828 ) | ( n10673 & n14828 ) ;
  assign n14834 = n8029 ^ n4021 ^ n1255 ;
  assign n14830 = n9526 & n10244 ;
  assign n14831 = n14830 ^ n11733 ^ 1'b0 ;
  assign n14832 = ~n3987 & n14831 ;
  assign n14833 = n3301 & ~n14832 ;
  assign n14835 = n14834 ^ n14833 ^ 1'b0 ;
  assign n14836 = ( n175 & ~n9441 ) | ( n175 & n14115 ) | ( ~n9441 & n14115 ) ;
  assign n14844 = ( n443 & n1559 ) | ( n443 & n2031 ) | ( n1559 & n2031 ) ;
  assign n14845 = n14844 ^ n4888 ^ n4247 ;
  assign n14841 = ( n3166 & n3905 ) | ( n3166 & ~n4640 ) | ( n3905 & ~n4640 ) ;
  assign n14838 = n8446 ^ n1280 ^ n859 ;
  assign n14839 = n14838 ^ n362 ^ n344 ;
  assign n14840 = n14839 ^ n10175 ^ n5182 ;
  assign n14842 = n14841 ^ n14840 ^ n6519 ;
  assign n14843 = n14842 ^ n14090 ^ 1'b0 ;
  assign n14837 = ( n4789 & ~n8905 ) | ( n4789 & n9817 ) | ( ~n8905 & n9817 ) ;
  assign n14846 = n14845 ^ n14843 ^ n14837 ;
  assign n14847 = n3019 ^ n1692 ^ n1291 ;
  assign n14848 = ( ~n2740 & n13619 ) | ( ~n2740 & n14847 ) | ( n13619 & n14847 ) ;
  assign n14849 = n8297 ^ n5285 ^ n1727 ;
  assign n14850 = ( n4015 & ~n14848 ) | ( n4015 & n14849 ) | ( ~n14848 & n14849 ) ;
  assign n14851 = n12687 ^ n9247 ^ n6241 ;
  assign n14852 = n14851 ^ n6993 ^ n2306 ;
  assign n14855 = n5567 ^ n2598 ^ n2132 ;
  assign n14856 = n14855 ^ n1655 ^ 1'b0 ;
  assign n14857 = n2848 | n14856 ;
  assign n14853 = n12661 ^ n10001 ^ n8538 ;
  assign n14854 = n14853 ^ n13299 ^ n625 ;
  assign n14858 = n14857 ^ n14854 ^ n3162 ;
  assign n14859 = n12429 ^ n2391 ^ 1'b0 ;
  assign n14860 = n5583 | n14859 ;
  assign n14861 = n8629 ^ n2747 ^ n1791 ;
  assign n14862 = n14861 ^ n5924 ^ n2978 ;
  assign n14863 = ( ~n3183 & n13689 ) | ( ~n3183 & n14862 ) | ( n13689 & n14862 ) ;
  assign n14864 = n14863 ^ n13529 ^ n3204 ;
  assign n14865 = n14860 & ~n14864 ;
  assign n14866 = n12014 ^ n2409 ^ n424 ;
  assign n14868 = n6591 ^ n5159 ^ n1080 ;
  assign n14869 = n14868 ^ n6985 ^ n6308 ;
  assign n14867 = ( ~n4408 & n7104 ) | ( ~n4408 & n8580 ) | ( n7104 & n8580 ) ;
  assign n14870 = n14869 ^ n14867 ^ n7905 ;
  assign n14871 = ( n5423 & n8900 ) | ( n5423 & n14870 ) | ( n8900 & n14870 ) ;
  assign n14872 = ( n3259 & ~n6374 ) | ( n3259 & n7488 ) | ( ~n6374 & n7488 ) ;
  assign n14874 = n2400 ^ n1584 ^ n296 ;
  assign n14873 = n11843 | n12102 ;
  assign n14875 = n14874 ^ n14873 ^ 1'b0 ;
  assign n14877 = n4037 & ~n6531 ;
  assign n14876 = n9503 ^ n3676 ^ n2840 ;
  assign n14878 = n14877 ^ n14876 ^ n5754 ;
  assign n14879 = n2932 & n6855 ;
  assign n14880 = n11916 & n14879 ;
  assign n14881 = n14880 ^ n10020 ^ n2246 ;
  assign n14882 = ( n152 & n1273 ) | ( n152 & n14881 ) | ( n1273 & n14881 ) ;
  assign n14883 = n7092 ^ n5685 ^ n343 ;
  assign n14884 = n4624 ^ n2113 ^ n1255 ;
  assign n14885 = n7961 ^ n4289 ^ n4008 ;
  assign n14886 = n4427 & ~n6061 ;
  assign n14887 = ~n14885 & n14886 ;
  assign n14888 = n14884 & ~n14887 ;
  assign n14889 = n522 & n14888 ;
  assign n14890 = ( ~n5262 & n7505 ) | ( ~n5262 & n14889 ) | ( n7505 & n14889 ) ;
  assign n14891 = ( n1129 & n2732 ) | ( n1129 & ~n6922 ) | ( n2732 & ~n6922 ) ;
  assign n14892 = ( ~n1024 & n11967 ) | ( ~n1024 & n14891 ) | ( n11967 & n14891 ) ;
  assign n14893 = n6723 ^ n4894 ^ 1'b0 ;
  assign n14904 = ( n2134 & n5535 ) | ( n2134 & n8585 ) | ( n5535 & n8585 ) ;
  assign n14902 = n9941 ^ n5682 ^ 1'b0 ;
  assign n14903 = ( n330 & n4408 ) | ( n330 & ~n14902 ) | ( n4408 & ~n14902 ) ;
  assign n14905 = n14904 ^ n14903 ^ n4615 ;
  assign n14894 = n2576 ^ n2557 ^ n226 ;
  assign n14895 = n14894 ^ n1822 ^ n176 ;
  assign n14896 = n11604 ^ n2513 ^ n288 ;
  assign n14897 = ( ~n633 & n5847 ) | ( ~n633 & n14896 ) | ( n5847 & n14896 ) ;
  assign n14898 = n14895 | n14897 ;
  assign n14899 = n14898 ^ n12938 ^ n12411 ;
  assign n14900 = n14116 ^ n7639 ^ n7382 ;
  assign n14901 = ( n2004 & n14899 ) | ( n2004 & ~n14900 ) | ( n14899 & ~n14900 ) ;
  assign n14906 = n14905 ^ n14901 ^ n7626 ;
  assign n14907 = n1069 & ~n5944 ;
  assign n14908 = ~n6919 & n14907 ;
  assign n14909 = n12112 | n14908 ;
  assign n14910 = n2496 | n14909 ;
  assign n14911 = n12895 ^ n7400 ^ n5395 ;
  assign n14915 = ( n6497 & n8198 ) | ( n6497 & n12811 ) | ( n8198 & n12811 ) ;
  assign n14912 = n6152 & ~n6409 ;
  assign n14913 = n6426 & n14912 ;
  assign n14914 = n14913 ^ n10336 ^ n364 ;
  assign n14916 = n14915 ^ n14914 ^ n6112 ;
  assign n14917 = n2608 & ~n14916 ;
  assign n14918 = n12586 ^ n5021 ^ n2419 ;
  assign n14919 = x46 & ~n14918 ;
  assign n14920 = n14919 ^ n5615 ^ 1'b0 ;
  assign n14921 = ~n13917 & n14920 ;
  assign n14922 = ~n6770 & n14921 ;
  assign n14923 = ( n6364 & n14917 ) | ( n6364 & n14922 ) | ( n14917 & n14922 ) ;
  assign n14924 = n11016 ^ n7180 ^ n4127 ;
  assign n14925 = ( n926 & n2453 ) | ( n926 & ~n5497 ) | ( n2453 & ~n5497 ) ;
  assign n14926 = ~n1976 & n9418 ;
  assign n14927 = ~n4392 & n14926 ;
  assign n14928 = n14927 ^ n11695 ^ 1'b0 ;
  assign n14929 = ~n6645 & n14928 ;
  assign n14930 = n14929 ^ n9510 ^ n7923 ;
  assign n14931 = ( n6287 & n7131 ) | ( n6287 & ~n14930 ) | ( n7131 & ~n14930 ) ;
  assign n14932 = ( n5193 & ~n8406 ) | ( n5193 & n14004 ) | ( ~n8406 & n14004 ) ;
  assign n14933 = n1568 | n14932 ;
  assign n14934 = n14931 & ~n14933 ;
  assign n14935 = ( n1105 & n6340 ) | ( n1105 & ~n13334 ) | ( n6340 & ~n13334 ) ;
  assign n14936 = ( ~n2759 & n6324 ) | ( ~n2759 & n8995 ) | ( n6324 & n8995 ) ;
  assign n14937 = n10012 ^ n7939 ^ n4057 ;
  assign n14938 = ( n7726 & n14936 ) | ( n7726 & n14937 ) | ( n14936 & n14937 ) ;
  assign n14939 = n14938 ^ n8648 ^ n4062 ;
  assign n14940 = ( n444 & n4423 ) | ( n444 & n11480 ) | ( n4423 & n11480 ) ;
  assign n14941 = n3229 & ~n14940 ;
  assign n14942 = n7805 ^ n3446 ^ 1'b0 ;
  assign n14943 = ( n2375 & n4730 ) | ( n2375 & ~n14942 ) | ( n4730 & ~n14942 ) ;
  assign n14944 = n946 & ~n2451 ;
  assign n14945 = n14944 ^ n12847 ^ 1'b0 ;
  assign n14946 = n14945 ^ n14703 ^ 1'b0 ;
  assign n14959 = n3854 ^ n2870 ^ n2320 ;
  assign n14958 = n14412 ^ n8275 ^ n5355 ;
  assign n14951 = n2100 ^ x18 ^ 1'b0 ;
  assign n14952 = n8933 & n14951 ;
  assign n14953 = n10271 ^ n8753 ^ n1727 ;
  assign n14954 = ( x80 & n4237 ) | ( x80 & n14953 ) | ( n4237 & n14953 ) ;
  assign n14955 = ( n13741 & n14952 ) | ( n13741 & n14954 ) | ( n14952 & n14954 ) ;
  assign n14956 = n14955 ^ n7016 ^ n2053 ;
  assign n14949 = n4063 ^ n2406 ^ n2100 ;
  assign n14947 = n1702 & ~n1758 ;
  assign n14948 = ~n3210 & n14947 ;
  assign n14950 = n14949 ^ n14948 ^ n5369 ;
  assign n14957 = n14956 ^ n14950 ^ n6719 ;
  assign n14960 = n14959 ^ n14958 ^ n14957 ;
  assign n14961 = n9669 ^ n4274 ^ 1'b0 ;
  assign n14962 = ~n12910 & n14961 ;
  assign n14968 = n4379 ^ n3688 ^ n1993 ;
  assign n14965 = ( ~n283 & n2645 ) | ( ~n283 & n3233 ) | ( n2645 & n3233 ) ;
  assign n14966 = n14965 ^ n9330 ^ n7737 ;
  assign n14963 = ~n1523 & n5149 ;
  assign n14964 = ( n211 & ~n2322 ) | ( n211 & n14963 ) | ( ~n2322 & n14963 ) ;
  assign n14967 = n14966 ^ n14964 ^ n1553 ;
  assign n14969 = n14968 ^ n14967 ^ n6570 ;
  assign n14970 = ( n3224 & n4540 ) | ( n3224 & ~n9324 ) | ( n4540 & ~n9324 ) ;
  assign n14971 = n14440 ^ n13756 ^ n2912 ;
  assign n14972 = ( n2616 & n11649 ) | ( n2616 & n14971 ) | ( n11649 & n14971 ) ;
  assign n14973 = ( ~n14006 & n14970 ) | ( ~n14006 & n14972 ) | ( n14970 & n14972 ) ;
  assign n14974 = ( n3180 & n14969 ) | ( n3180 & ~n14973 ) | ( n14969 & ~n14973 ) ;
  assign n14975 = n10979 ^ n3422 ^ n2905 ;
  assign n14977 = n14651 ^ n6555 ^ n2421 ;
  assign n14976 = n11569 ^ n5630 ^ n3841 ;
  assign n14978 = n14977 ^ n14976 ^ n7577 ;
  assign n14979 = n14978 ^ n14293 ^ n219 ;
  assign n14980 = ( n1062 & ~n3992 ) | ( n1062 & n10930 ) | ( ~n3992 & n10930 ) ;
  assign n14981 = n7416 ^ n6037 ^ n3178 ;
  assign n14982 = n14981 ^ n5110 ^ 1'b0 ;
  assign n14983 = n14215 & ~n14982 ;
  assign n14984 = n4770 & n14983 ;
  assign n14985 = n14984 ^ n13011 ^ 1'b0 ;
  assign n14986 = ( n1857 & n4880 ) | ( n1857 & n14259 ) | ( n4880 & n14259 ) ;
  assign n14987 = ( n694 & n7576 ) | ( n694 & ~n14986 ) | ( n7576 & ~n14986 ) ;
  assign n14988 = ( n7246 & n14985 ) | ( n7246 & n14987 ) | ( n14985 & n14987 ) ;
  assign n14989 = ( n13315 & n14980 ) | ( n13315 & ~n14988 ) | ( n14980 & ~n14988 ) ;
  assign n14990 = n13946 ^ n1255 ^ n917 ;
  assign n14991 = ( n3061 & ~n3503 ) | ( n3061 & n14990 ) | ( ~n3503 & n14990 ) ;
  assign n14992 = n14991 ^ n2328 ^ n400 ;
  assign n14993 = n8677 ^ n6479 ^ n1693 ;
  assign n14994 = n14993 ^ n2332 ^ n2062 ;
  assign n14995 = n14994 ^ n12267 ^ n4901 ;
  assign n14996 = ( n8857 & n10772 ) | ( n8857 & ~n11310 ) | ( n10772 & ~n11310 ) ;
  assign n14997 = n7418 ^ n6477 ^ n1706 ;
  assign n14998 = ( ~n14995 & n14996 ) | ( ~n14995 & n14997 ) | ( n14996 & n14997 ) ;
  assign n14999 = n14898 ^ n8886 ^ n6216 ;
  assign n15000 = n14999 ^ n6884 ^ n5477 ;
  assign n15001 = ( n1858 & ~n2436 ) | ( n1858 & n3762 ) | ( ~n2436 & n3762 ) ;
  assign n15002 = n15001 ^ n5197 ^ n2673 ;
  assign n15003 = n15002 ^ n4029 ^ n555 ;
  assign n15005 = ( n2507 & n3670 ) | ( n2507 & ~n5314 ) | ( n3670 & ~n5314 ) ;
  assign n15006 = ~n1597 & n15005 ;
  assign n15007 = n15006 ^ n11007 ^ 1'b0 ;
  assign n15004 = ( n3394 & n3412 ) | ( n3394 & n7192 ) | ( n3412 & n7192 ) ;
  assign n15008 = n15007 ^ n15004 ^ n11982 ;
  assign n15009 = n15008 ^ n9968 ^ n2904 ;
  assign n15010 = n14443 ^ n14275 ^ n6704 ;
  assign n15011 = ( n3685 & n4064 ) | ( n3685 & ~n15010 ) | ( n4064 & ~n15010 ) ;
  assign n15012 = ( n1738 & ~n3318 ) | ( n1738 & n6643 ) | ( ~n3318 & n6643 ) ;
  assign n15013 = n15012 ^ n10881 ^ 1'b0 ;
  assign n15014 = n15013 ^ n7459 ^ n6288 ;
  assign n15023 = n12216 ^ n5815 ^ 1'b0 ;
  assign n15024 = n8934 & n15023 ;
  assign n15015 = ( n4655 & n5364 ) | ( n4655 & ~n13382 ) | ( n5364 & ~n13382 ) ;
  assign n15016 = ( x17 & n3317 ) | ( x17 & ~n15015 ) | ( n3317 & ~n15015 ) ;
  assign n15019 = n3939 | n7685 ;
  assign n15020 = n13780 | n15019 ;
  assign n15017 = n4403 ^ n1995 ^ n1347 ;
  assign n15018 = n15017 ^ n11930 ^ n7234 ;
  assign n15021 = n15020 ^ n15018 ^ n14674 ;
  assign n15022 = ( n1103 & n15016 ) | ( n1103 & n15021 ) | ( n15016 & n15021 ) ;
  assign n15025 = n15024 ^ n15022 ^ n3683 ;
  assign n15026 = n4068 ^ n1544 ^ n384 ;
  assign n15027 = n15026 ^ n13635 ^ n1287 ;
  assign n15028 = n10012 ^ n8877 ^ 1'b0 ;
  assign n15029 = n15028 ^ n10623 ^ n2670 ;
  assign n15030 = ~n2332 & n10577 ;
  assign n15031 = n10326 & n15030 ;
  assign n15032 = n15031 ^ n12057 ^ n9709 ;
  assign n15042 = n13601 ^ n7141 ^ n4634 ;
  assign n15036 = n1597 ^ n1349 ^ 1'b0 ;
  assign n15037 = n15036 ^ n14159 ^ n11347 ;
  assign n15038 = n15037 ^ n9375 ^ n5022 ;
  assign n15039 = n7029 ^ n6258 ^ n6007 ;
  assign n15040 = ~n2653 & n15039 ;
  assign n15041 = ~n15038 & n15040 ;
  assign n15033 = n9247 ^ n4321 ^ n723 ;
  assign n15034 = n5939 | n15033 ;
  assign n15035 = n15034 ^ n12386 ^ n11458 ;
  assign n15043 = n15042 ^ n15041 ^ n15035 ;
  assign n15044 = n11662 ^ n10223 ^ n2200 ;
  assign n15045 = n15044 ^ n1546 ^ 1'b0 ;
  assign n15048 = ( n1693 & ~n3360 ) | ( n1693 & n5266 ) | ( ~n3360 & n5266 ) ;
  assign n15049 = n15048 ^ n8242 ^ n4015 ;
  assign n15046 = ( n759 & n5703 ) | ( n759 & ~n8628 ) | ( n5703 & ~n8628 ) ;
  assign n15047 = n15046 ^ n8703 ^ n4335 ;
  assign n15050 = n15049 ^ n15047 ^ n6104 ;
  assign n15051 = n9276 ^ n8370 ^ n814 ;
  assign n15052 = n11488 ^ n8242 ^ n5894 ;
  assign n15053 = ( ~n1770 & n7340 ) | ( ~n1770 & n15052 ) | ( n7340 & n15052 ) ;
  assign n15054 = n15053 ^ n11220 ^ 1'b0 ;
  assign n15055 = n7338 ^ n5027 ^ 1'b0 ;
  assign n15056 = ( n889 & n9857 ) | ( n889 & n14224 ) | ( n9857 & n14224 ) ;
  assign n15057 = ( ~n9084 & n15055 ) | ( ~n9084 & n15056 ) | ( n15055 & n15056 ) ;
  assign n15058 = ( n2613 & n6531 ) | ( n2613 & n15057 ) | ( n6531 & n15057 ) ;
  assign n15059 = ( n955 & n1334 ) | ( n955 & n6494 ) | ( n1334 & n6494 ) ;
  assign n15060 = ( ~n2021 & n8481 ) | ( ~n2021 & n15059 ) | ( n8481 & n15059 ) ;
  assign n15061 = n11515 ^ n4703 ^ n2204 ;
  assign n15062 = ( n5630 & n7448 ) | ( n5630 & ~n9960 ) | ( n7448 & ~n9960 ) ;
  assign n15063 = ( n15060 & n15061 ) | ( n15060 & n15062 ) | ( n15061 & n15062 ) ;
  assign n15064 = ( n8895 & ~n14848 ) | ( n8895 & n15063 ) | ( ~n14848 & n15063 ) ;
  assign n15065 = ( ~n9733 & n15058 ) | ( ~n9733 & n15064 ) | ( n15058 & n15064 ) ;
  assign n15066 = ( n5446 & n9476 ) | ( n5446 & n14904 ) | ( n9476 & n14904 ) ;
  assign n15067 = n15066 ^ n8946 ^ 1'b0 ;
  assign n15068 = n10310 | n15067 ;
  assign n15072 = n484 | n8015 ;
  assign n15073 = n15072 ^ n6701 ^ 1'b0 ;
  assign n15069 = n11333 ^ n2200 ^ 1'b0 ;
  assign n15070 = n6189 & ~n15069 ;
  assign n15071 = ~n4991 & n15070 ;
  assign n15074 = n15073 ^ n15071 ^ n12062 ;
  assign n15075 = ( n1135 & n6784 ) | ( n1135 & ~n15074 ) | ( n6784 & ~n15074 ) ;
  assign n15076 = n9303 | n13198 ;
  assign n15077 = n15076 ^ n14970 ^ n10112 ;
  assign n15078 = n5228 ^ n3743 ^ n1235 ;
  assign n15079 = n10971 | n15078 ;
  assign n15080 = n15079 ^ n11279 ^ 1'b0 ;
  assign n15081 = ~n715 & n15080 ;
  assign n15082 = ( ~n12316 & n15077 ) | ( ~n12316 & n15081 ) | ( n15077 & n15081 ) ;
  assign n15083 = n11580 ^ n5256 ^ n2769 ;
  assign n15084 = ( ~n2712 & n9270 ) | ( ~n2712 & n13335 ) | ( n9270 & n13335 ) ;
  assign n15085 = n4078 ^ n2485 ^ 1'b0 ;
  assign n15086 = n2741 | n8244 ;
  assign n15087 = n15086 ^ n2441 ^ 1'b0 ;
  assign n15088 = n15087 ^ n14002 ^ n3922 ;
  assign n15089 = ( n2917 & ~n15085 ) | ( n2917 & n15088 ) | ( ~n15085 & n15088 ) ;
  assign n15090 = ( n9299 & ~n10809 ) | ( n9299 & n13976 ) | ( ~n10809 & n13976 ) ;
  assign n15091 = ( n6145 & n15089 ) | ( n6145 & n15090 ) | ( n15089 & n15090 ) ;
  assign n15092 = n9079 ^ n1730 ^ n1129 ;
  assign n15093 = ( ~n5383 & n9915 ) | ( ~n5383 & n15092 ) | ( n9915 & n15092 ) ;
  assign n15094 = ( n2601 & n6539 ) | ( n2601 & n15093 ) | ( n6539 & n15093 ) ;
  assign n15095 = n15094 ^ x6 ^ 1'b0 ;
  assign n15096 = n5246 | n15095 ;
  assign n15097 = ( n647 & ~n14717 ) | ( n647 & n15096 ) | ( ~n14717 & n15096 ) ;
  assign n15098 = ~n3192 & n7733 ;
  assign n15099 = n15098 ^ n3422 ^ 1'b0 ;
  assign n15100 = ( n1809 & ~n15097 ) | ( n1809 & n15099 ) | ( ~n15097 & n15099 ) ;
  assign n15105 = ( n1596 & ~n4595 ) | ( n1596 & n9939 ) | ( ~n4595 & n9939 ) ;
  assign n15106 = ( n614 & n5525 ) | ( n614 & ~n15105 ) | ( n5525 & ~n15105 ) ;
  assign n15102 = n12008 ^ n1446 ^ n524 ;
  assign n15103 = ( n718 & n5153 ) | ( n718 & ~n15102 ) | ( n5153 & ~n15102 ) ;
  assign n15104 = n15103 ^ n12018 ^ n150 ;
  assign n15101 = n10819 & ~n14619 ;
  assign n15107 = n15106 ^ n15104 ^ n15101 ;
  assign n15108 = ( n3107 & n4468 ) | ( n3107 & n8910 ) | ( n4468 & n8910 ) ;
  assign n15109 = ( ~n6924 & n14129 ) | ( ~n6924 & n15108 ) | ( n14129 & n15108 ) ;
  assign n15110 = ( n3704 & n5375 ) | ( n3704 & n7459 ) | ( n5375 & n7459 ) ;
  assign n15111 = ( n2694 & n9604 ) | ( n2694 & ~n10444 ) | ( n9604 & ~n10444 ) ;
  assign n15112 = ( ~n10140 & n15110 ) | ( ~n10140 & n15111 ) | ( n15110 & n15111 ) ;
  assign n15113 = n790 & n10266 ;
  assign n15114 = n7151 & n15113 ;
  assign n15115 = ( n1403 & n2745 ) | ( n1403 & n11769 ) | ( n2745 & n11769 ) ;
  assign n15116 = ( n8199 & n12906 ) | ( n8199 & ~n15115 ) | ( n12906 & ~n15115 ) ;
  assign n15117 = n15116 ^ n9845 ^ n4131 ;
  assign n15118 = n13617 ^ n12232 ^ n9001 ;
  assign n15119 = ( n9268 & n10148 ) | ( n9268 & n15118 ) | ( n10148 & n15118 ) ;
  assign n15120 = n15119 ^ n3392 ^ n1013 ;
  assign n15121 = ( ~n1087 & n2563 ) | ( ~n1087 & n2820 ) | ( n2563 & n2820 ) ;
  assign n15122 = ~n4020 & n15121 ;
  assign n15123 = n8958 & n15122 ;
  assign n15124 = n15123 ^ n14164 ^ n5368 ;
  assign n15125 = ( x82 & n4517 ) | ( x82 & n7924 ) | ( n4517 & n7924 ) ;
  assign n15126 = n15125 ^ n6245 ^ n6111 ;
  assign n15129 = n1761 & n9391 ;
  assign n15130 = n4203 & n15129 ;
  assign n15127 = n13272 ^ n11064 ^ n7227 ;
  assign n15128 = ( n2640 & n5754 ) | ( n2640 & ~n15127 ) | ( n5754 & ~n15127 ) ;
  assign n15131 = n15130 ^ n15128 ^ n5386 ;
  assign n15132 = ( x9 & ~n5155 ) | ( x9 & n5320 ) | ( ~n5155 & n5320 ) ;
  assign n15133 = ( n3685 & n5601 ) | ( n3685 & ~n5877 ) | ( n5601 & ~n5877 ) ;
  assign n15134 = ( n9328 & n15132 ) | ( n9328 & ~n15133 ) | ( n15132 & ~n15133 ) ;
  assign n15135 = n15134 ^ n9053 ^ 1'b0 ;
  assign n15136 = n7766 & ~n15135 ;
  assign n15137 = ( n2024 & ~n3104 ) | ( n2024 & n8514 ) | ( ~n3104 & n8514 ) ;
  assign n15138 = n7961 ^ n3377 ^ n853 ;
  assign n15139 = ( n3611 & n15137 ) | ( n3611 & ~n15138 ) | ( n15137 & ~n15138 ) ;
  assign n15140 = n15139 ^ n5749 ^ n4411 ;
  assign n15141 = n6224 ^ n5922 ^ n4056 ;
  assign n15142 = ( ~n658 & n8301 ) | ( ~n658 & n9107 ) | ( n8301 & n9107 ) ;
  assign n15144 = ( n305 & n2930 ) | ( n305 & n7911 ) | ( n2930 & n7911 ) ;
  assign n15143 = ( n1470 & ~n5840 ) | ( n1470 & n13630 ) | ( ~n5840 & n13630 ) ;
  assign n15145 = n15144 ^ n15143 ^ n10551 ;
  assign n15146 = n15142 & n15145 ;
  assign n15147 = n10131 & n15146 ;
  assign n15149 = ( n3116 & ~n3293 ) | ( n3116 & n4311 ) | ( ~n3293 & n4311 ) ;
  assign n15150 = ~n8272 & n15149 ;
  assign n15151 = n15150 ^ n1267 ^ 1'b0 ;
  assign n15148 = ( ~n8034 & n8075 ) | ( ~n8034 & n9338 ) | ( n8075 & n9338 ) ;
  assign n15152 = n15151 ^ n15148 ^ n7818 ;
  assign n15153 = n8623 ^ n2836 ^ n2519 ;
  assign n15154 = n15153 ^ n4257 ^ 1'b0 ;
  assign n15155 = n15154 ^ n7540 ^ n2751 ;
  assign n15156 = ( n3631 & ~n7207 ) | ( n3631 & n13623 ) | ( ~n7207 & n13623 ) ;
  assign n15157 = n15092 ^ n13935 ^ n1940 ;
  assign n15158 = ( ~n10598 & n14248 ) | ( ~n10598 & n15157 ) | ( n14248 & n15157 ) ;
  assign n15161 = ~n792 & n13171 ;
  assign n15162 = n15161 ^ n2668 ^ 1'b0 ;
  assign n15159 = n3202 & n9096 ;
  assign n15160 = n15159 ^ n3283 ^ 1'b0 ;
  assign n15163 = n15162 ^ n15160 ^ n14399 ;
  assign n15164 = ( n1963 & n4799 ) | ( n1963 & n10941 ) | ( n4799 & n10941 ) ;
  assign n15165 = n2555 ^ n2179 ^ n1862 ;
  assign n15166 = ( ~n2226 & n11052 ) | ( ~n2226 & n15165 ) | ( n11052 & n15165 ) ;
  assign n15167 = n11042 ^ n906 ^ 1'b0 ;
  assign n15168 = n10611 & n15167 ;
  assign n15169 = n6038 ^ n381 ^ 1'b0 ;
  assign n15170 = ~n9905 & n15169 ;
  assign n15171 = n15170 ^ n2540 ^ n2193 ;
  assign n15172 = n8738 ^ n6904 ^ n4213 ;
  assign n15173 = ~n3750 & n8352 ;
  assign n15174 = n15173 ^ n8713 ^ 1'b0 ;
  assign n15175 = ( n2579 & n3044 ) | ( n2579 & n15174 ) | ( n3044 & n15174 ) ;
  assign n15176 = ( n5166 & ~n14608 ) | ( n5166 & n15175 ) | ( ~n14608 & n15175 ) ;
  assign n15177 = n13707 ^ n13352 ^ n3257 ;
  assign n15178 = ( x126 & n5886 ) | ( x126 & ~n12072 ) | ( n5886 & ~n12072 ) ;
  assign n15179 = n13827 ^ n5012 ^ n3972 ;
  assign n15180 = ( n4141 & n10787 ) | ( n4141 & n12697 ) | ( n10787 & n12697 ) ;
  assign n15187 = ( ~n2368 & n4497 ) | ( ~n2368 & n4884 ) | ( n4497 & n4884 ) ;
  assign n15188 = ( ~n4461 & n5157 ) | ( ~n4461 & n15187 ) | ( n5157 & n15187 ) ;
  assign n15189 = n15188 ^ n8992 ^ n2604 ;
  assign n15181 = n2002 | n3362 ;
  assign n15182 = n6428 | n15181 ;
  assign n15183 = ( n6491 & n9481 ) | ( n6491 & ~n15182 ) | ( n9481 & ~n15182 ) ;
  assign n15184 = ( n1431 & ~n1517 ) | ( n1431 & n15183 ) | ( ~n1517 & n15183 ) ;
  assign n15185 = n15184 ^ n12860 ^ n8074 ;
  assign n15186 = n9395 & ~n15185 ;
  assign n15190 = n15189 ^ n15186 ^ 1'b0 ;
  assign n15191 = n1331 ^ n867 ^ n670 ;
  assign n15192 = n15191 ^ n1219 ^ n883 ;
  assign n15193 = ( n2948 & n8614 ) | ( n2948 & ~n15192 ) | ( n8614 & ~n15192 ) ;
  assign n15194 = ( n4646 & n5978 ) | ( n4646 & ~n15193 ) | ( n5978 & ~n15193 ) ;
  assign n15195 = n10103 ^ n6871 ^ n5762 ;
  assign n15196 = n15195 ^ n10545 ^ n7792 ;
  assign n15197 = n15196 ^ n6582 ^ n4562 ;
  assign n15198 = n15197 ^ n12992 ^ n7860 ;
  assign n15199 = ~n3897 & n7562 ;
  assign n15200 = n15199 ^ n3977 ^ 1'b0 ;
  assign n15201 = n3327 ^ n2837 ^ n2501 ;
  assign n15202 = n6351 & ~n10447 ;
  assign n15203 = n13878 & n15202 ;
  assign n15204 = ( n12413 & n15201 ) | ( n12413 & ~n15203 ) | ( n15201 & ~n15203 ) ;
  assign n15210 = n9892 ^ n1743 ^ n373 ;
  assign n15205 = ( n390 & n478 ) | ( n390 & n9284 ) | ( n478 & n9284 ) ;
  assign n15206 = n13667 ^ n8267 ^ n1995 ;
  assign n15207 = ( n1672 & n3240 ) | ( n1672 & n5644 ) | ( n3240 & n5644 ) ;
  assign n15208 = ( n4066 & n15206 ) | ( n4066 & n15207 ) | ( n15206 & n15207 ) ;
  assign n15209 = ( ~n6158 & n15205 ) | ( ~n6158 & n15208 ) | ( n15205 & n15208 ) ;
  assign n15211 = n15210 ^ n15209 ^ n8255 ;
  assign n15212 = n9414 ^ n8050 ^ n2091 ;
  assign n15216 = n15206 ^ n14880 ^ 1'b0 ;
  assign n15213 = n14803 ^ n10472 ^ n591 ;
  assign n15214 = ~n8714 & n15213 ;
  assign n15215 = ~n7076 & n15214 ;
  assign n15217 = n15216 ^ n15215 ^ n2169 ;
  assign n15218 = n15201 ^ n8168 ^ 1'b0 ;
  assign n15219 = n10905 & ~n11416 ;
  assign n15220 = n15218 & n15219 ;
  assign n15221 = n11902 ^ n11177 ^ n2638 ;
  assign n15222 = n15221 ^ n7694 ^ n5398 ;
  assign n15223 = n10045 ^ n3264 ^ 1'b0 ;
  assign n15224 = ~n8967 & n15223 ;
  assign n15225 = n15224 ^ n575 ^ 1'b0 ;
  assign n15226 = n15225 ^ n7243 ^ n3303 ;
  assign n15227 = n10923 ^ n6195 ^ 1'b0 ;
  assign n15228 = n15226 & ~n15227 ;
  assign n15229 = ( n5093 & n10107 ) | ( n5093 & n15228 ) | ( n10107 & n15228 ) ;
  assign n15230 = ( ~n4269 & n6290 ) | ( ~n4269 & n15229 ) | ( n6290 & n15229 ) ;
  assign n15231 = ( n422 & ~n2615 ) | ( n422 & n4787 ) | ( ~n2615 & n4787 ) ;
  assign n15232 = ( n1246 & n11245 ) | ( n1246 & ~n15231 ) | ( n11245 & ~n15231 ) ;
  assign n15233 = ( n2037 & ~n11146 ) | ( n2037 & n13748 ) | ( ~n11146 & n13748 ) ;
  assign n15234 = ( ~n11474 & n15232 ) | ( ~n11474 & n15233 ) | ( n15232 & n15233 ) ;
  assign n15235 = n1557 | n5307 ;
  assign n15236 = n15235 ^ n11907 ^ n3554 ;
  assign n15237 = n14388 ^ n4176 ^ n4025 ;
  assign n15238 = n9564 ^ n6697 ^ n6590 ;
  assign n15239 = n1351 ^ n164 ^ 1'b0 ;
  assign n15240 = ~n7349 & n15239 ;
  assign n15241 = n15240 ^ n12229 ^ 1'b0 ;
  assign n15242 = ( n268 & ~n3364 ) | ( n268 & n15241 ) | ( ~n3364 & n15241 ) ;
  assign n15243 = ( n4122 & n7696 ) | ( n4122 & ~n15242 ) | ( n7696 & ~n15242 ) ;
  assign n15244 = n1592 ^ n1129 ^ 1'b0 ;
  assign n15245 = ~n683 & n15244 ;
  assign n15246 = ( n6340 & n11816 ) | ( n6340 & n15245 ) | ( n11816 & n15245 ) ;
  assign n15247 = n8885 ^ n2761 ^ n360 ;
  assign n15248 = ( n656 & ~n4645 ) | ( n656 & n15247 ) | ( ~n4645 & n15247 ) ;
  assign n15249 = ( n3753 & ~n6770 ) | ( n3753 & n15248 ) | ( ~n6770 & n15248 ) ;
  assign n15250 = n319 | n15249 ;
  assign n15251 = n5664 ^ n3370 ^ n876 ;
  assign n15252 = n11928 ^ n11064 ^ n5253 ;
  assign n15253 = ( n2050 & ~n15251 ) | ( n2050 & n15252 ) | ( ~n15251 & n15252 ) ;
  assign n15254 = ( n1134 & n1425 ) | ( n1134 & ~n7403 ) | ( n1425 & ~n7403 ) ;
  assign n15255 = ( n6320 & ~n10411 ) | ( n6320 & n15254 ) | ( ~n10411 & n15254 ) ;
  assign n15256 = n15255 ^ n7047 ^ n3543 ;
  assign n15257 = n15256 ^ n4034 ^ n3056 ;
  assign n15258 = ( n4471 & n12013 ) | ( n4471 & n15257 ) | ( n12013 & n15257 ) ;
  assign n15259 = n15258 ^ n8545 ^ n4766 ;
  assign n15261 = n11313 ^ n6329 ^ n2398 ;
  assign n15260 = n8712 & n10785 ;
  assign n15262 = n15261 ^ n15260 ^ 1'b0 ;
  assign n15268 = n14990 ^ n5193 ^ n1512 ;
  assign n15263 = ( ~n1166 & n4926 ) | ( ~n1166 & n10114 ) | ( n4926 & n10114 ) ;
  assign n15264 = n12899 ^ n12088 ^ 1'b0 ;
  assign n15265 = n15263 | n15264 ;
  assign n15266 = ( n6805 & n7000 ) | ( n6805 & ~n15265 ) | ( n7000 & ~n15265 ) ;
  assign n15267 = n1508 & ~n15266 ;
  assign n15269 = n15268 ^ n15267 ^ 1'b0 ;
  assign n15270 = n7342 ^ n3190 ^ n2833 ;
  assign n15271 = n15270 ^ n15059 ^ n13292 ;
  assign n15272 = n10749 ^ n6787 ^ 1'b0 ;
  assign n15273 = n15272 ^ n2358 ^ n853 ;
  assign n15274 = n917 ^ n900 ^ n396 ;
  assign n15275 = n15274 ^ n8286 ^ n484 ;
  assign n15276 = ( n1305 & n7581 ) | ( n1305 & ~n8206 ) | ( n7581 & ~n8206 ) ;
  assign n15277 = ( n1063 & n9312 ) | ( n1063 & ~n15276 ) | ( n9312 & ~n15276 ) ;
  assign n15278 = ( n5743 & n13509 ) | ( n5743 & ~n15277 ) | ( n13509 & ~n15277 ) ;
  assign n15283 = ( n1598 & n2519 ) | ( n1598 & ~n2848 ) | ( n2519 & ~n2848 ) ;
  assign n15280 = n12947 ^ n8412 ^ n193 ;
  assign n15281 = ( ~x48 & n6255 ) | ( ~x48 & n15280 ) | ( n6255 & n15280 ) ;
  assign n15279 = n14017 ^ n10795 ^ n5903 ;
  assign n15282 = n15281 ^ n15279 ^ n949 ;
  assign n15284 = n15283 ^ n15282 ^ n4641 ;
  assign n15288 = n9622 ^ n5921 ^ n1709 ;
  assign n15287 = n10107 ^ n4711 ^ n4602 ;
  assign n15285 = n6412 | n8686 ;
  assign n15286 = n15285 ^ x56 ^ 1'b0 ;
  assign n15289 = n15288 ^ n15287 ^ n15286 ;
  assign n15290 = ( x14 & ~n8828 ) | ( x14 & n10576 ) | ( ~n8828 & n10576 ) ;
  assign n15291 = n15290 ^ n7595 ^ n1179 ;
  assign n15292 = n13074 ^ n4974 ^ 1'b0 ;
  assign n15293 = n15292 ^ n7313 ^ n2537 ;
  assign n15301 = ( ~n2038 & n7090 ) | ( ~n2038 & n8294 ) | ( n7090 & n8294 ) ;
  assign n15294 = n6180 ^ n1624 ^ n511 ;
  assign n15295 = ( n1262 & ~n7229 ) | ( n1262 & n8392 ) | ( ~n7229 & n8392 ) ;
  assign n15296 = ( ~n2557 & n10522 ) | ( ~n2557 & n15295 ) | ( n10522 & n15295 ) ;
  assign n15297 = n15296 ^ n4497 ^ n1793 ;
  assign n15298 = n8873 & ~n15297 ;
  assign n15299 = ~n11760 & n15298 ;
  assign n15300 = ( n7692 & n15294 ) | ( n7692 & ~n15299 ) | ( n15294 & ~n15299 ) ;
  assign n15302 = n15301 ^ n15300 ^ n7722 ;
  assign n15304 = n4581 ^ n3484 ^ n1031 ;
  assign n15303 = n806 & n4039 ;
  assign n15305 = n15304 ^ n15303 ^ 1'b0 ;
  assign n15306 = ( ~n3289 & n9774 ) | ( ~n3289 & n15305 ) | ( n9774 & n15305 ) ;
  assign n15307 = ( ~n781 & n7046 ) | ( ~n781 & n10146 ) | ( n7046 & n10146 ) ;
  assign n15308 = ~n9012 & n9377 ;
  assign n15309 = n15308 ^ n510 ^ 1'b0 ;
  assign n15310 = n15307 | n15309 ;
  assign n15311 = n8416 ^ n3940 ^ n1815 ;
  assign n15312 = n15311 ^ n12073 ^ n978 ;
  assign n15313 = ~n4832 & n11844 ;
  assign n15314 = ~n11311 & n15313 ;
  assign n15315 = ~n5123 & n9036 ;
  assign n15316 = ~n4839 & n15315 ;
  assign n15317 = n13775 ^ n10029 ^ n8415 ;
  assign n15318 = n11424 ^ n7303 ^ n2466 ;
  assign n15319 = n12085 & n15318 ;
  assign n15320 = ( n4589 & n15317 ) | ( n4589 & ~n15319 ) | ( n15317 & ~n15319 ) ;
  assign n15321 = ( n2938 & n4835 ) | ( n2938 & ~n7044 ) | ( n4835 & ~n7044 ) ;
  assign n15322 = n13844 & n14401 ;
  assign n15323 = ~n9909 & n15322 ;
  assign n15324 = n11541 ^ n8089 ^ n7990 ;
  assign n15325 = n2267 ^ n2172 ^ x51 ;
  assign n15326 = n15325 ^ n12655 ^ n1515 ;
  assign n15327 = ( n15323 & n15324 ) | ( n15323 & ~n15326 ) | ( n15324 & ~n15326 ) ;
  assign n15336 = ( n722 & n4622 ) | ( n722 & n5196 ) | ( n4622 & n5196 ) ;
  assign n15334 = n1207 | n7382 ;
  assign n15335 = n8538 & ~n15334 ;
  assign n15337 = n15336 ^ n15335 ^ 1'b0 ;
  assign n15338 = n15337 ^ n6750 ^ 1'b0 ;
  assign n15339 = n9185 & ~n15338 ;
  assign n15328 = n6922 ^ n3575 ^ n1460 ;
  assign n15329 = ~n2638 & n15328 ;
  assign n15330 = n15329 ^ n575 ^ 1'b0 ;
  assign n15331 = ( n1056 & n12348 ) | ( n1056 & ~n15330 ) | ( n12348 & ~n15330 ) ;
  assign n15332 = ~n4797 & n15331 ;
  assign n15333 = n10829 & n15332 ;
  assign n15340 = n15339 ^ n15333 ^ n6135 ;
  assign n15341 = ( n2973 & n5249 ) | ( n2973 & ~n13930 ) | ( n5249 & ~n13930 ) ;
  assign n15345 = n6842 ^ n6288 ^ x28 ;
  assign n15346 = ( n1596 & n1788 ) | ( n1596 & ~n3803 ) | ( n1788 & ~n3803 ) ;
  assign n15347 = n15346 ^ n11666 ^ n9434 ;
  assign n15348 = ( n6891 & n15345 ) | ( n6891 & n15347 ) | ( n15345 & n15347 ) ;
  assign n15342 = ~n3919 & n11520 ;
  assign n15343 = ~n1438 & n15342 ;
  assign n15344 = n15343 ^ n12580 ^ n5023 ;
  assign n15349 = n15348 ^ n15344 ^ n13542 ;
  assign n15350 = n5149 ^ n2064 ^ 1'b0 ;
  assign n15351 = n7063 & n15350 ;
  assign n15352 = ( n2846 & n4329 ) | ( n2846 & n8430 ) | ( n4329 & n8430 ) ;
  assign n15353 = n15352 ^ n2186 ^ n994 ;
  assign n15354 = ( n2819 & n6450 ) | ( n2819 & ~n15353 ) | ( n6450 & ~n15353 ) ;
  assign n15355 = n15354 ^ n8642 ^ x107 ;
  assign n15356 = n1581 & n5316 ;
  assign n15357 = ~n8348 & n15356 ;
  assign n15358 = ( n6040 & ~n15283 ) | ( n6040 & n15357 ) | ( ~n15283 & n15357 ) ;
  assign n15359 = n14958 | n15358 ;
  assign n15360 = n12146 ^ n11319 ^ n5454 ;
  assign n15361 = ( ~n1786 & n3704 ) | ( ~n1786 & n15360 ) | ( n3704 & n15360 ) ;
  assign n15362 = n249 & ~n10673 ;
  assign n15365 = ( n1431 & ~n2833 ) | ( n1431 & n3797 ) | ( ~n2833 & n3797 ) ;
  assign n15363 = ( n1941 & ~n3011 ) | ( n1941 & n14082 ) | ( ~n3011 & n14082 ) ;
  assign n15364 = n15363 ^ n14682 ^ n838 ;
  assign n15366 = n15365 ^ n15364 ^ n5950 ;
  assign n15367 = n15366 ^ n8400 ^ n2908 ;
  assign n15368 = n8288 ^ n5218 ^ n4191 ;
  assign n15369 = ( ~n1080 & n12769 ) | ( ~n1080 & n13820 ) | ( n12769 & n13820 ) ;
  assign n15370 = n6651 ^ n4627 ^ n3809 ;
  assign n15371 = n15370 ^ n8250 ^ 1'b0 ;
  assign n15372 = ( ~n1353 & n6993 ) | ( ~n1353 & n15371 ) | ( n6993 & n15371 ) ;
  assign n15373 = n15372 ^ n10347 ^ n6227 ;
  assign n15374 = n11430 ^ n9450 ^ n2004 ;
  assign n15375 = n15374 ^ n14361 ^ n6170 ;
  assign n15376 = n11979 | n15375 ;
  assign n15377 = n15376 ^ n9552 ^ 1'b0 ;
  assign n15378 = n4203 & ~n15377 ;
  assign n15379 = ~n4306 & n15378 ;
  assign n15380 = n2507 ^ n1945 ^ n1662 ;
  assign n15381 = n3772 & ~n4399 ;
  assign n15382 = ~n258 & n15381 ;
  assign n15383 = ( n8016 & ~n10410 ) | ( n8016 & n15382 ) | ( ~n10410 & n15382 ) ;
  assign n15384 = ( n13895 & ~n15380 ) | ( n13895 & n15383 ) | ( ~n15380 & n15383 ) ;
  assign n15385 = ( ~n6598 & n9987 ) | ( ~n6598 & n10746 ) | ( n9987 & n10746 ) ;
  assign n15386 = n8703 ^ n5257 ^ n3929 ;
  assign n15387 = ( n8980 & ~n12928 ) | ( n8980 & n15386 ) | ( ~n12928 & n15386 ) ;
  assign n15389 = n9122 ^ n8764 ^ n6494 ;
  assign n15388 = x85 & ~n2424 ;
  assign n15390 = n15389 ^ n15388 ^ 1'b0 ;
  assign n15391 = ( n1541 & n10374 ) | ( n1541 & ~n15390 ) | ( n10374 & ~n15390 ) ;
  assign n15392 = ( ~n7624 & n9930 ) | ( ~n7624 & n14379 ) | ( n9930 & n14379 ) ;
  assign n15393 = n10482 & ~n13297 ;
  assign n15394 = n15393 ^ n4645 ^ 1'b0 ;
  assign n15395 = n15394 ^ n12591 ^ n7013 ;
  assign n15396 = ( n2010 & n4180 ) | ( n2010 & ~n11901 ) | ( n4180 & ~n11901 ) ;
  assign n15397 = n1460 | n15396 ;
  assign n15398 = n8006 | n15397 ;
  assign n15399 = n15398 ^ n10282 ^ n4817 ;
  assign n15400 = ( ~n4853 & n15395 ) | ( ~n4853 & n15399 ) | ( n15395 & n15399 ) ;
  assign n15401 = n5376 & n13578 ;
  assign n15402 = n15401 ^ n12092 ^ 1'b0 ;
  assign n15403 = n15402 ^ n11769 ^ n5128 ;
  assign n15408 = ( n462 & n6333 ) | ( n462 & n10947 ) | ( n6333 & n10947 ) ;
  assign n15404 = n12252 ^ n6924 ^ n4245 ;
  assign n15405 = ( ~n3007 & n6423 ) | ( ~n3007 & n13244 ) | ( n6423 & n13244 ) ;
  assign n15406 = ( n7249 & n15404 ) | ( n7249 & ~n15405 ) | ( n15404 & ~n15405 ) ;
  assign n15407 = n15406 ^ n12429 ^ n5533 ;
  assign n15409 = n15408 ^ n15407 ^ n12528 ;
  assign n15410 = ( ~n4297 & n5992 ) | ( ~n4297 & n6905 ) | ( n5992 & n6905 ) ;
  assign n15411 = n9562 ^ n2505 ^ 1'b0 ;
  assign n15412 = n6211 & ~n12469 ;
  assign n15413 = n1991 & ~n10874 ;
  assign n15414 = n2993 | n12734 ;
  assign n15415 = n15414 ^ n14559 ^ n1659 ;
  assign n15416 = ( n3204 & n6347 ) | ( n3204 & ~n7926 ) | ( n6347 & ~n7926 ) ;
  assign n15417 = n15416 ^ n3828 ^ n3297 ;
  assign n15418 = n11894 ^ n3972 ^ 1'b0 ;
  assign n15419 = ~n15417 & n15418 ;
  assign n15420 = ( n2428 & n3617 ) | ( n2428 & n15419 ) | ( n3617 & n15419 ) ;
  assign n15421 = n15185 ^ n7349 ^ n834 ;
  assign n15424 = ( x107 & n835 ) | ( x107 & n1377 ) | ( n835 & n1377 ) ;
  assign n15422 = ( n6122 & n12096 ) | ( n6122 & n15348 ) | ( n12096 & n15348 ) ;
  assign n15423 = ( n685 & ~n8974 ) | ( n685 & n15422 ) | ( ~n8974 & n15422 ) ;
  assign n15425 = n15424 ^ n15423 ^ n1374 ;
  assign n15431 = n3987 | n10630 ;
  assign n15432 = n15431 ^ n13251 ^ n6886 ;
  assign n15429 = n15055 ^ n12369 ^ n8397 ;
  assign n15426 = n8093 ^ n6026 ^ n5051 ;
  assign n15427 = n10595 & ~n15426 ;
  assign n15428 = n15427 ^ n4863 ^ 1'b0 ;
  assign n15430 = n15429 ^ n15428 ^ n11609 ;
  assign n15433 = n15432 ^ n15430 ^ 1'b0 ;
  assign n15434 = ( n357 & n801 ) | ( n357 & n10596 ) | ( n801 & n10596 ) ;
  assign n15435 = n15434 ^ n12459 ^ n1055 ;
  assign n15436 = n15435 ^ n3319 ^ n1941 ;
  assign n15437 = ( ~n2293 & n12258 ) | ( ~n2293 & n14493 ) | ( n12258 & n14493 ) ;
  assign n15438 = ( n14942 & n15436 ) | ( n14942 & n15437 ) | ( n15436 & n15437 ) ;
  assign n15439 = ( n3626 & n3734 ) | ( n3626 & ~n8483 ) | ( n3734 & ~n8483 ) ;
  assign n15440 = ( n739 & n12247 ) | ( n739 & ~n15439 ) | ( n12247 & ~n15439 ) ;
  assign n15441 = n5155 & n7323 ;
  assign n15442 = n15441 ^ n2770 ^ 1'b0 ;
  assign n15443 = n15442 ^ n6326 ^ n528 ;
  assign n15444 = n13653 ^ n704 ^ 1'b0 ;
  assign n15445 = n6764 | n15444 ;
  assign n15446 = n1437 | n15445 ;
  assign n15447 = n15443 & n15446 ;
  assign n15448 = ( n1896 & n3053 ) | ( n1896 & n4760 ) | ( n3053 & n4760 ) ;
  assign n15449 = n15448 ^ n4433 ^ n3374 ;
  assign n15450 = n15449 ^ n6579 ^ 1'b0 ;
  assign n15451 = ~n1391 & n15450 ;
  assign n15452 = ~n8242 & n15451 ;
  assign n15453 = n569 & n15452 ;
  assign n15457 = n2544 ^ n847 ^ 1'b0 ;
  assign n15458 = n6787 | n15457 ;
  assign n15459 = n15458 ^ n9495 ^ n6315 ;
  assign n15454 = ( n4334 & n10541 ) | ( n4334 & n14035 ) | ( n10541 & n14035 ) ;
  assign n15455 = n3728 ^ n2708 ^ n522 ;
  assign n15456 = ( n13943 & n15454 ) | ( n13943 & n15455 ) | ( n15454 & n15455 ) ;
  assign n15460 = n15459 ^ n15456 ^ n12414 ;
  assign n15461 = ( n2744 & n3885 ) | ( n2744 & ~n12562 ) | ( n3885 & ~n12562 ) ;
  assign n15462 = ( n1997 & n3194 ) | ( n1997 & ~n15461 ) | ( n3194 & ~n15461 ) ;
  assign n15463 = ( ~x125 & n2899 ) | ( ~x125 & n10295 ) | ( n2899 & n10295 ) ;
  assign n15464 = ( n354 & n4820 ) | ( n354 & ~n15463 ) | ( n4820 & ~n15463 ) ;
  assign n15465 = ( ~n8446 & n8715 ) | ( ~n8446 & n15464 ) | ( n8715 & n15464 ) ;
  assign n15466 = n3640 & n15465 ;
  assign n15467 = ( n2104 & n6870 ) | ( n2104 & ~n15466 ) | ( n6870 & ~n15466 ) ;
  assign n15468 = n11458 ^ n10107 ^ n924 ;
  assign n15469 = n15468 ^ n9790 ^ n1901 ;
  assign n15470 = ( n777 & ~n8862 ) | ( n777 & n12655 ) | ( ~n8862 & n12655 ) ;
  assign n15471 = n6114 & n15470 ;
  assign n15474 = n3639 ^ n2986 ^ n2831 ;
  assign n15475 = ~n3384 & n15474 ;
  assign n15476 = n15475 ^ n2834 ^ 1'b0 ;
  assign n15477 = n15476 ^ n4097 ^ 1'b0 ;
  assign n15478 = n5103 ^ n4129 ^ n2871 ;
  assign n15479 = n15478 ^ n8482 ^ n221 ;
  assign n15480 = ( n1151 & n15477 ) | ( n1151 & n15479 ) | ( n15477 & n15479 ) ;
  assign n15472 = n12743 ^ n5381 ^ n5362 ;
  assign n15473 = n15472 ^ n9859 ^ n6650 ;
  assign n15481 = n15480 ^ n15473 ^ n15464 ;
  assign n15482 = n12604 ^ n10657 ^ n9695 ;
  assign n15483 = ( n2620 & ~n7378 ) | ( n2620 & n7522 ) | ( ~n7378 & n7522 ) ;
  assign n15484 = ( ~n1316 & n1400 ) | ( ~n1316 & n3713 ) | ( n1400 & n3713 ) ;
  assign n15485 = n15484 ^ n10281 ^ n3236 ;
  assign n15486 = n7125 & n8288 ;
  assign n15487 = n15486 ^ n11560 ^ 1'b0 ;
  assign n15488 = ( x26 & n10013 ) | ( x26 & ~n12039 ) | ( n10013 & ~n12039 ) ;
  assign n15489 = n15488 ^ n333 ^ 1'b0 ;
  assign n15490 = n15246 ^ n5433 ^ n3070 ;
  assign n15491 = ( n3159 & ~n8182 ) | ( n3159 & n11552 ) | ( ~n8182 & n11552 ) ;
  assign n15492 = ( n2847 & n4790 ) | ( n2847 & n11050 ) | ( n4790 & n11050 ) ;
  assign n15494 = ( n1446 & ~n7324 ) | ( n1446 & n8938 ) | ( ~n7324 & n8938 ) ;
  assign n15495 = n15494 ^ n7030 ^ n5373 ;
  assign n15493 = ( n4275 & n6079 ) | ( n4275 & n14502 ) | ( n6079 & n14502 ) ;
  assign n15496 = n15495 ^ n15493 ^ n2262 ;
  assign n15497 = n15496 ^ n9043 ^ n9007 ;
  assign n15498 = n9504 ^ n870 ^ 1'b0 ;
  assign n15499 = n686 | n15498 ;
  assign n15500 = n915 & ~n6509 ;
  assign n15501 = ( ~n2572 & n6247 ) | ( ~n2572 & n15500 ) | ( n6247 & n15500 ) ;
  assign n15502 = n11807 ^ n6802 ^ n5437 ;
  assign n15503 = ~n6263 & n15502 ;
  assign n15504 = ( n5597 & n11412 ) | ( n5597 & ~n12851 ) | ( n11412 & ~n12851 ) ;
  assign n15505 = n4999 & n15504 ;
  assign n15506 = ~n5400 & n15505 ;
  assign n15507 = ( ~n679 & n13316 ) | ( ~n679 & n15506 ) | ( n13316 & n15506 ) ;
  assign n15508 = ~n8784 & n11460 ;
  assign n15509 = ( n6041 & n7685 ) | ( n6041 & ~n9339 ) | ( n7685 & ~n9339 ) ;
  assign n15510 = ( n285 & ~n9885 ) | ( n285 & n13727 ) | ( ~n9885 & n13727 ) ;
  assign n15511 = n10426 ^ n8422 ^ 1'b0 ;
  assign n15512 = n15510 | n15511 ;
  assign n15513 = n1790 | n1916 ;
  assign n15525 = n8355 ^ n3987 ^ n1337 ;
  assign n15516 = n5504 ^ n164 ^ 1'b0 ;
  assign n15517 = ( n2029 & ~n3378 ) | ( n2029 & n15516 ) | ( ~n3378 & n15516 ) ;
  assign n15518 = n3850 & ~n15517 ;
  assign n15519 = ( ~n624 & n3715 ) | ( ~n624 & n15518 ) | ( n3715 & n15518 ) ;
  assign n15520 = ( ~n3593 & n10458 ) | ( ~n3593 & n15519 ) | ( n10458 & n15519 ) ;
  assign n15521 = n8197 | n10127 ;
  assign n15522 = n15520 | n15521 ;
  assign n15514 = n5434 & ~n13858 ;
  assign n15515 = ( n1126 & n4898 ) | ( n1126 & ~n15514 ) | ( n4898 & ~n15514 ) ;
  assign n15523 = n15522 ^ n15515 ^ n7454 ;
  assign n15524 = n15523 ^ n15510 ^ n9609 ;
  assign n15526 = n15525 ^ n15524 ^ n1157 ;
  assign n15527 = ( ~n1274 & n15513 ) | ( ~n1274 & n15526 ) | ( n15513 & n15526 ) ;
  assign n15528 = ( x115 & n2444 ) | ( x115 & n3241 ) | ( n2444 & n3241 ) ;
  assign n15529 = n9528 ^ n7781 ^ n1742 ;
  assign n15530 = n15529 ^ n13187 ^ n594 ;
  assign n15531 = ( n8035 & ~n15528 ) | ( n8035 & n15530 ) | ( ~n15528 & n15530 ) ;
  assign n15532 = n15531 ^ n8420 ^ n2505 ;
  assign n15533 = n5079 ^ n4569 ^ n2122 ;
  assign n15534 = n15533 ^ n9257 ^ n3938 ;
  assign n15535 = n15534 ^ n9257 ^ n4978 ;
  assign n15536 = ( n11881 & n12481 ) | ( n11881 & ~n15535 ) | ( n12481 & ~n15535 ) ;
  assign n15537 = n15536 ^ n11063 ^ n7074 ;
  assign n15538 = n14123 ^ n10946 ^ n6053 ;
  assign n15542 = n4327 ^ n2318 ^ 1'b0 ;
  assign n15541 = n12576 ^ n6588 ^ n5196 ;
  assign n15539 = n3788 & ~n13360 ;
  assign n15540 = n417 & n15539 ;
  assign n15543 = n15542 ^ n15541 ^ n15540 ;
  assign n15545 = ( ~n2158 & n2622 ) | ( ~n2158 & n6743 ) | ( n2622 & n6743 ) ;
  assign n15544 = ~n6399 & n6992 ;
  assign n15546 = n15545 ^ n15544 ^ n1480 ;
  assign n15547 = ( n1394 & n3984 ) | ( n1394 & n5303 ) | ( n3984 & n5303 ) ;
  assign n15548 = n15547 ^ n12037 ^ n3274 ;
  assign n15549 = ~n3419 & n6650 ;
  assign n15550 = ( ~n2406 & n15548 ) | ( ~n2406 & n15549 ) | ( n15548 & n15549 ) ;
  assign n15551 = n5367 ^ n3970 ^ n3414 ;
  assign n15552 = n13688 ^ n12939 ^ x111 ;
  assign n15553 = ~n164 & n15552 ;
  assign n15559 = n9461 ^ n9182 ^ n4161 ;
  assign n15555 = n710 & ~n11847 ;
  assign n15556 = n1235 | n13259 ;
  assign n15557 = n15555 & ~n15556 ;
  assign n15558 = n15557 ^ n11970 ^ n5983 ;
  assign n15560 = n15559 ^ n15558 ^ n11017 ;
  assign n15554 = n7431 ^ n4351 ^ n3853 ;
  assign n15561 = n15560 ^ n15554 ^ n12344 ;
  assign n15562 = ( n15551 & ~n15553 ) | ( n15551 & n15561 ) | ( ~n15553 & n15561 ) ;
  assign n15563 = ( n10708 & ~n12388 ) | ( n10708 & n14143 ) | ( ~n12388 & n14143 ) ;
  assign n15564 = n7124 ^ n5864 ^ n5701 ;
  assign n15565 = n7966 ^ n4173 ^ n3199 ;
  assign n15566 = ( x48 & n2522 ) | ( x48 & n2700 ) | ( n2522 & n2700 ) ;
  assign n15567 = ( ~n4891 & n15565 ) | ( ~n4891 & n15566 ) | ( n15565 & n15566 ) ;
  assign n15568 = x125 & n9881 ;
  assign n15569 = n13627 & n15568 ;
  assign n15570 = ( n1703 & n4832 ) | ( n1703 & ~n15569 ) | ( n4832 & ~n15569 ) ;
  assign n15571 = ( n6044 & ~n7236 ) | ( n6044 & n15570 ) | ( ~n7236 & n15570 ) ;
  assign n15572 = ( n1270 & n8382 ) | ( n1270 & n11540 ) | ( n8382 & n11540 ) ;
  assign n15573 = n11048 | n15480 ;
  assign n15574 = n12633 ^ n9990 ^ n3853 ;
  assign n15575 = n12463 ^ n9811 ^ n8596 ;
  assign n15576 = n11068 ^ n10766 ^ n8639 ;
  assign n15577 = ( n15574 & n15575 ) | ( n15574 & n15576 ) | ( n15575 & n15576 ) ;
  assign n15579 = ( ~n1240 & n2520 ) | ( ~n1240 & n12676 ) | ( n2520 & n12676 ) ;
  assign n15578 = ( n4861 & n9658 ) | ( n4861 & n13493 ) | ( n9658 & n13493 ) ;
  assign n15580 = n15579 ^ n15578 ^ n6502 ;
  assign n15585 = ( n3695 & n3817 ) | ( n3695 & ~n12923 ) | ( n3817 & ~n12923 ) ;
  assign n15583 = ( ~n1953 & n4130 ) | ( ~n1953 & n8046 ) | ( n4130 & n8046 ) ;
  assign n15581 = n1757 ^ n687 ^ x12 ;
  assign n15582 = ( ~n9512 & n13605 ) | ( ~n9512 & n15581 ) | ( n13605 & n15581 ) ;
  assign n15584 = n15583 ^ n15582 ^ n2408 ;
  assign n15586 = n15585 ^ n15584 ^ n5274 ;
  assign n15587 = n14713 ^ n9316 ^ n5301 ;
  assign n15588 = n15587 ^ n12109 ^ 1'b0 ;
  assign n15589 = ~x86 & n15588 ;
  assign n15590 = n15589 ^ n7262 ^ n2460 ;
  assign n15591 = n5252 ^ n4231 ^ x99 ;
  assign n15592 = n15591 ^ n4866 ^ n4270 ;
  assign n15593 = n15590 & n15592 ;
  assign n15594 = n913 & n15593 ;
  assign n15595 = ( n3876 & n5940 ) | ( n3876 & ~n6455 ) | ( n5940 & ~n6455 ) ;
  assign n15596 = n15595 ^ n401 ^ 1'b0 ;
  assign n15597 = ( ~n3857 & n6998 ) | ( ~n3857 & n15596 ) | ( n6998 & n15596 ) ;
  assign n15598 = n15597 ^ n10702 ^ n9816 ;
  assign n15599 = ( n2098 & n2591 ) | ( n2098 & ~n15598 ) | ( n2591 & ~n15598 ) ;
  assign n15600 = ( ~n5531 & n6455 ) | ( ~n5531 & n7233 ) | ( n6455 & n7233 ) ;
  assign n15601 = n4857 & n7797 ;
  assign n15602 = n15601 ^ n12552 ^ 1'b0 ;
  assign n15603 = ( n2903 & ~n11714 ) | ( n2903 & n15602 ) | ( ~n11714 & n15602 ) ;
  assign n15604 = ( ~n1452 & n2501 ) | ( ~n1452 & n10760 ) | ( n2501 & n10760 ) ;
  assign n15605 = n15328 & n15604 ;
  assign n15606 = ~n9236 & n15605 ;
  assign n15607 = n15555 ^ n13626 ^ 1'b0 ;
  assign n15608 = ( ~n281 & n1042 ) | ( ~n281 & n7859 ) | ( n1042 & n7859 ) ;
  assign n15609 = ( ~n2446 & n5151 ) | ( ~n2446 & n15608 ) | ( n5151 & n15608 ) ;
  assign n15614 = n13627 ^ n9731 ^ n292 ;
  assign n15610 = n11569 ^ n1630 ^ n243 ;
  assign n15611 = n11088 ^ n7357 ^ n669 ;
  assign n15612 = n15611 ^ n15348 ^ n6861 ;
  assign n15613 = ( n4440 & ~n15610 ) | ( n4440 & n15612 ) | ( ~n15610 & n15612 ) ;
  assign n15615 = n15614 ^ n15613 ^ n2064 ;
  assign n15616 = n15615 ^ n13975 ^ n1476 ;
  assign n15622 = n14818 ^ n7156 ^ n4766 ;
  assign n15620 = ~n2640 & n6120 ;
  assign n15621 = n15620 ^ n3172 ^ 1'b0 ;
  assign n15623 = n15622 ^ n15621 ^ n939 ;
  assign n15617 = n791 | n817 ;
  assign n15618 = n15617 ^ n5035 ^ n558 ;
  assign n15619 = n15618 ^ n6050 ^ n4614 ;
  assign n15624 = n15623 ^ n15619 ^ n8274 ;
  assign n15625 = ( n6127 & n6962 ) | ( n6127 & ~n12889 ) | ( n6962 & ~n12889 ) ;
  assign n15626 = n15625 ^ n8869 ^ 1'b0 ;
  assign n15637 = ( n1765 & ~n3748 ) | ( n1765 & n4742 ) | ( ~n3748 & n4742 ) ;
  assign n15638 = n15637 ^ n12402 ^ n950 ;
  assign n15634 = ( ~n2060 & n8187 ) | ( ~n2060 & n11460 ) | ( n8187 & n11460 ) ;
  assign n15635 = ( n151 & n6139 ) | ( n151 & ~n15634 ) | ( n6139 & ~n15634 ) ;
  assign n15636 = ( n6076 & ~n13520 ) | ( n6076 & n15635 ) | ( ~n13520 & n15635 ) ;
  assign n15631 = n1061 ^ n773 ^ n730 ;
  assign n15629 = n10750 ^ n3859 ^ 1'b0 ;
  assign n15630 = n13635 | n15629 ;
  assign n15627 = n1896 & ~n13881 ;
  assign n15628 = ~n8867 & n15627 ;
  assign n15632 = n15631 ^ n15630 ^ n15628 ;
  assign n15633 = n15632 ^ n2428 ^ n243 ;
  assign n15639 = n15638 ^ n15636 ^ n15633 ;
  assign n15640 = ( ~n1153 & n6479 ) | ( ~n1153 & n14212 ) | ( n6479 & n14212 ) ;
  assign n15641 = n8550 & n15640 ;
  assign n15642 = n15641 ^ n7616 ^ 1'b0 ;
  assign n15643 = n15642 ^ n286 ^ 1'b0 ;
  assign n15644 = n7934 & n15643 ;
  assign n15645 = n1953 | n6166 ;
  assign n15646 = n15645 ^ n3644 ^ 1'b0 ;
  assign n15657 = ( ~n6633 & n7088 ) | ( ~n6633 & n9517 ) | ( n7088 & n9517 ) ;
  assign n15656 = n7717 ^ n5589 ^ n845 ;
  assign n15658 = n15657 ^ n15656 ^ n3194 ;
  assign n15659 = n15658 ^ n13940 ^ n12614 ;
  assign n15655 = n8249 ^ n7530 ^ 1'b0 ;
  assign n15650 = n7932 ^ n1744 ^ n815 ;
  assign n15647 = n4075 ^ n3249 ^ x3 ;
  assign n15648 = ~n3636 & n5161 ;
  assign n15649 = ( ~n1737 & n15647 ) | ( ~n1737 & n15648 ) | ( n15647 & n15648 ) ;
  assign n15651 = n15650 ^ n15649 ^ n8943 ;
  assign n15652 = ( n4006 & n5559 ) | ( n4006 & n8770 ) | ( n5559 & n8770 ) ;
  assign n15653 = ( n2342 & ~n6290 ) | ( n2342 & n15652 ) | ( ~n6290 & n15652 ) ;
  assign n15654 = ( n1164 & n15651 ) | ( n1164 & ~n15653 ) | ( n15651 & ~n15653 ) ;
  assign n15660 = n15659 ^ n15655 ^ n15654 ;
  assign n15661 = ( ~n4848 & n10025 ) | ( ~n4848 & n10613 ) | ( n10025 & n10613 ) ;
  assign n15662 = n15661 ^ n5133 ^ n4434 ;
  assign n15663 = n5384 ^ n4554 ^ n2178 ;
  assign n15664 = ( n707 & n13591 ) | ( n707 & ~n15663 ) | ( n13591 & ~n15663 ) ;
  assign n15665 = n15664 ^ n8150 ^ n3112 ;
  assign n15666 = n12350 ^ n11316 ^ n4476 ;
  assign n15667 = n15666 ^ n11124 ^ n9639 ;
  assign n15668 = ( ~n6594 & n15665 ) | ( ~n6594 & n15667 ) | ( n15665 & n15667 ) ;
  assign n15669 = ( x8 & n721 ) | ( x8 & n4812 ) | ( n721 & n4812 ) ;
  assign n15674 = n582 & ~n2899 ;
  assign n15675 = n15674 ^ n4396 ^ 1'b0 ;
  assign n15676 = n15675 ^ n11970 ^ n2344 ;
  assign n15671 = n1446 | n2793 ;
  assign n15672 = n6521 | n15671 ;
  assign n15670 = n3867 ^ n1551 ^ n1361 ;
  assign n15673 = n15672 ^ n15670 ^ n4967 ;
  assign n15677 = n15676 ^ n15673 ^ n4960 ;
  assign n15678 = n15677 ^ n5091 ^ 1'b0 ;
  assign n15679 = n15669 & ~n15678 ;
  assign n15683 = ( n611 & ~n3260 ) | ( n611 & n9278 ) | ( ~n3260 & n9278 ) ;
  assign n15684 = n15683 ^ n5997 ^ n3208 ;
  assign n15680 = n12636 ^ n8702 ^ n175 ;
  assign n15681 = n15680 ^ n8147 ^ n2022 ;
  assign n15682 = ( n2542 & n12177 ) | ( n2542 & n15681 ) | ( n12177 & n15681 ) ;
  assign n15685 = n15684 ^ n15682 ^ n14384 ;
  assign n15686 = ( n2791 & n13160 ) | ( n2791 & n14874 ) | ( n13160 & n14874 ) ;
  assign n15689 = n9658 ^ n8594 ^ n8020 ;
  assign n15687 = ~n840 & n14288 ;
  assign n15688 = n1635 & n15687 ;
  assign n15690 = n15689 ^ n15688 ^ n9874 ;
  assign n15691 = n5287 ^ n2967 ^ 1'b0 ;
  assign n15692 = n11147 ^ n5615 ^ n1368 ;
  assign n15693 = ( n11695 & n11907 ) | ( n11695 & n15692 ) | ( n11907 & n15692 ) ;
  assign n15694 = n15432 ^ n1527 ^ 1'b0 ;
  assign n15695 = n15694 ^ n7695 ^ n3709 ;
  assign n15703 = n5022 ^ n3028 ^ n1869 ;
  assign n15699 = n2845 & n11894 ;
  assign n15700 = n5861 & n15699 ;
  assign n15701 = n11264 & ~n15700 ;
  assign n15702 = n15701 ^ n13919 ^ n7172 ;
  assign n15696 = ( n390 & n1718 ) | ( n390 & ~n8482 ) | ( n1718 & ~n8482 ) ;
  assign n15697 = ( ~n8394 & n11963 ) | ( ~n8394 & n15696 ) | ( n11963 & n15696 ) ;
  assign n15698 = n7910 & n15697 ;
  assign n15704 = n15703 ^ n15702 ^ n15698 ;
  assign n15705 = n13842 ^ n9101 ^ n9051 ;
  assign n15706 = ( n1411 & ~n4409 ) | ( n1411 & n5026 ) | ( ~n4409 & n5026 ) ;
  assign n15707 = n7055 ^ n6674 ^ n1652 ;
  assign n15708 = n15707 ^ n15105 ^ n5052 ;
  assign n15709 = n11760 ^ n6374 ^ n3138 ;
  assign n15710 = ( n15162 & n15708 ) | ( n15162 & ~n15709 ) | ( n15708 & ~n15709 ) ;
  assign n15711 = ( n4711 & n15706 ) | ( n4711 & n15710 ) | ( n15706 & n15710 ) ;
  assign n15712 = ( n8797 & ~n15705 ) | ( n8797 & n15711 ) | ( ~n15705 & n15711 ) ;
  assign n15713 = n3013 ^ n2771 ^ n2306 ;
  assign n15714 = n2427 & ~n15713 ;
  assign n15715 = ( n4833 & ~n12485 ) | ( n4833 & n15714 ) | ( ~n12485 & n15714 ) ;
  assign n15716 = n3774 | n15715 ;
  assign n15717 = n15648 ^ n9825 ^ n2253 ;
  assign n15719 = n647 ^ n358 ^ n249 ;
  assign n15720 = n15719 ^ n8938 ^ n5414 ;
  assign n15718 = ( n339 & n6866 ) | ( n339 & ~n9658 ) | ( n6866 & ~n9658 ) ;
  assign n15721 = n15720 ^ n15718 ^ n11335 ;
  assign n15722 = ( ~n480 & n1213 ) | ( ~n480 & n1663 ) | ( n1213 & n1663 ) ;
  assign n15723 = n15722 ^ n12493 ^ n2400 ;
  assign n15726 = n12171 ^ n7966 ^ 1'b0 ;
  assign n15724 = n7723 ^ n4643 ^ n3934 ;
  assign n15725 = n13390 | n15724 ;
  assign n15727 = n15726 ^ n15725 ^ n7143 ;
  assign n15728 = n7580 ^ n4852 ^ 1'b0 ;
  assign n15729 = n4756 & n15728 ;
  assign n15730 = n1520 | n8566 ;
  assign n15731 = n10323 | n15730 ;
  assign n15740 = ( ~n5012 & n7210 ) | ( ~n5012 & n15123 ) | ( n7210 & n15123 ) ;
  assign n15736 = n11533 ^ n9441 ^ n1327 ;
  assign n15732 = ( n2124 & n4329 ) | ( n2124 & n6143 ) | ( n4329 & n6143 ) ;
  assign n15733 = n2870 | n3389 ;
  assign n15734 = ( n2457 & ~n15732 ) | ( n2457 & n15733 ) | ( ~n15732 & n15733 ) ;
  assign n15735 = n15734 ^ n990 ^ n792 ;
  assign n15737 = n15736 ^ n15735 ^ n10688 ;
  assign n15738 = n8598 | n10700 ;
  assign n15739 = n15737 & ~n15738 ;
  assign n15741 = n15740 ^ n15739 ^ n1868 ;
  assign n15742 = n7753 ^ n7604 ^ n5884 ;
  assign n15743 = n7808 ^ n6966 ^ n2587 ;
  assign n15744 = n1929 | n1947 ;
  assign n15745 = n15743 | n15744 ;
  assign n15748 = n2708 ^ n633 ^ 1'b0 ;
  assign n15749 = n15748 ^ n13045 ^ n7721 ;
  assign n15750 = n15749 ^ n8674 ^ 1'b0 ;
  assign n15751 = ~n881 & n15750 ;
  assign n15746 = ( n837 & ~n4429 ) | ( n837 & n5694 ) | ( ~n4429 & n5694 ) ;
  assign n15747 = ( n3570 & n4108 ) | ( n3570 & ~n15746 ) | ( n4108 & ~n15746 ) ;
  assign n15752 = n15751 ^ n15747 ^ n10750 ;
  assign n15753 = ( ~n15742 & n15745 ) | ( ~n15742 & n15752 ) | ( n15745 & n15752 ) ;
  assign n15754 = n15753 ^ n8623 ^ 1'b0 ;
  assign n15755 = ( n3446 & ~n4853 ) | ( n3446 & n11958 ) | ( ~n4853 & n11958 ) ;
  assign n15756 = n15755 ^ n3563 ^ n1116 ;
  assign n15757 = n13913 ^ n13776 ^ x111 ;
  assign n15758 = ( n991 & n4654 ) | ( n991 & ~n15757 ) | ( n4654 & ~n15757 ) ;
  assign n15759 = ( n1647 & n6401 ) | ( n1647 & ~n8097 ) | ( n6401 & ~n8097 ) ;
  assign n15760 = ( ~n7708 & n13443 ) | ( ~n7708 & n15759 ) | ( n13443 & n15759 ) ;
  assign n15761 = n10994 ^ n10006 ^ n1527 ;
  assign n15762 = n4010 ^ n1064 ^ n242 ;
  assign n15763 = ( n1450 & n5696 ) | ( n1450 & ~n15762 ) | ( n5696 & ~n15762 ) ;
  assign n15764 = ( n4488 & n6355 ) | ( n4488 & n13097 ) | ( n6355 & n13097 ) ;
  assign n15765 = n9505 ^ n5295 ^ n5197 ;
  assign n15766 = n11007 ^ n5359 ^ n1170 ;
  assign n15767 = ( n5371 & n7117 ) | ( n5371 & ~n15766 ) | ( n7117 & ~n15766 ) ;
  assign n15768 = n15767 ^ n7797 ^ n5106 ;
  assign n15771 = n5568 ^ n2583 ^ n1934 ;
  assign n15772 = ( ~n175 & n4362 ) | ( ~n175 & n15771 ) | ( n4362 & n15771 ) ;
  assign n15773 = ( n1628 & ~n9936 ) | ( n1628 & n15772 ) | ( ~n9936 & n15772 ) ;
  assign n15769 = n1331 | n5889 ;
  assign n15770 = n1240 & ~n15769 ;
  assign n15774 = n15773 ^ n15770 ^ n1146 ;
  assign n15775 = ( n751 & n2426 ) | ( n751 & n9894 ) | ( n2426 & n9894 ) ;
  assign n15776 = n15775 ^ n3920 ^ n1719 ;
  assign n15777 = n4304 & n5126 ;
  assign n15778 = ~n15776 & n15777 ;
  assign n15779 = ( n1727 & ~n1743 ) | ( n1727 & n6012 ) | ( ~n1743 & n6012 ) ;
  assign n15780 = ( ~n3352 & n4797 ) | ( ~n3352 & n15779 ) | ( n4797 & n15779 ) ;
  assign n15781 = ( n2301 & n15778 ) | ( n2301 & ~n15780 ) | ( n15778 & ~n15780 ) ;
  assign n15782 = ~n11147 & n12036 ;
  assign n15783 = ( n4152 & ~n8814 ) | ( n4152 & n14844 ) | ( ~n8814 & n14844 ) ;
  assign n15784 = n1137 | n3559 ;
  assign n15785 = n2286 | n15784 ;
  assign n15786 = n15785 ^ n11930 ^ n6330 ;
  assign n15787 = n1284 & ~n8884 ;
  assign n15788 = n10794 ^ n9247 ^ n3331 ;
  assign n15789 = ( n709 & n1429 ) | ( n709 & n4522 ) | ( n1429 & n4522 ) ;
  assign n15790 = n8187 ^ n6923 ^ 1'b0 ;
  assign n15791 = n3088 & n11013 ;
  assign n15792 = n15791 ^ n4869 ^ 1'b0 ;
  assign n15794 = ( ~n524 & n3864 ) | ( ~n524 & n11760 ) | ( n3864 & n11760 ) ;
  assign n15795 = n9461 & n15794 ;
  assign n15793 = ( n5039 & ~n11430 ) | ( n5039 & n15734 ) | ( ~n11430 & n15734 ) ;
  assign n15796 = n15795 ^ n15793 ^ 1'b0 ;
  assign n15797 = ( x81 & n2538 ) | ( x81 & ~n15796 ) | ( n2538 & ~n15796 ) ;
  assign n15798 = ( ~n1562 & n11440 ) | ( ~n1562 & n11941 ) | ( n11440 & n11941 ) ;
  assign n15799 = ( n5154 & ~n9772 ) | ( n5154 & n12019 ) | ( ~n9772 & n12019 ) ;
  assign n15800 = n8140 ^ n8072 ^ n7711 ;
  assign n15801 = ( ~n13600 & n14844 ) | ( ~n13600 & n15800 ) | ( n14844 & n15800 ) ;
  assign n15802 = ( ~n2522 & n15799 ) | ( ~n2522 & n15801 ) | ( n15799 & n15801 ) ;
  assign n15803 = n15802 ^ n11914 ^ n2416 ;
  assign n15804 = n12808 ^ n11371 ^ n10800 ;
  assign n15805 = ( n4314 & n11103 ) | ( n4314 & ~n15804 ) | ( n11103 & ~n15804 ) ;
  assign n15806 = n14028 ^ n6713 ^ n1197 ;
  assign n15807 = ~n644 & n8454 ;
  assign n15808 = ( n1449 & ~n1789 ) | ( n1449 & n6205 ) | ( ~n1789 & n6205 ) ;
  assign n15809 = n1860 ^ n1067 ^ 1'b0 ;
  assign n15810 = n614 | n15809 ;
  assign n15811 = n15810 ^ n10725 ^ n5331 ;
  assign n15812 = n15811 ^ n11225 ^ n8702 ;
  assign n15813 = n3559 | n15812 ;
  assign n15814 = n15808 & ~n15813 ;
  assign n15815 = ( n2241 & ~n15807 ) | ( n2241 & n15814 ) | ( ~n15807 & n15814 ) ;
  assign n15816 = ( n658 & ~n746 ) | ( n658 & n15174 ) | ( ~n746 & n15174 ) ;
  assign n15817 = n15816 ^ n9837 ^ n7087 ;
  assign n15818 = n5386 & n7858 ;
  assign n15819 = ( n5580 & n15817 ) | ( n5580 & n15818 ) | ( n15817 & n15818 ) ;
  assign n15820 = n13324 ^ n1565 ^ n716 ;
  assign n15821 = n15820 ^ n9694 ^ n1668 ;
  assign n15822 = n4547 & n6107 ;
  assign n15823 = n15822 ^ n10814 ^ 1'b0 ;
  assign n15824 = ~n15821 & n15823 ;
  assign n15825 = n2863 & ~n9966 ;
  assign n15826 = n15825 ^ n11542 ^ n2208 ;
  assign n15827 = ( ~n4349 & n8222 ) | ( ~n4349 & n15755 ) | ( n8222 & n15755 ) ;
  assign n15828 = ( n5913 & n7771 ) | ( n5913 & ~n15827 ) | ( n7771 & ~n15827 ) ;
  assign n15829 = n15828 ^ n13274 ^ n2079 ;
  assign n15830 = ( n2043 & ~n6624 ) | ( n2043 & n6698 ) | ( ~n6624 & n6698 ) ;
  assign n15831 = ( n7672 & n10199 ) | ( n7672 & n12720 ) | ( n10199 & n12720 ) ;
  assign n15832 = ( n6941 & n9568 ) | ( n6941 & n12809 ) | ( n9568 & n12809 ) ;
  assign n15833 = n15832 ^ n10085 ^ n1371 ;
  assign n15842 = n10874 ^ n3425 ^ 1'b0 ;
  assign n15843 = ( n6921 & n10929 ) | ( n6921 & ~n15842 ) | ( n10929 & ~n15842 ) ;
  assign n15834 = ( n1161 & ~n2347 ) | ( n1161 & n11944 ) | ( ~n2347 & n11944 ) ;
  assign n15835 = n15834 ^ n4955 ^ 1'b0 ;
  assign n15836 = n9330 & n15835 ;
  assign n15837 = ( ~n4278 & n12491 ) | ( ~n4278 & n15836 ) | ( n12491 & n15836 ) ;
  assign n15838 = n4477 & ~n15837 ;
  assign n15839 = n11614 ^ n8103 ^ n5885 ;
  assign n15840 = ( n1456 & n12019 ) | ( n1456 & n15839 ) | ( n12019 & n15839 ) ;
  assign n15841 = ( n8610 & n15838 ) | ( n8610 & n15840 ) | ( n15838 & n15840 ) ;
  assign n15844 = n15843 ^ n15841 ^ n4623 ;
  assign n15853 = n15555 ^ n5605 ^ n5189 ;
  assign n15851 = ( ~n1108 & n3632 ) | ( ~n1108 & n4640 ) | ( n3632 & n4640 ) ;
  assign n15852 = n15851 ^ n1474 ^ n900 ;
  assign n15846 = n7660 ^ n2917 ^ 1'b0 ;
  assign n15847 = n9054 | n15846 ;
  assign n15848 = n15847 ^ n8269 ^ n1086 ;
  assign n15845 = n7455 ^ n6378 ^ n3901 ;
  assign n15849 = n15848 ^ n15845 ^ n9310 ;
  assign n15850 = ( n4113 & n15814 ) | ( n4113 & ~n15849 ) | ( n15814 & ~n15849 ) ;
  assign n15854 = n15853 ^ n15852 ^ n15850 ;
  assign n15856 = n5985 | n8397 ;
  assign n15855 = n8548 ^ n5942 ^ n4816 ;
  assign n15857 = n15856 ^ n15855 ^ n14419 ;
  assign n15858 = n7676 ^ n2022 ^ n2004 ;
  assign n15859 = n211 & n15858 ;
  assign n15860 = n15859 ^ n744 ^ 1'b0 ;
  assign n15861 = n15650 ^ n8881 ^ 1'b0 ;
  assign n15864 = ( n4055 & n4201 ) | ( n4055 & ~n9554 ) | ( n4201 & ~n9554 ) ;
  assign n15863 = n6396 ^ n4474 ^ n3742 ;
  assign n15862 = ( ~n631 & n4591 ) | ( ~n631 & n7535 ) | ( n4591 & n7535 ) ;
  assign n15865 = n15864 ^ n15863 ^ n15862 ;
  assign n15866 = ( ~n380 & n3661 ) | ( ~n380 & n15865 ) | ( n3661 & n15865 ) ;
  assign n15867 = ( n6615 & n15861 ) | ( n6615 & n15866 ) | ( n15861 & n15866 ) ;
  assign n15868 = n8969 ^ n4414 ^ 1'b0 ;
  assign n15869 = ( ~x81 & n4943 ) | ( ~x81 & n15868 ) | ( n4943 & n15868 ) ;
  assign n15870 = n1650 ^ n1610 ^ n205 ;
  assign n15871 = ~n15810 & n15870 ;
  assign n15872 = ( n4020 & n6369 ) | ( n4020 & ~n12805 ) | ( n6369 & ~n12805 ) ;
  assign n15873 = n15872 ^ n13254 ^ 1'b0 ;
  assign n15874 = n15871 & n15873 ;
  assign n15875 = n3819 ^ n3742 ^ n2259 ;
  assign n15876 = ( n11103 & ~n11117 ) | ( n11103 & n15875 ) | ( ~n11117 & n15875 ) ;
  assign n15877 = ( n700 & n3821 ) | ( n700 & n14380 ) | ( n3821 & n14380 ) ;
  assign n15878 = ( n1939 & ~n2678 ) | ( n1939 & n5649 ) | ( ~n2678 & n5649 ) ;
  assign n15879 = n15878 ^ n2263 ^ n654 ;
  assign n15880 = n15879 ^ n7511 ^ n3417 ;
  assign n15881 = n14952 ^ n10505 ^ n3794 ;
  assign n15882 = ( n8253 & n15272 ) | ( n8253 & ~n15881 ) | ( n15272 & ~n15881 ) ;
  assign n15883 = ( n1878 & n15880 ) | ( n1878 & ~n15882 ) | ( n15880 & ~n15882 ) ;
  assign n15884 = ( n14813 & n15877 ) | ( n14813 & ~n15883 ) | ( n15877 & ~n15883 ) ;
  assign n15885 = ( n6060 & n9895 ) | ( n6060 & n15884 ) | ( n9895 & n15884 ) ;
  assign n15886 = n15876 | n15885 ;
  assign n15887 = n15886 ^ n5116 ^ 1'b0 ;
  assign n15888 = ( n10390 & ~n15874 ) | ( n10390 & n15887 ) | ( ~n15874 & n15887 ) ;
  assign n15891 = n3057 & n11355 ;
  assign n15892 = n15891 ^ n1291 ^ 1'b0 ;
  assign n15889 = ( n581 & ~n3198 ) | ( n581 & n5699 ) | ( ~n3198 & n5699 ) ;
  assign n15890 = ( n3351 & ~n7859 ) | ( n3351 & n15889 ) | ( ~n7859 & n15889 ) ;
  assign n15893 = n15892 ^ n15890 ^ 1'b0 ;
  assign n15894 = ( n6111 & ~n10307 ) | ( n6111 & n14920 ) | ( ~n10307 & n14920 ) ;
  assign n15895 = ( n6129 & n6395 ) | ( n6129 & n14484 ) | ( n6395 & n14484 ) ;
  assign n15896 = ( n7502 & n15894 ) | ( n7502 & n15895 ) | ( n15894 & n15895 ) ;
  assign n15897 = ( n3137 & n8320 ) | ( n3137 & ~n9118 ) | ( n8320 & ~n9118 ) ;
  assign n15898 = ( ~n10240 & n15055 ) | ( ~n10240 & n15897 ) | ( n15055 & n15897 ) ;
  assign n15899 = ( n7698 & ~n15896 ) | ( n7698 & n15898 ) | ( ~n15896 & n15898 ) ;
  assign n15900 = n14775 ^ n10929 ^ n3304 ;
  assign n15901 = ( n412 & ~n2088 ) | ( n412 & n5319 ) | ( ~n2088 & n5319 ) ;
  assign n15902 = n12917 ^ n4992 ^ n2000 ;
  assign n15903 = n1212 & n10567 ;
  assign n15904 = ( n599 & n9548 ) | ( n599 & n15903 ) | ( n9548 & n15903 ) ;
  assign n15905 = ( n15901 & n15902 ) | ( n15901 & n15904 ) | ( n15902 & n15904 ) ;
  assign n15906 = n15905 ^ n15044 ^ n7237 ;
  assign n15907 = n15208 ^ n7785 ^ 1'b0 ;
  assign n15908 = n15907 ^ n14331 ^ 1'b0 ;
  assign n15909 = n6557 & ~n15908 ;
  assign n15910 = n15909 ^ n6184 ^ n5933 ;
  assign n15911 = n15191 ^ n1401 ^ 1'b0 ;
  assign n15912 = n3971 | n15911 ;
  assign n15913 = n15912 ^ n11519 ^ 1'b0 ;
  assign n15914 = ( n7990 & n10883 ) | ( n7990 & ~n15913 ) | ( n10883 & ~n15913 ) ;
  assign n15915 = ( n1706 & n4238 ) | ( n1706 & n13582 ) | ( n4238 & n13582 ) ;
  assign n15916 = ( x101 & n10544 ) | ( x101 & n15915 ) | ( n10544 & n15915 ) ;
  assign n15917 = n6614 ^ n4563 ^ n2103 ;
  assign n15918 = n5937 ^ n5132 ^ n3306 ;
  assign n15919 = n5606 ^ n3919 ^ n1872 ;
  assign n15920 = ( n4965 & n8472 ) | ( n4965 & ~n15919 ) | ( n8472 & ~n15919 ) ;
  assign n15921 = ( x60 & n2459 ) | ( x60 & ~n2468 ) | ( n2459 & ~n2468 ) ;
  assign n15922 = n15921 ^ n10338 ^ n423 ;
  assign n15923 = n14030 ^ n13547 ^ n456 ;
  assign n15924 = n15923 ^ n2839 ^ n629 ;
  assign n15928 = n6459 ^ n5409 ^ n2814 ;
  assign n15929 = ( n3919 & ~n5078 ) | ( n3919 & n15928 ) | ( ~n5078 & n15928 ) ;
  assign n15925 = n8294 ^ n4730 ^ 1'b0 ;
  assign n15926 = n4846 & n15925 ;
  assign n15927 = ( n2345 & n7952 ) | ( n2345 & n15926 ) | ( n7952 & n15926 ) ;
  assign n15930 = n15929 ^ n15927 ^ n11917 ;
  assign n15931 = n6505 ^ n6075 ^ n3231 ;
  assign n15932 = ( n11018 & n15930 ) | ( n11018 & n15931 ) | ( n15930 & n15931 ) ;
  assign n15933 = n14206 ^ n10223 ^ n1550 ;
  assign n15934 = n15933 ^ n11939 ^ 1'b0 ;
  assign n15935 = n7186 & ~n15934 ;
  assign n15936 = n15935 ^ n12535 ^ n7536 ;
  assign n15937 = ( n3652 & n15932 ) | ( n3652 & ~n15936 ) | ( n15932 & ~n15936 ) ;
  assign n15938 = n15254 ^ n11017 ^ n6065 ;
  assign n15939 = ~n3643 & n9554 ;
  assign n15940 = n15939 ^ n6662 ^ 1'b0 ;
  assign n15941 = ( ~n4058 & n4993 ) | ( ~n4058 & n15940 ) | ( n4993 & n15940 ) ;
  assign n15942 = n7939 ^ n2054 ^ 1'b0 ;
  assign n15943 = n2519 & ~n12092 ;
  assign n15944 = ~n2194 & n15943 ;
  assign n15945 = ( n3734 & n15942 ) | ( n3734 & n15944 ) | ( n15942 & n15944 ) ;
  assign n15951 = n15825 ^ n1512 ^ n721 ;
  assign n15952 = n10655 ^ n3655 ^ n2704 ;
  assign n15953 = ( n272 & ~n6093 ) | ( n272 & n15952 ) | ( ~n6093 & n15952 ) ;
  assign n15954 = ( n6039 & n15951 ) | ( n6039 & ~n15953 ) | ( n15951 & ~n15953 ) ;
  assign n15955 = n15954 ^ n10527 ^ n610 ;
  assign n15946 = ~n290 & n3776 ;
  assign n15947 = n15946 ^ n219 ^ 1'b0 ;
  assign n15948 = ( n2574 & n4925 ) | ( n2574 & n15947 ) | ( n4925 & n15947 ) ;
  assign n15949 = ( n3264 & n4608 ) | ( n3264 & n8935 ) | ( n4608 & n8935 ) ;
  assign n15950 = ( n7938 & n15948 ) | ( n7938 & ~n15949 ) | ( n15948 & ~n15949 ) ;
  assign n15956 = n15955 ^ n15950 ^ n15795 ;
  assign n15957 = n10863 ^ n8624 ^ n1927 ;
  assign n15958 = ( n2731 & n15736 ) | ( n2731 & ~n15957 ) | ( n15736 & ~n15957 ) ;
  assign n15960 = n5566 ^ n4036 ^ n2701 ;
  assign n15959 = ( ~n4622 & n8403 ) | ( ~n4622 & n11604 ) | ( n8403 & n11604 ) ;
  assign n15961 = n15960 ^ n15959 ^ n819 ;
  assign n15966 = ( n1276 & n1461 ) | ( n1276 & n9435 ) | ( n1461 & n9435 ) ;
  assign n15967 = n15966 ^ n11305 ^ n9917 ;
  assign n15965 = n12267 ^ n10517 ^ n502 ;
  assign n15968 = n15967 ^ n15965 ^ n12475 ;
  assign n15962 = ~n543 & n4364 ;
  assign n15963 = n15962 ^ n1231 ^ 1'b0 ;
  assign n15964 = n8311 & ~n15963 ;
  assign n15969 = n15968 ^ n15964 ^ n5379 ;
  assign n15975 = ( n1617 & ~n1777 ) | ( n1617 & n15458 ) | ( ~n1777 & n15458 ) ;
  assign n15971 = ( n6864 & n9473 ) | ( n6864 & n10506 ) | ( n9473 & n10506 ) ;
  assign n15972 = n15971 ^ n5251 ^ n3677 ;
  assign n15973 = n1553 ^ n884 ^ 1'b0 ;
  assign n15974 = ( ~n664 & n15972 ) | ( ~n664 & n15973 ) | ( n15972 & n15973 ) ;
  assign n15970 = n8148 ^ n6262 ^ 1'b0 ;
  assign n15976 = n15975 ^ n15974 ^ n15970 ;
  assign n15977 = ( n3066 & n9232 ) | ( n3066 & ~n15132 ) | ( n9232 & ~n15132 ) ;
  assign n15978 = ( ~n9777 & n14990 ) | ( ~n9777 & n15977 ) | ( n14990 & n15977 ) ;
  assign n15979 = n8981 | n13340 ;
  assign n15980 = n5620 & ~n6537 ;
  assign n15981 = ( n4585 & n15979 ) | ( n4585 & ~n15980 ) | ( n15979 & ~n15980 ) ;
  assign n15982 = n6855 ^ n2549 ^ 1'b0 ;
  assign n15983 = ( n3351 & ~n10063 ) | ( n3351 & n15982 ) | ( ~n10063 & n15982 ) ;
  assign n15984 = n15983 ^ n7691 ^ 1'b0 ;
  assign n15985 = ( n1884 & n5495 ) | ( n1884 & n14884 ) | ( n5495 & n14884 ) ;
  assign n15986 = ( n3439 & ~n3905 ) | ( n3439 & n15985 ) | ( ~n3905 & n15985 ) ;
  assign n15987 = ( n8791 & n14426 ) | ( n8791 & ~n14760 ) | ( n14426 & ~n14760 ) ;
  assign n15988 = ~n15986 & n15987 ;
  assign n15989 = ~n2168 & n15988 ;
  assign n15990 = ( n2429 & ~n6963 ) | ( n2429 & n7248 ) | ( ~n6963 & n7248 ) ;
  assign n15991 = ( n2671 & n9447 ) | ( n2671 & n14978 ) | ( n9447 & n14978 ) ;
  assign n15993 = n4150 | n9575 ;
  assign n15994 = ( n2853 & n15494 ) | ( n2853 & ~n15993 ) | ( n15494 & ~n15993 ) ;
  assign n15992 = ~n1961 & n12491 ;
  assign n15995 = n15994 ^ n15992 ^ 1'b0 ;
  assign n15996 = n7059 & n7739 ;
  assign n15997 = ( n2195 & n3060 ) | ( n2195 & ~n4415 ) | ( n3060 & ~n4415 ) ;
  assign n15998 = ( n4354 & n13694 ) | ( n4354 & n15997 ) | ( n13694 & n15997 ) ;
  assign n15999 = ( ~n7292 & n9896 ) | ( ~n7292 & n15998 ) | ( n9896 & n15998 ) ;
  assign n16000 = ( n420 & ~n821 ) | ( n420 & n1840 ) | ( ~n821 & n1840 ) ;
  assign n16001 = n16000 ^ n3890 ^ 1'b0 ;
  assign n16002 = ( ~n3675 & n5183 ) | ( ~n3675 & n8463 ) | ( n5183 & n8463 ) ;
  assign n16003 = n16002 ^ n15977 ^ n6646 ;
  assign n16004 = ( n442 & n1934 ) | ( n442 & n4766 ) | ( n1934 & n4766 ) ;
  assign n16005 = n16004 ^ n5742 ^ n5169 ;
  assign n16006 = ( ~n218 & n879 ) | ( ~n218 & n6104 ) | ( n879 & n6104 ) ;
  assign n16007 = ( n1553 & ~n15707 ) | ( n1553 & n16006 ) | ( ~n15707 & n16006 ) ;
  assign n16008 = n16007 ^ n5949 ^ n4830 ;
  assign n16009 = ( n852 & ~n7522 ) | ( n852 & n16008 ) | ( ~n7522 & n16008 ) ;
  assign n16010 = n16009 ^ n1130 ^ 1'b0 ;
  assign n16011 = ~n3053 & n16010 ;
  assign n16012 = n9340 ^ n4050 ^ n448 ;
  assign n16013 = n16012 ^ n10828 ^ n7309 ;
  assign n16014 = n16013 ^ n8194 ^ n5491 ;
  assign n16015 = ( n1529 & n6143 ) | ( n1529 & ~n16014 ) | ( n6143 & ~n16014 ) ;
  assign n16016 = n14271 ^ n1729 ^ 1'b0 ;
  assign n16017 = n16015 & ~n16016 ;
  assign n16018 = n880 | n5119 ;
  assign n16019 = n5497 & ~n16018 ;
  assign n16020 = n237 & ~n16019 ;
  assign n16021 = n5805 ^ n3410 ^ n155 ;
  assign n16022 = ( ~n2592 & n4133 ) | ( ~n2592 & n5974 ) | ( n4133 & n5974 ) ;
  assign n16023 = n16022 ^ n1075 ^ n981 ;
  assign n16024 = ( n7644 & n16021 ) | ( n7644 & ~n16023 ) | ( n16021 & ~n16023 ) ;
  assign n16025 = ( n7708 & ~n16020 ) | ( n7708 & n16024 ) | ( ~n16020 & n16024 ) ;
  assign n16026 = n16025 ^ n10788 ^ n3528 ;
  assign n16027 = n13140 ^ n6188 ^ n3834 ;
  assign n16028 = ( n623 & n14061 ) | ( n623 & n16027 ) | ( n14061 & n16027 ) ;
  assign n16029 = n16028 ^ n15523 ^ n11250 ;
  assign n16030 = n4536 ^ n4015 ^ n698 ;
  assign n16031 = ( n735 & n8100 ) | ( n735 & ~n10630 ) | ( n8100 & ~n10630 ) ;
  assign n16032 = n6026 | n12321 ;
  assign n16033 = n16031 & ~n16032 ;
  assign n16034 = ( n6514 & n16030 ) | ( n6514 & ~n16033 ) | ( n16030 & ~n16033 ) ;
  assign n16035 = n10674 ^ n7598 ^ n411 ;
  assign n16036 = n16035 ^ n14690 ^ n4954 ;
  assign n16037 = n1388 & ~n11521 ;
  assign n16038 = ~n13046 & n16037 ;
  assign n16039 = ( n5834 & ~n6258 ) | ( n5834 & n14482 ) | ( ~n6258 & n14482 ) ;
  assign n16044 = ( n3537 & n4447 ) | ( n3537 & n9392 ) | ( n4447 & n9392 ) ;
  assign n16045 = ( n8162 & ~n13668 ) | ( n8162 & n16044 ) | ( ~n13668 & n16044 ) ;
  assign n16040 = ( n4602 & n5101 ) | ( n4602 & n11715 ) | ( n5101 & n11715 ) ;
  assign n16041 = ( n7273 & n14045 ) | ( n7273 & ~n16040 ) | ( n14045 & ~n16040 ) ;
  assign n16042 = n6729 | n16041 ;
  assign n16043 = n16042 ^ n10665 ^ n4833 ;
  assign n16046 = n16045 ^ n16043 ^ n3941 ;
  assign n16047 = n13316 ^ n6606 ^ n4597 ;
  assign n16048 = ( n2069 & n5669 ) | ( n2069 & ~n16047 ) | ( n5669 & ~n16047 ) ;
  assign n16049 = n6954 ^ n2613 ^ n1968 ;
  assign n16050 = n16049 ^ n9431 ^ 1'b0 ;
  assign n16052 = ( n2429 & n2552 ) | ( n2429 & ~n7797 ) | ( n2552 & ~n7797 ) ;
  assign n16053 = n14076 | n16052 ;
  assign n16054 = n6366 & ~n16053 ;
  assign n16051 = n5636 & ~n5852 ;
  assign n16055 = n16054 ^ n16051 ^ 1'b0 ;
  assign n16056 = n5882 ^ n3112 ^ n2247 ;
  assign n16057 = n16056 ^ n14817 ^ n6288 ;
  assign n16058 = ( n2563 & n3811 ) | ( n2563 & ~n16057 ) | ( n3811 & ~n16057 ) ;
  assign n16059 = ( n1304 & n16055 ) | ( n1304 & ~n16058 ) | ( n16055 & ~n16058 ) ;
  assign n16066 = n5313 ^ n3032 ^ 1'b0 ;
  assign n16063 = n4602 & n6189 ;
  assign n16064 = n16063 ^ n2737 ^ 1'b0 ;
  assign n16065 = n16064 ^ n7964 ^ n2935 ;
  assign n16060 = n6491 ^ n4362 ^ n3096 ;
  assign n16061 = ( ~n5188 & n14383 ) | ( ~n5188 & n16060 ) | ( n14383 & n16060 ) ;
  assign n16062 = ( n10355 & n13645 ) | ( n10355 & n16061 ) | ( n13645 & n16061 ) ;
  assign n16067 = n16066 ^ n16065 ^ n16062 ;
  assign n16068 = n8148 ^ n4372 ^ n4194 ;
  assign n16069 = ( n373 & n4746 ) | ( n373 & n16068 ) | ( n4746 & n16068 ) ;
  assign n16070 = n16069 ^ n10905 ^ n8539 ;
  assign n16071 = ( n5007 & ~n11799 ) | ( n5007 & n16070 ) | ( ~n11799 & n16070 ) ;
  assign n16073 = ( n408 & ~n7358 ) | ( n408 & n10203 ) | ( ~n7358 & n10203 ) ;
  assign n16072 = ( x26 & ~n6204 ) | ( x26 & n9173 ) | ( ~n6204 & n9173 ) ;
  assign n16074 = n16073 ^ n16072 ^ 1'b0 ;
  assign n16075 = n5137 & n11216 ;
  assign n16076 = ( ~n16071 & n16074 ) | ( ~n16071 & n16075 ) | ( n16074 & n16075 ) ;
  assign n16080 = n1538 & n2712 ;
  assign n16081 = ~n15517 & n16080 ;
  assign n16077 = n8075 ^ n261 ^ 1'b0 ;
  assign n16078 = n8495 & ~n16077 ;
  assign n16079 = n16078 ^ n4769 ^ n807 ;
  assign n16082 = n16081 ^ n16079 ^ n9260 ;
  assign n16083 = n10921 & n16082 ;
  assign n16084 = n13520 ^ n6243 ^ n5835 ;
  assign n16085 = n16084 ^ n7822 ^ n4039 ;
  assign n16086 = ( n8565 & n11099 ) | ( n8565 & n16085 ) | ( n11099 & n16085 ) ;
  assign n16087 = ( n4322 & n9556 ) | ( n4322 & n16086 ) | ( n9556 & n16086 ) ;
  assign n16088 = ( n5365 & n16083 ) | ( n5365 & n16087 ) | ( n16083 & n16087 ) ;
  assign n16089 = n13876 ^ n3650 ^ n194 ;
  assign n16090 = n16089 ^ n14526 ^ n11462 ;
  assign n16093 = ~n1525 & n7543 ;
  assign n16094 = n16093 ^ n14119 ^ 1'b0 ;
  assign n16091 = ~n1955 & n14307 ;
  assign n16092 = n16091 ^ n12075 ^ n5551 ;
  assign n16095 = n16094 ^ n16092 ^ n11555 ;
  assign n16096 = ( ~n5835 & n6727 ) | ( ~n5835 & n9643 ) | ( n6727 & n9643 ) ;
  assign n16097 = n2975 | n7948 ;
  assign n16098 = ( ~n5866 & n8221 ) | ( ~n5866 & n10652 ) | ( n8221 & n10652 ) ;
  assign n16099 = ( n549 & n16097 ) | ( n549 & n16098 ) | ( n16097 & n16098 ) ;
  assign n16100 = ~n1426 & n13775 ;
  assign n16101 = ~n2510 & n16100 ;
  assign n16102 = ( n1056 & n11162 ) | ( n1056 & ~n16101 ) | ( n11162 & ~n16101 ) ;
  assign n16103 = n16102 ^ n13045 ^ n4966 ;
  assign n16104 = n4755 & ~n10136 ;
  assign n16105 = n16103 & n16104 ;
  assign n16106 = n16105 ^ n13534 ^ n11897 ;
  assign n16107 = ~n9246 & n16102 ;
  assign n16108 = n16107 ^ n6103 ^ 1'b0 ;
  assign n16109 = ( n5080 & n7264 ) | ( n5080 & n15651 ) | ( n7264 & n15651 ) ;
  assign n16110 = n16109 ^ n1712 ^ n744 ;
  assign n16111 = n6008 ^ n2403 ^ n2082 ;
  assign n16112 = n4840 | n16111 ;
  assign n16113 = n6789 & ~n16112 ;
  assign n16114 = ( n2213 & n3241 ) | ( n2213 & n16113 ) | ( n3241 & n16113 ) ;
  assign n16115 = n5477 | n8420 ;
  assign n16116 = n1486 & ~n16115 ;
  assign n16117 = n6627 ^ n5514 ^ n237 ;
  assign n16118 = ( ~n3533 & n3547 ) | ( ~n3533 & n4042 ) | ( n3547 & n4042 ) ;
  assign n16119 = ( n13119 & n15080 ) | ( n13119 & n16118 ) | ( n15080 & n16118 ) ;
  assign n16120 = n4204 | n8690 ;
  assign n16121 = n4410 | n16120 ;
  assign n16122 = n16121 ^ n9568 ^ n2956 ;
  assign n16123 = ( ~n3777 & n7988 ) | ( ~n3777 & n9098 ) | ( n7988 & n9098 ) ;
  assign n16124 = ( n176 & n3721 ) | ( n176 & n9714 ) | ( n3721 & n9714 ) ;
  assign n16125 = ~n10510 & n16124 ;
  assign n16126 = ~n13357 & n16125 ;
  assign n16127 = n11081 ^ n9211 ^ n5061 ;
  assign n16128 = n16127 ^ n12231 ^ 1'b0 ;
  assign n16129 = n16126 | n16128 ;
  assign n16130 = n10314 ^ n310 ^ 1'b0 ;
  assign n16131 = n4969 | n16130 ;
  assign n16133 = ( ~n949 & n10039 ) | ( ~n949 & n10314 ) | ( n10039 & n10314 ) ;
  assign n16132 = n9584 ^ n1094 ^ 1'b0 ;
  assign n16134 = n16133 ^ n16132 ^ n6884 ;
  assign n16135 = n15274 ^ n5802 ^ n1846 ;
  assign n16136 = ( ~n1529 & n9426 ) | ( ~n1529 & n16135 ) | ( n9426 & n16135 ) ;
  assign n16137 = ( n16131 & ~n16134 ) | ( n16131 & n16136 ) | ( ~n16134 & n16136 ) ;
  assign n16139 = ( n626 & ~n4775 ) | ( n626 & n9976 ) | ( ~n4775 & n9976 ) ;
  assign n16140 = ( n3736 & n10366 ) | ( n3736 & n16139 ) | ( n10366 & n16139 ) ;
  assign n16138 = n10995 ^ n6312 ^ n4378 ;
  assign n16141 = n16140 ^ n16138 ^ n2525 ;
  assign n16142 = n15630 ^ n12512 ^ n4218 ;
  assign n16143 = n14895 ^ n11439 ^ n11317 ;
  assign n16144 = ( n2316 & ~n16142 ) | ( n2316 & n16143 ) | ( ~n16142 & n16143 ) ;
  assign n16145 = n16144 ^ n3317 ^ 1'b0 ;
  assign n16146 = n4541 | n16145 ;
  assign n16147 = n3111 ^ n3033 ^ n233 ;
  assign n16148 = ( n5706 & ~n12899 ) | ( n5706 & n16147 ) | ( ~n12899 & n16147 ) ;
  assign n16149 = n16148 ^ n9182 ^ n6295 ;
  assign n16150 = ~n9524 & n16149 ;
  assign n16151 = n16150 ^ n12379 ^ 1'b0 ;
  assign n16152 = n16151 ^ n9314 ^ 1'b0 ;
  assign n16153 = n11873 ^ n4940 ^ n3332 ;
  assign n16154 = ( n1048 & ~n8861 ) | ( n1048 & n13357 ) | ( ~n8861 & n13357 ) ;
  assign n16155 = ( ~n12857 & n16153 ) | ( ~n12857 & n16154 ) | ( n16153 & n16154 ) ;
  assign n16156 = n10348 ^ n7762 ^ n2910 ;
  assign n16157 = n16155 | n16156 ;
  assign n16158 = n16157 ^ n9066 ^ 1'b0 ;
  assign n16159 = ( n9152 & ~n13209 ) | ( n9152 & n16158 ) | ( ~n13209 & n16158 ) ;
  assign n16161 = ( n709 & n2119 ) | ( n709 & ~n9258 ) | ( n2119 & ~n9258 ) ;
  assign n16160 = ( n170 & ~n7465 ) | ( n170 & n11961 ) | ( ~n7465 & n11961 ) ;
  assign n16162 = n16161 ^ n16160 ^ n2465 ;
  assign n16163 = n16162 ^ n7133 ^ n1197 ;
  assign n16164 = ( n15875 & n15998 ) | ( n15875 & n16163 ) | ( n15998 & n16163 ) ;
  assign n16165 = n8516 ^ n2324 ^ n1293 ;
  assign n16166 = ( n2186 & n9396 ) | ( n2186 & ~n14567 ) | ( n9396 & ~n14567 ) ;
  assign n16167 = ( x121 & n3899 ) | ( x121 & ~n16166 ) | ( n3899 & ~n16166 ) ;
  assign n16169 = n4721 ^ n1958 ^ n891 ;
  assign n16168 = n10788 ^ n5156 ^ n2168 ;
  assign n16170 = n16169 ^ n16168 ^ n4499 ;
  assign n16171 = n3942 ^ n2320 ^ x48 ;
  assign n16172 = ( n5380 & n15719 ) | ( n5380 & n16171 ) | ( n15719 & n16171 ) ;
  assign n16173 = n8671 ^ n6759 ^ n5195 ;
  assign n16174 = n16173 ^ n15647 ^ n3251 ;
  assign n16175 = n16174 ^ n7041 ^ 1'b0 ;
  assign n16176 = ~n16172 & n16175 ;
  assign n16177 = ~n6789 & n13410 ;
  assign n16178 = n12078 ^ n11939 ^ 1'b0 ;
  assign n16179 = n3379 & ~n16178 ;
  assign n16180 = ~n640 & n16179 ;
  assign n16181 = n10959 ^ n10680 ^ n7229 ;
  assign n16182 = n3461 & ~n13493 ;
  assign n16183 = n16182 ^ n1588 ^ 1'b0 ;
  assign n16184 = ( n1077 & n2940 ) | ( n1077 & n6374 ) | ( n2940 & n6374 ) ;
  assign n16185 = n5893 ^ n5266 ^ n2552 ;
  assign n16186 = ( n16183 & n16184 ) | ( n16183 & n16185 ) | ( n16184 & n16185 ) ;
  assign n16187 = ( n4401 & ~n16181 ) | ( n4401 & n16186 ) | ( ~n16181 & n16186 ) ;
  assign n16188 = ( ~n2850 & n3239 ) | ( ~n2850 & n3637 ) | ( n3239 & n3637 ) ;
  assign n16189 = n16188 ^ n14639 ^ n7420 ;
  assign n16190 = ~n1451 & n16189 ;
  assign n16191 = ( n12745 & n16068 ) | ( n12745 & ~n16190 ) | ( n16068 & ~n16190 ) ;
  assign n16192 = ~n4876 & n13254 ;
  assign n16193 = ( n13174 & n14117 ) | ( n13174 & ~n16192 ) | ( n14117 & ~n16192 ) ;
  assign n16194 = ( ~n1355 & n3214 ) | ( ~n1355 & n4838 ) | ( n3214 & n4838 ) ;
  assign n16195 = ( n3781 & n9087 ) | ( n3781 & ~n16194 ) | ( n9087 & ~n16194 ) ;
  assign n16196 = n16195 ^ n13966 ^ n3133 ;
  assign n16197 = n16196 ^ n6676 ^ n3416 ;
  assign n16198 = n12501 ^ n7687 ^ n1459 ;
  assign n16199 = n11238 ^ n4684 ^ n2988 ;
  assign n16200 = ~n1680 & n16199 ;
  assign n16201 = ~n16198 & n16200 ;
  assign n16202 = n2906 ^ n546 ^ 1'b0 ;
  assign n16203 = n6031 & ~n16202 ;
  assign n16204 = ( n3731 & n3924 ) | ( n3731 & ~n9324 ) | ( n3924 & ~n9324 ) ;
  assign n16205 = n16204 ^ n6094 ^ 1'b0 ;
  assign n16206 = n16205 ^ n11689 ^ n1297 ;
  assign n16207 = n12497 ^ n8079 ^ n5544 ;
  assign n16208 = ~n3708 & n4742 ;
  assign n16209 = ~n16207 & n16208 ;
  assign n16210 = ( n3042 & ~n5783 ) | ( n3042 & n5882 ) | ( ~n5783 & n5882 ) ;
  assign n16211 = n15281 ^ n1251 ^ 1'b0 ;
  assign n16212 = n9434 | n16211 ;
  assign n16213 = ( ~n4922 & n16210 ) | ( ~n4922 & n16212 ) | ( n16210 & n16212 ) ;
  assign n16218 = n3544 ^ n3367 ^ 1'b0 ;
  assign n16219 = ( n10175 & ~n14066 ) | ( n10175 & n16218 ) | ( ~n14066 & n16218 ) ;
  assign n16214 = ( ~n2062 & n6036 ) | ( ~n2062 & n6592 ) | ( n6036 & n6592 ) ;
  assign n16215 = ( n4476 & n8034 ) | ( n4476 & n16214 ) | ( n8034 & n16214 ) ;
  assign n16216 = n16215 ^ n9142 ^ n7279 ;
  assign n16217 = n16216 ^ n4978 ^ x24 ;
  assign n16220 = n16219 ^ n16217 ^ n12957 ;
  assign n16221 = n12656 ^ n8962 ^ n761 ;
  assign n16222 = n9673 ^ n2276 ^ n2241 ;
  assign n16223 = ( ~x6 & n1629 ) | ( ~x6 & n11135 ) | ( n1629 & n11135 ) ;
  assign n16224 = ( n12873 & n14696 ) | ( n12873 & n16223 ) | ( n14696 & n16223 ) ;
  assign n16225 = n13865 | n16224 ;
  assign n16226 = n16225 ^ n6090 ^ 1'b0 ;
  assign n16227 = n6767 ^ n2364 ^ 1'b0 ;
  assign n16228 = x39 & n16227 ;
  assign n16229 = ( n1541 & n4676 ) | ( n1541 & ~n16228 ) | ( n4676 & ~n16228 ) ;
  assign n16230 = ( n16222 & n16226 ) | ( n16222 & ~n16229 ) | ( n16226 & ~n16229 ) ;
  assign n16237 = ( n6668 & ~n7635 ) | ( n6668 & n12969 ) | ( ~n7635 & n12969 ) ;
  assign n16238 = n16237 ^ n7607 ^ n4754 ;
  assign n16235 = ( n4154 & n8866 ) | ( n4154 & n15078 ) | ( n8866 & n15078 ) ;
  assign n16231 = ( n1486 & n8036 ) | ( n1486 & n13741 ) | ( n8036 & n13741 ) ;
  assign n16232 = ( n872 & n15426 ) | ( n872 & ~n16231 ) | ( n15426 & ~n16231 ) ;
  assign n16233 = n13086 | n16232 ;
  assign n16234 = n10729 | n16233 ;
  assign n16236 = n16235 ^ n16234 ^ n7094 ;
  assign n16239 = n16238 ^ n16236 ^ n15583 ;
  assign n16240 = n5808 & ~n13185 ;
  assign n16241 = n16240 ^ n4458 ^ 1'b0 ;
  assign n16242 = ( ~n1907 & n5014 ) | ( ~n1907 & n5914 ) | ( n5014 & n5914 ) ;
  assign n16243 = ( ~n3528 & n3679 ) | ( ~n3528 & n8566 ) | ( n3679 & n8566 ) ;
  assign n16244 = ( n6088 & ~n16242 ) | ( n6088 & n16243 ) | ( ~n16242 & n16243 ) ;
  assign n16245 = n10254 ^ n5272 ^ n3476 ;
  assign n16246 = n16244 | n16245 ;
  assign n16247 = n9712 ^ n4496 ^ n1617 ;
  assign n16248 = ( n1295 & n5695 ) | ( n1295 & ~n16247 ) | ( n5695 & ~n16247 ) ;
  assign n16249 = n13367 & ~n15670 ;
  assign n16250 = n1190 | n5463 ;
  assign n16251 = n16249 & ~n16250 ;
  assign n16252 = ( n5192 & n16248 ) | ( n5192 & n16251 ) | ( n16248 & n16251 ) ;
  assign n16253 = n1537 & n2767 ;
  assign n16254 = ( n6801 & ~n9035 ) | ( n6801 & n16253 ) | ( ~n9035 & n16253 ) ;
  assign n16255 = n775 ^ n288 ^ 1'b0 ;
  assign n16256 = ~n2884 & n12921 ;
  assign n16257 = ~n10178 & n16256 ;
  assign n16258 = ( n15484 & n16255 ) | ( n15484 & ~n16257 ) | ( n16255 & ~n16257 ) ;
  assign n16260 = n3204 ^ n2310 ^ 1'b0 ;
  assign n16261 = ( ~n11601 & n13023 ) | ( ~n11601 & n16260 ) | ( n13023 & n16260 ) ;
  assign n16259 = n9085 ^ n8643 ^ 1'b0 ;
  assign n16262 = n16261 ^ n16259 ^ n3860 ;
  assign n16263 = ( n2188 & ~n7408 ) | ( n2188 & n10764 ) | ( ~n7408 & n10764 ) ;
  assign n16264 = n16263 ^ n7069 ^ n6452 ;
  assign n16265 = n16264 ^ n14470 ^ n3086 ;
  assign n16266 = ( n11375 & n11564 ) | ( n11375 & n13990 ) | ( n11564 & n13990 ) ;
  assign n16267 = n16266 ^ n3203 ^ n596 ;
  assign n16273 = ( ~n4225 & n8611 ) | ( ~n4225 & n13198 ) | ( n8611 & n13198 ) ;
  assign n16270 = n7665 ^ n2727 ^ n2283 ;
  assign n16268 = n2253 & n4072 ;
  assign n16269 = n16268 ^ n2834 ^ 1'b0 ;
  assign n16271 = n16270 ^ n16269 ^ 1'b0 ;
  assign n16272 = ( n4557 & ~n10143 ) | ( n4557 & n16271 ) | ( ~n10143 & n16271 ) ;
  assign n16274 = n16273 ^ n16272 ^ n15183 ;
  assign n16275 = ( ~x16 & n1140 ) | ( ~x16 & n14416 ) | ( n1140 & n14416 ) ;
  assign n16276 = n210 & ~n1459 ;
  assign n16277 = n3005 & n16276 ;
  assign n16278 = ( n5844 & n6593 ) | ( n5844 & n16277 ) | ( n6593 & n16277 ) ;
  assign n16279 = n12342 & ~n16278 ;
  assign n16280 = n16279 ^ n14688 ^ 1'b0 ;
  assign n16281 = ( n3004 & ~n16275 ) | ( n3004 & n16280 ) | ( ~n16275 & n16280 ) ;
  assign n16286 = n9016 ^ n708 ^ 1'b0 ;
  assign n16282 = ( n5475 & ~n6674 ) | ( n5475 & n8281 ) | ( ~n6674 & n8281 ) ;
  assign n16283 = ( n1333 & n4874 ) | ( n1333 & n15346 ) | ( n4874 & n15346 ) ;
  assign n16284 = ( ~n10808 & n11840 ) | ( ~n10808 & n16283 ) | ( n11840 & n16283 ) ;
  assign n16285 = ( n9820 & n16282 ) | ( n9820 & ~n16284 ) | ( n16282 & ~n16284 ) ;
  assign n16287 = n16286 ^ n16285 ^ n9493 ;
  assign n16288 = ( n506 & n1578 ) | ( n506 & ~n5553 ) | ( n1578 & ~n5553 ) ;
  assign n16289 = n14097 | n16288 ;
  assign n16290 = n11156 | n16289 ;
  assign n16291 = n6698 ^ n5831 ^ 1'b0 ;
  assign n16292 = n16290 & ~n16291 ;
  assign n16293 = n16292 ^ n3375 ^ n2074 ;
  assign n16294 = n9610 ^ n9465 ^ n6712 ;
  assign n16297 = ( n454 & ~n6586 ) | ( n454 & n7879 ) | ( ~n6586 & n7879 ) ;
  assign n16298 = ( ~n7558 & n8221 ) | ( ~n7558 & n12277 ) | ( n8221 & n12277 ) ;
  assign n16299 = n16298 ^ n14902 ^ n612 ;
  assign n16300 = ( n9471 & ~n16297 ) | ( n9471 & n16299 ) | ( ~n16297 & n16299 ) ;
  assign n16295 = n4440 & ~n5010 ;
  assign n16296 = n4348 & n16295 ;
  assign n16301 = n16300 ^ n16296 ^ n654 ;
  assign n16302 = ~n3156 & n16301 ;
  assign n16303 = ~n16294 & n16302 ;
  assign n16304 = n11807 ^ n2043 ^ n1795 ;
  assign n16305 = n7219 & ~n16304 ;
  assign n16306 = n5623 ^ n2066 ^ 1'b0 ;
  assign n16307 = ( ~n9704 & n15372 ) | ( ~n9704 & n16306 ) | ( n15372 & n16306 ) ;
  assign n16308 = n14945 ^ n14762 ^ n13119 ;
  assign n16309 = ( ~n268 & n10176 ) | ( ~n268 & n12899 ) | ( n10176 & n12899 ) ;
  assign n16310 = ( n768 & n1655 ) | ( n768 & n16309 ) | ( n1655 & n16309 ) ;
  assign n16311 = n3833 ^ n3757 ^ n2157 ;
  assign n16312 = n14535 ^ n3402 ^ n2528 ;
  assign n16313 = ( n2947 & n5489 ) | ( n2947 & ~n9510 ) | ( n5489 & ~n9510 ) ;
  assign n16314 = n396 & ~n16313 ;
  assign n16315 = ~n9399 & n16314 ;
  assign n16316 = n13666 ^ n10083 ^ n2212 ;
  assign n16317 = n10375 ^ n4019 ^ 1'b0 ;
  assign n16318 = n16317 ^ n1324 ^ n259 ;
  assign n16319 = ( ~n7562 & n16316 ) | ( ~n7562 & n16318 ) | ( n16316 & n16318 ) ;
  assign n16320 = n16319 ^ n4381 ^ n2872 ;
  assign n16321 = n13883 ^ n11579 ^ n10822 ;
  assign n16322 = n5289 ^ n2788 ^ n2038 ;
  assign n16323 = ( n2410 & ~n6317 ) | ( n2410 & n12386 ) | ( ~n6317 & n12386 ) ;
  assign n16324 = n16323 ^ n14071 ^ n2193 ;
  assign n16325 = ( n10860 & n16322 ) | ( n10860 & ~n16324 ) | ( n16322 & ~n16324 ) ;
  assign n16326 = n9504 ^ n2481 ^ n2005 ;
  assign n16327 = n16326 ^ n12132 ^ n2498 ;
  assign n16328 = ( n10240 & n12637 ) | ( n10240 & ~n16327 ) | ( n12637 & ~n16327 ) ;
  assign n16329 = ( n528 & n8515 ) | ( n528 & ~n9712 ) | ( n8515 & ~n9712 ) ;
  assign n16330 = n16329 ^ n10664 ^ n6461 ;
  assign n16331 = ( n8036 & ~n8820 ) | ( n8036 & n10472 ) | ( ~n8820 & n10472 ) ;
  assign n16332 = n10728 ^ n9700 ^ n2553 ;
  assign n16333 = n10205 ^ x75 ^ 1'b0 ;
  assign n16334 = n16333 ^ n9000 ^ n1790 ;
  assign n16335 = n8901 ^ n8142 ^ n5049 ;
  assign n16336 = n4959 ^ n2250 ^ 1'b0 ;
  assign n16337 = n16335 & ~n16336 ;
  assign n16339 = n758 & n7532 ;
  assign n16340 = ~n13800 & n16339 ;
  assign n16338 = n13249 ^ n12561 ^ n6870 ;
  assign n16341 = n16340 ^ n16338 ^ n7234 ;
  assign n16342 = n2324 ^ n1267 ^ x108 ;
  assign n16343 = n16342 ^ n4002 ^ n2943 ;
  assign n16344 = n11178 ^ n1942 ^ n1577 ;
  assign n16345 = n8114 ^ n3356 ^ 1'b0 ;
  assign n16346 = n12712 & ~n16345 ;
  assign n16347 = ( n5359 & n6715 ) | ( n5359 & n16346 ) | ( n6715 & n16346 ) ;
  assign n16348 = ( ~n5387 & n6543 ) | ( ~n5387 & n8406 ) | ( n6543 & n8406 ) ;
  assign n16349 = n3219 & n16348 ;
  assign n16350 = ( n16344 & ~n16347 ) | ( n16344 & n16349 ) | ( ~n16347 & n16349 ) ;
  assign n16351 = n8643 ^ n5395 ^ 1'b0 ;
  assign n16352 = n4074 & ~n7161 ;
  assign n16353 = n13990 ^ n10639 ^ n7314 ;
  assign n16354 = n1822 ^ n132 ^ 1'b0 ;
  assign n16355 = n3686 | n16354 ;
  assign n16356 = n16353 | n16355 ;
  assign n16357 = n16356 ^ n10738 ^ 1'b0 ;
  assign n16358 = ( ~n16351 & n16352 ) | ( ~n16351 & n16357 ) | ( n16352 & n16357 ) ;
  assign n16359 = n15688 ^ n7857 ^ n7519 ;
  assign n16363 = ( n3402 & n6541 ) | ( n3402 & ~n10002 ) | ( n6541 & ~n10002 ) ;
  assign n16362 = n183 & n9222 ;
  assign n16364 = n16363 ^ n16362 ^ n11411 ;
  assign n16360 = ( n3129 & n8803 ) | ( n3129 & n13242 ) | ( n8803 & n13242 ) ;
  assign n16361 = ( n1957 & n2120 ) | ( n1957 & ~n16360 ) | ( n2120 & ~n16360 ) ;
  assign n16365 = n16364 ^ n16361 ^ n1442 ;
  assign n16368 = n9435 ^ n3043 ^ n2159 ;
  assign n16369 = n5977 ^ n5281 ^ n1663 ;
  assign n16370 = ( n8796 & n16368 ) | ( n8796 & ~n16369 ) | ( n16368 & ~n16369 ) ;
  assign n16367 = n9764 & n14000 ;
  assign n16371 = n16370 ^ n16367 ^ 1'b0 ;
  assign n16366 = n11057 ^ n7015 ^ n637 ;
  assign n16372 = n16371 ^ n16366 ^ n15134 ;
  assign n16373 = n4156 ^ n2740 ^ n2155 ;
  assign n16374 = n16373 ^ n7139 ^ n3198 ;
  assign n16375 = ( n2737 & ~n2876 ) | ( n2737 & n16374 ) | ( ~n2876 & n16374 ) ;
  assign n16376 = n16375 ^ n12922 ^ n2934 ;
  assign n16377 = n2941 & n16376 ;
  assign n16378 = n13753 ^ n6121 ^ 1'b0 ;
  assign n16379 = x24 & n16378 ;
  assign n16380 = ( n4087 & n7980 ) | ( n4087 & n16379 ) | ( n7980 & n16379 ) ;
  assign n16381 = n10332 & ~n16380 ;
  assign n16382 = n16381 ^ n5960 ^ 1'b0 ;
  assign n16386 = ~n2913 & n6543 ;
  assign n16387 = n16386 ^ n3784 ^ 1'b0 ;
  assign n16383 = n6712 ^ n3266 ^ 1'b0 ;
  assign n16384 = n3499 & ~n16383 ;
  assign n16385 = n16384 ^ n11970 ^ n3820 ;
  assign n16388 = n16387 ^ n16385 ^ n12463 ;
  assign n16389 = n2596 ^ n1713 ^ n495 ;
  assign n16390 = n1063 ^ x86 ^ 1'b0 ;
  assign n16391 = ( n6633 & ~n7699 ) | ( n6633 & n16390 ) | ( ~n7699 & n16390 ) ;
  assign n16392 = n16391 ^ n10819 ^ n6349 ;
  assign n16393 = ( ~n1612 & n1815 ) | ( ~n1612 & n1943 ) | ( n1815 & n1943 ) ;
  assign n16394 = n16393 ^ n15456 ^ n462 ;
  assign n16395 = n7722 | n9453 ;
  assign n16396 = ( n4393 & n11725 ) | ( n4393 & n12630 ) | ( n11725 & n12630 ) ;
  assign n16397 = n16395 | n16396 ;
  assign n16398 = n15177 ^ n811 ^ 1'b0 ;
  assign n16399 = n10272 & n16398 ;
  assign n16400 = n4042 ^ n2633 ^ n805 ;
  assign n16403 = n304 ^ x81 ^ 1'b0 ;
  assign n16404 = n16403 ^ n13919 ^ n6253 ;
  assign n16401 = n12833 & n14009 ;
  assign n16402 = n16401 ^ n8645 ^ 1'b0 ;
  assign n16405 = n16404 ^ n16402 ^ n2189 ;
  assign n16406 = ( n9855 & n16400 ) | ( n9855 & ~n16405 ) | ( n16400 & ~n16405 ) ;
  assign n16407 = n12123 ^ n1887 ^ 1'b0 ;
  assign n16408 = ( n4930 & n8147 ) | ( n4930 & ~n12422 ) | ( n8147 & ~n12422 ) ;
  assign n16409 = n16408 ^ n11840 ^ n8191 ;
  assign n16410 = n16409 ^ n13546 ^ n3787 ;
  assign n16411 = ( ~n3152 & n10460 ) | ( ~n3152 & n15799 ) | ( n10460 & n15799 ) ;
  assign n16412 = ( n6798 & n7069 ) | ( n6798 & n9434 ) | ( n7069 & n9434 ) ;
  assign n16413 = ( n8369 & ~n11422 ) | ( n8369 & n16412 ) | ( ~n11422 & n16412 ) ;
  assign n16414 = ( n11224 & ~n16411 ) | ( n11224 & n16413 ) | ( ~n16411 & n16413 ) ;
  assign n16415 = ( n1926 & ~n5695 ) | ( n1926 & n7778 ) | ( ~n5695 & n7778 ) ;
  assign n16416 = n16415 ^ n9171 ^ n6429 ;
  assign n16417 = n7258 ^ n3378 ^ n2245 ;
  assign n16422 = ( n962 & ~n3346 ) | ( n962 & n10955 ) | ( ~n3346 & n10955 ) ;
  assign n16423 = n4201 & n16422 ;
  assign n16420 = ( n4582 & n6961 ) | ( n4582 & n7149 ) | ( n6961 & n7149 ) ;
  assign n16418 = n7077 ^ n5753 ^ 1'b0 ;
  assign n16419 = n15255 & ~n16418 ;
  assign n16421 = n16420 ^ n16419 ^ n14315 ;
  assign n16424 = n16423 ^ n16421 ^ n1275 ;
  assign n16425 = n15831 ^ n8890 ^ n4322 ;
  assign n16426 = ( n563 & ~n11942 ) | ( n563 & n14116 ) | ( ~n11942 & n14116 ) ;
  assign n16427 = n16426 ^ n13959 ^ n884 ;
  assign n16428 = ( ~n6444 & n8759 ) | ( ~n6444 & n16427 ) | ( n8759 & n16427 ) ;
  assign n16429 = n5917 ^ n4073 ^ n3324 ;
  assign n16430 = ( n280 & n1271 ) | ( n280 & n5793 ) | ( n1271 & n5793 ) ;
  assign n16431 = ( ~n4954 & n9076 ) | ( ~n4954 & n16430 ) | ( n9076 & n16430 ) ;
  assign n16432 = n16431 ^ n13273 ^ n10371 ;
  assign n16433 = n16429 | n16432 ;
  assign n16434 = n16433 ^ n762 ^ 1'b0 ;
  assign n16435 = n4572 & ~n6016 ;
  assign n16436 = n16435 ^ n6417 ^ 1'b0 ;
  assign n16437 = ( ~n827 & n5632 ) | ( ~n827 & n16436 ) | ( n5632 & n16436 ) ;
  assign n16438 = ( n3679 & n9206 ) | ( n3679 & n10981 ) | ( n9206 & n10981 ) ;
  assign n16439 = n12032 ^ n11082 ^ n1610 ;
  assign n16440 = n5154 ^ n2833 ^ n1275 ;
  assign n16441 = n6088 ^ n5675 ^ 1'b0 ;
  assign n16442 = n16440 | n16441 ;
  assign n16443 = ~n2170 & n5627 ;
  assign n16444 = n16442 & n16443 ;
  assign n16445 = ( n762 & ~n8285 ) | ( n762 & n13316 ) | ( ~n8285 & n13316 ) ;
  assign n16446 = ( n2342 & n4451 ) | ( n2342 & n16445 ) | ( n4451 & n16445 ) ;
  assign n16447 = n10298 | n13220 ;
  assign n16448 = n16447 ^ n2522 ^ n594 ;
  assign n16449 = n16448 ^ n14145 ^ n9189 ;
  assign n16450 = ( ~n3034 & n3281 ) | ( ~n3034 & n4614 ) | ( n3281 & n4614 ) ;
  assign n16452 = n12095 ^ n11164 ^ n6900 ;
  assign n16451 = n9652 ^ n1995 ^ n510 ;
  assign n16453 = n16452 ^ n16451 ^ n11077 ;
  assign n16454 = ( n4822 & n4876 ) | ( n4822 & n9189 ) | ( n4876 & n9189 ) ;
  assign n16455 = n16454 ^ n10156 ^ 1'b0 ;
  assign n16456 = n2630 & ~n13305 ;
  assign n16457 = ~n16455 & n16456 ;
  assign n16459 = n3133 ^ n1814 ^ 1'b0 ;
  assign n16460 = ~n1288 & n16459 ;
  assign n16458 = n14273 ^ n10106 ^ n2295 ;
  assign n16461 = n16460 ^ n16458 ^ n11382 ;
  assign n16462 = ( ~n1160 & n4846 ) | ( ~n1160 & n11694 ) | ( n4846 & n11694 ) ;
  assign n16463 = n7217 & n16462 ;
  assign n16464 = n10586 ^ n7660 ^ n2443 ;
  assign n16465 = ( ~n199 & n2143 ) | ( ~n199 & n16464 ) | ( n2143 & n16464 ) ;
  assign n16466 = ( n9827 & n16463 ) | ( n9827 & ~n16465 ) | ( n16463 & ~n16465 ) ;
  assign n16467 = ( n3488 & n8075 ) | ( n3488 & ~n14969 ) | ( n8075 & ~n14969 ) ;
  assign n16468 = n4569 & ~n7443 ;
  assign n16469 = n2270 & n16468 ;
  assign n16470 = n16469 ^ n7211 ^ n1835 ;
  assign n16471 = ( n8496 & ~n10742 ) | ( n8496 & n16470 ) | ( ~n10742 & n16470 ) ;
  assign n16472 = n16471 ^ n2164 ^ 1'b0 ;
  assign n16473 = n16467 & n16472 ;
  assign n16478 = ( n854 & n1794 ) | ( n854 & n10359 ) | ( n1794 & n10359 ) ;
  assign n16474 = ( n385 & n1558 ) | ( n385 & ~n10051 ) | ( n1558 & ~n10051 ) ;
  assign n16475 = ( n950 & n2874 ) | ( n950 & n8607 ) | ( n2874 & n8607 ) ;
  assign n16476 = n16474 | n16475 ;
  assign n16477 = n7919 | n16476 ;
  assign n16479 = n16478 ^ n16477 ^ n4783 ;
  assign n16480 = ( ~n1630 & n6096 ) | ( ~n1630 & n8383 ) | ( n6096 & n8383 ) ;
  assign n16481 = n16480 ^ n12150 ^ n8541 ;
  assign n16487 = n14789 ^ n13652 ^ n365 ;
  assign n16482 = n5745 & ~n11703 ;
  assign n16483 = n16482 ^ n6103 ^ 1'b0 ;
  assign n16484 = ( ~n5976 & n10397 ) | ( ~n5976 & n16483 ) | ( n10397 & n16483 ) ;
  assign n16485 = n16484 ^ n9058 ^ n751 ;
  assign n16486 = n16485 ^ n4021 ^ n876 ;
  assign n16488 = n16487 ^ n16486 ^ n3494 ;
  assign n16489 = ( n1715 & n8016 ) | ( n1715 & n15347 ) | ( n8016 & n15347 ) ;
  assign n16490 = n4093 ^ n2217 ^ n909 ;
  assign n16491 = ( n5727 & ~n6439 ) | ( n5727 & n16490 ) | ( ~n6439 & n16490 ) ;
  assign n16492 = ( ~n11012 & n12570 ) | ( ~n11012 & n16491 ) | ( n12570 & n16491 ) ;
  assign n16493 = ( ~n2583 & n5377 ) | ( ~n2583 & n9795 ) | ( n5377 & n9795 ) ;
  assign n16494 = n16493 ^ n9373 ^ n1577 ;
  assign n16495 = n16494 ^ n5753 ^ n1815 ;
  assign n16496 = ( n4554 & ~n8090 ) | ( n4554 & n16495 ) | ( ~n8090 & n16495 ) ;
  assign n16497 = ( n13932 & n16492 ) | ( n13932 & n16496 ) | ( n16492 & n16496 ) ;
  assign n16498 = n14326 ^ n4948 ^ n1594 ;
  assign n16500 = ( ~n302 & n3011 ) | ( ~n302 & n14040 ) | ( n3011 & n14040 ) ;
  assign n16499 = n10087 ^ n5982 ^ n2029 ;
  assign n16501 = n16500 ^ n16499 ^ n13953 ;
  assign n16502 = ( n646 & ~n4440 ) | ( n646 & n11926 ) | ( ~n4440 & n11926 ) ;
  assign n16503 = n12486 ^ n8652 ^ n3101 ;
  assign n16504 = n16503 ^ n11572 ^ n3560 ;
  assign n16505 = ( n6194 & ~n13617 ) | ( n6194 & n16504 ) | ( ~n13617 & n16504 ) ;
  assign n16506 = n13627 ^ n3332 ^ n2453 ;
  assign n16507 = n16506 ^ n12044 ^ n5038 ;
  assign n16508 = n13880 ^ n3629 ^ n3568 ;
  assign n16509 = ( ~n9236 & n15855 ) | ( ~n9236 & n16508 ) | ( n15855 & n16508 ) ;
  assign n16510 = ( n1789 & ~n5741 ) | ( n1789 & n16509 ) | ( ~n5741 & n16509 ) ;
  assign n16511 = n12402 ^ n12319 ^ n2910 ;
  assign n16512 = n16511 ^ n9244 ^ 1'b0 ;
  assign n16513 = ( n3796 & ~n9872 ) | ( n3796 & n14567 ) | ( ~n9872 & n14567 ) ;
  assign n16515 = n10052 ^ n2589 ^ n747 ;
  assign n16514 = n5903 ^ n2361 ^ n1566 ;
  assign n16516 = n16515 ^ n16514 ^ n513 ;
  assign n16517 = ( ~n974 & n6899 ) | ( ~n974 & n9558 ) | ( n6899 & n9558 ) ;
  assign n16518 = ( ~x62 & n3597 ) | ( ~x62 & n10573 ) | ( n3597 & n10573 ) ;
  assign n16519 = n16518 ^ n10250 ^ 1'b0 ;
  assign n16520 = n16517 & ~n16519 ;
  assign n16521 = ( n5615 & n11483 ) | ( n5615 & n14258 ) | ( n11483 & n14258 ) ;
  assign n16522 = n16521 ^ n10323 ^ 1'b0 ;
  assign n16523 = n16522 ^ n13971 ^ n7287 ;
  assign n16524 = n9596 ^ n8939 ^ 1'b0 ;
  assign n16525 = ~n5790 & n16524 ;
  assign n16526 = n16525 ^ n6269 ^ n2213 ;
  assign n16530 = n10626 ^ n6240 ^ n2034 ;
  assign n16528 = ( n7217 & ~n11724 ) | ( n7217 & n15528 ) | ( ~n11724 & n15528 ) ;
  assign n16529 = ( n11839 & n16266 ) | ( n11839 & ~n16528 ) | ( n16266 & ~n16528 ) ;
  assign n16527 = n11037 ^ n6697 ^ 1'b0 ;
  assign n16531 = n16530 ^ n16529 ^ n16527 ;
  assign n16532 = ( ~n8300 & n16526 ) | ( ~n8300 & n16531 ) | ( n16526 & n16531 ) ;
  assign n16533 = n8406 ^ n3952 ^ n2919 ;
  assign n16534 = ( n10157 & n16189 ) | ( n10157 & n16533 ) | ( n16189 & n16533 ) ;
  assign n16535 = ( n1253 & n1813 ) | ( n1253 & n4121 ) | ( n1813 & n4121 ) ;
  assign n16536 = n16535 ^ n5504 ^ n5410 ;
  assign n16537 = n10454 & ~n16536 ;
  assign n16538 = n2275 & ~n9818 ;
  assign n16539 = ( ~n2705 & n5079 ) | ( ~n2705 & n16538 ) | ( n5079 & n16538 ) ;
  assign n16540 = n16539 ^ n12154 ^ n7616 ;
  assign n16541 = n4764 | n5286 ;
  assign n16542 = ( ~x19 & n2124 ) | ( ~x19 & n3527 ) | ( n2124 & n3527 ) ;
  assign n16543 = ( n3107 & n7210 ) | ( n3107 & n10640 ) | ( n7210 & n10640 ) ;
  assign n16544 = ~n1645 & n16543 ;
  assign n16545 = ~n16542 & n16544 ;
  assign n16546 = ~n16541 & n16545 ;
  assign n16554 = ( n471 & n11349 ) | ( n471 & ~n13337 ) | ( n11349 & ~n13337 ) ;
  assign n16555 = n16554 ^ n6416 ^ n5777 ;
  assign n16556 = n129 & n16181 ;
  assign n16557 = ~n7583 & n16556 ;
  assign n16558 = ( n8505 & ~n16555 ) | ( n8505 & n16557 ) | ( ~n16555 & n16557 ) ;
  assign n16549 = ( ~n2892 & n10063 ) | ( ~n2892 & n14045 ) | ( n10063 & n14045 ) ;
  assign n16550 = n1820 ^ n1148 ^ n193 ;
  assign n16551 = ( n1521 & ~n2834 ) | ( n1521 & n8064 ) | ( ~n2834 & n8064 ) ;
  assign n16552 = ( ~n16549 & n16550 ) | ( ~n16549 & n16551 ) | ( n16550 & n16551 ) ;
  assign n16547 = n7129 ^ n6801 ^ n3574 ;
  assign n16548 = n3780 | n16547 ;
  assign n16553 = n16552 ^ n16548 ^ 1'b0 ;
  assign n16559 = n16558 ^ n16553 ^ n15858 ;
  assign n16560 = n11595 ^ n7951 ^ n6417 ;
  assign n16561 = n13104 ^ n4394 ^ n2908 ;
  assign n16562 = n16561 ^ n9571 ^ 1'b0 ;
  assign n16563 = n9869 ^ n5480 ^ n4437 ;
  assign n16564 = n16563 ^ n12264 ^ n3429 ;
  assign n16565 = n11809 ^ n11489 ^ n7920 ;
  assign n16566 = n10339 ^ n7336 ^ n3881 ;
  assign n16567 = n10990 ^ n4362 ^ n3316 ;
  assign n16568 = ( ~n224 & n5850 ) | ( ~n224 & n16567 ) | ( n5850 & n16567 ) ;
  assign n16569 = ( n2400 & n4541 ) | ( n2400 & n4567 ) | ( n4541 & n4567 ) ;
  assign n16570 = ~n9852 & n16569 ;
  assign n16571 = ~n16568 & n16570 ;
  assign n16572 = ( n8953 & n11431 ) | ( n8953 & ~n16571 ) | ( n11431 & ~n16571 ) ;
  assign n16574 = ( ~n4933 & n6915 ) | ( ~n4933 & n11038 ) | ( n6915 & n11038 ) ;
  assign n16573 = ~n1260 & n5741 ;
  assign n16575 = n16574 ^ n16573 ^ n10072 ;
  assign n16576 = n16326 ^ n9435 ^ n2232 ;
  assign n16577 = ( x71 & n11728 ) | ( x71 & n16576 ) | ( n11728 & n16576 ) ;
  assign n16578 = ( n5171 & n7393 ) | ( n5171 & n16577 ) | ( n7393 & n16577 ) ;
  assign n16580 = n2946 ^ n1348 ^ n321 ;
  assign n16579 = ( ~n2041 & n4263 ) | ( ~n2041 & n10481 ) | ( n4263 & n10481 ) ;
  assign n16581 = n16580 ^ n16579 ^ n11182 ;
  assign n16582 = n14491 ^ n8715 ^ n2048 ;
  assign n16583 = n1169 | n15235 ;
  assign n16584 = n16582 & ~n16583 ;
  assign n16592 = ( n1436 & ~n6040 ) | ( n1436 & n7210 ) | ( ~n6040 & n7210 ) ;
  assign n16585 = ( ~n625 & n1114 ) | ( ~n625 & n3136 ) | ( n1114 & n3136 ) ;
  assign n16587 = n1849 ^ n1478 ^ n832 ;
  assign n16586 = n12156 ^ n1468 ^ n1392 ;
  assign n16588 = n16587 ^ n16586 ^ n3410 ;
  assign n16589 = n16585 | n16588 ;
  assign n16590 = n16589 ^ n5369 ^ 1'b0 ;
  assign n16591 = ~n3153 & n16590 ;
  assign n16593 = n16592 ^ n16591 ^ n5737 ;
  assign n16595 = n5036 ^ n4693 ^ 1'b0 ;
  assign n16596 = ( n4473 & ~n4879 ) | ( n4473 & n16595 ) | ( ~n4879 & n16595 ) ;
  assign n16594 = ( n3260 & n5343 ) | ( n3260 & ~n10655 ) | ( n5343 & ~n10655 ) ;
  assign n16597 = n16596 ^ n16594 ^ n1385 ;
  assign n16598 = ( n2041 & n12355 ) | ( n2041 & n16597 ) | ( n12355 & n16597 ) ;
  assign n16599 = n9851 ^ n3757 ^ 1'b0 ;
  assign n16600 = ( n13702 & n15466 ) | ( n13702 & ~n16599 ) | ( n15466 & ~n16599 ) ;
  assign n16601 = ( n2514 & n8646 ) | ( n2514 & ~n11462 ) | ( n8646 & ~n11462 ) ;
  assign n16602 = n16601 ^ n11041 ^ n3129 ;
  assign n16603 = n16602 ^ n7226 ^ n6924 ;
  assign n16604 = ( n4061 & ~n4949 ) | ( n4061 & n16603 ) | ( ~n4949 & n16603 ) ;
  assign n16605 = n15778 ^ n7333 ^ 1'b0 ;
  assign n16606 = ( n4309 & ~n4562 ) | ( n4309 & n9205 ) | ( ~n4562 & n9205 ) ;
  assign n16607 = ( n3708 & n6937 ) | ( n3708 & ~n11467 ) | ( n6937 & ~n11467 ) ;
  assign n16608 = n15971 ^ n4822 ^ 1'b0 ;
  assign n16609 = ~n16607 & n16608 ;
  assign n16611 = n14884 ^ n7156 ^ n4204 ;
  assign n16612 = n16611 ^ n9808 ^ n2048 ;
  assign n16610 = ( n2220 & n4764 ) | ( n2220 & ~n14986 ) | ( n4764 & ~n14986 ) ;
  assign n16613 = n16612 ^ n16610 ^ n4516 ;
  assign n16614 = n10235 ^ n6620 ^ 1'b0 ;
  assign n16615 = n3029 & ~n16614 ;
  assign n16616 = ( n7053 & n7908 ) | ( n7053 & n10988 ) | ( n7908 & n10988 ) ;
  assign n16617 = n1282 | n2123 ;
  assign n16618 = n16617 ^ n3415 ^ 1'b0 ;
  assign n16619 = ( n16615 & n16616 ) | ( n16615 & n16618 ) | ( n16616 & n16618 ) ;
  assign n16622 = n12865 ^ n10115 ^ n4306 ;
  assign n16620 = n3163 ^ n2765 ^ n1421 ;
  assign n16621 = ( n1753 & n11347 ) | ( n1753 & ~n16620 ) | ( n11347 & ~n16620 ) ;
  assign n16623 = n16622 ^ n16621 ^ n5949 ;
  assign n16624 = n14739 ^ n6311 ^ n1500 ;
  assign n16625 = ( n7006 & ~n8653 ) | ( n7006 & n15514 ) | ( ~n8653 & n15514 ) ;
  assign n16626 = n16625 ^ n2221 ^ n234 ;
  assign n16629 = n15442 ^ n3895 ^ n2804 ;
  assign n16627 = ( n9732 & n10656 ) | ( n9732 & n11636 ) | ( n10656 & n11636 ) ;
  assign n16628 = ( n4192 & ~n9714 ) | ( n4192 & n16627 ) | ( ~n9714 & n16627 ) ;
  assign n16630 = n16629 ^ n16628 ^ n12449 ;
  assign n16631 = n14351 ^ n5101 ^ n3415 ;
  assign n16632 = ( n1672 & ~n5095 ) | ( n1672 & n5470 ) | ( ~n5095 & n5470 ) ;
  assign n16636 = n14708 ^ n8212 ^ 1'b0 ;
  assign n16633 = n5358 & ~n6340 ;
  assign n16634 = n16633 ^ n716 ^ 1'b0 ;
  assign n16635 = ( n1869 & n11731 ) | ( n1869 & ~n16634 ) | ( n11731 & ~n16634 ) ;
  assign n16637 = n16636 ^ n16635 ^ n8897 ;
  assign n16639 = ( ~n3883 & n5552 ) | ( ~n3883 & n11842 ) | ( n5552 & n11842 ) ;
  assign n16640 = ( n4074 & n9122 ) | ( n4074 & n16639 ) | ( n9122 & n16639 ) ;
  assign n16638 = n4783 | n14117 ;
  assign n16641 = n16640 ^ n16638 ^ 1'b0 ;
  assign n16642 = n5597 ^ n4695 ^ n2233 ;
  assign n16643 = n10060 ^ n8490 ^ 1'b0 ;
  assign n16644 = n10750 & ~n16643 ;
  assign n16645 = ( ~n7262 & n15426 ) | ( ~n7262 & n16644 ) | ( n15426 & n16644 ) ;
  assign n16646 = ( n10675 & ~n16642 ) | ( n10675 & n16645 ) | ( ~n16642 & n16645 ) ;
  assign n16647 = n3762 | n5108 ;
  assign n16648 = n16647 ^ n15575 ^ 1'b0 ;
  assign n16649 = n5390 & n8056 ;
  assign n16650 = n16649 ^ n1213 ^ 1'b0 ;
  assign n16651 = n16650 ^ n12331 ^ n2510 ;
  assign n16652 = ( n1893 & n13055 ) | ( n1893 & n16651 ) | ( n13055 & n16651 ) ;
  assign n16658 = ( n3971 & n4735 ) | ( n3971 & ~n13037 ) | ( n4735 & ~n13037 ) ;
  assign n16656 = n1419 & n3751 ;
  assign n16657 = ( n1834 & n5036 ) | ( n1834 & ~n16656 ) | ( n5036 & ~n16656 ) ;
  assign n16653 = ( n3748 & n6400 ) | ( n3748 & ~n11917 ) | ( n6400 & ~n11917 ) ;
  assign n16654 = n3271 | n16653 ;
  assign n16655 = n16654 ^ n3957 ^ 1'b0 ;
  assign n16659 = n16658 ^ n16657 ^ n16655 ;
  assign n16660 = ( n4258 & n9128 ) | ( n4258 & ~n14132 ) | ( n9128 & ~n14132 ) ;
  assign n16661 = x61 & n14614 ;
  assign n16662 = ~n277 & n16661 ;
  assign n16663 = ( ~n8681 & n16660 ) | ( ~n8681 & n16662 ) | ( n16660 & n16662 ) ;
  assign n16664 = n7740 ^ n6044 ^ 1'b0 ;
  assign n16665 = n6269 ^ n4388 ^ n1462 ;
  assign n16666 = ( n1842 & n8854 ) | ( n1842 & ~n16665 ) | ( n8854 & ~n16665 ) ;
  assign n16668 = n15549 ^ n10247 ^ n2749 ;
  assign n16667 = ( n3597 & n5412 ) | ( n3597 & n11499 ) | ( n5412 & n11499 ) ;
  assign n16669 = n16668 ^ n16667 ^ n1203 ;
  assign n16670 = n13423 ^ n6425 ^ n4870 ;
  assign n16671 = n8576 ^ n5263 ^ n2691 ;
  assign n16672 = n16671 ^ n12001 ^ n10363 ;
  assign n16673 = ( n2866 & ~n3676 ) | ( n2866 & n15137 ) | ( ~n3676 & n15137 ) ;
  assign n16674 = n16673 ^ n5315 ^ n1262 ;
  assign n16675 = n6524 ^ n3524 ^ n1939 ;
  assign n16676 = n4263 ^ n595 ^ 1'b0 ;
  assign n16677 = ( ~n4540 & n16675 ) | ( ~n4540 & n16676 ) | ( n16675 & n16676 ) ;
  assign n16678 = ( n5515 & ~n16674 ) | ( n5515 & n16677 ) | ( ~n16674 & n16677 ) ;
  assign n16679 = ( n8711 & n9299 ) | ( n8711 & ~n13355 ) | ( n9299 & ~n13355 ) ;
  assign n16680 = n5008 & n6960 ;
  assign n16681 = ( n3767 & n3902 ) | ( n3767 & n15610 ) | ( n3902 & n15610 ) ;
  assign n16682 = ( n14948 & n16680 ) | ( n14948 & n16681 ) | ( n16680 & n16681 ) ;
  assign n16686 = n7500 ^ n6806 ^ n5299 ;
  assign n16687 = n16686 ^ n9543 ^ n8795 ;
  assign n16683 = n5472 ^ n4394 ^ n680 ;
  assign n16684 = n16683 ^ n6981 ^ n4916 ;
  assign n16685 = ( n1667 & ~n11061 ) | ( n1667 & n16684 ) | ( ~n11061 & n16684 ) ;
  assign n16688 = n16687 ^ n16685 ^ n6061 ;
  assign n16689 = ( ~n2686 & n10001 ) | ( ~n2686 & n11255 ) | ( n10001 & n11255 ) ;
  assign n16690 = ( n14131 & n16370 ) | ( n14131 & n16689 ) | ( n16370 & n16689 ) ;
  assign n16691 = n2083 ^ n303 ^ 1'b0 ;
  assign n16692 = n9239 & ~n15363 ;
  assign n16693 = n4232 & n16692 ;
  assign n16694 = ( n4850 & ~n16691 ) | ( n4850 & n16693 ) | ( ~n16691 & n16693 ) ;
  assign n16695 = ( n903 & n10815 ) | ( n903 & ~n13266 ) | ( n10815 & ~n13266 ) ;
  assign n16696 = n16695 ^ n8496 ^ n5742 ;
  assign n16697 = ( n1264 & n2382 ) | ( n1264 & n14153 ) | ( n2382 & n14153 ) ;
  assign n16698 = ( n7391 & ~n7916 ) | ( n7391 & n16697 ) | ( ~n7916 & n16697 ) ;
  assign n16699 = ~n6698 & n16698 ;
  assign n16700 = n16699 ^ n8622 ^ n5434 ;
  assign n16701 = ~n4006 & n14100 ;
  assign n16702 = n15949 & n16701 ;
  assign n16703 = ( n2617 & ~n6877 ) | ( n2617 & n16702 ) | ( ~n6877 & n16702 ) ;
  assign n16704 = ( n2174 & ~n4356 ) | ( n2174 & n10037 ) | ( ~n4356 & n10037 ) ;
  assign n16705 = ( n6056 & ~n7420 ) | ( n6056 & n15232 ) | ( ~n7420 & n15232 ) ;
  assign n16706 = ~n12062 & n16705 ;
  assign n16707 = n9883 & n16706 ;
  assign n16708 = n14412 ^ n7611 ^ n3520 ;
  assign n16709 = ( ~n524 & n5885 ) | ( ~n524 & n14388 ) | ( n5885 & n14388 ) ;
  assign n16710 = ( n1290 & n2881 ) | ( n1290 & ~n11216 ) | ( n2881 & ~n11216 ) ;
  assign n16711 = n9129 ^ n6162 ^ n2076 ;
  assign n16712 = ( ~n13017 & n16710 ) | ( ~n13017 & n16711 ) | ( n16710 & n16711 ) ;
  assign n16713 = ( n906 & ~n3919 ) | ( n906 & n7546 ) | ( ~n3919 & n7546 ) ;
  assign n16714 = n5716 ^ n1329 ^ 1'b0 ;
  assign n16715 = ( ~n10681 & n15828 ) | ( ~n10681 & n16714 ) | ( n15828 & n16714 ) ;
  assign n16716 = ( n11552 & n16713 ) | ( n11552 & ~n16715 ) | ( n16713 & ~n16715 ) ;
  assign n16717 = ( x90 & ~n9168 ) | ( x90 & n13504 ) | ( ~n9168 & n13504 ) ;
  assign n16718 = n16717 ^ n5982 ^ n5705 ;
  assign n16719 = n13440 ^ n9894 ^ n5340 ;
  assign n16720 = ( n7654 & n12148 ) | ( n7654 & n16719 ) | ( n12148 & n16719 ) ;
  assign n16723 = n11887 ^ n6669 ^ 1'b0 ;
  assign n16724 = n11088 & n16723 ;
  assign n16721 = ( n242 & n1457 ) | ( n242 & ~n2862 ) | ( n1457 & ~n2862 ) ;
  assign n16722 = ( ~n1544 & n6642 ) | ( ~n1544 & n16721 ) | ( n6642 & n16721 ) ;
  assign n16725 = n16724 ^ n16722 ^ n5960 ;
  assign n16726 = n3734 ^ n2930 ^ n871 ;
  assign n16727 = n16726 ^ n13676 ^ n6443 ;
  assign n16728 = ( ~n13400 & n16725 ) | ( ~n13400 & n16727 ) | ( n16725 & n16727 ) ;
  assign n16731 = ( n2680 & n3459 ) | ( n2680 & n3471 ) | ( n3459 & n3471 ) ;
  assign n16732 = ( n6094 & n6404 ) | ( n6094 & n16731 ) | ( n6404 & n16731 ) ;
  assign n16729 = n5819 ^ n2001 ^ 1'b0 ;
  assign n16730 = n16729 ^ n10304 ^ n10179 ;
  assign n16733 = n16732 ^ n16730 ^ n3494 ;
  assign n16735 = ( n3371 & n7412 ) | ( n3371 & n11543 ) | ( n7412 & n11543 ) ;
  assign n16734 = ( x55 & n1148 ) | ( x55 & ~n6978 ) | ( n1148 & ~n6978 ) ;
  assign n16736 = n16735 ^ n16734 ^ n1857 ;
  assign n16737 = ( ~n6662 & n16629 ) | ( ~n6662 & n16736 ) | ( n16629 & n16736 ) ;
  assign n16738 = n145 | n9481 ;
  assign n16739 = n16738 ^ n14522 ^ n5188 ;
  assign n16740 = ( ~n2824 & n6407 ) | ( ~n2824 & n16739 ) | ( n6407 & n16739 ) ;
  assign n16741 = ( ~n3721 & n9269 ) | ( ~n3721 & n12708 ) | ( n9269 & n12708 ) ;
  assign n16742 = n11380 ^ n9538 ^ n1690 ;
  assign n16743 = n16742 ^ n12095 ^ n3988 ;
  assign n16744 = n16743 ^ n4142 ^ x12 ;
  assign n16745 = ( ~n5112 & n10023 ) | ( ~n5112 & n16744 ) | ( n10023 & n16744 ) ;
  assign n16746 = ( n15967 & ~n16741 ) | ( n15967 & n16745 ) | ( ~n16741 & n16745 ) ;
  assign n16747 = ( n1095 & ~n1655 ) | ( n1095 & n5257 ) | ( ~n1655 & n5257 ) ;
  assign n16748 = ( n856 & n8881 ) | ( n856 & n16747 ) | ( n8881 & n16747 ) ;
  assign n16749 = ( ~n1119 & n11499 ) | ( ~n1119 & n13564 ) | ( n11499 & n13564 ) ;
  assign n16750 = n5185 ^ n335 ^ 1'b0 ;
  assign n16751 = n6567 & ~n16750 ;
  assign n16752 = ( n7905 & ~n15502 ) | ( n7905 & n16751 ) | ( ~n15502 & n16751 ) ;
  assign n16753 = ( n3111 & n3463 ) | ( n3111 & ~n5389 ) | ( n3463 & ~n5389 ) ;
  assign n16754 = n16753 ^ n12576 ^ n9425 ;
  assign n16755 = n16754 ^ n5304 ^ 1'b0 ;
  assign n16756 = ( n8385 & ~n16752 ) | ( n8385 & n16755 ) | ( ~n16752 & n16755 ) ;
  assign n16757 = n16756 ^ n9238 ^ n843 ;
  assign n16758 = n7249 ^ n5961 ^ n2360 ;
  assign n16759 = n16758 ^ n12226 ^ n440 ;
  assign n16760 = n6361 & ~n14805 ;
  assign n16761 = n16760 ^ n3628 ^ 1'b0 ;
  assign n16762 = ( n578 & n7909 ) | ( n578 & n15587 ) | ( n7909 & n15587 ) ;
  assign n16764 = ( n3349 & ~n8304 ) | ( n3349 & n11661 ) | ( ~n8304 & n11661 ) ;
  assign n16763 = n1628 ^ n740 ^ 1'b0 ;
  assign n16765 = n16764 ^ n16763 ^ n596 ;
  assign n16766 = n6618 ^ n1985 ^ 1'b0 ;
  assign n16767 = n7282 | n16766 ;
  assign n16768 = n16767 ^ n6604 ^ 1'b0 ;
  assign n16769 = n6378 | n12165 ;
  assign n16770 = n1863 ^ n1102 ^ n550 ;
  assign n16771 = n16770 ^ n7435 ^ n953 ;
  assign n16772 = n16771 ^ n7124 ^ n4756 ;
  assign n16773 = n14795 ^ n14142 ^ n11071 ;
  assign n16774 = ( n2638 & n10261 ) | ( n2638 & ~n16773 ) | ( n10261 & ~n16773 ) ;
  assign n16776 = n6415 ^ n4403 ^ 1'b0 ;
  assign n16777 = n4728 | n16776 ;
  assign n16775 = n14338 ^ n6922 ^ n427 ;
  assign n16778 = n16777 ^ n16775 ^ n5102 ;
  assign n16779 = n6459 ^ n5755 ^ n2368 ;
  assign n16780 = n16779 ^ n12757 ^ n6614 ;
  assign n16781 = n2504 ^ n264 ^ 1'b0 ;
  assign n16782 = n5919 ^ n2179 ^ n1154 ;
  assign n16783 = n14347 ^ n13657 ^ n461 ;
  assign n16784 = ( n6289 & ~n16022 ) | ( n6289 & n16783 ) | ( ~n16022 & n16783 ) ;
  assign n16785 = ( n8626 & n16782 ) | ( n8626 & n16784 ) | ( n16782 & n16784 ) ;
  assign n16786 = ~n11933 & n14292 ;
  assign n16787 = n8424 & n16786 ;
  assign n16788 = ( n12448 & n16785 ) | ( n12448 & n16787 ) | ( n16785 & n16787 ) ;
  assign n16789 = ( n5734 & n16781 ) | ( n5734 & ~n16788 ) | ( n16781 & ~n16788 ) ;
  assign n16790 = ( n7879 & ~n10586 ) | ( n7879 & n13423 ) | ( ~n10586 & n13423 ) ;
  assign n16791 = n10305 ^ n7097 ^ n6947 ;
  assign n16792 = ( n16669 & ~n16790 ) | ( n16669 & n16791 ) | ( ~n16790 & n16791 ) ;
  assign n16793 = n8988 ^ n4019 ^ 1'b0 ;
  assign n16794 = n15276 ^ n12418 ^ n10099 ;
  assign n16795 = n16794 ^ n11375 ^ n10816 ;
  assign n16796 = ~n4996 & n15463 ;
  assign n16797 = ( n629 & ~n7309 ) | ( n629 & n16796 ) | ( ~n7309 & n16796 ) ;
  assign n16798 = n14173 & n16797 ;
  assign n16799 = ( ~n1907 & n6492 ) | ( ~n1907 & n12946 ) | ( n6492 & n12946 ) ;
  assign n16800 = n8968 ^ n2472 ^ n1056 ;
  assign n16801 = ( n1785 & ~n5409 ) | ( n1785 & n10884 ) | ( ~n5409 & n10884 ) ;
  assign n16802 = ( n9727 & ~n10759 ) | ( n9727 & n16801 ) | ( ~n10759 & n16801 ) ;
  assign n16804 = n11350 ^ n290 ^ 1'b0 ;
  assign n16805 = ( n6751 & n13493 ) | ( n6751 & ~n16804 ) | ( n13493 & ~n16804 ) ;
  assign n16806 = ( n3008 & n13107 ) | ( n3008 & n16805 ) | ( n13107 & n16805 ) ;
  assign n16803 = n5288 | n11060 ;
  assign n16807 = n16806 ^ n16803 ^ 1'b0 ;
  assign n16808 = n16475 ^ n12808 ^ n7927 ;
  assign n16809 = n16808 ^ n8883 ^ n3416 ;
  assign n16810 = n15085 ^ n13278 ^ n8485 ;
  assign n16811 = n16810 ^ n10879 ^ n10747 ;
  assign n16812 = n4755 ^ n4645 ^ n3447 ;
  assign n16813 = ( n9574 & n12660 ) | ( n9574 & n16812 ) | ( n12660 & n16812 ) ;
  assign n16814 = ( n5773 & ~n7328 ) | ( n5773 & n9847 ) | ( ~n7328 & n9847 ) ;
  assign n16815 = n5754 | n16814 ;
  assign n16817 = ( n3288 & n4356 ) | ( n3288 & ~n5550 ) | ( n4356 & ~n5550 ) ;
  assign n16816 = n9634 ^ n8381 ^ n3676 ;
  assign n16818 = n16817 ^ n16816 ^ 1'b0 ;
  assign n16819 = ( n11810 & n12142 ) | ( n11810 & n16818 ) | ( n12142 & n16818 ) ;
  assign n16820 = n11643 ^ n5974 ^ 1'b0 ;
  assign n16821 = ( n894 & ~n2355 ) | ( n894 & n9810 ) | ( ~n2355 & n9810 ) ;
  assign n16822 = n6748 ^ n6165 ^ n1797 ;
  assign n16823 = n16822 ^ n4834 ^ n2903 ;
  assign n16824 = ( n1334 & ~n1787 ) | ( n1334 & n13324 ) | ( ~n1787 & n13324 ) ;
  assign n16825 = ( n639 & n6098 ) | ( n639 & ~n16824 ) | ( n6098 & ~n16824 ) ;
  assign n16826 = ( n11531 & ~n12734 ) | ( n11531 & n16825 ) | ( ~n12734 & n16825 ) ;
  assign n16827 = ( n772 & ~n7310 ) | ( n772 & n9451 ) | ( ~n7310 & n9451 ) ;
  assign n16828 = ( n506 & n13124 ) | ( n506 & n16827 ) | ( n13124 & n16827 ) ;
  assign n16829 = ( n4001 & ~n11689 ) | ( n4001 & n16828 ) | ( ~n11689 & n16828 ) ;
  assign n16830 = ( ~n5482 & n14333 ) | ( ~n5482 & n16829 ) | ( n14333 & n16829 ) ;
  assign n16831 = ( n5675 & n11805 ) | ( n5675 & n13760 ) | ( n11805 & n13760 ) ;
  assign n16832 = n4942 ^ n2726 ^ n1907 ;
  assign n16833 = n10408 ^ n5039 ^ x126 ;
  assign n16834 = ( x20 & ~n5136 ) | ( x20 & n16833 ) | ( ~n5136 & n16833 ) ;
  assign n16835 = n10937 ^ n6294 ^ n5931 ;
  assign n16836 = n16835 ^ n13394 ^ n3692 ;
  assign n16837 = ( n4313 & ~n16834 ) | ( n4313 & n16836 ) | ( ~n16834 & n16836 ) ;
  assign n16838 = n16837 ^ n13843 ^ n4139 ;
  assign n16839 = n649 & n16838 ;
  assign n16840 = n16839 ^ n16494 ^ 1'b0 ;
  assign n16841 = ( ~n16831 & n16832 ) | ( ~n16831 & n16840 ) | ( n16832 & n16840 ) ;
  assign n16842 = ( ~n2256 & n7325 ) | ( ~n2256 & n16223 ) | ( n7325 & n16223 ) ;
  assign n16843 = ( n1462 & n4454 ) | ( n1462 & ~n16842 ) | ( n4454 & ~n16842 ) ;
  assign n16844 = ( x110 & ~n1060 ) | ( x110 & n4288 ) | ( ~n1060 & n4288 ) ;
  assign n16845 = n16844 ^ n7431 ^ n4508 ;
  assign n16846 = n13625 & ~n16845 ;
  assign n16847 = ~n8617 & n16846 ;
  assign n16848 = n16847 ^ n7669 ^ n3783 ;
  assign n16849 = n12242 ^ n9895 ^ n6165 ;
  assign n16850 = n8663 & n16849 ;
  assign n16851 = ~n13133 & n16850 ;
  assign n16852 = n16851 ^ n13136 ^ n1665 ;
  assign n16854 = n6296 ^ n2377 ^ 1'b0 ;
  assign n16853 = ( ~n2197 & n2276 ) | ( ~n2197 & n3250 ) | ( n2276 & n3250 ) ;
  assign n16855 = n16854 ^ n16853 ^ n4454 ;
  assign n16856 = ( ~n2755 & n15566 ) | ( ~n2755 & n16855 ) | ( n15566 & n16855 ) ;
  assign n16857 = n6897 ^ n4624 ^ n3009 ;
  assign n16858 = n12448 ^ n4702 ^ 1'b0 ;
  assign n16859 = n16857 & n16858 ;
  assign n16860 = n16859 ^ n12857 ^ n1826 ;
  assign n16861 = n14436 ^ n2908 ^ n1954 ;
  assign n16862 = n3175 ^ n1938 ^ 1'b0 ;
  assign n16863 = n6066 & n16862 ;
  assign n16864 = ( n4652 & n15770 ) | ( n4652 & ~n16863 ) | ( n15770 & ~n16863 ) ;
  assign n16865 = ( n1387 & ~n16861 ) | ( n1387 & n16864 ) | ( ~n16861 & n16864 ) ;
  assign n16866 = ( n3830 & n16860 ) | ( n3830 & ~n16865 ) | ( n16860 & ~n16865 ) ;
  assign n16867 = n16866 ^ n6055 ^ n256 ;
  assign n16870 = ~n3716 & n14842 ;
  assign n16868 = n7323 ^ n5971 ^ n641 ;
  assign n16869 = ~n8514 & n16868 ;
  assign n16871 = n16870 ^ n16869 ^ 1'b0 ;
  assign n16872 = n16118 ^ n3366 ^ 1'b0 ;
  assign n16873 = n16871 & n16872 ;
  assign n16874 = ( n2757 & n3859 ) | ( n2757 & ~n9258 ) | ( n3859 & ~n9258 ) ;
  assign n16875 = n16368 ^ n12759 ^ n5696 ;
  assign n16876 = n16875 ^ n6681 ^ n5564 ;
  assign n16877 = n9864 ^ n6965 ^ n6079 ;
  assign n16878 = n10461 ^ n9610 ^ n8718 ;
  assign n16880 = ( ~n263 & n3855 ) | ( ~n263 & n10060 ) | ( n3855 & n10060 ) ;
  assign n16881 = n14250 ^ n6965 ^ 1'b0 ;
  assign n16882 = ~n16880 & n16881 ;
  assign n16879 = n12072 ^ n5620 ^ n3091 ;
  assign n16883 = n16882 ^ n16879 ^ n14008 ;
  assign n16884 = ( n7443 & n11442 ) | ( n7443 & n13855 ) | ( n11442 & n13855 ) ;
  assign n16885 = n11885 ^ n6361 ^ n1532 ;
  assign n16886 = n9749 & n16885 ;
  assign n16887 = ~n10699 & n16886 ;
  assign n16888 = ( n2283 & n4438 ) | ( n2283 & ~n16887 ) | ( n4438 & ~n16887 ) ;
  assign n16889 = ~n16884 & n16888 ;
  assign n16890 = ~n10753 & n16889 ;
  assign n16891 = n2143 | n10658 ;
  assign n16892 = n16891 ^ n6770 ^ n3725 ;
  assign n16893 = ( n2143 & n5012 ) | ( n2143 & n13855 ) | ( n5012 & n13855 ) ;
  assign n16894 = ( n5677 & ~n10464 ) | ( n5677 & n16893 ) | ( ~n10464 & n16893 ) ;
  assign n16895 = n6616 ^ n2269 ^ n1008 ;
  assign n16896 = ( ~n7377 & n15555 ) | ( ~n7377 & n16895 ) | ( n15555 & n16895 ) ;
  assign n16897 = ( ~n11043 & n11570 ) | ( ~n11043 & n16896 ) | ( n11570 & n16896 ) ;
  assign n16898 = n5122 ^ n1917 ^ 1'b0 ;
  assign n16899 = n14361 ^ n11569 ^ n10513 ;
  assign n16900 = ( n3133 & n16898 ) | ( n3133 & ~n16899 ) | ( n16898 & ~n16899 ) ;
  assign n16906 = ( ~n612 & n3698 ) | ( ~n612 & n16814 ) | ( n3698 & n16814 ) ;
  assign n16904 = n5239 ^ n4846 ^ n4684 ;
  assign n16901 = n13059 ^ n3362 ^ n1678 ;
  assign n16902 = ( n2201 & n3261 ) | ( n2201 & ~n16901 ) | ( n3261 & ~n16901 ) ;
  assign n16903 = ( ~n10099 & n11725 ) | ( ~n10099 & n16902 ) | ( n11725 & n16902 ) ;
  assign n16905 = n16904 ^ n16903 ^ n8191 ;
  assign n16907 = n16906 ^ n16905 ^ 1'b0 ;
  assign n16908 = n7600 & ~n16907 ;
  assign n16909 = ~n6583 & n16908 ;
  assign n16913 = n6894 ^ n1566 ^ n948 ;
  assign n16910 = n16525 ^ n9491 ^ n4996 ;
  assign n16911 = ( ~x120 & n6546 ) | ( ~x120 & n16910 ) | ( n6546 & n16910 ) ;
  assign n16912 = n16911 ^ n8193 ^ n3725 ;
  assign n16914 = n16913 ^ n16912 ^ n14061 ;
  assign n16915 = ( n6613 & n11618 ) | ( n6613 & n15642 ) | ( n11618 & n15642 ) ;
  assign n16916 = ( n4201 & n6211 ) | ( n4201 & n10095 ) | ( n6211 & n10095 ) ;
  assign n16917 = n16916 ^ n14249 ^ n4812 ;
  assign n16918 = ( ~n13415 & n14751 ) | ( ~n13415 & n16917 ) | ( n14751 & n16917 ) ;
  assign n16919 = n16918 ^ n5154 ^ 1'b0 ;
  assign n16920 = ( ~n1790 & n2353 ) | ( ~n1790 & n14716 ) | ( n2353 & n14716 ) ;
  assign n16921 = x6 & n7144 ;
  assign n16922 = n16921 ^ n7739 ^ 1'b0 ;
  assign n16923 = n16922 ^ n14931 ^ n3517 ;
  assign n16924 = n16923 ^ n11135 ^ n9101 ;
  assign n16927 = ( ~n5693 & n7924 ) | ( ~n5693 & n8754 ) | ( n7924 & n8754 ) ;
  assign n16926 = n10929 ^ n9178 ^ n137 ;
  assign n16925 = ( ~n670 & n5934 ) | ( ~n670 & n7515 ) | ( n5934 & n7515 ) ;
  assign n16928 = n16927 ^ n16926 ^ n16925 ;
  assign n16929 = n5349 | n16928 ;
  assign n16930 = ( n817 & n6177 ) | ( n817 & n7155 ) | ( n6177 & n7155 ) ;
  assign n16931 = ( n3493 & n6972 ) | ( n3493 & n16930 ) | ( n6972 & n16930 ) ;
  assign n16932 = n2004 & ~n16931 ;
  assign n16933 = ~n15020 & n16932 ;
  assign n16934 = n16933 ^ n10572 ^ n8626 ;
  assign n16935 = ( n493 & n10886 ) | ( n493 & ~n16934 ) | ( n10886 & ~n16934 ) ;
  assign n16936 = ( n625 & n11222 ) | ( n625 & ~n16393 ) | ( n11222 & ~n16393 ) ;
  assign n16937 = n8704 ^ n5733 ^ n3425 ;
  assign n16938 = ( n5900 & n6668 ) | ( n5900 & n16031 ) | ( n6668 & n16031 ) ;
  assign n16939 = ( n9905 & n16937 ) | ( n9905 & ~n16938 ) | ( n16937 & ~n16938 ) ;
  assign n16940 = n250 & ~n16939 ;
  assign n16941 = ~n181 & n16199 ;
  assign n16942 = ~n10929 & n16941 ;
  assign n16943 = ( n7311 & ~n7337 ) | ( n7311 & n14968 ) | ( ~n7337 & n14968 ) ;
  assign n16944 = n11541 ^ n11132 ^ n6579 ;
  assign n16945 = n16944 ^ n10199 ^ n2976 ;
  assign n16946 = ( n1496 & n16943 ) | ( n1496 & ~n16945 ) | ( n16943 & ~n16945 ) ;
  assign n16947 = ( n12784 & ~n13412 ) | ( n12784 & n14688 ) | ( ~n13412 & n14688 ) ;
  assign n16948 = ( n1298 & n9237 ) | ( n1298 & n16947 ) | ( n9237 & n16947 ) ;
  assign n16950 = ( n623 & n1964 ) | ( n623 & ~n3416 ) | ( n1964 & ~n3416 ) ;
  assign n16951 = n16950 ^ n12702 ^ n6313 ;
  assign n16949 = ( n2748 & n7266 ) | ( n2748 & n12229 ) | ( n7266 & n12229 ) ;
  assign n16952 = n16951 ^ n16949 ^ n12275 ;
  assign n16953 = n15348 ^ n4650 ^ n4242 ;
  assign n16954 = n7233 & ~n16953 ;
  assign n16955 = n16954 ^ n5113 ^ n1435 ;
  assign n16956 = n4112 ^ n3777 ^ 1'b0 ;
  assign n16957 = ~n3035 & n13171 ;
  assign n16958 = n16957 ^ n4870 ^ 1'b0 ;
  assign n16959 = ( ~n15103 & n15737 ) | ( ~n15103 & n16585 ) | ( n15737 & n16585 ) ;
  assign n16960 = ( n11193 & ~n11731 ) | ( n11193 & n16959 ) | ( ~n11731 & n16959 ) ;
  assign n16961 = n11460 ^ n1747 ^ n1732 ;
  assign n16962 = ( x98 & n9339 ) | ( x98 & ~n16961 ) | ( n9339 & ~n16961 ) ;
  assign n16963 = n16962 ^ n1680 ^ n541 ;
  assign n16964 = ( n997 & n10716 ) | ( n997 & ~n12413 ) | ( n10716 & ~n12413 ) ;
  assign n16966 = n473 & n1796 ;
  assign n16967 = n16966 ^ n2089 ^ 1'b0 ;
  assign n16968 = n16967 ^ n4807 ^ n1737 ;
  assign n16965 = n3195 & ~n8689 ;
  assign n16969 = n16968 ^ n16965 ^ 1'b0 ;
  assign n16970 = n16057 & n16969 ;
  assign n16971 = n16970 ^ n14887 ^ 1'b0 ;
  assign n16972 = n11861 ^ n9069 ^ n8398 ;
  assign n16973 = ( n14521 & n16971 ) | ( n14521 & ~n16972 ) | ( n16971 & ~n16972 ) ;
  assign n16975 = n11804 ^ n10969 ^ 1'b0 ;
  assign n16976 = n3252 & ~n16975 ;
  assign n16974 = n12463 ^ n1406 ^ n1241 ;
  assign n16977 = n16976 ^ n16974 ^ n14456 ;
  assign n16978 = ( n4488 & n4953 ) | ( n4488 & ~n11636 ) | ( n4953 & ~n11636 ) ;
  assign n16979 = n8240 | n16978 ;
  assign n16980 = n13023 ^ n7242 ^ n5420 ;
  assign n16981 = ( n10365 & n16979 ) | ( n10365 & ~n16980 ) | ( n16979 & ~n16980 ) ;
  assign n16982 = ~n5197 & n7218 ;
  assign n16983 = ( n2227 & n10886 ) | ( n2227 & ~n16982 ) | ( n10886 & ~n16982 ) ;
  assign n16984 = ( ~n2679 & n10441 ) | ( ~n2679 & n16983 ) | ( n10441 & n16983 ) ;
  assign n16985 = n626 | n3390 ;
  assign n16986 = n3789 | n16985 ;
  assign n16987 = ( n3757 & n9079 ) | ( n3757 & n16052 ) | ( n9079 & n16052 ) ;
  assign n16988 = ( ~n1340 & n2645 ) | ( ~n1340 & n3297 ) | ( n2645 & n3297 ) ;
  assign n16989 = n16988 ^ n3547 ^ n3449 ;
  assign n16990 = n16989 ^ n11323 ^ n4043 ;
  assign n16991 = ( ~n9953 & n16987 ) | ( ~n9953 & n16990 ) | ( n16987 & n16990 ) ;
  assign n16992 = ( n4097 & n4230 ) | ( n4097 & ~n15089 ) | ( n4230 & ~n15089 ) ;
  assign n16993 = n16992 ^ n14651 ^ n3127 ;
  assign n16994 = ( ~n2889 & n11466 ) | ( ~n2889 & n15656 ) | ( n11466 & n15656 ) ;
  assign n16995 = n13770 ^ n7088 ^ n2283 ;
  assign n16996 = n10893 ^ n8896 ^ n3703 ;
  assign n16997 = ( n16223 & ~n16995 ) | ( n16223 & n16996 ) | ( ~n16995 & n16996 ) ;
  assign n16998 = ~n5608 & n16997 ;
  assign n16999 = n14007 ^ n6436 ^ n2531 ;
  assign n17000 = n11318 ^ n9588 ^ n910 ;
  assign n17001 = n17000 ^ n1523 ^ n705 ;
  assign n17002 = ( n3908 & n16999 ) | ( n3908 & n17001 ) | ( n16999 & n17001 ) ;
  assign n17003 = n9135 ^ n8959 ^ n8287 ;
  assign n17004 = n17003 ^ n11914 ^ n855 ;
  assign n17006 = n8096 ^ n7639 ^ n2505 ;
  assign n17005 = n1569 & ~n14332 ;
  assign n17007 = n17006 ^ n17005 ^ n4423 ;
  assign n17008 = n6765 & n8070 ;
  assign n17011 = n8710 ^ n5133 ^ 1'b0 ;
  assign n17009 = n7465 | n14348 ;
  assign n17010 = n6092 & ~n17009 ;
  assign n17012 = n17011 ^ n17010 ^ n13411 ;
  assign n17013 = ( n5566 & n17008 ) | ( n5566 & n17012 ) | ( n17008 & n17012 ) ;
  assign n17014 = ( ~x15 & n10127 ) | ( ~x15 & n10812 ) | ( n10127 & n10812 ) ;
  assign n17015 = n5088 ^ n1893 ^ 1'b0 ;
  assign n17016 = n17015 ^ n9532 ^ n3137 ;
  assign n17017 = ( n4113 & n4158 ) | ( n4113 & ~n17016 ) | ( n4158 & ~n17016 ) ;
  assign n17020 = n5398 ^ n4782 ^ n2612 ;
  assign n17018 = ( n2175 & n2472 ) | ( n2175 & n13828 ) | ( n2472 & n13828 ) ;
  assign n17019 = ( ~n927 & n16547 ) | ( ~n927 & n17018 ) | ( n16547 & n17018 ) ;
  assign n17021 = n17020 ^ n17019 ^ n11864 ;
  assign n17022 = n15396 ^ n14632 ^ 1'b0 ;
  assign n17023 = n17022 ^ n15522 ^ n3267 ;
  assign n17024 = n14039 ^ n6036 ^ n3218 ;
  assign n17025 = ( ~n2461 & n7292 ) | ( ~n2461 & n17024 ) | ( n7292 & n17024 ) ;
  assign n17026 = ( ~n8742 & n12132 ) | ( ~n8742 & n17025 ) | ( n12132 & n17025 ) ;
  assign n17027 = ( n619 & n16596 ) | ( n619 & ~n17026 ) | ( n16596 & ~n17026 ) ;
  assign n17028 = n11267 ^ n4764 ^ n848 ;
  assign n17029 = ( n3893 & n5704 ) | ( n3893 & n17028 ) | ( n5704 & n17028 ) ;
  assign n17030 = n6638 & ~n17029 ;
  assign n17031 = n17030 ^ n2987 ^ 1'b0 ;
  assign n17032 = n17031 ^ n16997 ^ n1334 ;
  assign n17033 = n10111 ^ n2327 ^ 1'b0 ;
  assign n17034 = n8138 | n17033 ;
  assign n17036 = ( n3519 & n3761 ) | ( n3519 & ~n5835 ) | ( n3761 & ~n5835 ) ;
  assign n17035 = n6219 | n13741 ;
  assign n17037 = n17036 ^ n17035 ^ n1871 ;
  assign n17038 = ~n5621 & n17037 ;
  assign n17039 = ( n564 & ~n3476 ) | ( n564 & n9316 ) | ( ~n3476 & n9316 ) ;
  assign n17040 = n17039 ^ n11543 ^ n7351 ;
  assign n17041 = ( n2855 & ~n4510 ) | ( n2855 & n17040 ) | ( ~n4510 & n17040 ) ;
  assign n17042 = n17041 ^ n10861 ^ n6238 ;
  assign n17043 = ( n10467 & n12195 ) | ( n10467 & n15036 ) | ( n12195 & n15036 ) ;
  assign n17044 = ( n6922 & ~n8886 ) | ( n6922 & n10689 ) | ( ~n8886 & n10689 ) ;
  assign n17045 = n17044 ^ n16891 ^ n14307 ;
  assign n17046 = ( ~n13943 & n14653 ) | ( ~n13943 & n17045 ) | ( n14653 & n17045 ) ;
  assign n17047 = n12095 ^ n9091 ^ n4933 ;
  assign n17048 = n2170 & n17047 ;
  assign n17049 = ~n4327 & n4519 ;
  assign n17050 = n17049 ^ n15288 ^ n5536 ;
  assign n17052 = n9077 ^ n4587 ^ n1377 ;
  assign n17051 = n14069 ^ n8996 ^ 1'b0 ;
  assign n17053 = n17052 ^ n17051 ^ n11418 ;
  assign n17054 = n8872 ^ n4447 ^ n492 ;
  assign n17055 = ( n245 & n3694 ) | ( n245 & ~n17054 ) | ( n3694 & ~n17054 ) ;
  assign n17056 = n4294 & n17055 ;
  assign n17057 = n11506 & n17056 ;
  assign n17058 = ~n6799 & n17057 ;
  assign n17059 = n5738 ^ n3652 ^ 1'b0 ;
  assign n17060 = n2790 & n17059 ;
  assign n17061 = n17060 ^ n9519 ^ n7909 ;
  assign n17062 = n17061 ^ n14153 ^ n11043 ;
  assign n17063 = n17062 ^ n11016 ^ n2206 ;
  assign n17066 = ( n608 & n3801 ) | ( n608 & ~n8343 ) | ( n3801 & ~n8343 ) ;
  assign n17064 = n9682 ^ n4848 ^ 1'b0 ;
  assign n17065 = n2730 | n17064 ;
  assign n17067 = n17066 ^ n17065 ^ n8850 ;
  assign n17068 = ( ~n3356 & n5737 ) | ( ~n3356 & n8159 ) | ( n5737 & n8159 ) ;
  assign n17069 = n17068 ^ n12355 ^ n3247 ;
  assign n17071 = ( n2268 & ~n8587 ) | ( n2268 & n10503 ) | ( ~n8587 & n10503 ) ;
  assign n17070 = n8839 ^ n7556 ^ n1175 ;
  assign n17072 = n17071 ^ n17070 ^ n2250 ;
  assign n17073 = n1968 | n5545 ;
  assign n17074 = n17073 ^ n9360 ^ 1'b0 ;
  assign n17075 = ( n5659 & ~n5919 ) | ( n5659 & n17074 ) | ( ~n5919 & n17074 ) ;
  assign n17076 = n17075 ^ n13965 ^ n3648 ;
  assign n17077 = ( n2316 & n2509 ) | ( n2316 & ~n17076 ) | ( n2509 & ~n17076 ) ;
  assign n17078 = ( n3274 & n10848 ) | ( n3274 & ~n17077 ) | ( n10848 & ~n17077 ) ;
  assign n17079 = n11187 ^ n10319 ^ n5195 ;
  assign n17080 = n10829 ^ n1354 ^ n297 ;
  assign n17081 = n13483 ^ n12898 ^ n5182 ;
  assign n17082 = n17081 ^ n16927 ^ n1797 ;
  assign n17083 = n14710 ^ n7064 ^ n4530 ;
  assign n17084 = ~n2819 & n5090 ;
  assign n17085 = n14006 & n17084 ;
  assign n17086 = ( n6499 & n13263 ) | ( n6499 & n15795 ) | ( n13263 & n15795 ) ;
  assign n17087 = ( n1614 & n4183 ) | ( n1614 & ~n17086 ) | ( n4183 & ~n17086 ) ;
  assign n17088 = n2671 & n17087 ;
  assign n17089 = n17085 & n17088 ;
  assign n17092 = n16012 ^ n1434 ^ n223 ;
  assign n17090 = n3430 ^ n1455 ^ n1064 ;
  assign n17091 = n17090 ^ n14320 ^ n4637 ;
  assign n17093 = n17092 ^ n17091 ^ n811 ;
  assign n17094 = ( x102 & n5611 ) | ( x102 & n17049 ) | ( n5611 & n17049 ) ;
  assign n17097 = n12472 ^ n4641 ^ n3669 ;
  assign n17096 = n10881 ^ n9020 ^ n3044 ;
  assign n17095 = n2913 | n9486 ;
  assign n17098 = n17097 ^ n17096 ^ n17095 ;
  assign n17099 = n1267 | n7617 ;
  assign n17100 = n17099 ^ n7743 ^ 1'b0 ;
  assign n17101 = n15847 ^ n3533 ^ n2288 ;
  assign n17102 = ~n3090 & n7938 ;
  assign n17103 = n3244 & ~n17102 ;
  assign n17104 = ~n17101 & n17103 ;
  assign n17105 = n8514 ^ n6896 ^ n764 ;
  assign n17106 = n17105 ^ n4101 ^ n3975 ;
  assign n17107 = n1232 & ~n2826 ;
  assign n17108 = n17107 ^ n7937 ^ 1'b0 ;
  assign n17109 = n17108 ^ n15651 ^ n4445 ;
  assign n17110 = ( n9964 & n10432 ) | ( n9964 & ~n16342 ) | ( n10432 & ~n16342 ) ;
  assign n17111 = n17110 ^ n16547 ^ 1'b0 ;
  assign n17112 = n9091 ^ n2310 ^ 1'b0 ;
  assign n17113 = n17112 ^ n11479 ^ n1162 ;
  assign n17114 = n17113 ^ n825 ^ n339 ;
  assign n17115 = n15885 ^ n7925 ^ n4055 ;
  assign n17116 = ( n644 & n2082 ) | ( n644 & ~n7109 ) | ( n2082 & ~n7109 ) ;
  assign n17117 = n17116 ^ n6915 ^ 1'b0 ;
  assign n17118 = n13217 | n17117 ;
  assign n17119 = ( n2801 & n3343 ) | ( n2801 & n10068 ) | ( n3343 & n10068 ) ;
  assign n17120 = ( ~n1154 & n15442 ) | ( ~n1154 & n17119 ) | ( n15442 & n17119 ) ;
  assign n17121 = n7226 ^ n3695 ^ n2378 ;
  assign n17122 = n17121 ^ n8859 ^ 1'b0 ;
  assign n17123 = n5047 | n17122 ;
  assign n17124 = ( n4520 & n5514 ) | ( n4520 & ~n17123 ) | ( n5514 & ~n17123 ) ;
  assign n17125 = n5885 ^ n3233 ^ x74 ;
  assign n17126 = ( n9593 & ~n16452 ) | ( n9593 & n17125 ) | ( ~n16452 & n17125 ) ;
  assign n17127 = n13710 ^ n9447 ^ n5189 ;
  assign n17128 = n3572 & ~n6197 ;
  assign n17129 = n17128 ^ n744 ^ x6 ;
  assign n17130 = n17129 ^ n5154 ^ n5005 ;
  assign n17131 = n17130 ^ n13339 ^ 1'b0 ;
  assign n17132 = ( n3722 & n5939 ) | ( n3722 & n8677 ) | ( n5939 & n8677 ) ;
  assign n17133 = n17092 ^ n15380 ^ n3073 ;
  assign n17134 = ( n8622 & n9307 ) | ( n8622 & ~n17133 ) | ( n9307 & ~n17133 ) ;
  assign n17135 = n17134 ^ n7118 ^ n1476 ;
  assign n17136 = ( n15558 & n17132 ) | ( n15558 & ~n17135 ) | ( n17132 & ~n17135 ) ;
  assign n17137 = ( n7481 & n10234 ) | ( n7481 & ~n15667 ) | ( n10234 & ~n15667 ) ;
  assign n17138 = n15614 ^ n4796 ^ 1'b0 ;
  assign n17139 = n17138 ^ n4344 ^ n3493 ;
  assign n17140 = n8932 ^ n7822 ^ n3938 ;
  assign n17141 = n8530 | n11093 ;
  assign n17142 = n12921 ^ n4861 ^ n782 ;
  assign n17143 = ( n692 & n1566 ) | ( n692 & n2228 ) | ( n1566 & n2228 ) ;
  assign n17144 = ( n1452 & n17142 ) | ( n1452 & ~n17143 ) | ( n17142 & ~n17143 ) ;
  assign n17145 = n11730 ^ n6974 ^ n5748 ;
  assign n17146 = ( n11959 & ~n15848 ) | ( n11959 & n17145 ) | ( ~n15848 & n17145 ) ;
  assign n17147 = n12655 & n12676 ;
  assign n17148 = n17147 ^ n13688 ^ 1'b0 ;
  assign n17149 = n17148 ^ n16734 ^ n7607 ;
  assign n17151 = ( n3571 & ~n6685 ) | ( n3571 & n7717 ) | ( ~n6685 & n7717 ) ;
  assign n17150 = n13249 ^ n11924 ^ n8595 ;
  assign n17152 = n17151 ^ n17150 ^ n4414 ;
  assign n17154 = n9029 ^ n658 ^ x29 ;
  assign n17155 = n17154 ^ n6669 ^ 1'b0 ;
  assign n17153 = ( n1392 & ~n5917 ) | ( n1392 & n12085 ) | ( ~n5917 & n12085 ) ;
  assign n17156 = n17155 ^ n17153 ^ n13250 ;
  assign n17157 = n17156 ^ n4876 ^ 1'b0 ;
  assign n17158 = ( n3019 & n7553 ) | ( n3019 & n14063 ) | ( n7553 & n14063 ) ;
  assign n17159 = n17158 ^ n13397 ^ 1'b0 ;
  assign n17160 = ( ~n4796 & n8283 ) | ( ~n4796 & n17000 ) | ( n8283 & n17000 ) ;
  assign n17161 = n11785 ^ n2937 ^ 1'b0 ;
  assign n17162 = n11576 ^ n8853 ^ n7469 ;
  assign n17163 = n17162 ^ n13493 ^ 1'b0 ;
  assign n17164 = ( x101 & n2392 ) | ( x101 & ~n9939 ) | ( n2392 & ~n9939 ) ;
  assign n17165 = n11211 & n17164 ;
  assign n17166 = ~n1088 & n17165 ;
  assign n17167 = n17166 ^ n3822 ^ n3284 ;
  assign n17168 = ( ~n8513 & n12379 ) | ( ~n8513 & n17167 ) | ( n12379 & n17167 ) ;
  assign n17169 = n9366 ^ n5742 ^ n1836 ;
  assign n17170 = n11912 ^ n9128 ^ n3392 ;
  assign n17171 = ~n2256 & n17170 ;
  assign n17172 = n17171 ^ n7445 ^ 1'b0 ;
  assign n17173 = ( n2737 & n17169 ) | ( n2737 & n17172 ) | ( n17169 & n17172 ) ;
  assign n17175 = ( n2124 & n3185 ) | ( n2124 & n3226 ) | ( n3185 & n3226 ) ;
  assign n17176 = n17175 ^ n9769 ^ n7679 ;
  assign n17174 = n8099 & ~n9437 ;
  assign n17177 = n17176 ^ n17174 ^ 1'b0 ;
  assign n17178 = n5385 ^ n4609 ^ n4108 ;
  assign n17179 = n9056 & n17178 ;
  assign n17180 = ( n8514 & n13849 ) | ( n8514 & n14149 ) | ( n13849 & n14149 ) ;
  assign n17181 = ( n528 & n1026 ) | ( n528 & ~n15378 ) | ( n1026 & ~n15378 ) ;
  assign n17182 = n17181 ^ n9948 ^ n9316 ;
  assign n17183 = n3891 ^ n752 ^ x1 ;
  assign n17184 = ( n6649 & n7847 ) | ( n6649 & n17183 ) | ( n7847 & n17183 ) ;
  assign n17185 = n566 | n3898 ;
  assign n17186 = n17184 & ~n17185 ;
  assign n17187 = n3990 & n7687 ;
  assign n17191 = n15858 ^ n13382 ^ n9480 ;
  assign n17192 = n17191 ^ n10970 ^ 1'b0 ;
  assign n17193 = ( ~n9333 & n12982 ) | ( ~n9333 & n17192 ) | ( n12982 & n17192 ) ;
  assign n17188 = ( n1779 & n6315 ) | ( n1779 & ~n9090 ) | ( n6315 & ~n9090 ) ;
  assign n17189 = n7998 ^ n2951 ^ 1'b0 ;
  assign n17190 = ( ~n1816 & n17188 ) | ( ~n1816 & n17189 ) | ( n17188 & n17189 ) ;
  assign n17194 = n17193 ^ n17190 ^ n11671 ;
  assign n17195 = n4480 ^ n3154 ^ n2657 ;
  assign n17196 = ( n7619 & n10077 ) | ( n7619 & n17195 ) | ( n10077 & n17195 ) ;
  assign n17197 = n4392 ^ n3333 ^ n958 ;
  assign n17198 = n9846 ^ n2831 ^ n694 ;
  assign n17199 = n17197 & ~n17198 ;
  assign n17200 = ~n1894 & n17199 ;
  assign n17201 = n17200 ^ n11623 ^ 1'b0 ;
  assign n17202 = n17045 & n17201 ;
  assign n17203 = n9458 ^ n3411 ^ n2191 ;
  assign n17204 = ( n6087 & ~n15590 ) | ( n6087 & n17203 ) | ( ~n15590 & n17203 ) ;
  assign n17205 = n1619 & ~n5145 ;
  assign n17206 = n7395 & n17205 ;
  assign n17207 = n17206 ^ n10218 ^ n2188 ;
  assign n17208 = ( n1466 & n5118 ) | ( n1466 & ~n8117 ) | ( n5118 & ~n8117 ) ;
  assign n17209 = n17208 ^ n5385 ^ 1'b0 ;
  assign n17210 = n10875 | n17209 ;
  assign n17211 = ( ~n3987 & n13267 ) | ( ~n3987 & n17210 ) | ( n13267 & n17210 ) ;
  assign n17212 = ( n10904 & n17207 ) | ( n10904 & ~n17211 ) | ( n17207 & ~n17211 ) ;
  assign n17219 = n16901 ^ n10803 ^ 1'b0 ;
  assign n17220 = n3815 | n17219 ;
  assign n17213 = n15928 ^ n9909 ^ 1'b0 ;
  assign n17214 = n15904 ^ n9951 ^ n8884 ;
  assign n17215 = n17214 ^ n8796 ^ 1'b0 ;
  assign n17216 = n13209 | n17215 ;
  assign n17217 = n15579 & ~n17216 ;
  assign n17218 = n17213 & n17217 ;
  assign n17221 = n17220 ^ n17218 ^ n6366 ;
  assign n17222 = n7054 ^ n6100 ^ n197 ;
  assign n17223 = n17222 ^ n16022 ^ n2421 ;
  assign n17224 = n17223 ^ n2686 ^ n2515 ;
  assign n17225 = ( n6289 & ~n15213 ) | ( n6289 & n17224 ) | ( ~n15213 & n17224 ) ;
  assign n17226 = n10449 ^ n6570 ^ n5219 ;
  assign n17227 = n17226 ^ n10982 ^ n5450 ;
  assign n17228 = n250 & ~n576 ;
  assign n17229 = ~n14443 & n17228 ;
  assign n17230 = n12570 ^ n10541 ^ n7146 ;
  assign n17231 = n17230 ^ n15251 ^ n4157 ;
  assign n17234 = n1336 | n1824 ;
  assign n17235 = ( ~n8697 & n15069 ) | ( ~n8697 & n17234 ) | ( n15069 & n17234 ) ;
  assign n17232 = n5137 ^ n1705 ^ n1482 ;
  assign n17233 = ( n3171 & ~n11519 ) | ( n3171 & n17232 ) | ( ~n11519 & n17232 ) ;
  assign n17236 = n17235 ^ n17233 ^ n11093 ;
  assign n17242 = n4581 ^ n1331 ^ n380 ;
  assign n17240 = n1649 & n8996 ;
  assign n17241 = n17240 ^ n14356 ^ 1'b0 ;
  assign n17243 = n17242 ^ n17241 ^ n12511 ;
  assign n17238 = n11925 ^ n8117 ^ n1256 ;
  assign n17237 = n6738 ^ n3473 ^ n576 ;
  assign n17239 = n17238 ^ n17237 ^ n13180 ;
  assign n17244 = n17243 ^ n17239 ^ n7431 ;
  assign n17245 = n12421 ^ n5236 ^ 1'b0 ;
  assign n17246 = ( n10936 & n14207 ) | ( n10936 & ~n17245 ) | ( n14207 & ~n17245 ) ;
  assign n17247 = n9876 ^ n9138 ^ n796 ;
  assign n17248 = ( n9259 & n10913 ) | ( n9259 & n13252 ) | ( n10913 & n13252 ) ;
  assign n17249 = n2840 ^ n490 ^ x12 ;
  assign n17250 = ( n5105 & n6700 ) | ( n5105 & n13496 ) | ( n6700 & n13496 ) ;
  assign n17251 = ( n9385 & n17249 ) | ( n9385 & n17250 ) | ( n17249 & n17250 ) ;
  assign n17254 = n2196 ^ n1079 ^ n858 ;
  assign n17253 = n5457 & ~n7284 ;
  assign n17255 = n17254 ^ n17253 ^ n220 ;
  assign n17252 = ( n282 & ~n6861 ) | ( n282 & n12795 ) | ( ~n6861 & n12795 ) ;
  assign n17256 = n17255 ^ n17252 ^ n893 ;
  assign n17257 = n13126 ^ n6673 ^ n5277 ;
  assign n17258 = n17257 ^ n13683 ^ n1554 ;
  assign n17259 = ( n3097 & n7563 ) | ( n3097 & n11234 ) | ( n7563 & n11234 ) ;
  assign n17260 = n11689 ^ n4996 ^ 1'b0 ;
  assign n17261 = n6855 ^ n4569 ^ n1991 ;
  assign n17262 = n17261 ^ n9622 ^ n8339 ;
  assign n17263 = ( ~n3310 & n10412 ) | ( ~n3310 & n17262 ) | ( n10412 & n17262 ) ;
  assign n17264 = n17263 ^ n3431 ^ 1'b0 ;
  assign n17265 = n17163 ^ n1413 ^ 1'b0 ;
  assign n17267 = ( n1867 & ~n5737 ) | ( n1867 & n12733 ) | ( ~n5737 & n12733 ) ;
  assign n17266 = ( ~n1967 & n10310 ) | ( ~n1967 & n16554 ) | ( n10310 & n16554 ) ;
  assign n17268 = n17267 ^ n17266 ^ n10026 ;
  assign n17269 = ( ~n416 & n704 ) | ( ~n416 & n5991 ) | ( n704 & n5991 ) ;
  assign n17270 = n17269 ^ n13478 ^ n3387 ;
  assign n17271 = n12667 ^ n10680 ^ n6217 ;
  assign n17272 = ( n17268 & n17270 ) | ( n17268 & ~n17271 ) | ( n17270 & ~n17271 ) ;
  assign n17273 = n17272 ^ n3105 ^ 1'b0 ;
  assign n17274 = n2608 & n10237 ;
  assign n17275 = n8065 ^ n882 ^ n192 ;
  assign n17276 = ( ~n6274 & n11687 ) | ( ~n6274 & n17275 ) | ( n11687 & n17275 ) ;
  assign n17277 = ( n1960 & ~n2147 ) | ( n1960 & n17276 ) | ( ~n2147 & n17276 ) ;
  assign n17278 = n9517 ^ n8971 ^ n6984 ;
  assign n17279 = n4577 & n9990 ;
  assign n17280 = n15110 & ~n17279 ;
  assign n17281 = n17280 ^ n3278 ^ 1'b0 ;
  assign n17282 = ( n3420 & n9019 ) | ( n3420 & n11226 ) | ( n9019 & n11226 ) ;
  assign n17283 = ( n4063 & ~n14457 ) | ( n4063 & n17282 ) | ( ~n14457 & n17282 ) ;
  assign n17284 = n5151 ^ n1287 ^ n1094 ;
  assign n17294 = n10408 ^ n2525 ^ 1'b0 ;
  assign n17295 = n15073 & ~n17294 ;
  assign n17287 = ( ~n3603 & n3821 ) | ( ~n3603 & n5463 ) | ( n3821 & n5463 ) ;
  assign n17288 = n3232 ^ n1801 ^ n1603 ;
  assign n17289 = ( n2004 & n2989 ) | ( n2004 & ~n12280 ) | ( n2989 & ~n12280 ) ;
  assign n17290 = n17289 ^ n11807 ^ n8256 ;
  assign n17291 = ( n11649 & n17288 ) | ( n11649 & ~n17290 ) | ( n17288 & ~n17290 ) ;
  assign n17292 = ( n9145 & n17287 ) | ( n9145 & n17291 ) | ( n17287 & n17291 ) ;
  assign n17285 = n3940 | n7525 ;
  assign n17286 = n17285 ^ n7980 ^ 1'b0 ;
  assign n17293 = n17292 ^ n17286 ^ n9429 ;
  assign n17296 = n17295 ^ n17293 ^ n3331 ;
  assign n17297 = n17296 ^ n14141 ^ n940 ;
  assign n17298 = ( n10623 & n17284 ) | ( n10623 & ~n17297 ) | ( n17284 & ~n17297 ) ;
  assign n17299 = n17298 ^ n9259 ^ n1576 ;
  assign n17300 = n13292 ^ n4780 ^ n390 ;
  assign n17301 = n7471 ^ n3939 ^ n2138 ;
  assign n17302 = ( ~n3160 & n9330 ) | ( ~n3160 & n17301 ) | ( n9330 & n17301 ) ;
  assign n17303 = ( ~n2138 & n10419 ) | ( ~n2138 & n17302 ) | ( n10419 & n17302 ) ;
  assign n17304 = n9466 ^ n4298 ^ 1'b0 ;
  assign n17305 = ( n17300 & ~n17303 ) | ( n17300 & n17304 ) | ( ~n17303 & n17304 ) ;
  assign n17306 = n9203 ^ n4890 ^ n4779 ;
  assign n17307 = n17306 ^ n15451 ^ n10632 ;
  assign n17308 = ( n6212 & ~n6242 ) | ( n6212 & n10979 ) | ( ~n6242 & n10979 ) ;
  assign n17309 = n4571 & ~n17308 ;
  assign n17310 = n17309 ^ n11639 ^ 1'b0 ;
  assign n17311 = ( n3039 & n3396 ) | ( n3039 & n5101 ) | ( n3396 & n5101 ) ;
  assign n17312 = n17311 ^ n9720 ^ 1'b0 ;
  assign n17313 = ( n9717 & n12373 ) | ( n9717 & n17312 ) | ( n12373 & n17312 ) ;
  assign n17314 = ( n2977 & n4386 ) | ( n2977 & n4400 ) | ( n4386 & n4400 ) ;
  assign n17315 = n17314 ^ n12041 ^ n6089 ;
  assign n17316 = n17315 ^ n11015 ^ n920 ;
  assign n17317 = n17316 ^ n14342 ^ n12157 ;
  assign n17318 = n7288 & ~n8941 ;
  assign n17319 = n2314 ^ n972 ^ 1'b0 ;
  assign n17320 = ~n4949 & n17319 ;
  assign n17321 = n8719 ^ n7447 ^ n2768 ;
  assign n17322 = ( n4666 & n17320 ) | ( n4666 & ~n17321 ) | ( n17320 & ~n17321 ) ;
  assign n17323 = n2919 | n9646 ;
  assign n17324 = n10998 ^ n4602 ^ 1'b0 ;
  assign n17325 = n17323 | n17324 ;
  assign n17326 = n1419 & ~n3683 ;
  assign n17327 = n17326 ^ n16049 ^ n198 ;
  assign n17331 = ( n6710 & n7671 ) | ( n6710 & n16040 ) | ( n7671 & n16040 ) ;
  assign n17332 = ( n1024 & n9395 ) | ( n1024 & ~n17331 ) | ( n9395 & ~n17331 ) ;
  assign n17333 = n17332 ^ n10016 ^ n9212 ;
  assign n17328 = n4774 & ~n5293 ;
  assign n17329 = n17328 ^ n9194 ^ 1'b0 ;
  assign n17330 = n2155 & n17329 ;
  assign n17334 = n17333 ^ n17330 ^ n9718 ;
  assign n17335 = ( ~n974 & n14646 ) | ( ~n974 & n17334 ) | ( n14646 & n17334 ) ;
  assign n17337 = n9208 ^ n467 ^ 1'b0 ;
  assign n17338 = n301 & n787 ;
  assign n17339 = n16814 & n17338 ;
  assign n17340 = ( n5348 & n17337 ) | ( n5348 & n17339 ) | ( n17337 & n17339 ) ;
  assign n17336 = ( n1002 & ~n10177 ) | ( n1002 & n14860 ) | ( ~n10177 & n14860 ) ;
  assign n17341 = n17340 ^ n17336 ^ n8084 ;
  assign n17342 = ( n8139 & n9608 ) | ( n8139 & ~n13128 ) | ( n9608 & ~n13128 ) ;
  assign n17343 = n13141 ^ n4081 ^ n2180 ;
  assign n17344 = n14539 ^ n4559 ^ n780 ;
  assign n17345 = n17344 ^ n1055 ^ n319 ;
  assign n17346 = ( n10436 & ~n11119 ) | ( n10436 & n17345 ) | ( ~n11119 & n17345 ) ;
  assign n17347 = ~n2230 & n17346 ;
  assign n17348 = n7538 ^ n4045 ^ n1426 ;
  assign n17349 = ( n371 & ~n5554 ) | ( n371 & n8492 ) | ( ~n5554 & n8492 ) ;
  assign n17350 = n17349 ^ n13671 ^ n13527 ;
  assign n17351 = n5796 ^ n1821 ^ 1'b0 ;
  assign n17352 = n17350 | n17351 ;
  assign n17353 = ~n3686 & n5231 ;
  assign n17354 = n16674 & n17353 ;
  assign n17361 = n9450 ^ n7880 ^ n3926 ;
  assign n17358 = n13808 ^ n11245 ^ n2478 ;
  assign n17355 = n10686 ^ n9837 ^ n2864 ;
  assign n17356 = ( ~n6722 & n15810 ) | ( ~n6722 & n17355 ) | ( n15810 & n17355 ) ;
  assign n17357 = n17356 ^ n3070 ^ n206 ;
  assign n17359 = n17358 ^ n17357 ^ n2940 ;
  assign n17360 = n17359 ^ n14213 ^ n5649 ;
  assign n17362 = n17361 ^ n17360 ^ n11936 ;
  assign n17363 = n10659 ^ n1335 ^ n325 ;
  assign n17364 = n17363 ^ n7885 ^ n499 ;
  assign n17365 = ( ~n482 & n6784 ) | ( ~n482 & n14090 ) | ( n6784 & n14090 ) ;
  assign n17366 = ~n6078 & n10238 ;
  assign n17367 = ~n11317 & n17366 ;
  assign n17368 = ( ~n6802 & n14592 ) | ( ~n6802 & n17367 ) | ( n14592 & n17367 ) ;
  assign n17369 = ( n16689 & ~n17365 ) | ( n16689 & n17368 ) | ( ~n17365 & n17368 ) ;
  assign n17370 = ( x62 & ~n9651 ) | ( x62 & n13203 ) | ( ~n9651 & n13203 ) ;
  assign n17371 = n17370 ^ n12695 ^ 1'b0 ;
  assign n17372 = n4543 ^ n2409 ^ 1'b0 ;
  assign n17373 = n17371 & n17372 ;
  assign n17374 = ( ~n1603 & n3300 ) | ( ~n1603 & n17373 ) | ( n3300 & n17373 ) ;
  assign n17375 = ( n4151 & ~n6363 ) | ( n4151 & n14035 ) | ( ~n6363 & n14035 ) ;
  assign n17376 = ( n383 & n15464 ) | ( n383 & n17375 ) | ( n15464 & n17375 ) ;
  assign n17379 = ( n1895 & n5566 ) | ( n1895 & n16169 ) | ( n5566 & n16169 ) ;
  assign n17377 = n9752 ^ n8064 ^ n4590 ;
  assign n17378 = ( n9487 & n13999 ) | ( n9487 & n17377 ) | ( n13999 & n17377 ) ;
  assign n17380 = n17379 ^ n17378 ^ n358 ;
  assign n17381 = n15422 ^ n13520 ^ n8889 ;
  assign n17385 = n15317 ^ n7138 ^ n5749 ;
  assign n17386 = n17385 ^ n13855 ^ n3564 ;
  assign n17382 = n7785 ^ n6021 ^ n730 ;
  assign n17383 = n17382 ^ n13653 ^ 1'b0 ;
  assign n17384 = ~n7639 & n17383 ;
  assign n17387 = n17386 ^ n17384 ^ n9450 ;
  assign n17388 = ( n6792 & ~n17381 ) | ( n6792 & n17387 ) | ( ~n17381 & n17387 ) ;
  assign n17389 = n3377 & n11237 ;
  assign n17390 = n17389 ^ n9434 ^ 1'b0 ;
  assign n17395 = n697 & n3977 ;
  assign n17396 = n17395 ^ n4236 ^ 1'b0 ;
  assign n17391 = n9937 ^ n9337 ^ 1'b0 ;
  assign n17392 = ~n8361 & n17391 ;
  assign n17393 = n1122 & n17392 ;
  assign n17394 = n17393 ^ n4131 ^ 1'b0 ;
  assign n17397 = n17396 ^ n17394 ^ n10663 ;
  assign n17398 = n6449 ^ n5621 ^ n3285 ;
  assign n17399 = n17398 ^ n3813 ^ 1'b0 ;
  assign n17400 = n12270 ^ n5522 ^ n1769 ;
  assign n17401 = ( n3426 & ~n7083 ) | ( n3426 & n17400 ) | ( ~n7083 & n17400 ) ;
  assign n17407 = ( n5302 & ~n6200 ) | ( n5302 & n8259 ) | ( ~n6200 & n8259 ) ;
  assign n17408 = ( ~n5793 & n7665 ) | ( ~n5793 & n17407 ) | ( n7665 & n17407 ) ;
  assign n17406 = n4519 & n16148 ;
  assign n17402 = n7218 ^ n7117 ^ n4447 ;
  assign n17403 = n10926 ^ n6665 ^ 1'b0 ;
  assign n17404 = ( n129 & n17402 ) | ( n129 & ~n17403 ) | ( n17402 & ~n17403 ) ;
  assign n17405 = n17404 ^ n6863 ^ n1378 ;
  assign n17409 = n17408 ^ n17406 ^ n17405 ;
  assign n17411 = n1711 ^ n240 ^ 1'b0 ;
  assign n17412 = n5132 & ~n17411 ;
  assign n17410 = ( n7224 & ~n10235 ) | ( n7224 & n11027 ) | ( ~n10235 & n11027 ) ;
  assign n17413 = n17412 ^ n17410 ^ n8791 ;
  assign n17414 = n7143 & n14608 ;
  assign n17415 = n3501 & n17414 ;
  assign n17416 = n6485 ^ n5619 ^ n430 ;
  assign n17417 = n6887 & ~n17416 ;
  assign n17418 = ~n11985 & n17417 ;
  assign n17419 = n14076 ^ n5458 ^ n4379 ;
  assign n17420 = n5834 ^ n5745 ^ n3934 ;
  assign n17421 = n17420 ^ n15402 ^ n13240 ;
  assign n17422 = n17232 & ~n17421 ;
  assign n17424 = n6747 ^ n1810 ^ x10 ;
  assign n17423 = n2394 | n7195 ;
  assign n17425 = n17424 ^ n17423 ^ 1'b0 ;
  assign n17426 = n17425 ^ n13930 ^ n5355 ;
  assign n17429 = n14759 ^ n12475 ^ n3241 ;
  assign n17427 = n12631 ^ n5112 ^ n486 ;
  assign n17428 = n13204 | n17427 ;
  assign n17430 = n17429 ^ n17428 ^ n3107 ;
  assign n17431 = ( ~n366 & n8275 ) | ( ~n366 & n13605 ) | ( n8275 & n13605 ) ;
  assign n17433 = ~n2031 & n3075 ;
  assign n17434 = n9549 ^ n3976 ^ n3523 ;
  assign n17435 = n17434 ^ n1718 ^ 1'b0 ;
  assign n17436 = ( n4016 & n17433 ) | ( n4016 & ~n17435 ) | ( n17433 & ~n17435 ) ;
  assign n17432 = n5091 ^ n4586 ^ n2090 ;
  assign n17437 = n17436 ^ n17432 ^ n4172 ;
  assign n17438 = ( ~n5050 & n6849 ) | ( ~n5050 & n14703 ) | ( n6849 & n14703 ) ;
  assign n17439 = n5898 & ~n12059 ;
  assign n17440 = n15479 ^ n11907 ^ n463 ;
  assign n17441 = ~n1449 & n17440 ;
  assign n17442 = n8981 ^ n7401 ^ 1'b0 ;
  assign n17443 = n17442 ^ n9906 ^ n7173 ;
  assign n17444 = ( n2770 & ~n9134 ) | ( n2770 & n17443 ) | ( ~n9134 & n17443 ) ;
  assign n17445 = n15618 ^ n1457 ^ 1'b0 ;
  assign n17446 = ( n11421 & ~n15594 ) | ( n11421 & n17105 ) | ( ~n15594 & n17105 ) ;
  assign n17447 = n10006 ^ n3440 ^ 1'b0 ;
  assign n17448 = ~n6051 & n17447 ;
  assign n17449 = n17448 ^ n15632 ^ n7665 ;
  assign n17450 = n16500 ^ n4418 ^ n3889 ;
  assign n17451 = n17450 ^ n9598 ^ n6210 ;
  assign n17452 = n6333 | n17451 ;
  assign n17453 = n4016 | n17452 ;
  assign n17454 = ( n4087 & ~n7043 ) | ( n4087 & n16288 ) | ( ~n7043 & n16288 ) ;
  assign n17455 = n17454 ^ n14380 ^ n4306 ;
  assign n17456 = ( n13182 & ~n17453 ) | ( n13182 & n17455 ) | ( ~n17453 & n17455 ) ;
  assign n17457 = ( ~n5456 & n7985 ) | ( ~n5456 & n11925 ) | ( n7985 & n11925 ) ;
  assign n17461 = n10968 ^ n1884 ^ n211 ;
  assign n17460 = ( n475 & n2565 ) | ( n475 & n3815 ) | ( n2565 & n3815 ) ;
  assign n17462 = n17461 ^ n17460 ^ n738 ;
  assign n17463 = n17462 ^ n11419 ^ n10609 ;
  assign n17459 = ( n992 & n1712 ) | ( n992 & ~n13220 ) | ( n1712 & ~n13220 ) ;
  assign n17458 = n8445 ^ n7106 ^ n2777 ;
  assign n17464 = n17463 ^ n17459 ^ n17458 ;
  assign n17465 = ( ~n465 & n5619 ) | ( ~n465 & n17256 ) | ( n5619 & n17256 ) ;
  assign n17466 = n7758 & n15753 ;
  assign n17470 = ( n556 & n1468 ) | ( n556 & ~n6247 ) | ( n1468 & ~n6247 ) ;
  assign n17467 = n2910 ^ n2363 ^ n1507 ;
  assign n17468 = n13534 ^ n4018 ^ n1760 ;
  assign n17469 = ( n1736 & n17467 ) | ( n1736 & n17468 ) | ( n17467 & n17468 ) ;
  assign n17471 = n17470 ^ n17469 ^ n14632 ;
  assign n17472 = ( ~n499 & n2236 ) | ( ~n499 & n15853 ) | ( n2236 & n15853 ) ;
  assign n17473 = ( n1376 & n11091 ) | ( n1376 & ~n17472 ) | ( n11091 & ~n17472 ) ;
  assign n17474 = n6335 ^ n5821 ^ n696 ;
  assign n17475 = n5966 | n13023 ;
  assign n17476 = n14969 & ~n17475 ;
  assign n17477 = n17476 ^ n9733 ^ n3917 ;
  assign n17478 = n17474 & n17477 ;
  assign n17479 = n17478 ^ n15480 ^ 1'b0 ;
  assign n17481 = ( n234 & n2182 ) | ( n234 & n2853 ) | ( n2182 & n2853 ) ;
  assign n17480 = ( n8613 & n9173 ) | ( n8613 & ~n16136 ) | ( n9173 & ~n16136 ) ;
  assign n17482 = n17481 ^ n17480 ^ n15965 ;
  assign n17483 = n15845 ^ n10545 ^ n8644 ;
  assign n17484 = n7648 ^ n1377 ^ n1079 ;
  assign n17485 = n17484 ^ n1157 ^ n586 ;
  assign n17486 = n17485 ^ n5053 ^ n2243 ;
  assign n17487 = n12292 ^ n5214 ^ 1'b0 ;
  assign n17488 = ~n3392 & n5420 ;
  assign n17489 = ~n3556 & n17488 ;
  assign n17490 = n11843 ^ n10505 ^ 1'b0 ;
  assign n17491 = ( n2449 & n11181 ) | ( n2449 & ~n11566 ) | ( n11181 & ~n11566 ) ;
  assign n17492 = ( n17489 & ~n17490 ) | ( n17489 & n17491 ) | ( ~n17490 & n17491 ) ;
  assign n17494 = ( n9415 & n10388 ) | ( n9415 & ~n15042 ) | ( n10388 & ~n15042 ) ;
  assign n17493 = n8443 ^ n1303 ^ n207 ;
  assign n17495 = n17494 ^ n17493 ^ n5299 ;
  assign n17497 = n13481 ^ n11237 ^ n4061 ;
  assign n17496 = ( n6049 & n7642 ) | ( n6049 & n7899 ) | ( n7642 & n7899 ) ;
  assign n17498 = n17497 ^ n17496 ^ n3274 ;
  assign n17499 = ( n3173 & n6611 ) | ( n3173 & n17468 ) | ( n6611 & n17468 ) ;
  assign n17500 = n3530 ^ n1871 ^ n1569 ;
  assign n17501 = n17500 ^ n5487 ^ n5192 ;
  assign n17502 = ( n3678 & ~n10875 ) | ( n3678 & n17501 ) | ( ~n10875 & n17501 ) ;
  assign n17503 = n17142 ^ n3621 ^ n2896 ;
  assign n17504 = ( n1590 & n3303 ) | ( n1590 & n17503 ) | ( n3303 & n17503 ) ;
  assign n17505 = n17504 ^ n15292 ^ n12966 ;
  assign n17506 = ( ~n12518 & n17502 ) | ( ~n12518 & n17505 ) | ( n17502 & n17505 ) ;
  assign n17507 = n16147 ^ n13263 ^ 1'b0 ;
  assign n17508 = ( ~n8047 & n8946 ) | ( ~n8047 & n17507 ) | ( n8946 & n17507 ) ;
  assign n17510 = ( n944 & n12182 ) | ( n944 & ~n13143 ) | ( n12182 & ~n13143 ) ;
  assign n17509 = n3494 & ~n9095 ;
  assign n17511 = n17510 ^ n17509 ^ 1'b0 ;
  assign n17512 = n518 | n17511 ;
  assign n17513 = n17512 ^ n4888 ^ 1'b0 ;
  assign n17514 = n5308 ^ n3806 ^ n801 ;
  assign n17515 = n17514 ^ n8016 ^ n3531 ;
  assign n17516 = ( n5740 & ~n10927 ) | ( n5740 & n14570 ) | ( ~n10927 & n14570 ) ;
  assign n17519 = n12107 ^ n7260 ^ n819 ;
  assign n17517 = n12672 ^ n4778 ^ n1887 ;
  assign n17518 = ( ~n15596 & n16934 ) | ( ~n15596 & n17517 ) | ( n16934 & n17517 ) ;
  assign n17520 = n17519 ^ n17518 ^ n10235 ;
  assign n17521 = n6566 ^ n5934 ^ n5551 ;
  assign n17522 = n17521 ^ n7389 ^ n6430 ;
  assign n17523 = ~n5903 & n8013 ;
  assign n17524 = n17523 ^ n10044 ^ n7874 ;
  assign n17525 = n16374 ^ n10726 ^ n1775 ;
  assign n17526 = n1809 & ~n9391 ;
  assign n17527 = ( n788 & ~n1778 ) | ( n788 & n2382 ) | ( ~n1778 & n2382 ) ;
  assign n17528 = n17527 ^ n14715 ^ 1'b0 ;
  assign n17529 = n17528 ^ n15714 ^ n1217 ;
  assign n17530 = n15101 ^ n2101 ^ 1'b0 ;
  assign n17531 = ~n17529 & n17530 ;
  assign n17532 = n10610 ^ n4888 ^ n3866 ;
  assign n17533 = n17532 ^ n4493 ^ 1'b0 ;
  assign n17534 = ( n4400 & ~n5978 ) | ( n4400 & n11880 ) | ( ~n5978 & n11880 ) ;
  assign n17535 = ( n7787 & n17533 ) | ( n7787 & ~n17534 ) | ( n17533 & ~n17534 ) ;
  assign n17536 = n10573 ^ n5719 ^ n3994 ;
  assign n17537 = n17536 ^ n10206 ^ 1'b0 ;
  assign n17538 = ( ~n3789 & n16969 ) | ( ~n3789 & n17537 ) | ( n16969 & n17537 ) ;
  assign n17539 = ( n8942 & n13297 ) | ( n8942 & n17538 ) | ( n13297 & n17538 ) ;
  assign n17541 = n1320 ^ n758 ^ 1'b0 ;
  assign n17540 = n6767 ^ n6076 ^ n4054 ;
  assign n17542 = n17541 ^ n17540 ^ n580 ;
  assign n17543 = ( n1277 & ~n6719 ) | ( n1277 & n17542 ) | ( ~n6719 & n17542 ) ;
  assign n17544 = ( n3356 & ~n11256 ) | ( n3356 & n17543 ) | ( ~n11256 & n17543 ) ;
  assign n17546 = n4780 ^ n3411 ^ n3020 ;
  assign n17545 = n15405 ^ n14222 ^ n4174 ;
  assign n17547 = n17546 ^ n17545 ^ n12149 ;
  assign n17551 = n7948 ^ n4455 ^ n411 ;
  assign n17552 = ~n1298 & n17551 ;
  assign n17553 = ~n4430 & n5386 ;
  assign n17554 = n17552 & n17553 ;
  assign n17548 = ( ~n594 & n620 ) | ( ~n594 & n6048 ) | ( n620 & n6048 ) ;
  assign n17549 = n12995 ^ n9986 ^ n3383 ;
  assign n17550 = ( n11934 & n17548 ) | ( n11934 & n17549 ) | ( n17548 & n17549 ) ;
  assign n17555 = n17554 ^ n17550 ^ n6362 ;
  assign n17556 = ( n797 & n7530 ) | ( n797 & n15795 ) | ( n7530 & n15795 ) ;
  assign n17557 = n17556 ^ n15325 ^ 1'b0 ;
  assign n17558 = n12565 & n17557 ;
  assign n17559 = n2196 | n6860 ;
  assign n17560 = ( n4391 & ~n8907 ) | ( n4391 & n12511 ) | ( ~n8907 & n12511 ) ;
  assign n17561 = ( ~n17484 & n17559 ) | ( ~n17484 & n17560 ) | ( n17559 & n17560 ) ;
  assign n17562 = n3433 & n11174 ;
  assign n17563 = ( n12116 & n15663 ) | ( n12116 & n15823 ) | ( n15663 & n15823 ) ;
  assign n17564 = n7997 ^ n5078 ^ n2967 ;
  assign n17565 = ( n4557 & n14243 ) | ( n4557 & n17564 ) | ( n14243 & n17564 ) ;
  assign n17566 = n17565 ^ n15247 ^ n12035 ;
  assign n17567 = n6257 ^ n3055 ^ n2422 ;
  assign n17568 = n9838 ^ n6364 ^ n6041 ;
  assign n17571 = n2432 ^ n467 ^ x29 ;
  assign n17569 = n3554 & ~n4585 ;
  assign n17570 = ~n4871 & n17569 ;
  assign n17572 = n17571 ^ n17570 ^ n922 ;
  assign n17573 = ( n1093 & n8096 ) | ( n1093 & n15569 ) | ( n8096 & n15569 ) ;
  assign n17574 = ( n5363 & n8864 ) | ( n5363 & ~n11473 ) | ( n8864 & ~n11473 ) ;
  assign n17575 = ( n2091 & n17573 ) | ( n2091 & ~n17574 ) | ( n17573 & ~n17574 ) ;
  assign n17586 = n4683 & n8933 ;
  assign n17587 = ~n2888 & n17586 ;
  assign n17588 = n17587 ^ n16770 ^ n9547 ;
  assign n17589 = ( n9017 & ~n9830 ) | ( n9017 & n17588 ) | ( ~n9830 & n17588 ) ;
  assign n17590 = ( n3643 & n8501 ) | ( n3643 & ~n17589 ) | ( n8501 & ~n17589 ) ;
  assign n17576 = n13111 ^ n3184 ^ n2679 ;
  assign n17577 = n5696 & ~n17576 ;
  assign n17578 = n17577 ^ n3763 ^ 1'b0 ;
  assign n17579 = n17578 ^ n16214 ^ n12784 ;
  assign n17580 = n6449 ^ n1946 ^ 1'b0 ;
  assign n17581 = n5936 & ~n17580 ;
  assign n17582 = ( n874 & ~n1929 ) | ( n874 & n10670 ) | ( ~n1929 & n10670 ) ;
  assign n17583 = n17582 ^ n13109 ^ n6236 ;
  assign n17584 = ( n12382 & n17581 ) | ( n12382 & n17583 ) | ( n17581 & n17583 ) ;
  assign n17585 = n17579 & n17584 ;
  assign n17591 = n17590 ^ n17585 ^ 1'b0 ;
  assign n17592 = n17503 ^ n7581 ^ n246 ;
  assign n17593 = n7088 ^ n1834 ^ n565 ;
  assign n17594 = ( n640 & ~n987 ) | ( n640 & n17593 ) | ( ~n987 & n17593 ) ;
  assign n17595 = ~n7204 & n17594 ;
  assign n17596 = ( n4846 & n8946 ) | ( n4846 & n16134 ) | ( n8946 & n16134 ) ;
  assign n17598 = n8717 ^ n7657 ^ 1'b0 ;
  assign n17597 = n12958 ^ n8253 ^ n2805 ;
  assign n17599 = n17598 ^ n17597 ^ n1062 ;
  assign n17600 = n17599 ^ n15073 ^ n1335 ;
  assign n17601 = ( n3808 & n10649 ) | ( n3808 & n17218 ) | ( n10649 & n17218 ) ;
  assign n17602 = ~n11047 & n17076 ;
  assign n17603 = n575 & n8729 ;
  assign n17604 = n2458 ^ n2029 ^ n335 ;
  assign n17605 = n17604 ^ n2112 ^ n1964 ;
  assign n17606 = ( n1476 & n5431 ) | ( n1476 & ~n17605 ) | ( n5431 & ~n17605 ) ;
  assign n17607 = ( n5010 & n7937 ) | ( n5010 & ~n9793 ) | ( n7937 & ~n9793 ) ;
  assign n17608 = ( n3916 & n7385 ) | ( n3916 & ~n17607 ) | ( n7385 & ~n17607 ) ;
  assign n17609 = ( n6754 & ~n9901 ) | ( n6754 & n17608 ) | ( ~n9901 & n17608 ) ;
  assign n17610 = n10250 ^ n4869 ^ n1839 ;
  assign n17611 = n13067 & n17610 ;
  assign n17612 = ~n17609 & n17611 ;
  assign n17613 = ( n17603 & n17606 ) | ( n17603 & ~n17612 ) | ( n17606 & ~n17612 ) ;
  assign n17614 = n10224 ^ n6713 ^ 1'b0 ;
  assign n17615 = ~n4369 & n17614 ;
  assign n17616 = ~n10356 & n16753 ;
  assign n17617 = n6430 & n17616 ;
  assign n17618 = ~n2554 & n3145 ;
  assign n17619 = ~n4767 & n17618 ;
  assign n17620 = n10549 ^ n7550 ^ n6289 ;
  assign n17621 = n9512 ^ n8472 ^ n1955 ;
  assign n17622 = ( ~n2875 & n6023 ) | ( ~n2875 & n6572 ) | ( n6023 & n6572 ) ;
  assign n17623 = n17622 ^ n16323 ^ n7054 ;
  assign n17624 = ( n13607 & n17621 ) | ( n13607 & ~n17623 ) | ( n17621 & ~n17623 ) ;
  assign n17625 = n13193 ^ n12236 ^ n2449 ;
  assign n17626 = ( n10821 & n16653 ) | ( n10821 & ~n17625 ) | ( n16653 & ~n17625 ) ;
  assign n17627 = ( ~n17620 & n17624 ) | ( ~n17620 & n17626 ) | ( n17624 & n17626 ) ;
  assign n17628 = n17619 | n17627 ;
  assign n17629 = n17617 & ~n17628 ;
  assign n17630 = n16072 ^ n8900 ^ n1697 ;
  assign n17631 = ( ~n9392 & n17589 ) | ( ~n9392 & n17630 ) | ( n17589 & n17630 ) ;
  assign n17632 = n14159 ^ n3949 ^ n3677 ;
  assign n17633 = n16442 ^ n4833 ^ n2275 ;
  assign n17634 = n13058 & ~n17633 ;
  assign n17635 = n6412 ^ n2364 ^ n664 ;
  assign n17636 = n687 & n1661 ;
  assign n17637 = n5470 & n17636 ;
  assign n17638 = n17637 ^ n17605 ^ n8748 ;
  assign n17639 = n17635 | n17638 ;
  assign n17640 = n15967 ^ n7756 ^ 1'b0 ;
  assign n17641 = ( ~n5191 & n17639 ) | ( ~n5191 & n17640 ) | ( n17639 & n17640 ) ;
  assign n17642 = ( ~n6452 & n10050 ) | ( ~n6452 & n11752 ) | ( n10050 & n11752 ) ;
  assign n17643 = n17642 ^ n3457 ^ 1'b0 ;
  assign n17644 = n5827 ^ n2557 ^ n1195 ;
  assign n17645 = ( n6171 & ~n7539 ) | ( n6171 & n12109 ) | ( ~n7539 & n12109 ) ;
  assign n17646 = n5863 & ~n13627 ;
  assign n17647 = n17645 & n17646 ;
  assign n17648 = ( n2181 & ~n4403 ) | ( n2181 & n17647 ) | ( ~n4403 & n17647 ) ;
  assign n17649 = n4852 ^ n3893 ^ n3378 ;
  assign n17650 = n17649 ^ n9028 ^ n3865 ;
  assign n17651 = n17650 ^ n14320 ^ n11994 ;
  assign n17652 = n6796 ^ n6243 ^ n4955 ;
  assign n17667 = n9007 ^ n5077 ^ n418 ;
  assign n17668 = n17667 ^ n4876 ^ n1429 ;
  assign n17663 = ( n4351 & n6828 ) | ( n4351 & n10003 ) | ( n6828 & n10003 ) ;
  assign n17664 = ( n4959 & n6847 ) | ( n4959 & ~n17663 ) | ( n6847 & ~n17663 ) ;
  assign n17665 = ( n1667 & n2085 ) | ( n1667 & ~n10596 ) | ( n2085 & ~n10596 ) ;
  assign n17666 = ( n7367 & ~n17664 ) | ( n7367 & n17665 ) | ( ~n17664 & n17665 ) ;
  assign n17669 = n17668 ^ n17666 ^ n13023 ;
  assign n17653 = ( n1016 & ~n4079 ) | ( n1016 & n10436 ) | ( ~n4079 & n10436 ) ;
  assign n17654 = n17653 ^ n2650 ^ 1'b0 ;
  assign n17655 = n4224 & ~n17654 ;
  assign n17656 = n4281 ^ n4210 ^ 1'b0 ;
  assign n17657 = ( n8314 & n17655 ) | ( n8314 & n17656 ) | ( n17655 & n17656 ) ;
  assign n17658 = ( n381 & ~n1935 ) | ( n381 & n7532 ) | ( ~n1935 & n7532 ) ;
  assign n17659 = n15443 & n17658 ;
  assign n17660 = ~n17657 & n17659 ;
  assign n17661 = x87 & ~n17660 ;
  assign n17662 = n17661 ^ n11927 ^ n201 ;
  assign n17670 = n17669 ^ n17662 ^ n13383 ;
  assign n17671 = ( ~n8354 & n17652 ) | ( ~n8354 & n17670 ) | ( n17652 & n17670 ) ;
  assign n17672 = ~n11325 & n13566 ;
  assign n17673 = n4655 & n5225 ;
  assign n17674 = n7798 & n17673 ;
  assign n17675 = ~n7864 & n17674 ;
  assign n17676 = ( n2416 & n3752 ) | ( n2416 & ~n8147 ) | ( n3752 & ~n8147 ) ;
  assign n17677 = n11391 ^ n5253 ^ 1'b0 ;
  assign n17678 = ( n14073 & n17676 ) | ( n14073 & n17677 ) | ( n17676 & n17677 ) ;
  assign n17679 = ( n289 & ~n1955 ) | ( n289 & n6008 ) | ( ~n1955 & n6008 ) ;
  assign n17680 = n17679 ^ n11571 ^ n2971 ;
  assign n17681 = n13297 ^ n12437 ^ n5155 ;
  assign n17682 = n17681 ^ n9222 ^ n4074 ;
  assign n17683 = ( ~n14284 & n15276 ) | ( ~n14284 & n17682 ) | ( n15276 & n17682 ) ;
  assign n17686 = n6434 & ~n8043 ;
  assign n17687 = n7364 & n17686 ;
  assign n17688 = n17687 ^ n8208 ^ n1519 ;
  assign n17684 = n12480 ^ n3561 ^ n959 ;
  assign n17685 = n17684 ^ n16973 ^ n2342 ;
  assign n17689 = n17688 ^ n17685 ^ n11928 ;
  assign n17690 = ( n7332 & n9683 ) | ( n7332 & n13800 ) | ( n9683 & n13800 ) ;
  assign n17691 = n17690 ^ n5888 ^ 1'b0 ;
  assign n17692 = ~n16506 & n17691 ;
  assign n17693 = n17692 ^ n1680 ^ n1377 ;
  assign n17695 = n4129 ^ n2386 ^ n606 ;
  assign n17694 = n13021 ^ n10178 ^ n3008 ;
  assign n17696 = n17695 ^ n17694 ^ n11981 ;
  assign n17697 = ( n2770 & ~n8473 ) | ( n2770 & n17696 ) | ( ~n8473 & n17696 ) ;
  assign n17698 = ( n1662 & ~n3080 ) | ( n1662 & n3330 ) | ( ~n3080 & n3330 ) ;
  assign n17699 = n17698 ^ n4233 ^ n3030 ;
  assign n17700 = ( ~n6236 & n11965 ) | ( ~n6236 & n12457 ) | ( n11965 & n12457 ) ;
  assign n17701 = ( n3600 & n10057 ) | ( n3600 & n11953 ) | ( n10057 & n11953 ) ;
  assign n17702 = ( n10073 & n14160 ) | ( n10073 & ~n17701 ) | ( n14160 & ~n17701 ) ;
  assign n17703 = n3389 & n17702 ;
  assign n17704 = ( n5921 & n17700 ) | ( n5921 & ~n17703 ) | ( n17700 & ~n17703 ) ;
  assign n17706 = ( n1116 & ~n3683 ) | ( n1116 & n4162 ) | ( ~n3683 & n4162 ) ;
  assign n17705 = n14880 ^ n10407 ^ n1401 ;
  assign n17707 = n17706 ^ n17705 ^ n4251 ;
  assign n17709 = ( n8453 & ~n9446 ) | ( n8453 & n15611 ) | ( ~n9446 & n15611 ) ;
  assign n17708 = ( ~n2765 & n6277 ) | ( ~n2765 & n10161 ) | ( n6277 & n10161 ) ;
  assign n17710 = n17709 ^ n17708 ^ n14399 ;
  assign n17711 = n7680 & ~n14521 ;
  assign n17712 = n17711 ^ n7008 ^ 1'b0 ;
  assign n17713 = n17712 ^ n10373 ^ n8563 ;
  assign n17714 = ( n1672 & n5485 ) | ( n1672 & n17713 ) | ( n5485 & n17713 ) ;
  assign n17715 = n6407 ^ n2900 ^ n929 ;
  assign n17716 = n17715 ^ n12795 ^ n12050 ;
  assign n17718 = ( n13010 & n14315 ) | ( n13010 & ~n15911 ) | ( n14315 & ~n15911 ) ;
  assign n17717 = n13762 ^ n8299 ^ n4704 ;
  assign n17719 = n17718 ^ n17717 ^ n9542 ;
  assign n17720 = ~n9786 & n13078 ;
  assign n17721 = ( n5058 & n12150 ) | ( n5058 & n17720 ) | ( n12150 & n17720 ) ;
  assign n17723 = ( ~n6743 & n7330 ) | ( ~n6743 & n13598 ) | ( n7330 & n13598 ) ;
  assign n17724 = n17723 ^ n7486 ^ n1288 ;
  assign n17722 = n668 | n3549 ;
  assign n17725 = n17724 ^ n17722 ^ 1'b0 ;
  assign n17726 = n4249 ^ n3950 ^ 1'b0 ;
  assign n17727 = ( n6612 & n6701 ) | ( n6612 & ~n17726 ) | ( n6701 & ~n17726 ) ;
  assign n17728 = n17727 ^ n10333 ^ n3762 ;
  assign n17729 = n15808 ^ n6372 ^ n3909 ;
  assign n17730 = n1410 & ~n2443 ;
  assign n17731 = n17730 ^ n1538 ^ 1'b0 ;
  assign n17732 = n17731 ^ n13480 ^ n8127 ;
  assign n17733 = ( n10429 & ~n17729 ) | ( n10429 & n17732 ) | ( ~n17729 & n17732 ) ;
  assign n17734 = n6031 & n9073 ;
  assign n17735 = n17734 ^ n5664 ^ 1'b0 ;
  assign n17738 = n2105 ^ n1858 ^ 1'b0 ;
  assign n17739 = n17738 ^ n2509 ^ n2203 ;
  assign n17736 = n16184 ^ n10943 ^ 1'b0 ;
  assign n17737 = n17736 ^ n14920 ^ n9926 ;
  assign n17740 = n17739 ^ n17737 ^ n804 ;
  assign n17741 = ( n250 & n4001 ) | ( n250 & ~n9003 ) | ( n4001 & ~n9003 ) ;
  assign n17742 = n10101 ^ n3375 ^ n1524 ;
  assign n17743 = ( n4165 & n6582 ) | ( n4165 & ~n14151 ) | ( n6582 & ~n14151 ) ;
  assign n17744 = ( n7425 & ~n9181 ) | ( n7425 & n13047 ) | ( ~n9181 & n13047 ) ;
  assign n17745 = n1669 & ~n17744 ;
  assign n17746 = n17745 ^ n16422 ^ n7101 ;
  assign n17747 = n17746 ^ n12581 ^ x100 ;
  assign n17748 = n8943 ^ n7525 ^ n3587 ;
  assign n17749 = n15154 ^ n14570 ^ n2609 ;
  assign n17750 = ( n4030 & ~n17748 ) | ( n4030 & n17749 ) | ( ~n17748 & n17749 ) ;
  assign n17751 = ( n2358 & ~n7499 ) | ( n2358 & n9171 ) | ( ~n7499 & n9171 ) ;
  assign n17752 = ( n5969 & ~n13167 ) | ( n5969 & n17751 ) | ( ~n13167 & n17751 ) ;
  assign n17753 = n4537 ^ n4132 ^ n3294 ;
  assign n17754 = n16148 & n17753 ;
  assign n17755 = n15225 ^ n1485 ^ n756 ;
  assign n17756 = ~n5118 & n17755 ;
  assign n17757 = ~n1718 & n17756 ;
  assign n17758 = n6228 ^ n5327 ^ n1355 ;
  assign n17759 = n5791 ^ n5755 ^ n2419 ;
  assign n17760 = n17759 ^ n17529 ^ n9399 ;
  assign n17761 = n17760 ^ n16072 ^ n3148 ;
  assign n17762 = n10610 ^ n1336 ^ 1'b0 ;
  assign n17763 = n17762 ^ n3271 ^ x75 ;
  assign n17764 = n9702 & n16222 ;
  assign n17765 = n2029 & n17764 ;
  assign n17766 = n11576 ^ n4367 ^ n635 ;
  assign n17767 = n17766 ^ n13294 ^ n5024 ;
  assign n17768 = ( n17763 & n17765 ) | ( n17763 & ~n17767 ) | ( n17765 & ~n17767 ) ;
  assign n17769 = n12751 ^ n12348 ^ n8331 ;
  assign n17771 = ( n1178 & n11559 ) | ( n1178 & ~n11896 ) | ( n11559 & ~n11896 ) ;
  assign n17770 = n15836 ^ n5414 ^ n5378 ;
  assign n17772 = n17771 ^ n17770 ^ n14757 ;
  assign n17773 = n17772 ^ n4516 ^ n1562 ;
  assign n17774 = n17773 ^ n7375 ^ n6054 ;
  assign n17775 = ( n945 & ~n15272 ) | ( n945 & n17500 ) | ( ~n15272 & n17500 ) ;
  assign n17776 = n17775 ^ n16906 ^ n2633 ;
  assign n17777 = n17776 ^ n9686 ^ 1'b0 ;
  assign n17778 = n16547 ^ n6799 ^ n3098 ;
  assign n17779 = ( n1883 & n11348 ) | ( n1883 & n17642 ) | ( n11348 & n17642 ) ;
  assign n17780 = ~n17778 & n17779 ;
  assign n17781 = ( ~n3443 & n8759 ) | ( ~n3443 & n11499 ) | ( n8759 & n11499 ) ;
  assign n17782 = ~n5463 & n17781 ;
  assign n17783 = n6183 ^ n5331 ^ 1'b0 ;
  assign n17784 = ( ~n1497 & n2510 ) | ( ~n1497 & n5385 ) | ( n2510 & n5385 ) ;
  assign n17785 = n17784 ^ n6230 ^ n1280 ;
  assign n17786 = n7693 ^ n3945 ^ n1392 ;
  assign n17787 = n2576 ^ n1042 ^ n234 ;
  assign n17788 = n1323 | n17787 ;
  assign n17789 = ( n1104 & n17786 ) | ( n1104 & n17788 ) | ( n17786 & n17788 ) ;
  assign n17790 = n1183 ^ n876 ^ 1'b0 ;
  assign n17791 = ( ~n313 & n393 ) | ( ~n313 & n5423 ) | ( n393 & n5423 ) ;
  assign n17792 = n17791 ^ n3308 ^ 1'b0 ;
  assign n17793 = n2745 & ~n17792 ;
  assign n17794 = ( n324 & n1258 ) | ( n324 & ~n2327 ) | ( n1258 & ~n2327 ) ;
  assign n17795 = n17794 ^ n14035 ^ 1'b0 ;
  assign n17796 = n17795 ^ n16198 ^ n5738 ;
  assign n17797 = ( n3099 & ~n17793 ) | ( n3099 & n17796 ) | ( ~n17793 & n17796 ) ;
  assign n17798 = n17797 ^ n14978 ^ n8420 ;
  assign n17801 = ( ~n2524 & n3429 ) | ( ~n2524 & n15947 ) | ( n3429 & n15947 ) ;
  assign n17799 = n7702 & ~n13941 ;
  assign n17800 = n17799 ^ n6749 ^ 1'b0 ;
  assign n17802 = n17801 ^ n17800 ^ n15496 ;
  assign n17803 = n2109 & n3884 ;
  assign n17808 = n13623 ^ n1571 ^ 1'b0 ;
  assign n17809 = ~n1285 & n17808 ;
  assign n17804 = n6884 ^ n3248 ^ n2613 ;
  assign n17805 = n11032 ^ n10461 ^ 1'b0 ;
  assign n17806 = n14973 & ~n17805 ;
  assign n17807 = ( n16620 & ~n17804 ) | ( n16620 & n17806 ) | ( ~n17804 & n17806 ) ;
  assign n17810 = n17809 ^ n17807 ^ n10207 ;
  assign n17811 = n16783 ^ n9452 ^ 1'b0 ;
  assign n17812 = ~n645 & n17811 ;
  assign n17813 = ( x28 & ~n1405 ) | ( x28 & n7100 ) | ( ~n1405 & n7100 ) ;
  assign n17814 = ~n480 & n13411 ;
  assign n17815 = ~n843 & n17814 ;
  assign n17816 = ( n3588 & n5638 ) | ( n3588 & n7979 ) | ( n5638 & n7979 ) ;
  assign n17817 = n17815 | n17816 ;
  assign n17818 = n2001 | n17817 ;
  assign n17819 = ( n4724 & n17813 ) | ( n4724 & ~n17818 ) | ( n17813 & ~n17818 ) ;
  assign n17820 = ( x68 & n587 ) | ( x68 & ~n4041 ) | ( n587 & ~n4041 ) ;
  assign n17821 = n17820 ^ n4949 ^ n3931 ;
  assign n17822 = n17821 ^ n7688 ^ n3645 ;
  assign n17823 = n7228 | n17822 ;
  assign n17824 = n17461 ^ n11513 ^ x114 ;
  assign n17825 = n17824 ^ n15370 ^ n4718 ;
  assign n17826 = ( n588 & n3277 ) | ( n588 & n12758 ) | ( n3277 & n12758 ) ;
  assign n17827 = ( n1164 & n12825 ) | ( n1164 & n17826 ) | ( n12825 & n17826 ) ;
  assign n17828 = n14274 & ~n14666 ;
  assign n17829 = ( n1681 & n8482 ) | ( n1681 & n10376 ) | ( n8482 & n10376 ) ;
  assign n17830 = ( n858 & ~n1240 ) | ( n858 & n6461 ) | ( ~n1240 & n6461 ) ;
  assign n17831 = ( n9593 & n13547 ) | ( n9593 & ~n13994 ) | ( n13547 & ~n13994 ) ;
  assign n17832 = ( n9591 & n17830 ) | ( n9591 & ~n17831 ) | ( n17830 & ~n17831 ) ;
  assign n17833 = ( n14697 & n16683 ) | ( n14697 & ~n17832 ) | ( n16683 & ~n17832 ) ;
  assign n17834 = n6152 ^ n5217 ^ n2051 ;
  assign n17835 = ( n2419 & n9530 ) | ( n2419 & ~n12663 ) | ( n9530 & ~n12663 ) ;
  assign n17836 = n2502 & n9367 ;
  assign n17837 = ~n2045 & n17836 ;
  assign n17838 = n137 | n17837 ;
  assign n17839 = n17838 ^ n8530 ^ 1'b0 ;
  assign n17840 = ( ~n5060 & n9440 ) | ( ~n5060 & n10652 ) | ( n9440 & n10652 ) ;
  assign n17841 = n17840 ^ n3137 ^ 1'b0 ;
  assign n17842 = ( n1887 & ~n17839 ) | ( n1887 & n17841 ) | ( ~n17839 & n17841 ) ;
  assign n17843 = ( n3197 & ~n6992 ) | ( n3197 & n15402 ) | ( ~n6992 & n15402 ) ;
  assign n17844 = ( n11981 & n13327 ) | ( n11981 & n13493 ) | ( n13327 & n13493 ) ;
  assign n17845 = ~n2545 & n9365 ;
  assign n17846 = ~n5005 & n17845 ;
  assign n17847 = n17846 ^ n8343 ^ 1'b0 ;
  assign n17848 = n17847 ^ n5355 ^ n3678 ;
  assign n17849 = n11332 & ~n15330 ;
  assign n17850 = n17849 ^ n1056 ^ 1'b0 ;
  assign n17851 = ~n10252 & n17850 ;
  assign n17852 = ~n4141 & n17851 ;
  assign n17853 = n17848 & ~n17852 ;
  assign n17854 = n17853 ^ n10476 ^ 1'b0 ;
  assign n17855 = n12089 | n14090 ;
  assign n17856 = n12708 & ~n17855 ;
  assign n17857 = ( n7208 & n8535 ) | ( n7208 & n9423 ) | ( n8535 & n9423 ) ;
  assign n17858 = n845 & ~n10118 ;
  assign n17859 = n17858 ^ n8870 ^ 1'b0 ;
  assign n17860 = n17859 ^ n14401 ^ n1566 ;
  assign n17861 = n7481 ^ n3414 ^ n915 ;
  assign n17862 = n17861 ^ n4715 ^ 1'b0 ;
  assign n17863 = n13974 ^ n7391 ^ n7014 ;
  assign n17864 = n11709 ^ n2519 ^ x33 ;
  assign n17865 = ( n3150 & ~n4231 ) | ( n3150 & n17864 ) | ( ~n4231 & n17864 ) ;
  assign n17866 = ( n4996 & n14058 ) | ( n4996 & n17865 ) | ( n14058 & n17865 ) ;
  assign n17867 = n5189 ^ n3762 ^ n891 ;
  assign n17868 = ( ~n845 & n12396 ) | ( ~n845 & n17867 ) | ( n12396 & n17867 ) ;
  assign n17871 = ( n1081 & ~n2992 ) | ( n1081 & n8150 ) | ( ~n2992 & n8150 ) ;
  assign n17869 = ( n2309 & n7176 ) | ( n2309 & n9418 ) | ( n7176 & n9418 ) ;
  assign n17870 = n372 | n17869 ;
  assign n17872 = n17871 ^ n17870 ^ 1'b0 ;
  assign n17873 = n15127 ^ n14841 ^ n2401 ;
  assign n17874 = n15111 ^ n9855 ^ 1'b0 ;
  assign n17875 = ~n11220 & n17874 ;
  assign n17876 = ( n3854 & n17873 ) | ( n3854 & n17875 ) | ( n17873 & n17875 ) ;
  assign n17877 = ( n4742 & n10925 ) | ( n4742 & n14596 ) | ( n10925 & n14596 ) ;
  assign n17878 = n14778 ^ n5207 ^ n4679 ;
  assign n17879 = n205 & ~n17878 ;
  assign n17880 = n17877 & n17879 ;
  assign n17881 = ( ~n3782 & n14523 ) | ( ~n3782 & n17880 ) | ( n14523 & n17880 ) ;
  assign n17882 = n12630 | n17250 ;
  assign n17883 = ( ~n5201 & n8454 ) | ( ~n5201 & n17142 ) | ( n8454 & n17142 ) ;
  assign n17884 = n17883 ^ n13965 ^ n13327 ;
  assign n17885 = ( n5887 & n8762 ) | ( n5887 & ~n15836 ) | ( n8762 & ~n15836 ) ;
  assign n17886 = n17885 ^ n9028 ^ n8033 ;
  assign n17887 = n17886 ^ n11703 ^ n4623 ;
  assign n17888 = n10408 ^ n4794 ^ n1298 ;
  assign n17889 = n17888 ^ n3362 ^ n2541 ;
  assign n17890 = ( n6816 & n10373 ) | ( n6816 & n14061 ) | ( n10373 & n14061 ) ;
  assign n17891 = ( ~n10557 & n17889 ) | ( ~n10557 & n17890 ) | ( n17889 & n17890 ) ;
  assign n17892 = n12051 ^ n1241 ^ n975 ;
  assign n17893 = n8856 ^ n7794 ^ n2821 ;
  assign n17894 = n9292 ^ n7615 ^ n7323 ;
  assign n17895 = n12551 ^ n4658 ^ n1349 ;
  assign n17896 = ~n17894 & n17895 ;
  assign n17897 = ( n5111 & n17893 ) | ( n5111 & n17896 ) | ( n17893 & n17896 ) ;
  assign n17898 = ~n2930 & n12466 ;
  assign n17899 = n1447 & n17898 ;
  assign n17900 = ( n11762 & n16384 ) | ( n11762 & ~n17899 ) | ( n16384 & ~n17899 ) ;
  assign n17901 = n17900 ^ n14957 ^ n1316 ;
  assign n17902 = ( n2803 & n8155 ) | ( n2803 & ~n15305 ) | ( n8155 & ~n15305 ) ;
  assign n17903 = n17902 ^ n10908 ^ n2847 ;
  assign n17904 = ( n341 & n8480 ) | ( n341 & ~n9367 ) | ( n8480 & ~n9367 ) ;
  assign n17905 = n410 ^ n382 ^ 1'b0 ;
  assign n17906 = n17904 | n17905 ;
  assign n17907 = n3114 | n17906 ;
  assign n17908 = ( n1181 & n3983 ) | ( n1181 & n12707 ) | ( n3983 & n12707 ) ;
  assign n17909 = ( n9265 & ~n14138 ) | ( n9265 & n17908 ) | ( ~n14138 & n17908 ) ;
  assign n17910 = ( n5260 & n11649 ) | ( n5260 & n14215 ) | ( n11649 & n14215 ) ;
  assign n17911 = n3401 ^ n3125 ^ 1'b0 ;
  assign n17912 = n6966 & ~n17911 ;
  assign n17913 = ( n4198 & ~n17910 ) | ( n4198 & n17912 ) | ( ~n17910 & n17912 ) ;
  assign n17914 = ( n4415 & n6915 ) | ( n4415 & ~n7550 ) | ( n6915 & ~n7550 ) ;
  assign n17915 = ( ~n3516 & n6891 ) | ( ~n3516 & n7488 ) | ( n6891 & n7488 ) ;
  assign n17916 = n17914 & n17915 ;
  assign n17917 = n17916 ^ n4479 ^ 1'b0 ;
  assign n17918 = ( n4635 & n8716 ) | ( n4635 & ~n17917 ) | ( n8716 & ~n17917 ) ;
  assign n17919 = ( n1282 & n2387 ) | ( n1282 & n14493 ) | ( n2387 & n14493 ) ;
  assign n17920 = n11731 ^ n8016 ^ 1'b0 ;
  assign n17921 = ( n6079 & n12924 ) | ( n6079 & ~n17920 ) | ( n12924 & ~n17920 ) ;
  assign n17922 = ( ~n924 & n4118 ) | ( ~n924 & n14616 ) | ( n4118 & n14616 ) ;
  assign n17923 = n3854 ^ n2924 ^ 1'b0 ;
  assign n17924 = n6754 & n17923 ;
  assign n17925 = n14106 ^ n10940 ^ n3164 ;
  assign n17926 = n17925 ^ n15595 ^ 1'b0 ;
  assign n17927 = n851 | n9643 ;
  assign n17928 = n17927 ^ n653 ^ 1'b0 ;
  assign n17929 = n17037 ^ n13413 ^ 1'b0 ;
  assign n17930 = n17928 & ~n17929 ;
  assign n17931 = n12530 | n13463 ;
  assign n17932 = n17931 ^ n8022 ^ 1'b0 ;
  assign n17933 = n5500 & n7748 ;
  assign n17934 = n1753 & n17933 ;
  assign n17935 = ( n5685 & n6154 ) | ( n5685 & ~n17934 ) | ( n6154 & ~n17934 ) ;
  assign n17936 = n8223 ^ n5959 ^ n1297 ;
  assign n17937 = n17936 ^ n13471 ^ n12284 ;
  assign n17938 = ( n917 & n2129 ) | ( n917 & ~n7604 ) | ( n2129 & ~n7604 ) ;
  assign n17939 = ( x3 & n14578 ) | ( x3 & ~n17938 ) | ( n14578 & ~n17938 ) ;
  assign n17943 = n3828 & ~n11965 ;
  assign n17944 = ~n780 & n17943 ;
  assign n17945 = ~n3435 & n17944 ;
  assign n17940 = n9392 ^ n2136 ^ n1799 ;
  assign n17941 = n17940 ^ n14714 ^ 1'b0 ;
  assign n17942 = n361 | n17941 ;
  assign n17946 = n17945 ^ n17942 ^ n10134 ;
  assign n17947 = ~n4413 & n10404 ;
  assign n17948 = n17947 ^ n12189 ^ n5539 ;
  assign n17949 = n17948 ^ n14488 ^ n5130 ;
  assign n17950 = n9722 ^ n4386 ^ n1963 ;
  assign n17951 = n247 | n8006 ;
  assign n17952 = ( n5338 & n17950 ) | ( n5338 & n17951 ) | ( n17950 & n17951 ) ;
  assign n17955 = n1289 & ~n2460 ;
  assign n17956 = n7308 & n17955 ;
  assign n17953 = n8110 ^ n7578 ^ 1'b0 ;
  assign n17954 = n13943 | n17953 ;
  assign n17957 = n17956 ^ n17954 ^ n3971 ;
  assign n17958 = n10510 & n17957 ;
  assign n17959 = n17958 ^ n13203 ^ n8268 ;
  assign n17962 = n2770 & n6437 ;
  assign n17960 = n6533 ^ n1695 ^ 1'b0 ;
  assign n17961 = n17960 ^ n13157 ^ n3787 ;
  assign n17963 = n17962 ^ n17961 ^ n6448 ;
  assign n17964 = ( n3804 & n5977 ) | ( n3804 & n17963 ) | ( n5977 & n17963 ) ;
  assign n17966 = n3899 ^ n2148 ^ n1776 ;
  assign n17965 = n13011 ^ n11763 ^ n4338 ;
  assign n17967 = n17966 ^ n17965 ^ n1421 ;
  assign n17968 = n17485 ^ n9922 ^ n6297 ;
  assign n17969 = ~n15707 & n17968 ;
  assign n17970 = n17967 & n17969 ;
  assign n17971 = n2555 ^ n1679 ^ 1'b0 ;
  assign n17972 = n12379 & n17971 ;
  assign n17973 = n16309 ^ n8795 ^ n953 ;
  assign n17974 = n17973 ^ n14198 ^ n4451 ;
  assign n17975 = n130 & n2705 ;
  assign n17976 = n7244 & n17975 ;
  assign n17977 = n9507 ^ n8009 ^ n3588 ;
  assign n17978 = ( n435 & ~n17976 ) | ( n435 & n17977 ) | ( ~n17976 & n17977 ) ;
  assign n17979 = ( n612 & n1723 ) | ( n612 & n16371 ) | ( n1723 & n16371 ) ;
  assign n17980 = ( n9122 & n10375 ) | ( n9122 & ~n15077 ) | ( n10375 & ~n15077 ) ;
  assign n17981 = n891 & n16632 ;
  assign n17982 = n17981 ^ n12053 ^ 1'b0 ;
  assign n17983 = n12604 ^ n2553 ^ n2485 ;
  assign n17984 = n17983 ^ n11939 ^ n4642 ;
  assign n17985 = n17984 ^ n11329 ^ n6177 ;
  assign n17986 = ~n16006 & n17985 ;
  assign n17987 = ( ~n2914 & n3767 ) | ( ~n2914 & n17986 ) | ( n3767 & n17986 ) ;
  assign n17988 = n16832 ^ n14554 ^ n7207 ;
  assign n17989 = n3947 ^ n2372 ^ 1'b0 ;
  assign n17990 = n10560 | n17989 ;
  assign n17991 = n9290 | n14592 ;
  assign n17992 = ( n2936 & n17990 ) | ( n2936 & n17991 ) | ( n17990 & n17991 ) ;
  assign n17993 = ( n2662 & n17988 ) | ( n2662 & ~n17992 ) | ( n17988 & ~n17992 ) ;
  assign n17999 = ( n950 & ~n1429 ) | ( n950 & n9645 ) | ( ~n1429 & n9645 ) ;
  assign n18000 = ( n3044 & n8774 ) | ( n3044 & ~n16660 ) | ( n8774 & ~n16660 ) ;
  assign n18001 = ( n3020 & n8187 ) | ( n3020 & n18000 ) | ( n8187 & n18000 ) ;
  assign n18002 = ( n6606 & n17999 ) | ( n6606 & ~n18001 ) | ( n17999 & ~n18001 ) ;
  assign n17994 = n14689 ^ n657 ^ 1'b0 ;
  assign n17995 = ~n14307 & n17994 ;
  assign n17996 = n17995 ^ n7066 ^ n1742 ;
  assign n17997 = ( n4624 & n7672 ) | ( n4624 & n17996 ) | ( n7672 & n17996 ) ;
  assign n17998 = ( ~n11888 & n12093 ) | ( ~n11888 & n17997 ) | ( n12093 & n17997 ) ;
  assign n18003 = n18002 ^ n17998 ^ 1'b0 ;
  assign n18004 = ~n11166 & n18003 ;
  assign n18005 = n11103 ^ n10242 ^ n5860 ;
  assign n18006 = ( n1209 & ~n8356 ) | ( n1209 & n9070 ) | ( ~n8356 & n9070 ) ;
  assign n18007 = ( n11394 & n18005 ) | ( n11394 & ~n18006 ) | ( n18005 & ~n18006 ) ;
  assign n18008 = n11912 ^ n7405 ^ n2752 ;
  assign n18009 = n18008 ^ n5605 ^ n1354 ;
  assign n18010 = ( n6681 & ~n10142 ) | ( n6681 & n11498 ) | ( ~n10142 & n11498 ) ;
  assign n18011 = n3168 ^ n1514 ^ n1290 ;
  assign n18012 = n11515 ^ n9292 ^ n1674 ;
  assign n18013 = n3114 | n10360 ;
  assign n18014 = n18012 | n18013 ;
  assign n18015 = ( n1457 & ~n4153 ) | ( n1457 & n13038 ) | ( ~n4153 & n13038 ) ;
  assign n18016 = ( ~n5195 & n18014 ) | ( ~n5195 & n18015 ) | ( n18014 & n18015 ) ;
  assign n18017 = n18016 ^ n7765 ^ n6130 ;
  assign n18018 = n1262 | n18017 ;
  assign n18019 = n18011 | n18018 ;
  assign n18020 = ( ~n8731 & n11688 ) | ( ~n8731 & n12017 ) | ( n11688 & n12017 ) ;
  assign n18021 = ( n2875 & n10472 ) | ( n2875 & n18020 ) | ( n10472 & n18020 ) ;
  assign n18022 = n823 | n18021 ;
  assign n18023 = ( n521 & n7697 ) | ( n521 & ~n8598 ) | ( n7697 & ~n8598 ) ;
  assign n18024 = n18023 ^ n2138 ^ n1660 ;
  assign n18025 = ( n5697 & n6178 ) | ( n5697 & ~n6465 ) | ( n6178 & ~n6465 ) ;
  assign n18026 = ( ~n1465 & n8407 ) | ( ~n1465 & n10655 ) | ( n8407 & n10655 ) ;
  assign n18027 = ( n1485 & ~n17736 ) | ( n1485 & n18026 ) | ( ~n17736 & n18026 ) ;
  assign n18028 = ( n7614 & ~n18025 ) | ( n7614 & n18027 ) | ( ~n18025 & n18027 ) ;
  assign n18029 = n12132 ^ n11885 ^ n1594 ;
  assign n18030 = n8886 ^ n4766 ^ n480 ;
  assign n18031 = ( n1231 & ~n1710 ) | ( n1231 & n2826 ) | ( ~n1710 & n2826 ) ;
  assign n18032 = ( ~n510 & n3381 ) | ( ~n510 & n18031 ) | ( n3381 & n18031 ) ;
  assign n18033 = n17885 | n18032 ;
  assign n18034 = n4311 & ~n18033 ;
  assign n18035 = ( n723 & n5903 ) | ( n723 & n18034 ) | ( n5903 & n18034 ) ;
  assign n18036 = ( ~n6913 & n9780 ) | ( ~n6913 & n10588 ) | ( n9780 & n10588 ) ;
  assign n18037 = ~n9395 & n12984 ;
  assign n18038 = ( n1522 & n18036 ) | ( n1522 & ~n18037 ) | ( n18036 & ~n18037 ) ;
  assign n18039 = n3365 & n4066 ;
  assign n18040 = n18039 ^ n13592 ^ n2884 ;
  assign n18041 = ~n3500 & n18040 ;
  assign n18042 = n1495 & n18041 ;
  assign n18043 = ~n4361 & n12966 ;
  assign n18046 = n3783 & ~n15828 ;
  assign n18044 = ( ~n2492 & n8229 ) | ( ~n2492 & n15670 ) | ( n8229 & n15670 ) ;
  assign n18045 = n18044 ^ n12039 ^ n8669 ;
  assign n18047 = n18046 ^ n18045 ^ n13777 ;
  assign n18048 = ( n872 & n8028 ) | ( n872 & ~n10515 ) | ( n8028 & ~n10515 ) ;
  assign n18049 = n18048 ^ n10659 ^ n3871 ;
  assign n18050 = ( ~n521 & n6520 ) | ( ~n521 & n18049 ) | ( n6520 & n18049 ) ;
  assign n18051 = ( n1081 & n9748 ) | ( n1081 & n18050 ) | ( n9748 & n18050 ) ;
  assign n18052 = n3682 ^ n850 ^ n235 ;
  assign n18053 = n5804 & n8054 ;
  assign n18054 = ~n15952 & n18053 ;
  assign n18055 = ( ~n5407 & n13571 ) | ( ~n5407 & n18054 ) | ( n13571 & n18054 ) ;
  assign n18056 = n10218 ^ n8672 ^ n810 ;
  assign n18057 = n18056 ^ n12845 ^ 1'b0 ;
  assign n18058 = ( ~n4440 & n5419 ) | ( ~n4440 & n8383 ) | ( n5419 & n8383 ) ;
  assign n18059 = n11797 ^ n8633 ^ n4978 ;
  assign n18063 = ( ~n150 & n1917 ) | ( ~n150 & n6843 ) | ( n1917 & n6843 ) ;
  assign n18061 = n5263 ^ n4078 ^ n751 ;
  assign n18060 = n10347 ^ n3762 ^ n2164 ;
  assign n18062 = n18061 ^ n18060 ^ n6966 ;
  assign n18064 = n18063 ^ n18062 ^ n15608 ;
  assign n18066 = n6774 ^ n5618 ^ 1'b0 ;
  assign n18065 = ( ~n1625 & n4722 ) | ( ~n1625 & n7317 ) | ( n4722 & n7317 ) ;
  assign n18067 = n18066 ^ n18065 ^ n8908 ;
  assign n18068 = ( n5743 & n8518 ) | ( n5743 & n10698 ) | ( n8518 & n10698 ) ;
  assign n18069 = n6943 ^ n1906 ^ n1782 ;
  assign n18070 = n230 & ~n17533 ;
  assign n18071 = n8308 & n18070 ;
  assign n18072 = n18071 ^ n9029 ^ 1'b0 ;
  assign n18073 = ~n12472 & n14716 ;
  assign n18074 = ~n7014 & n18073 ;
  assign n18075 = n2690 & ~n18074 ;
  assign n18076 = ( n2353 & n4274 ) | ( n2353 & n10878 ) | ( n4274 & n10878 ) ;
  assign n18077 = n8782 ^ n3556 ^ n2484 ;
  assign n18078 = ( n2320 & n13493 ) | ( n2320 & ~n18077 ) | ( n13493 & ~n18077 ) ;
  assign n18079 = ( n13248 & ~n13294 ) | ( n13248 & n18078 ) | ( ~n13294 & n18078 ) ;
  assign n18080 = ( ~n1818 & n2969 ) | ( ~n1818 & n16054 ) | ( n2969 & n16054 ) ;
  assign n18081 = ~n4257 & n10882 ;
  assign n18082 = n2216 & n18081 ;
  assign n18083 = ( ~n8256 & n11085 ) | ( ~n8256 & n11992 ) | ( n11085 & n11992 ) ;
  assign n18084 = n7372 & ~n12528 ;
  assign n18085 = ( ~n7939 & n16379 ) | ( ~n7939 & n18084 ) | ( n16379 & n18084 ) ;
  assign n18087 = ( ~n3503 & n3560 ) | ( ~n3503 & n8628 ) | ( n3560 & n8628 ) ;
  assign n18086 = n15970 ^ n2609 ^ n1913 ;
  assign n18088 = n18087 ^ n18086 ^ n5805 ;
  assign n18089 = n3463 | n6859 ;
  assign n18090 = n13173 ^ n5602 ^ n3788 ;
  assign n18091 = ( n1122 & ~n3363 ) | ( n1122 & n9817 ) | ( ~n3363 & n9817 ) ;
  assign n18092 = n18091 ^ n16622 ^ n1887 ;
  assign n18093 = n18092 ^ n9821 ^ 1'b0 ;
  assign n18094 = n18090 & n18093 ;
  assign n18098 = n1722 & ~n2919 ;
  assign n18099 = ~n572 & n18098 ;
  assign n18100 = n18099 ^ n13520 ^ n2399 ;
  assign n18101 = n18100 ^ n10981 ^ n10671 ;
  assign n18096 = ( n5830 & n6029 ) | ( n5830 & ~n12685 ) | ( n6029 & ~n12685 ) ;
  assign n18095 = ( ~n4146 & n10560 ) | ( ~n4146 & n11580 ) | ( n10560 & n11580 ) ;
  assign n18097 = n18096 ^ n18095 ^ n6068 ;
  assign n18102 = n18101 ^ n18097 ^ 1'b0 ;
  assign n18103 = ( ~n7533 & n13607 ) | ( ~n7533 & n16938 ) | ( n13607 & n16938 ) ;
  assign n18104 = ( ~n3199 & n4444 ) | ( ~n3199 & n13089 ) | ( n4444 & n13089 ) ;
  assign n18105 = n18104 ^ n15597 ^ n4364 ;
  assign n18106 = ( n14096 & ~n18103 ) | ( n14096 & n18105 ) | ( ~n18103 & n18105 ) ;
  assign n18109 = n3101 ^ n957 ^ x43 ;
  assign n18107 = ( n5029 & n8259 ) | ( n5029 & ~n15997 ) | ( n8259 & ~n15997 ) ;
  assign n18108 = ( n4082 & n7763 ) | ( n4082 & ~n18107 ) | ( n7763 & ~n18107 ) ;
  assign n18110 = n18109 ^ n18108 ^ 1'b0 ;
  assign n18111 = ( n1014 & n3679 ) | ( n1014 & ~n6630 ) | ( n3679 & ~n6630 ) ;
  assign n18112 = n15220 ^ n4637 ^ n1094 ;
  assign n18125 = ( ~n845 & n2245 ) | ( ~n845 & n5137 ) | ( n2245 & n5137 ) ;
  assign n18123 = n3501 | n13162 ;
  assign n18124 = n18123 ^ n2262 ^ 1'b0 ;
  assign n18126 = n18125 ^ n18124 ^ n9044 ;
  assign n18115 = ~n4333 & n9496 ;
  assign n18117 = n1986 ^ n1793 ^ n1690 ;
  assign n18118 = ( n1878 & ~n4338 ) | ( n1878 & n18117 ) | ( ~n4338 & n18117 ) ;
  assign n18116 = n16639 ^ n4077 ^ n1285 ;
  assign n18119 = n18118 ^ n18116 ^ n4897 ;
  assign n18120 = ( ~n4068 & n18115 ) | ( ~n4068 & n18119 ) | ( n18115 & n18119 ) ;
  assign n18121 = n9370 ^ n8510 ^ 1'b0 ;
  assign n18122 = n18120 & ~n18121 ;
  assign n18127 = n18126 ^ n18122 ^ n2494 ;
  assign n18113 = ( ~n7144 & n7478 ) | ( ~n7144 & n8694 ) | ( n7478 & n8694 ) ;
  assign n18114 = n18113 ^ n6581 ^ 1'b0 ;
  assign n18128 = n18127 ^ n18114 ^ n15973 ;
  assign n18129 = ( n6775 & n10468 ) | ( n6775 & n10809 ) | ( n10468 & n10809 ) ;
  assign n18130 = n12024 ^ n8472 ^ 1'b0 ;
  assign n18131 = n15724 ^ n14258 ^ 1'b0 ;
  assign n18132 = n15130 | n18131 ;
  assign n18133 = ~n5632 & n9098 ;
  assign n18134 = n18132 & n18133 ;
  assign n18135 = n18130 & ~n18134 ;
  assign n18136 = n8718 | n17144 ;
  assign n18137 = n18136 ^ n10487 ^ 1'b0 ;
  assign n18138 = ( n8811 & ~n16071 ) | ( n8811 & n17965 ) | ( ~n16071 & n17965 ) ;
  assign n18139 = n6243 | n18138 ;
  assign n18140 = n12769 ^ n1671 ^ 1'b0 ;
  assign n18141 = n18139 & n18140 ;
  assign n18142 = ( n919 & n2779 ) | ( n919 & n11721 ) | ( n2779 & n11721 ) ;
  assign n18143 = ( n227 & n2370 ) | ( n227 & n6501 ) | ( n2370 & n6501 ) ;
  assign n18144 = ( n369 & n3503 ) | ( n369 & n9190 ) | ( n3503 & n9190 ) ;
  assign n18151 = n7841 ^ n5248 ^ n3723 ;
  assign n18152 = n7224 | n18151 ;
  assign n18153 = n18152 ^ n2784 ^ n1843 ;
  assign n18154 = n17321 & ~n18153 ;
  assign n18155 = n18154 ^ n6275 ^ 1'b0 ;
  assign n18156 = n14977 ^ n10854 ^ n1281 ;
  assign n18157 = ( n643 & ~n18155 ) | ( n643 & n18156 ) | ( ~n18155 & n18156 ) ;
  assign n18158 = ( n6727 & n16594 ) | ( n6727 & n18157 ) | ( n16594 & n18157 ) ;
  assign n18148 = n1485 ^ n1432 ^ x5 ;
  assign n18146 = n15647 ^ n4807 ^ n3825 ;
  assign n18147 = n3841 | n18146 ;
  assign n18149 = n18148 ^ n18147 ^ n16680 ;
  assign n18150 = n18149 ^ n9972 ^ n3000 ;
  assign n18145 = ( n1102 & n9465 ) | ( n1102 & n10071 ) | ( n9465 & n10071 ) ;
  assign n18159 = n18158 ^ n18150 ^ n18145 ;
  assign n18160 = n11027 | n13668 ;
  assign n18161 = n18160 ^ n14418 ^ 1'b0 ;
  assign n18162 = n18161 ^ n10587 ^ n9607 ;
  assign n18163 = n16237 ^ n749 ^ 1'b0 ;
  assign n18171 = ( n715 & ~n2254 ) | ( n715 & n2633 ) | ( ~n2254 & n2633 ) ;
  assign n18172 = n18171 ^ n5739 ^ n685 ;
  assign n18167 = n14287 ^ n9717 ^ n5340 ;
  assign n18168 = ( n11252 & n14440 ) | ( n11252 & n18167 ) | ( n14440 & n18167 ) ;
  assign n18169 = n18168 ^ n14287 ^ n6312 ;
  assign n18170 = n18169 ^ n6672 ^ n2839 ;
  assign n18164 = n8358 ^ n3619 ^ x90 ;
  assign n18165 = ( ~n905 & n3261 ) | ( ~n905 & n18164 ) | ( n3261 & n18164 ) ;
  assign n18166 = ( n8992 & n14827 ) | ( n8992 & n18165 ) | ( n14827 & n18165 ) ;
  assign n18173 = n18172 ^ n18170 ^ n18166 ;
  assign n18174 = n16642 ^ n11814 ^ n9563 ;
  assign n18175 = ( n3230 & n13398 ) | ( n3230 & ~n14072 ) | ( n13398 & ~n14072 ) ;
  assign n18176 = n2381 ^ n1932 ^ n377 ;
  assign n18177 = n18176 ^ n5452 ^ n3561 ;
  assign n18178 = n8844 & n18177 ;
  assign n18179 = n18178 ^ n10209 ^ n3922 ;
  assign n18180 = n14442 ^ n11868 ^ n183 ;
  assign n18181 = ( n6667 & n14473 ) | ( n6667 & ~n18180 ) | ( n14473 & ~n18180 ) ;
  assign n18182 = ( n2200 & n3325 ) | ( n2200 & n10407 ) | ( n3325 & n10407 ) ;
  assign n18183 = ( ~x43 & n7401 ) | ( ~x43 & n18182 ) | ( n7401 & n18182 ) ;
  assign n18184 = n7267 ^ n5879 ^ n2449 ;
  assign n18185 = n18184 ^ n3593 ^ n2386 ;
  assign n18186 = ( n1521 & ~n16224 ) | ( n1521 & n18185 ) | ( ~n16224 & n18185 ) ;
  assign n18187 = n8663 ^ n6922 ^ n5942 ;
  assign n18188 = n18187 ^ n14654 ^ n8295 ;
  assign n18190 = n17755 ^ n9858 ^ n1294 ;
  assign n18191 = n18190 ^ n2607 ^ n1776 ;
  assign n18189 = ( n7576 & ~n13649 ) | ( n7576 & n15726 ) | ( ~n13649 & n15726 ) ;
  assign n18192 = n18191 ^ n18189 ^ n5442 ;
  assign n18193 = ( n7555 & n8184 ) | ( n7555 & ~n13339 ) | ( n8184 & ~n13339 ) ;
  assign n18194 = n8398 ^ n4711 ^ n4027 ;
  assign n18195 = ( n12136 & n18193 ) | ( n12136 & ~n18194 ) | ( n18193 & ~n18194 ) ;
  assign n18196 = n11375 ^ n9731 ^ n9321 ;
  assign n18198 = n12032 ^ n3707 ^ 1'b0 ;
  assign n18199 = n18198 ^ n17213 ^ 1'b0 ;
  assign n18197 = n12313 ^ n947 ^ 1'b0 ;
  assign n18200 = n18199 ^ n18197 ^ n6173 ;
  assign n18201 = ( n1278 & n4464 ) | ( n1278 & n9505 ) | ( n4464 & n9505 ) ;
  assign n18202 = ( n4163 & n15021 ) | ( n4163 & n18201 ) | ( n15021 & n18201 ) ;
  assign n18204 = ( n3404 & ~n3715 ) | ( n3404 & n5610 ) | ( ~n3715 & n5610 ) ;
  assign n18205 = ( n4274 & n15552 ) | ( n4274 & ~n18204 ) | ( n15552 & ~n18204 ) ;
  assign n18203 = n17995 ^ n13451 ^ n3941 ;
  assign n18206 = n18205 ^ n18203 ^ n5174 ;
  assign n18207 = n18206 ^ n1682 ^ 1'b0 ;
  assign n18208 = n18207 ^ n6555 ^ 1'b0 ;
  assign n18213 = n8528 ^ n3407 ^ 1'b0 ;
  assign n18212 = n7737 ^ n7467 ^ n837 ;
  assign n18209 = n14462 ^ n12365 ^ n4814 ;
  assign n18210 = n16582 ^ n12605 ^ n1936 ;
  assign n18211 = ( n13267 & n18209 ) | ( n13267 & n18210 ) | ( n18209 & n18210 ) ;
  assign n18214 = n18213 ^ n18212 ^ n18211 ;
  assign n18215 = ( ~n3138 & n12235 ) | ( ~n3138 & n17147 ) | ( n12235 & n17147 ) ;
  assign n18216 = ( ~n10996 & n11476 ) | ( ~n10996 & n18215 ) | ( n11476 & n18215 ) ;
  assign n18217 = n17200 ^ n14646 ^ n11563 ;
  assign n18218 = ( ~n797 & n1760 ) | ( ~n797 & n2912 ) | ( n1760 & n2912 ) ;
  assign n18219 = n9115 ^ n7745 ^ n3550 ;
  assign n18220 = n9305 & ~n9538 ;
  assign n18221 = n18219 & n18220 ;
  assign n18222 = n10154 ^ n7423 ^ 1'b0 ;
  assign n18223 = ( n18218 & ~n18221 ) | ( n18218 & n18222 ) | ( ~n18221 & n18222 ) ;
  assign n18227 = ( ~n6168 & n8594 ) | ( ~n6168 & n12959 ) | ( n8594 & n12959 ) ;
  assign n18224 = n6922 ^ n4965 ^ 1'b0 ;
  assign n18225 = n12445 ^ n6105 ^ n280 ;
  assign n18226 = ( n13354 & n18224 ) | ( n13354 & ~n18225 ) | ( n18224 & ~n18225 ) ;
  assign n18228 = n18227 ^ n18226 ^ n7056 ;
  assign n18229 = n5546 & ~n18228 ;
  assign n18230 = ( n377 & n7282 ) | ( n377 & n9245 ) | ( n7282 & n9245 ) ;
  assign n18231 = n18230 ^ n3420 ^ n3400 ;
  assign n18232 = n17011 ^ n12226 ^ n8804 ;
  assign n18233 = n4397 & ~n18232 ;
  assign n18234 = ( ~n5520 & n11205 ) | ( ~n5520 & n13554 ) | ( n11205 & n13554 ) ;
  assign n18235 = ( n3389 & n6228 ) | ( n3389 & ~n7888 ) | ( n6228 & ~n7888 ) ;
  assign n18237 = ( n5019 & n7308 ) | ( n5019 & n12423 ) | ( n7308 & n12423 ) ;
  assign n18236 = ( n4627 & n14041 ) | ( n4627 & n16393 ) | ( n14041 & n16393 ) ;
  assign n18238 = n18237 ^ n18236 ^ n9696 ;
  assign n18239 = ( n18234 & n18235 ) | ( n18234 & n18238 ) | ( n18235 & n18238 ) ;
  assign n18240 = ( ~n6065 & n8811 ) | ( ~n6065 & n18239 ) | ( n8811 & n18239 ) ;
  assign n18241 = n18240 ^ n4234 ^ n3788 ;
  assign n18245 = n7991 | n9707 ;
  assign n18243 = ( ~n6231 & n8489 ) | ( ~n6231 & n9607 ) | ( n8489 & n9607 ) ;
  assign n18244 = ~n2842 & n18243 ;
  assign n18246 = n18245 ^ n18244 ^ 1'b0 ;
  assign n18242 = n168 & ~n9936 ;
  assign n18247 = n18246 ^ n18242 ^ 1'b0 ;
  assign n18248 = n15395 ^ n8509 ^ n6782 ;
  assign n18249 = n18006 ^ n3107 ^ n1056 ;
  assign n18250 = ( n7315 & n12548 ) | ( n7315 & n18249 ) | ( n12548 & n18249 ) ;
  assign n18251 = ( n1732 & n2420 ) | ( n1732 & n4176 ) | ( n2420 & n4176 ) ;
  assign n18252 = n2582 & ~n18251 ;
  assign n18253 = n18252 ^ n8234 ^ 1'b0 ;
  assign n18254 = n18253 ^ n7794 ^ 1'b0 ;
  assign n18255 = ( n18248 & n18250 ) | ( n18248 & ~n18254 ) | ( n18250 & ~n18254 ) ;
  assign n18256 = ~n2812 & n6304 ;
  assign n18257 = n4393 | n11554 ;
  assign n18258 = n18256 | n18257 ;
  assign n18259 = n14788 ^ n11775 ^ n8599 ;
  assign n18260 = ( n5106 & ~n9716 ) | ( n5106 & n18259 ) | ( ~n9716 & n18259 ) ;
  assign n18261 = ( n5547 & n18258 ) | ( n5547 & ~n18260 ) | ( n18258 & ~n18260 ) ;
  assign n18262 = n7076 & ~n8223 ;
  assign n18263 = n18262 ^ n7386 ^ 1'b0 ;
  assign n18264 = ~n7194 & n8315 ;
  assign n18265 = n3293 | n9178 ;
  assign n18266 = n18264 & ~n18265 ;
  assign n18270 = n11891 ^ n5530 ^ n403 ;
  assign n18267 = ~n2379 & n3788 ;
  assign n18268 = n18267 ^ n6354 ^ 1'b0 ;
  assign n18269 = ( ~n683 & n11858 ) | ( ~n683 & n18268 ) | ( n11858 & n18268 ) ;
  assign n18271 = n18270 ^ n18269 ^ n15300 ;
  assign n18272 = ( ~n4709 & n6045 ) | ( ~n4709 & n11336 ) | ( n6045 & n11336 ) ;
  assign n18273 = n13582 ^ n8829 ^ n7349 ;
  assign n18274 = n13775 ^ n3630 ^ n630 ;
  assign n18275 = ( n666 & n18273 ) | ( n666 & ~n18274 ) | ( n18273 & ~n18274 ) ;
  assign n18276 = n4687 ^ n674 ^ n580 ;
  assign n18277 = n18276 ^ n9793 ^ n3195 ;
  assign n18278 = n18277 ^ n9445 ^ n7875 ;
  assign n18279 = n17537 ^ n15604 ^ 1'b0 ;
  assign n18280 = n13799 ^ n13544 ^ n3230 ;
  assign n18281 = ( n3791 & ~n17665 ) | ( n3791 & n18280 ) | ( ~n17665 & n18280 ) ;
  assign n18282 = ( n1442 & ~n8817 ) | ( n1442 & n11356 ) | ( ~n8817 & n11356 ) ;
  assign n18283 = n18282 ^ n8853 ^ 1'b0 ;
  assign n18284 = n4888 ^ x27 ^ 1'b0 ;
  assign n18285 = n2046 & n18284 ;
  assign n18287 = n8079 ^ n7392 ^ n1597 ;
  assign n18288 = n18287 ^ n2590 ^ 1'b0 ;
  assign n18289 = n14738 & ~n18288 ;
  assign n18286 = n5439 ^ n4574 ^ n1623 ;
  assign n18290 = n18289 ^ n18286 ^ n3136 ;
  assign n18295 = ( n909 & ~n4075 ) | ( n909 & n6159 ) | ( ~n4075 & n6159 ) ;
  assign n18293 = n15966 ^ n4782 ^ 1'b0 ;
  assign n18294 = n6176 & ~n18293 ;
  assign n18296 = n18295 ^ n18294 ^ n2843 ;
  assign n18291 = ( ~n3714 & n15395 ) | ( ~n3714 & n17300 ) | ( n15395 & n17300 ) ;
  assign n18292 = ( n5115 & n15670 ) | ( n5115 & ~n18291 ) | ( n15670 & ~n18291 ) ;
  assign n18297 = n18296 ^ n18292 ^ n4566 ;
  assign n18298 = n18297 ^ n18251 ^ n1943 ;
  assign n18299 = ( ~n1795 & n3440 ) | ( ~n1795 & n6039 ) | ( n3440 & n6039 ) ;
  assign n18300 = n10117 ^ n9231 ^ n4961 ;
  assign n18303 = n7645 ^ n4582 ^ n190 ;
  assign n18301 = n10910 ^ n8614 ^ n2073 ;
  assign n18302 = ( ~n8211 & n10604 ) | ( ~n8211 & n18301 ) | ( n10604 & n18301 ) ;
  assign n18304 = n18303 ^ n18302 ^ n8645 ;
  assign n18305 = n14580 | n18304 ;
  assign n18306 = n18305 ^ n1790 ^ 1'b0 ;
  assign n18307 = ( n18299 & n18300 ) | ( n18299 & n18306 ) | ( n18300 & n18306 ) ;
  assign n18311 = ( n5484 & n8250 ) | ( n5484 & n9334 ) | ( n8250 & n9334 ) ;
  assign n18312 = n18311 ^ n9767 ^ n1333 ;
  assign n18310 = ~n3042 & n8151 ;
  assign n18308 = n11026 ^ n8314 ^ n2478 ;
  assign n18309 = n18308 ^ n3365 ^ 1'b0 ;
  assign n18313 = n18312 ^ n18310 ^ n18309 ;
  assign n18316 = ( x0 & n6542 ) | ( x0 & n8089 ) | ( n6542 & n8089 ) ;
  assign n18317 = n18316 ^ n7541 ^ n5746 ;
  assign n18318 = n5300 & n12260 ;
  assign n18319 = n18318 ^ n2724 ^ 1'b0 ;
  assign n18320 = n18319 ^ n7573 ^ n879 ;
  assign n18321 = n4770 & ~n18320 ;
  assign n18322 = n18321 ^ n12795 ^ n9877 ;
  assign n18323 = ( n3176 & n18317 ) | ( n3176 & n18322 ) | ( n18317 & n18322 ) ;
  assign n18314 = n4392 & ~n9957 ;
  assign n18315 = ~x82 & n18314 ;
  assign n18324 = n18323 ^ n18315 ^ n4096 ;
  assign n18325 = n14834 ^ n10447 ^ n2941 ;
  assign n18326 = ( ~n1151 & n9891 ) | ( ~n1151 & n18325 ) | ( n9891 & n18325 ) ;
  assign n18327 = n9920 ^ n9212 ^ 1'b0 ;
  assign n18328 = ~n18326 & n18327 ;
  assign n18329 = n5348 ^ n1006 ^ 1'b0 ;
  assign n18330 = n2082 | n18329 ;
  assign n18331 = ( n429 & n5504 ) | ( n429 & ~n7522 ) | ( n5504 & ~n7522 ) ;
  assign n18332 = n15058 ^ n7359 ^ n5668 ;
  assign n18333 = ( ~n3636 & n7411 ) | ( ~n3636 & n18332 ) | ( n7411 & n18332 ) ;
  assign n18334 = n10779 ^ n8739 ^ n4620 ;
  assign n18335 = n9042 ^ n4021 ^ 1'b0 ;
  assign n18336 = n12617 ^ n9174 ^ n3253 ;
  assign n18337 = ( ~n13324 & n18335 ) | ( ~n13324 & n18336 ) | ( n18335 & n18336 ) ;
  assign n18338 = n7187 ^ n3804 ^ 1'b0 ;
  assign n18339 = n4510 & n18338 ;
  assign n18340 = n4313 & n18339 ;
  assign n18341 = n4494 & n18340 ;
  assign n18342 = n7191 & ~n8936 ;
  assign n18343 = n18342 ^ n966 ^ n959 ;
  assign n18344 = n1912 & ~n3500 ;
  assign n18345 = n18344 ^ n11691 ^ 1'b0 ;
  assign n18346 = n18345 ^ n7877 ^ n1310 ;
  assign n18347 = n15555 ^ n9217 ^ n4939 ;
  assign n18348 = ( n1662 & n16028 ) | ( n1662 & n18347 ) | ( n16028 & n18347 ) ;
  assign n18349 = n11715 ^ n9274 ^ n3849 ;
  assign n18350 = n15464 ^ n1300 ^ 1'b0 ;
  assign n18351 = ~n18349 & n18350 ;
  assign n18352 = ( x17 & ~n14002 ) | ( x17 & n18351 ) | ( ~n14002 & n18351 ) ;
  assign n18353 = ( ~n988 & n4646 ) | ( ~n988 & n18352 ) | ( n4646 & n18352 ) ;
  assign n18354 = ( n1480 & n3457 ) | ( n1480 & n13080 ) | ( n3457 & n13080 ) ;
  assign n18355 = n5776 & n7602 ;
  assign n18356 = n18355 ^ n1579 ^ 1'b0 ;
  assign n18357 = n11165 & ~n18356 ;
  assign n18358 = n1174 & ~n18357 ;
  assign n18359 = ~n859 & n18358 ;
  assign n18360 = ( n4068 & n7087 ) | ( n4068 & n16572 ) | ( n7087 & n16572 ) ;
  assign n18361 = n9507 ^ n8486 ^ n247 ;
  assign n18362 = n18361 ^ n10200 ^ n4457 ;
  assign n18363 = n7833 ^ n3211 ^ n1941 ;
  assign n18364 = n16834 ^ n3828 ^ 1'b0 ;
  assign n18369 = n9645 ^ n4733 ^ n2463 ;
  assign n18366 = ( n627 & n1938 ) | ( n627 & n11187 ) | ( n1938 & n11187 ) ;
  assign n18367 = n18366 ^ n1891 ^ n1371 ;
  assign n18368 = ( n6988 & n12015 ) | ( n6988 & n18367 ) | ( n12015 & n18367 ) ;
  assign n18365 = ( n2569 & n3277 ) | ( n2569 & ~n6633 ) | ( n3277 & ~n6633 ) ;
  assign n18370 = n18369 ^ n18368 ^ n18365 ;
  assign n18371 = n2830 & n15395 ;
  assign n18372 = ( n4381 & ~n6116 ) | ( n4381 & n6845 ) | ( ~n6116 & n6845 ) ;
  assign n18373 = ( n2153 & ~n15656 ) | ( n2153 & n18372 ) | ( ~n15656 & n18372 ) ;
  assign n18374 = n18373 ^ n3141 ^ n1121 ;
  assign n18375 = n3536 & n8340 ;
  assign n18376 = n18375 ^ n7168 ^ 1'b0 ;
  assign n18377 = ( n1789 & ~n3113 ) | ( n1789 & n18376 ) | ( ~n3113 & n18376 ) ;
  assign n18378 = n10523 ^ n451 ^ 1'b0 ;
  assign n18379 = n4195 ^ n3320 ^ n847 ;
  assign n18380 = ( n11737 & ~n14448 ) | ( n11737 & n18379 ) | ( ~n14448 & n18379 ) ;
  assign n18381 = ( n8369 & ~n18378 ) | ( n8369 & n18380 ) | ( ~n18378 & n18380 ) ;
  assign n18382 = ~n1374 & n4213 ;
  assign n18383 = ( n3120 & n13128 ) | ( n3120 & n18382 ) | ( n13128 & n18382 ) ;
  assign n18384 = ( n1862 & n9643 ) | ( n1862 & ~n18383 ) | ( n9643 & ~n18383 ) ;
  assign n18385 = ( ~n14168 & n18002 ) | ( ~n14168 & n18384 ) | ( n18002 & n18384 ) ;
  assign n18386 = n5361 & n14762 ;
  assign n18387 = n18385 & n18386 ;
  assign n18388 = n11986 ^ n2357 ^ n2123 ;
  assign n18389 = ( n7735 & ~n14098 ) | ( n7735 & n18388 ) | ( ~n14098 & n18388 ) ;
  assign n18390 = n18164 ^ n16160 ^ 1'b0 ;
  assign n18391 = ~n3281 & n18390 ;
  assign n18395 = n4794 ^ n3008 ^ 1'b0 ;
  assign n18393 = n7938 ^ n6265 ^ 1'b0 ;
  assign n18394 = ( ~n6900 & n12226 ) | ( ~n6900 & n18393 ) | ( n12226 & n18393 ) ;
  assign n18396 = n18395 ^ n18394 ^ n11594 ;
  assign n18392 = ~n1105 & n7903 ;
  assign n18397 = n18396 ^ n18392 ^ 1'b0 ;
  assign n18398 = ( ~n8229 & n18391 ) | ( ~n8229 & n18397 ) | ( n18391 & n18397 ) ;
  assign n18399 = ( n9906 & n14249 ) | ( n9906 & n18398 ) | ( n14249 & n18398 ) ;
  assign n18400 = n340 | n4140 ;
  assign n18401 = ( n8611 & ~n11574 ) | ( n8611 & n18400 ) | ( ~n11574 & n18400 ) ;
  assign n18402 = n18401 ^ n13457 ^ n1937 ;
  assign n18403 = n4062 ^ n2966 ^ n2913 ;
  assign n18404 = n18403 ^ n9556 ^ n4046 ;
  assign n18405 = ( n3496 & n13746 ) | ( n3496 & ~n18404 ) | ( n13746 & ~n18404 ) ;
  assign n18406 = ( n3800 & n4400 ) | ( n3800 & ~n14489 ) | ( n4400 & ~n14489 ) ;
  assign n18407 = ( n1211 & ~n6954 ) | ( n1211 & n18406 ) | ( ~n6954 & n18406 ) ;
  assign n18408 = ( n15838 & n18405 ) | ( n15838 & n18407 ) | ( n18405 & n18407 ) ;
  assign n18409 = n5980 ^ n3374 ^ n1558 ;
  assign n18421 = n12529 ^ n4721 ^ 1'b0 ;
  assign n18417 = ( n3682 & ~n6268 ) | ( n3682 & n10347 ) | ( ~n6268 & n10347 ) ;
  assign n18415 = n5731 & ~n7283 ;
  assign n18416 = n8858 & n18415 ;
  assign n18418 = n18417 ^ n18416 ^ n2047 ;
  assign n18419 = ( n345 & n2985 ) | ( n345 & n18418 ) | ( n2985 & n18418 ) ;
  assign n18411 = n11829 ^ n3144 ^ n1217 ;
  assign n18412 = ( n2853 & n7332 ) | ( n2853 & ~n18411 ) | ( n7332 & ~n18411 ) ;
  assign n18410 = n7484 ^ n5318 ^ n3701 ;
  assign n18413 = n18412 ^ n18410 ^ n6284 ;
  assign n18414 = ~n12700 & n18413 ;
  assign n18420 = n18419 ^ n18414 ^ n2902 ;
  assign n18422 = n18421 ^ n18420 ^ n17039 ;
  assign n18423 = n10197 ^ n8921 ^ n3653 ;
  assign n18424 = n14318 ^ n1652 ^ 1'b0 ;
  assign n18425 = n18423 | n18424 ;
  assign n18431 = n6663 ^ n3897 ^ n1993 ;
  assign n18432 = n4569 | n18431 ;
  assign n18426 = n653 & ~n9412 ;
  assign n18427 = n18300 ^ n8044 ^ n3166 ;
  assign n18428 = n18427 ^ n3169 ^ 1'b0 ;
  assign n18429 = n18426 | n18428 ;
  assign n18430 = n18429 ^ n9727 ^ n8630 ;
  assign n18433 = n18432 ^ n18430 ^ n15203 ;
  assign n18434 = n11439 ^ n9115 ^ n6230 ;
  assign n18435 = ( n14314 & ~n16015 ) | ( n14314 & n17826 ) | ( ~n16015 & n17826 ) ;
  assign n18439 = ( n374 & n2286 ) | ( n374 & ~n2355 ) | ( n2286 & ~n2355 ) ;
  assign n18436 = ( n5096 & n7157 ) | ( n5096 & ~n8924 ) | ( n7157 & ~n8924 ) ;
  assign n18437 = n18436 ^ n3826 ^ n390 ;
  assign n18438 = ( n2966 & ~n5062 ) | ( n2966 & n18437 ) | ( ~n5062 & n18437 ) ;
  assign n18440 = n18439 ^ n18438 ^ n6784 ;
  assign n18441 = ( n3889 & n11191 ) | ( n3889 & ~n17652 ) | ( n11191 & ~n17652 ) ;
  assign n18442 = ( n5253 & n9721 ) | ( n5253 & ~n18441 ) | ( n9721 & ~n18441 ) ;
  assign n18443 = ( n1558 & ~n4794 ) | ( n1558 & n11816 ) | ( ~n4794 & n11816 ) ;
  assign n18444 = ( n6279 & n17915 ) | ( n6279 & ~n18443 ) | ( n17915 & ~n18443 ) ;
  assign n18445 = n7293 ^ n7129 ^ n412 ;
  assign n18446 = n18445 ^ n6633 ^ x27 ;
  assign n18447 = n14813 ^ n1700 ^ 1'b0 ;
  assign n18448 = n18447 ^ n396 ^ 1'b0 ;
  assign n18449 = ( n1414 & ~n15929 ) | ( n1414 & n18448 ) | ( ~n15929 & n18448 ) ;
  assign n18450 = n5836 ^ n1753 ^ n294 ;
  assign n18451 = ( n492 & ~n8061 ) | ( n492 & n18245 ) | ( ~n8061 & n18245 ) ;
  assign n18452 = ( n1185 & n18450 ) | ( n1185 & ~n18451 ) | ( n18450 & ~n18451 ) ;
  assign n18453 = ( n8550 & ~n10288 ) | ( n8550 & n10394 ) | ( ~n10288 & n10394 ) ;
  assign n18454 = ( n3135 & ~n4768 ) | ( n3135 & n18453 ) | ( ~n4768 & n18453 ) ;
  assign n18455 = n9591 ^ n7148 ^ n2980 ;
  assign n18456 = n7490 & n18455 ;
  assign n18457 = n18456 ^ x91 ^ 1'b0 ;
  assign n18458 = ( n1055 & n1587 ) | ( n1055 & ~n18457 ) | ( n1587 & ~n18457 ) ;
  assign n18459 = n6416 ^ n5538 ^ n1762 ;
  assign n18460 = ( n8621 & n10479 ) | ( n8621 & ~n18459 ) | ( n10479 & ~n18459 ) ;
  assign n18461 = ( n4141 & n7057 ) | ( n4141 & ~n18460 ) | ( n7057 & ~n18460 ) ;
  assign n18462 = ( ~n7987 & n18458 ) | ( ~n7987 & n18461 ) | ( n18458 & n18461 ) ;
  assign n18463 = ( n14869 & ~n18454 ) | ( n14869 & n18462 ) | ( ~n18454 & n18462 ) ;
  assign n18464 = n15623 ^ n15347 ^ n9662 ;
  assign n18466 = n6636 ^ n5869 ^ n2790 ;
  assign n18467 = ( n6629 & ~n9284 ) | ( n6629 & n14894 ) | ( ~n9284 & n14894 ) ;
  assign n18468 = ~n9518 & n18467 ;
  assign n18469 = ( n7144 & ~n18466 ) | ( n7144 & n18468 ) | ( ~n18466 & n18468 ) ;
  assign n18470 = n3217 | n18469 ;
  assign n18471 = n10469 & ~n18470 ;
  assign n18465 = n514 & n2777 ;
  assign n18472 = n18471 ^ n18465 ^ 1'b0 ;
  assign n18473 = ( n2308 & n13585 ) | ( n2308 & n16484 ) | ( n13585 & n16484 ) ;
  assign n18474 = ( n3779 & n10257 ) | ( n3779 & ~n18473 ) | ( n10257 & ~n18473 ) ;
  assign n18476 = n12751 ^ n8836 ^ n517 ;
  assign n18475 = n15048 ^ n11200 ^ n10961 ;
  assign n18477 = n18476 ^ n18475 ^ n18455 ;
  assign n18481 = n6169 ^ n2734 ^ n1930 ;
  assign n18482 = ( n2605 & n6362 ) | ( n2605 & n18481 ) | ( n6362 & n18481 ) ;
  assign n18483 = ( n5038 & ~n6230 ) | ( n5038 & n18482 ) | ( ~n6230 & n18482 ) ;
  assign n18478 = n13133 ^ n7988 ^ n1606 ;
  assign n18479 = ( ~n524 & n7181 ) | ( ~n524 & n18478 ) | ( n7181 & n18478 ) ;
  assign n18480 = n18479 ^ n16447 ^ n8877 ;
  assign n18484 = n18483 ^ n18480 ^ 1'b0 ;
  assign n18485 = n18199 & ~n18484 ;
  assign n18488 = n6069 | n7251 ;
  assign n18486 = n13370 ^ n3775 ^ n1459 ;
  assign n18487 = n18486 ^ n17378 ^ n8059 ;
  assign n18489 = n18488 ^ n18487 ^ n1684 ;
  assign n18491 = ( n1283 & ~n1365 ) | ( n1283 & n17607 ) | ( ~n1365 & n17607 ) ;
  assign n18490 = ( n3630 & n6511 ) | ( n3630 & ~n14889 ) | ( n6511 & ~n14889 ) ;
  assign n18492 = n18491 ^ n18490 ^ n5908 ;
  assign n18493 = n2211 & n18492 ;
  assign n18494 = ( n5625 & ~n18224 ) | ( n5625 & n18493 ) | ( ~n18224 & n18493 ) ;
  assign n18496 = n10067 ^ n6263 ^ n5052 ;
  assign n18495 = n9558 ^ n7767 ^ n2251 ;
  assign n18497 = n18496 ^ n18495 ^ n18391 ;
  assign n18498 = n9303 & ~n18497 ;
  assign n18499 = ( n950 & n2888 ) | ( n950 & n3229 ) | ( n2888 & n3229 ) ;
  assign n18500 = n18499 ^ n13226 ^ n4297 ;
  assign n18501 = n18287 ^ n14654 ^ 1'b0 ;
  assign n18502 = ( n14364 & ~n18500 ) | ( n14364 & n18501 ) | ( ~n18500 & n18501 ) ;
  assign n18505 = n7961 ^ n7541 ^ n1240 ;
  assign n18506 = n18505 ^ n5865 ^ n5002 ;
  assign n18507 = ( ~n5985 & n8458 ) | ( ~n5985 & n18506 ) | ( n8458 & n18506 ) ;
  assign n18508 = n18507 ^ n9670 ^ 1'b0 ;
  assign n18503 = ( n138 & ~n2039 ) | ( n138 & n11842 ) | ( ~n2039 & n11842 ) ;
  assign n18504 = ( n6961 & ~n9494 ) | ( n6961 & n18503 ) | ( ~n9494 & n18503 ) ;
  assign n18509 = n18508 ^ n18504 ^ n9634 ;
  assign n18510 = ~n2528 & n5594 ;
  assign n18511 = n2977 ^ n1680 ^ x58 ;
  assign n18512 = n18511 ^ n9249 ^ 1'b0 ;
  assign n18513 = ~n8730 & n18512 ;
  assign n18514 = n6271 ^ n6083 ^ n839 ;
  assign n18515 = n6709 & n18514 ;
  assign n18516 = n18515 ^ n12342 ^ 1'b0 ;
  assign n18517 = ( n232 & ~n2557 ) | ( n232 & n12533 ) | ( ~n2557 & n12533 ) ;
  assign n18518 = n18517 ^ n12244 ^ n5122 ;
  assign n18519 = n10083 & n18518 ;
  assign n18520 = ~n2269 & n18519 ;
  assign n18521 = n5278 & ~n10380 ;
  assign n18522 = n5223 ^ n2019 ^ 1'b0 ;
  assign n18523 = n10557 ^ n10125 ^ n1210 ;
  assign n18524 = n2458 & ~n2704 ;
  assign n18525 = n18523 & n18524 ;
  assign n18526 = ( n12604 & n18522 ) | ( n12604 & ~n18525 ) | ( n18522 & ~n18525 ) ;
  assign n18527 = n18526 ^ n9103 ^ n6010 ;
  assign n18528 = ( ~n15021 & n17337 ) | ( ~n15021 & n17787 ) | ( n17337 & n17787 ) ;
  assign n18529 = ( ~n9140 & n13802 ) | ( ~n9140 & n18528 ) | ( n13802 & n18528 ) ;
  assign n18530 = n11925 ^ n2597 ^ 1'b0 ;
  assign n18531 = n18530 ^ n16987 ^ n6563 ;
  assign n18532 = n4663 ^ n1545 ^ 1'b0 ;
  assign n18533 = n18531 | n18532 ;
  assign n18534 = n18533 ^ n8748 ^ 1'b0 ;
  assign n18535 = n14082 ^ n9568 ^ n9425 ;
  assign n18536 = n18535 ^ n557 ^ n207 ;
  assign n18537 = n16521 ^ n2642 ^ n750 ;
  assign n18539 = n542 & n5476 ;
  assign n18538 = ( n10356 & ~n12800 ) | ( n10356 & n17101 ) | ( ~n12800 & n17101 ) ;
  assign n18540 = n18539 ^ n18538 ^ n4120 ;
  assign n18541 = n8528 ^ n8309 ^ n1262 ;
  assign n18542 = ( n804 & ~n16781 ) | ( n804 & n18541 ) | ( ~n16781 & n18541 ) ;
  assign n18543 = ( n5551 & ~n18540 ) | ( n5551 & n18542 ) | ( ~n18540 & n18542 ) ;
  assign n18544 = ~n2934 & n18543 ;
  assign n18545 = ~n18537 & n18544 ;
  assign n18546 = ~n1817 & n3407 ;
  assign n18547 = n18546 ^ n11286 ^ 1'b0 ;
  assign n18548 = n8046 ^ n4470 ^ n2775 ;
  assign n18549 = n18548 ^ n12541 ^ n10150 ;
  assign n18550 = ~n7829 & n8343 ;
  assign n18551 = n3702 & n12988 ;
  assign n18552 = n7176 ^ n3711 ^ n3275 ;
  assign n18553 = n18552 ^ n10516 ^ n3708 ;
  assign n18554 = n18553 ^ n10460 ^ n2209 ;
  assign n18555 = n18554 ^ n8451 ^ n1805 ;
  assign n18556 = ( n1511 & ~n8006 ) | ( n1511 & n11564 ) | ( ~n8006 & n11564 ) ;
  assign n18557 = ( n671 & n3561 ) | ( n671 & ~n18556 ) | ( n3561 & ~n18556 ) ;
  assign n18558 = n18250 ^ n1330 ^ n947 ;
  assign n18559 = ( ~n12370 & n18557 ) | ( ~n12370 & n18558 ) | ( n18557 & n18558 ) ;
  assign n18560 = n4733 & ~n18559 ;
  assign n18561 = n18560 ^ n14416 ^ 1'b0 ;
  assign n18562 = n7556 ^ n4052 ^ n1874 ;
  assign n18563 = ( ~n1273 & n12615 ) | ( ~n1273 & n18562 ) | ( n12615 & n18562 ) ;
  assign n18564 = n18563 ^ n14158 ^ n4055 ;
  assign n18566 = ( n1874 & n7311 ) | ( n1874 & n15892 ) | ( n7311 & n15892 ) ;
  assign n18565 = n6090 ^ n2342 ^ n780 ;
  assign n18567 = n18566 ^ n18565 ^ n3661 ;
  assign n18568 = n8594 ^ n2553 ^ n1077 ;
  assign n18569 = n18568 ^ n7608 ^ 1'b0 ;
  assign n18570 = n4178 & ~n10557 ;
  assign n18571 = n18570 ^ n4110 ^ 1'b0 ;
  assign n18572 = n14640 | n18571 ;
  assign n18573 = ( ~n6921 & n18569 ) | ( ~n6921 & n18572 ) | ( n18569 & n18572 ) ;
  assign n18574 = ( n14809 & n18567 ) | ( n14809 & n18573 ) | ( n18567 & n18573 ) ;
  assign n18575 = n2038 | n6282 ;
  assign n18576 = ( ~n1939 & n5983 ) | ( ~n1939 & n18575 ) | ( n5983 & n18575 ) ;
  assign n18577 = n7130 | n18576 ;
  assign n18578 = n18577 ^ n6886 ^ n3206 ;
  assign n18579 = ( n9004 & ~n11798 ) | ( n9004 & n18578 ) | ( ~n11798 & n18578 ) ;
  assign n18580 = n18579 ^ n6436 ^ n5284 ;
  assign n18581 = ( n3266 & ~n3267 ) | ( n3266 & n8986 ) | ( ~n3267 & n8986 ) ;
  assign n18582 = ~n4501 & n18581 ;
  assign n18583 = n18582 ^ n14068 ^ 1'b0 ;
  assign n18584 = n10955 & n18583 ;
  assign n18585 = ~n18580 & n18584 ;
  assign n18586 = n14098 & n18585 ;
  assign n18587 = ( ~n6789 & n7981 ) | ( ~n6789 & n10643 ) | ( n7981 & n10643 ) ;
  assign n18588 = n4482 ^ n4220 ^ n1269 ;
  assign n18589 = n8602 ^ n3226 ^ 1'b0 ;
  assign n18590 = ( ~n6754 & n18588 ) | ( ~n6754 & n18589 ) | ( n18588 & n18589 ) ;
  assign n18591 = n13876 ^ n5328 ^ 1'b0 ;
  assign n18592 = n4425 & ~n4446 ;
  assign n18593 = ~n4071 & n18592 ;
  assign n18594 = n18593 ^ n18451 ^ n3680 ;
  assign n18595 = n571 | n5833 ;
  assign n18596 = n18595 ^ n10904 ^ 1'b0 ;
  assign n18597 = ( n8416 & ~n13478 ) | ( n8416 & n14513 ) | ( ~n13478 & n14513 ) ;
  assign n18598 = ( n7011 & ~n11323 ) | ( n7011 & n18597 ) | ( ~n11323 & n18597 ) ;
  assign n18599 = n18598 ^ n10516 ^ n2293 ;
  assign n18600 = n18599 ^ n12170 ^ n4367 ;
  assign n18601 = ( n4354 & n17237 ) | ( n4354 & n18600 ) | ( n17237 & n18600 ) ;
  assign n18602 = n14656 ^ n5326 ^ n2541 ;
  assign n18603 = ( n5853 & ~n7607 ) | ( n5853 & n18602 ) | ( ~n7607 & n18602 ) ;
  assign n18604 = n16832 ^ n10599 ^ n10219 ;
  assign n18605 = n18604 ^ n14783 ^ n8086 ;
  assign n18606 = n1143 & n4397 ;
  assign n18607 = ( ~n2417 & n12423 ) | ( ~n2417 & n18606 ) | ( n12423 & n18606 ) ;
  assign n18608 = n1515 ^ n812 ^ 1'b0 ;
  assign n18609 = ~n11138 & n18608 ;
  assign n18610 = ( n3244 & n12923 ) | ( n3244 & ~n18609 ) | ( n12923 & ~n18609 ) ;
  assign n18611 = ( x28 & ~n6869 ) | ( x28 & n8408 ) | ( ~n6869 & n8408 ) ;
  assign n18612 = n18611 ^ n3956 ^ n3505 ;
  assign n18613 = n18612 ^ n7133 ^ n408 ;
  assign n18614 = n18613 ^ n4565 ^ 1'b0 ;
  assign n18615 = ~n10675 & n18614 ;
  assign n18616 = n10328 & ~n11439 ;
  assign n18617 = n18616 ^ n17257 ^ n17092 ;
  assign n18618 = n18617 ^ n7513 ^ 1'b0 ;
  assign n18619 = n18481 ^ n12708 ^ n5021 ;
  assign n18620 = ( n3710 & ~n6757 ) | ( n3710 & n11244 ) | ( ~n6757 & n11244 ) ;
  assign n18621 = n18620 ^ n2940 ^ n626 ;
  assign n18622 = ( ~n442 & n8845 ) | ( ~n442 & n18621 ) | ( n8845 & n18621 ) ;
  assign n18623 = ( n2630 & n9793 ) | ( n2630 & n15517 ) | ( n9793 & n15517 ) ;
  assign n18624 = ( n18619 & n18622 ) | ( n18619 & ~n18623 ) | ( n18622 & ~n18623 ) ;
  assign n18625 = ( n1574 & n11064 ) | ( n1574 & n18624 ) | ( n11064 & n18624 ) ;
  assign n18626 = ( n2334 & n5423 ) | ( n2334 & ~n18625 ) | ( n5423 & ~n18625 ) ;
  assign n18627 = n10067 ^ n7072 ^ n6388 ;
  assign n18628 = n18627 ^ n16272 ^ n537 ;
  assign n18629 = n18558 ^ n16054 ^ n14868 ;
  assign n18630 = ( n908 & n2874 ) | ( n908 & ~n4929 ) | ( n2874 & ~n4929 ) ;
  assign n18631 = n6306 ^ n1433 ^ 1'b0 ;
  assign n18632 = n5444 & n18631 ;
  assign n18633 = n18632 ^ n17534 ^ n14258 ;
  assign n18634 = ( n10315 & n18630 ) | ( n10315 & ~n18633 ) | ( n18630 & ~n18633 ) ;
  assign n18635 = n647 & ~n11195 ;
  assign n18636 = n17701 ^ n10643 ^ n4251 ;
  assign n18637 = ( n13976 & n15609 ) | ( n13976 & ~n18636 ) | ( n15609 & ~n18636 ) ;
  assign n18638 = ( n10242 & ~n11570 ) | ( n10242 & n11722 ) | ( ~n11570 & n11722 ) ;
  assign n18639 = n18638 ^ n8472 ^ n2221 ;
  assign n18640 = n4343 | n4838 ;
  assign n18641 = ( n8748 & ~n13633 ) | ( n8748 & n18640 ) | ( ~n13633 & n18640 ) ;
  assign n18642 = n1713 & n17060 ;
  assign n18643 = ( n2604 & n11387 ) | ( n2604 & ~n18642 ) | ( n11387 & ~n18642 ) ;
  assign n18645 = n2456 ^ n1753 ^ n622 ;
  assign n18644 = ( ~n8966 & n9878 ) | ( ~n8966 & n11847 ) | ( n9878 & n11847 ) ;
  assign n18646 = n18645 ^ n18644 ^ n11254 ;
  assign n18647 = n1289 & n18646 ;
  assign n18648 = n18647 ^ n4118 ^ 1'b0 ;
  assign n18649 = n14029 ^ n4322 ^ n3743 ;
  assign n18650 = ~n4569 & n18649 ;
  assign n18651 = ( n11308 & n15630 ) | ( n11308 & ~n18650 ) | ( n15630 & ~n18650 ) ;
  assign n18652 = ( n3224 & n4772 ) | ( n3224 & n9568 ) | ( n4772 & n9568 ) ;
  assign n18653 = n5062 & n18652 ;
  assign n18654 = n17288 ^ n7553 ^ x1 ;
  assign n18655 = ~n16950 & n18654 ;
  assign n18656 = ( n1462 & n15928 ) | ( n1462 & ~n18655 ) | ( n15928 & ~n18655 ) ;
  assign n18657 = n18656 ^ n14725 ^ n13266 ;
  assign n18658 = n18657 ^ n9685 ^ n3287 ;
  assign n18662 = ( n638 & n4644 ) | ( n638 & n8830 ) | ( n4644 & n8830 ) ;
  assign n18659 = n7665 ^ n5969 ^ n2498 ;
  assign n18660 = ~n3009 & n18659 ;
  assign n18661 = ( ~n8450 & n8733 ) | ( ~n8450 & n18660 ) | ( n8733 & n18660 ) ;
  assign n18663 = n18662 ^ n18661 ^ 1'b0 ;
  assign n18664 = n18663 ^ n4557 ^ n4136 ;
  assign n18673 = n12668 ^ n4598 ^ n3988 ;
  assign n18672 = ( n567 & n4250 ) | ( n567 & ~n4466 ) | ( n4250 & ~n4466 ) ;
  assign n18674 = n18673 ^ n18672 ^ n5202 ;
  assign n18665 = n10307 ^ n5296 ^ n2397 ;
  assign n18666 = n18665 ^ n12734 ^ n11499 ;
  assign n18668 = ( n863 & ~n3892 ) | ( n863 & n10886 ) | ( ~n3892 & n10886 ) ;
  assign n18667 = n10790 ^ n7669 ^ n6706 ;
  assign n18669 = n18668 ^ n18667 ^ n10790 ;
  assign n18670 = n15858 & ~n18669 ;
  assign n18671 = ~n18666 & n18670 ;
  assign n18675 = n18674 ^ n18671 ^ n5468 ;
  assign n18676 = n15610 ^ n2900 ^ n2451 ;
  assign n18677 = n16790 ^ n2680 ^ n1519 ;
  assign n18678 = n18677 ^ n6636 ^ 1'b0 ;
  assign n18679 = n18676 & ~n18678 ;
  assign n18680 = n18679 ^ n8762 ^ 1'b0 ;
  assign n18681 = ~n14590 & n18680 ;
  assign n18683 = ( n1882 & n3270 ) | ( n1882 & ~n5220 ) | ( n3270 & ~n5220 ) ;
  assign n18684 = n5241 ^ n3018 ^ 1'b0 ;
  assign n18685 = n18683 & n18684 ;
  assign n18686 = ( n5881 & n17394 ) | ( n5881 & n18685 ) | ( n17394 & n18685 ) ;
  assign n18682 = n17542 ^ n13058 ^ n10774 ;
  assign n18687 = n18686 ^ n18682 ^ n7109 ;
  assign n18688 = ( n3781 & ~n5454 ) | ( n3781 & n18394 ) | ( ~n5454 & n18394 ) ;
  assign n18689 = ( n3547 & ~n6658 ) | ( n3547 & n11147 ) | ( ~n6658 & n11147 ) ;
  assign n18690 = n18689 ^ n11460 ^ n1482 ;
  assign n18691 = ( n4801 & n7683 ) | ( n4801 & ~n18690 ) | ( n7683 & ~n18690 ) ;
  assign n18692 = n8624 ^ n4059 ^ 1'b0 ;
  assign n18693 = n7626 & n18692 ;
  assign n18694 = ( n13267 & n18691 ) | ( n13267 & ~n18693 ) | ( n18691 & ~n18693 ) ;
  assign n18695 = n18694 ^ n5193 ^ 1'b0 ;
  assign n18696 = n1175 & ~n18695 ;
  assign n18697 = ~n15069 & n18696 ;
  assign n18698 = n10331 ^ n4467 ^ 1'b0 ;
  assign n18699 = n12985 ^ n415 ^ 1'b0 ;
  assign n18700 = ( n15549 & n18698 ) | ( n15549 & n18699 ) | ( n18698 & n18699 ) ;
  assign n18702 = n13779 ^ n8529 ^ n7838 ;
  assign n18701 = ( ~n3484 & n7649 ) | ( ~n3484 & n9934 ) | ( n7649 & n9934 ) ;
  assign n18703 = n18702 ^ n18701 ^ n16195 ;
  assign n18704 = n8089 ^ n2791 ^ n1247 ;
  assign n18705 = n10080 ^ n3672 ^ n707 ;
  assign n18706 = n14819 ^ n14583 ^ n4216 ;
  assign n18707 = n18706 ^ n17045 ^ n11838 ;
  assign n18708 = n4843 & ~n16315 ;
  assign n18709 = n18708 ^ n420 ^ 1'b0 ;
  assign n18710 = n11620 ^ n10211 ^ n9015 ;
  assign n18717 = n4949 & n6919 ;
  assign n18718 = ( n4445 & n6917 ) | ( n4445 & ~n18717 ) | ( n6917 & ~n18717 ) ;
  assign n18719 = ( n805 & ~n8988 ) | ( n805 & n12027 ) | ( ~n8988 & n12027 ) ;
  assign n18720 = ( n3482 & n18718 ) | ( n3482 & n18719 ) | ( n18718 & n18719 ) ;
  assign n18721 = n3536 & ~n18720 ;
  assign n18722 = n18721 ^ n3194 ^ 1'b0 ;
  assign n18723 = ( n4996 & ~n13668 ) | ( n4996 & n18722 ) | ( ~n13668 & n18722 ) ;
  assign n18712 = n13686 ^ n2148 ^ n234 ;
  assign n18713 = ( n894 & n16671 ) | ( n894 & n18712 ) | ( n16671 & n18712 ) ;
  assign n18711 = n7969 ^ n1891 ^ n1697 ;
  assign n18714 = n18713 ^ n18711 ^ n12995 ;
  assign n18715 = n8161 | n18714 ;
  assign n18716 = n18715 ^ n1379 ^ 1'b0 ;
  assign n18724 = n18723 ^ n18716 ^ n8541 ;
  assign n18725 = n5905 ^ n5147 ^ 1'b0 ;
  assign n18726 = n18725 ^ n4469 ^ n1524 ;
  assign n18727 = ( n10150 & n10982 ) | ( n10150 & n18726 ) | ( n10982 & n18726 ) ;
  assign n18728 = n8096 ^ n3381 ^ n1801 ;
  assign n18729 = ( ~n9151 & n11299 ) | ( ~n9151 & n18728 ) | ( n11299 & n18728 ) ;
  assign n18730 = ( ~n8929 & n9950 ) | ( ~n8929 & n14397 ) | ( n9950 & n14397 ) ;
  assign n18731 = ( n1044 & n18056 ) | ( n1044 & ~n18730 ) | ( n18056 & ~n18730 ) ;
  assign n18732 = ( n6061 & n18729 ) | ( n6061 & n18731 ) | ( n18729 & n18731 ) ;
  assign n18733 = ( n3658 & n11293 ) | ( n3658 & n17826 ) | ( n11293 & n17826 ) ;
  assign n18735 = ( ~x38 & n4441 ) | ( ~x38 & n5512 ) | ( n4441 & n5512 ) ;
  assign n18736 = ( ~n1725 & n4811 ) | ( ~n1725 & n18735 ) | ( n4811 & n18735 ) ;
  assign n18737 = n17947 & ~n18736 ;
  assign n18734 = n7087 ^ n6812 ^ n1355 ;
  assign n18738 = n18737 ^ n18734 ^ n18130 ;
  assign n18739 = ( n904 & ~n3435 ) | ( n904 & n9901 ) | ( ~n3435 & n9901 ) ;
  assign n18740 = ( n2001 & n8373 ) | ( n2001 & n18739 ) | ( n8373 & n18739 ) ;
  assign n18741 = n11178 & ~n18740 ;
  assign n18742 = n18741 ^ n11830 ^ 1'b0 ;
  assign n18743 = n13002 ^ n9145 ^ n7372 ;
  assign n18745 = n8398 ^ n5552 ^ n950 ;
  assign n18744 = ( n6497 & n9161 ) | ( n6497 & n13059 ) | ( n9161 & n13059 ) ;
  assign n18746 = n18745 ^ n18744 ^ 1'b0 ;
  assign n18747 = ( ~n198 & n6029 ) | ( ~n198 & n6407 ) | ( n6029 & n6407 ) ;
  assign n18748 = n18747 ^ n9682 ^ n599 ;
  assign n18749 = ( n1291 & n9719 ) | ( n1291 & n17197 ) | ( n9719 & n17197 ) ;
  assign n18750 = n18749 ^ n14222 ^ n7074 ;
  assign n18751 = ( ~n17326 & n18748 ) | ( ~n17326 & n18750 ) | ( n18748 & n18750 ) ;
  assign n18753 = n13603 ^ n1134 ^ 1'b0 ;
  assign n18752 = n17518 ^ n17197 ^ n880 ;
  assign n18754 = n18753 ^ n18752 ^ 1'b0 ;
  assign n18755 = n6358 & ~n18754 ;
  assign n18756 = n1410 & ~n6952 ;
  assign n18757 = ~n8849 & n18756 ;
  assign n18758 = n18757 ^ n3438 ^ 1'b0 ;
  assign n18759 = ( n12994 & ~n14004 ) | ( n12994 & n18758 ) | ( ~n14004 & n18758 ) ;
  assign n18760 = n11142 ^ n5579 ^ n5050 ;
  assign n18761 = n5874 & n18760 ;
  assign n18762 = n18761 ^ n6125 ^ 1'b0 ;
  assign n18763 = n18762 ^ n1429 ^ 1'b0 ;
  assign n18764 = ~n4247 & n18763 ;
  assign n18765 = ( n2483 & ~n10713 ) | ( n2483 & n18764 ) | ( ~n10713 & n18764 ) ;
  assign n18766 = n16070 ^ n9895 ^ n3587 ;
  assign n18767 = ( ~x46 & n3461 ) | ( ~x46 & n18766 ) | ( n3461 & n18766 ) ;
  assign n18768 = n15191 ^ n8166 ^ n1212 ;
  assign n18769 = n18768 ^ n14344 ^ n11218 ;
  assign n18770 = n6216 ^ n1684 ^ 1'b0 ;
  assign n18771 = n9588 | n16264 ;
  assign n18772 = n10825 ^ n7153 ^ n2343 ;
  assign n18778 = ( n244 & ~n1762 ) | ( n244 & n8613 ) | ( ~n1762 & n8613 ) ;
  assign n18777 = ~n5947 & n11155 ;
  assign n18779 = n18778 ^ n18777 ^ 1'b0 ;
  assign n18773 = n7897 | n10612 ;
  assign n18774 = n15858 ^ n6201 ^ n4104 ;
  assign n18775 = ( n3047 & n8337 ) | ( n3047 & ~n18774 ) | ( n8337 & ~n18774 ) ;
  assign n18776 = ( n3646 & ~n18773 ) | ( n3646 & n18775 ) | ( ~n18773 & n18775 ) ;
  assign n18780 = n18779 ^ n18776 ^ n2743 ;
  assign n18781 = ( n3022 & n7208 ) | ( n3022 & ~n18165 ) | ( n7208 & ~n18165 ) ;
  assign n18782 = n18781 ^ n15188 ^ n475 ;
  assign n18783 = ~n17541 & n18782 ;
  assign n18784 = n2763 | n8946 ;
  assign n18785 = n15323 & ~n18784 ;
  assign n18786 = ( ~n5476 & n5748 ) | ( ~n5476 & n15325 ) | ( n5748 & n15325 ) ;
  assign n18787 = ( n5850 & n15703 ) | ( n5850 & n18786 ) | ( n15703 & n18786 ) ;
  assign n18788 = n8848 & ~n18787 ;
  assign n18794 = ( n2428 & n5183 ) | ( n2428 & ~n10413 ) | ( n5183 & ~n10413 ) ;
  assign n18790 = n7961 ^ n1853 ^ 1'b0 ;
  assign n18789 = n15092 ^ n10880 ^ n5091 ;
  assign n18791 = n18790 ^ n18789 ^ n13949 ;
  assign n18792 = ~n9062 & n18791 ;
  assign n18793 = n18792 ^ n5041 ^ 1'b0 ;
  assign n18795 = n18794 ^ n18793 ^ n15683 ;
  assign n18796 = n11364 ^ n7027 ^ n5892 ;
  assign n18797 = n18796 ^ n7162 ^ n4168 ;
  assign n18799 = ( ~n3570 & n7756 ) | ( ~n3570 & n11687 ) | ( n7756 & n11687 ) ;
  assign n18798 = n6358 & n14245 ;
  assign n18800 = n18799 ^ n18798 ^ 1'b0 ;
  assign n18801 = n11439 ^ n8163 ^ n1715 ;
  assign n18802 = n18801 ^ n2113 ^ 1'b0 ;
  assign n18803 = ( n16522 & n18287 ) | ( n16522 & n18802 ) | ( n18287 & n18802 ) ;
  assign n18804 = n13281 ^ n7208 ^ n1179 ;
  assign n18805 = x84 & n7797 ;
  assign n18806 = ~n9236 & n18805 ;
  assign n18807 = ( n2335 & n7474 ) | ( n2335 & n11873 ) | ( n7474 & n11873 ) ;
  assign n18808 = n5291 & n18807 ;
  assign n18809 = n18808 ^ n4101 ^ 1'b0 ;
  assign n18810 = n14398 ^ n12238 ^ n3434 ;
  assign n18811 = ( n3035 & n4317 ) | ( n3035 & ~n11511 ) | ( n4317 & ~n11511 ) ;
  assign n18812 = ( n5191 & n11234 ) | ( n5191 & n15658 ) | ( n11234 & n15658 ) ;
  assign n18813 = ( ~n1758 & n7767 ) | ( ~n1758 & n7773 ) | ( n7767 & n7773 ) ;
  assign n18814 = ( ~n9402 & n18812 ) | ( ~n9402 & n18813 ) | ( n18812 & n18813 ) ;
  assign n18815 = n17992 ^ n9327 ^ 1'b0 ;
  assign n18816 = n15613 ^ n12403 ^ n1488 ;
  assign n18817 = n18815 & n18816 ;
  assign n18818 = n9300 ^ n3556 ^ n1068 ;
  assign n18819 = ( ~n3150 & n15751 ) | ( ~n3150 & n18818 ) | ( n15751 & n18818 ) ;
  assign n18820 = ( ~n9737 & n16413 ) | ( ~n9737 & n18819 ) | ( n16413 & n18819 ) ;
  assign n18821 = n15336 ^ n10472 ^ 1'b0 ;
  assign n18822 = n9500 ^ n5987 ^ n946 ;
  assign n18823 = ( n5728 & n16056 ) | ( n5728 & ~n18822 ) | ( n16056 & ~n18822 ) ;
  assign n18824 = n18717 ^ n11146 ^ n640 ;
  assign n18825 = ( ~n641 & n7500 ) | ( ~n641 & n9847 ) | ( n7500 & n9847 ) ;
  assign n18826 = n18825 ^ n795 ^ n591 ;
  assign n18827 = ( ~n10775 & n18824 ) | ( ~n10775 & n18826 ) | ( n18824 & n18826 ) ;
  assign n18828 = n16580 ^ n12478 ^ n9701 ;
  assign n18829 = n5406 & n12702 ;
  assign n18830 = ~n5141 & n14293 ;
  assign n18831 = n4922 & n18830 ;
  assign n18832 = n18506 ^ n8080 ^ n5632 ;
  assign n18833 = n16863 ^ n13352 ^ n1030 ;
  assign n18834 = ( n2408 & n12859 ) | ( n2408 & n18378 ) | ( n12859 & n18378 ) ;
  assign n18835 = n4329 ^ n1727 ^ n777 ;
  assign n18836 = n18835 ^ n7563 ^ 1'b0 ;
  assign n18837 = n5884 & ~n18836 ;
  assign n18838 = ( n1917 & n2962 ) | ( n1917 & n3473 ) | ( n2962 & n3473 ) ;
  assign n18839 = n18838 ^ n15534 ^ 1'b0 ;
  assign n18840 = n18511 ^ n17701 ^ n9817 ;
  assign n18841 = n9659 ^ n8190 ^ 1'b0 ;
  assign n18842 = n6797 & ~n18841 ;
  assign n18843 = ( ~x86 & n9285 ) | ( ~x86 & n18842 ) | ( n9285 & n18842 ) ;
  assign n18844 = n6221 ^ n3548 ^ n1450 ;
  assign n18845 = n893 | n18844 ;
  assign n18846 = n8002 | n18845 ;
  assign n18847 = ( ~n2076 & n4776 ) | ( ~n2076 & n9222 ) | ( n4776 & n9222 ) ;
  assign n18848 = n8985 & ~n17470 ;
  assign n18849 = ( n687 & n1552 ) | ( n687 & n13730 ) | ( n1552 & n13730 ) ;
  assign n18850 = n8198 ^ n6531 ^ n3033 ;
  assign n18851 = n18850 ^ n11327 ^ n4793 ;
  assign n18852 = ( n6007 & ~n6146 ) | ( n6007 & n6333 ) | ( ~n6146 & n6333 ) ;
  assign n18853 = n18852 ^ n6931 ^ n4444 ;
  assign n18854 = ( n2357 & ~n4624 ) | ( n2357 & n15842 ) | ( ~n4624 & n15842 ) ;
  assign n18855 = n12085 ^ n7746 ^ n2924 ;
  assign n18856 = ( ~n9168 & n18854 ) | ( ~n9168 & n18855 ) | ( n18854 & n18855 ) ;
  assign n18857 = n17796 ^ n4062 ^ n2774 ;
  assign n18858 = n18857 ^ n11192 ^ n4122 ;
  assign n18859 = ( n4559 & ~n4711 ) | ( n4559 & n11979 ) | ( ~n4711 & n11979 ) ;
  assign n18860 = n18859 ^ n13642 ^ n9582 ;
  assign n18861 = ( n854 & ~n5548 ) | ( n854 & n18860 ) | ( ~n5548 & n18860 ) ;
  assign n18862 = n10442 ^ n2420 ^ 1'b0 ;
  assign n18863 = x68 & n11476 ;
  assign n18864 = n1059 & n18863 ;
  assign n18865 = n15057 ^ n12467 ^ n10712 ;
  assign n18866 = n563 | n9502 ;
  assign n18867 = n6476 ^ n330 ^ 1'b0 ;
  assign n18868 = n18749 ^ n8568 ^ n5507 ;
  assign n18869 = ( n9174 & ~n18867 ) | ( n9174 & n18868 ) | ( ~n18867 & n18868 ) ;
  assign n18870 = n16002 ^ n1896 ^ n918 ;
  assign n18871 = ( n11583 & ~n13741 ) | ( n11583 & n18870 ) | ( ~n13741 & n18870 ) ;
  assign n18872 = n18871 ^ n13460 ^ n3197 ;
  assign n18873 = n1712 & ~n1846 ;
  assign n18874 = ( n2374 & ~n11060 ) | ( n2374 & n18873 ) | ( ~n11060 & n18873 ) ;
  assign n18875 = n1682 & n18874 ;
  assign n18876 = ( n500 & n508 ) | ( n500 & n5304 ) | ( n508 & n5304 ) ;
  assign n18877 = n18825 & n18876 ;
  assign n18878 = n18877 ^ n5496 ^ n870 ;
  assign n18879 = n18878 ^ n18219 ^ x62 ;
  assign n18882 = n10465 ^ n4483 ^ 1'b0 ;
  assign n18880 = n15718 ^ n1701 ^ 1'b0 ;
  assign n18881 = n2158 & ~n18880 ;
  assign n18883 = n18882 ^ n18881 ^ n5758 ;
  assign n18884 = n1889 & ~n6829 ;
  assign n18885 = n18884 ^ n4537 ^ 1'b0 ;
  assign n18886 = ( n2432 & n3141 ) | ( n2432 & n18885 ) | ( n3141 & n18885 ) ;
  assign n18887 = ( n5358 & n6928 ) | ( n5358 & n18886 ) | ( n6928 & n18886 ) ;
  assign n18888 = ( n13458 & n18883 ) | ( n13458 & ~n18887 ) | ( n18883 & ~n18887 ) ;
  assign n18889 = n5834 ^ n2378 ^ n1286 ;
  assign n18890 = n5981 & n18889 ;
  assign n18891 = ~n16825 & n18890 ;
  assign n18892 = n18891 ^ n18407 ^ n14626 ;
  assign n18893 = n17292 ^ n15374 ^ n14205 ;
  assign n18894 = ( n2106 & n6757 ) | ( n2106 & n8240 ) | ( n6757 & n8240 ) ;
  assign n18895 = n18894 ^ n17809 ^ n5951 ;
  assign n18896 = n18895 ^ n1035 ^ 1'b0 ;
  assign n18897 = n16031 ^ n10222 ^ 1'b0 ;
  assign n18898 = n18897 ^ n6558 ^ n3825 ;
  assign n18899 = ( n3075 & ~n7898 ) | ( n3075 & n18898 ) | ( ~n7898 & n18898 ) ;
  assign n18900 = n11019 | n13025 ;
  assign n18901 = n1844 & ~n18900 ;
  assign n18902 = n16572 | n18901 ;
  assign n18903 = n6587 & ~n18902 ;
  assign n18904 = ( n680 & n3969 ) | ( n680 & n12924 ) | ( n3969 & n12924 ) ;
  assign n18905 = n18904 ^ n13341 ^ n4578 ;
  assign n18906 = n8093 ^ n6619 ^ n3457 ;
  assign n18907 = n18906 ^ n5318 ^ n278 ;
  assign n18908 = ( n9209 & n16430 ) | ( n9209 & n18907 ) | ( n16430 & n18907 ) ;
  assign n18913 = n4660 ^ n4122 ^ n811 ;
  assign n18914 = ( n8921 & n8929 ) | ( n8921 & ~n18913 ) | ( n8929 & ~n18913 ) ;
  assign n18911 = ~n2129 & n8951 ;
  assign n18909 = n1540 & n3056 ;
  assign n18910 = n18909 ^ n12312 ^ 1'b0 ;
  assign n18912 = n18911 ^ n18910 ^ n1067 ;
  assign n18915 = n18914 ^ n18912 ^ n18020 ;
  assign n18916 = n18349 ^ n4376 ^ 1'b0 ;
  assign n18917 = n18916 ^ n6064 ^ n2178 ;
  assign n18918 = ( n2674 & n2850 ) | ( n2674 & n3172 ) | ( n2850 & n3172 ) ;
  assign n18919 = n16298 & ~n18918 ;
  assign n18920 = ~n18917 & n18919 ;
  assign n18925 = ( n3624 & ~n4216 ) | ( n3624 & n12211 ) | ( ~n4216 & n12211 ) ;
  assign n18924 = n14964 ^ n5222 ^ n683 ;
  assign n18926 = n18925 ^ n18924 ^ n10174 ;
  assign n18922 = n5284 ^ n1863 ^ n1017 ;
  assign n18923 = n18922 ^ n3097 ^ n367 ;
  assign n18927 = n18926 ^ n18923 ^ n13104 ;
  assign n18921 = ( n3188 & ~n11691 ) | ( n3188 & n12789 ) | ( ~n11691 & n12789 ) ;
  assign n18928 = n18927 ^ n18921 ^ n3789 ;
  assign n18929 = n18928 ^ n15875 ^ 1'b0 ;
  assign n18930 = n11507 ^ n10357 ^ n3357 ;
  assign n18931 = ( n967 & n5058 ) | ( n967 & n11249 ) | ( n5058 & n11249 ) ;
  assign n18932 = n18931 ^ n16304 ^ n12375 ;
  assign n18933 = ( ~n2298 & n4839 ) | ( ~n2298 & n4939 ) | ( n4839 & n4939 ) ;
  assign n18934 = ( n7558 & n11769 ) | ( n7558 & n18933 ) | ( n11769 & n18933 ) ;
  assign n18935 = ( n1846 & ~n3148 ) | ( n1846 & n3261 ) | ( ~n3148 & n3261 ) ;
  assign n18936 = ( n7539 & n16796 ) | ( n7539 & ~n18935 ) | ( n16796 & ~n18935 ) ;
  assign n18937 = ( ~n1424 & n17597 ) | ( ~n1424 & n18936 ) | ( n17597 & n18936 ) ;
  assign n18938 = n18571 ^ n4195 ^ n1509 ;
  assign n18939 = n4340 & ~n18938 ;
  assign n18940 = ~n18937 & n18939 ;
  assign n18941 = ( ~n12279 & n18934 ) | ( ~n12279 & n18940 ) | ( n18934 & n18940 ) ;
  assign n18942 = ( n6792 & n7994 ) | ( n6792 & ~n18066 ) | ( n7994 & ~n18066 ) ;
  assign n18943 = n18942 ^ n17287 ^ 1'b0 ;
  assign n18944 = ~n1768 & n18943 ;
  assign n18945 = n15266 ^ n13777 ^ n12287 ;
  assign n18946 = n18642 ^ n4230 ^ n1473 ;
  assign n18947 = ~n1957 & n6430 ;
  assign n18948 = n14660 ^ n9938 ^ n8415 ;
  assign n18949 = n10676 | n13796 ;
  assign n18950 = ( n18947 & ~n18948 ) | ( n18947 & n18949 ) | ( ~n18948 & n18949 ) ;
  assign n18951 = n12166 ^ n11290 ^ 1'b0 ;
  assign n18952 = ( n2389 & n5378 ) | ( n2389 & n18951 ) | ( n5378 & n18951 ) ;
  assign n18953 = n11170 ^ n6957 ^ n1645 ;
  assign n18954 = n18953 ^ n18382 ^ n4304 ;
  assign n18955 = ( n6362 & n10823 ) | ( n6362 & n18954 ) | ( n10823 & n18954 ) ;
  assign n18956 = n4040 & ~n17751 ;
  assign n18957 = ( n412 & n8774 ) | ( n412 & n9785 ) | ( n8774 & n9785 ) ;
  assign n18958 = n3757 & ~n9674 ;
  assign n18959 = n6343 & ~n18958 ;
  assign n18960 = ( n10734 & ~n12479 ) | ( n10734 & n18959 ) | ( ~n12479 & n18959 ) ;
  assign n18961 = n9612 & n18960 ;
  assign n18962 = n18957 & n18961 ;
  assign n18963 = ( n2455 & ~n4515 ) | ( n2455 & n5680 ) | ( ~n4515 & n5680 ) ;
  assign n18964 = n18963 ^ n11749 ^ n8626 ;
  assign n18965 = ( n4496 & ~n11809 ) | ( n4496 & n18964 ) | ( ~n11809 & n18964 ) ;
  assign n18966 = ~n2439 & n8439 ;
  assign n18967 = ~n10280 & n18966 ;
  assign n18968 = n8642 ^ n6227 ^ n3525 ;
  assign n18969 = ( ~n16105 & n18967 ) | ( ~n16105 & n18968 ) | ( n18967 & n18968 ) ;
  assign n18970 = n5787 ^ n4871 ^ n1060 ;
  assign n18971 = n7985 | n13074 ;
  assign n18972 = ( ~n10257 & n18970 ) | ( ~n10257 & n18971 ) | ( n18970 & n18971 ) ;
  assign n18973 = ( ~n1020 & n17154 ) | ( ~n1020 & n18972 ) | ( n17154 & n18972 ) ;
  assign n18974 = n18973 ^ n151 ^ 1'b0 ;
  assign n18977 = ( n5191 & n9444 ) | ( n5191 & n10562 ) | ( n9444 & n10562 ) ;
  assign n18975 = n17556 ^ n14870 ^ n4241 ;
  assign n18976 = n18975 ^ n13733 ^ n4668 ;
  assign n18978 = n18977 ^ n18976 ^ n2321 ;
  assign n18979 = n10961 ^ n4712 ^ n4094 ;
  assign n18980 = n18979 ^ n15581 ^ 1'b0 ;
  assign n18981 = ~n694 & n18980 ;
  assign n18982 = n18981 ^ n17074 ^ n15700 ;
  assign n18983 = n2732 & ~n4360 ;
  assign n18984 = n18983 ^ n571 ^ 1'b0 ;
  assign n18985 = ( ~n7651 & n10333 ) | ( ~n7651 & n18984 ) | ( n10333 & n18984 ) ;
  assign n18986 = ( n10912 & n16945 ) | ( n10912 & n18985 ) | ( n16945 & n18985 ) ;
  assign n18987 = n18982 | n18986 ;
  assign n18988 = ( n8294 & ~n17065 ) | ( n8294 & n17529 ) | ( ~n17065 & n17529 ) ;
  assign n18989 = n5838 | n7627 ;
  assign n18990 = n18989 ^ n14426 ^ n6531 ;
  assign n18991 = ( ~n5905 & n13551 ) | ( ~n5905 & n18990 ) | ( n13551 & n18990 ) ;
  assign n18992 = n6657 & ~n17885 ;
  assign n18993 = n10239 ^ n7746 ^ n824 ;
  assign n18994 = ( ~n4640 & n5880 ) | ( ~n4640 & n7040 ) | ( n5880 & n7040 ) ;
  assign n18995 = n18994 ^ n14443 ^ n10930 ;
  assign n18996 = ( n6913 & ~n9413 ) | ( n6913 & n11624 ) | ( ~n9413 & n11624 ) ;
  assign n18997 = ( n470 & ~n8642 ) | ( n470 & n18996 ) | ( ~n8642 & n18996 ) ;
  assign n18998 = n13585 ^ n13006 ^ n2963 ;
  assign n18999 = n6302 ^ n4673 ^ n2624 ;
  assign n19000 = n18999 ^ n5407 ^ n5349 ;
  assign n19001 = n19000 ^ n9228 ^ n3794 ;
  assign n19002 = ( n5619 & n10871 ) | ( n5619 & n17676 ) | ( n10871 & n17676 ) ;
  assign n19003 = ( n3066 & n16352 ) | ( n3066 & ~n19002 ) | ( n16352 & ~n19002 ) ;
  assign n19004 = ( n2871 & ~n6633 ) | ( n2871 & n15637 ) | ( ~n6633 & n15637 ) ;
  assign n19005 = n19004 ^ n8405 ^ n1017 ;
  assign n19006 = n13106 & ~n19005 ;
  assign n19007 = ( n358 & n8873 ) | ( n358 & ~n15279 ) | ( n8873 & ~n15279 ) ;
  assign n19008 = ( n5998 & n17540 ) | ( n5998 & ~n19007 ) | ( n17540 & ~n19007 ) ;
  assign n19009 = ( n2322 & n2712 ) | ( n2322 & n15555 ) | ( n2712 & n15555 ) ;
  assign n19010 = n19009 ^ n9001 ^ n1039 ;
  assign n19011 = ( n2575 & n3617 ) | ( n2575 & ~n11800 ) | ( n3617 & ~n11800 ) ;
  assign n19012 = ( ~n1443 & n1887 ) | ( ~n1443 & n7787 ) | ( n1887 & n7787 ) ;
  assign n19013 = n19012 ^ n14222 ^ n11286 ;
  assign n19014 = n13389 ^ n10187 ^ n7622 ;
  assign n19015 = ( n16903 & n19013 ) | ( n16903 & n19014 ) | ( n19013 & n19014 ) ;
  assign n19016 = ( ~n303 & n3770 ) | ( ~n303 & n4102 ) | ( n3770 & n4102 ) ;
  assign n19017 = n19016 ^ n16596 ^ n13590 ;
  assign n19018 = n19017 ^ n14293 ^ n5623 ;
  assign n19021 = n11462 ^ n4998 ^ n4680 ;
  assign n19020 = ( n2946 & n3907 ) | ( n2946 & n5433 ) | ( n3907 & n5433 ) ;
  assign n19019 = n16917 ^ n12419 ^ n1593 ;
  assign n19022 = n19021 ^ n19020 ^ n19019 ;
  assign n19023 = n5831 ^ n4191 ^ n3094 ;
  assign n19025 = n2059 | n7472 ;
  assign n19026 = n3961 | n19025 ;
  assign n19024 = n17311 ^ n5497 ^ 1'b0 ;
  assign n19027 = n19026 ^ n19024 ^ n15700 ;
  assign n19028 = n19027 ^ n16042 ^ n3095 ;
  assign n19029 = ( n1896 & n5236 ) | ( n1896 & n9749 ) | ( n5236 & n9749 ) ;
  assign n19030 = ( n3714 & n5588 ) | ( n3714 & ~n15982 ) | ( n5588 & ~n15982 ) ;
  assign n19031 = n17450 ^ n10103 ^ 1'b0 ;
  assign n19032 = n16440 ^ n7710 ^ n3040 ;
  assign n19033 = ( n668 & ~n2527 ) | ( n668 & n19032 ) | ( ~n2527 & n19032 ) ;
  assign n19034 = n19033 ^ n168 ^ 1'b0 ;
  assign n19035 = ( n3931 & n16212 ) | ( n3931 & n19034 ) | ( n16212 & n19034 ) ;
  assign n19038 = n6445 | n12872 ;
  assign n19036 = n6496 ^ n5450 ^ n3601 ;
  assign n19037 = ( n6789 & ~n6948 ) | ( n6789 & n19036 ) | ( ~n6948 & n19036 ) ;
  assign n19039 = n19038 ^ n19037 ^ 1'b0 ;
  assign n19040 = n18436 ^ n14449 ^ n5442 ;
  assign n19041 = n1729 & ~n9429 ;
  assign n19042 = n19040 & n19041 ;
  assign n19043 = n8463 ^ n2831 ^ n540 ;
  assign n19044 = ( ~n4009 & n10426 ) | ( ~n4009 & n19043 ) | ( n10426 & n19043 ) ;
  assign n19045 = n14579 ^ n2518 ^ 1'b0 ;
  assign n19046 = n6366 ^ n2699 ^ 1'b0 ;
  assign n19047 = n8539 ^ n4511 ^ 1'b0 ;
  assign n19048 = ( n4423 & n12639 ) | ( n4423 & n19047 ) | ( n12639 & n19047 ) ;
  assign n19049 = n10442 ^ n1494 ^ n1421 ;
  assign n19050 = ~n5134 & n15776 ;
  assign n19051 = n906 & n6210 ;
  assign n19053 = ( n601 & ~n2541 ) | ( n601 & n2851 ) | ( ~n2541 & n2851 ) ;
  assign n19052 = n10063 ^ n1022 ^ n377 ;
  assign n19054 = n19053 ^ n19052 ^ n12578 ;
  assign n19055 = n2521 & n6417 ;
  assign n19056 = n19055 ^ n1532 ^ 1'b0 ;
  assign n19057 = ( n4895 & n15240 ) | ( n4895 & n18203 ) | ( n15240 & n18203 ) ;
  assign n19058 = ( n5677 & ~n19056 ) | ( n5677 & n19057 ) | ( ~n19056 & n19057 ) ;
  assign n19059 = n3220 & n8688 ;
  assign n19060 = ( n3043 & ~n17360 ) | ( n3043 & n19059 ) | ( ~n17360 & n19059 ) ;
  assign n19061 = ( n15185 & n19058 ) | ( n15185 & n19060 ) | ( n19058 & n19060 ) ;
  assign n19062 = ( n859 & n1475 ) | ( n859 & n5454 ) | ( n1475 & n5454 ) ;
  assign n19063 = ( n1742 & n14490 ) | ( n1742 & ~n19062 ) | ( n14490 & ~n19062 ) ;
  assign n19064 = n16738 ^ n13810 ^ n4860 ;
  assign n19065 = n19063 & n19064 ;
  assign n19066 = ( n6465 & n7035 ) | ( n6465 & ~n12166 ) | ( n7035 & ~n12166 ) ;
  assign n19067 = ( n6853 & n15343 ) | ( n6853 & ~n16726 ) | ( n15343 & ~n16726 ) ;
  assign n19068 = n4991 & ~n18321 ;
  assign n19069 = n19068 ^ n7854 ^ 1'b0 ;
  assign n19070 = n18690 ^ n11691 ^ 1'b0 ;
  assign n19071 = ~n18852 & n19070 ;
  assign n19072 = ( ~n1522 & n15097 ) | ( ~n1522 & n19071 ) | ( n15097 & n19071 ) ;
  assign n19076 = n5222 & ~n11959 ;
  assign n19077 = ~n1134 & n19076 ;
  assign n19073 = n18427 ^ n14407 ^ n1403 ;
  assign n19074 = n19073 ^ n3543 ^ 1'b0 ;
  assign n19075 = n19074 ^ n15496 ^ n623 ;
  assign n19078 = n19077 ^ n19075 ^ n12897 ;
  assign n19079 = ( ~n2795 & n6486 ) | ( ~n2795 & n8807 ) | ( n6486 & n8807 ) ;
  assign n19080 = n12015 ^ n9092 ^ n5058 ;
  assign n19081 = ( n7094 & n19057 ) | ( n7094 & ~n19080 ) | ( n19057 & ~n19080 ) ;
  assign n19082 = n17845 & ~n18380 ;
  assign n19083 = n973 & ~n19082 ;
  assign n19084 = n19083 ^ n17991 ^ n10112 ;
  assign n19086 = ( n2693 & ~n8297 ) | ( n2693 & n9097 ) | ( ~n8297 & n9097 ) ;
  assign n19085 = n11017 ^ n6962 ^ n4099 ;
  assign n19087 = n19086 ^ n19085 ^ n6614 ;
  assign n19088 = n7602 & n19087 ;
  assign n19095 = ( n1790 & ~n2798 ) | ( n1790 & n5454 ) | ( ~n2798 & n5454 ) ;
  assign n19096 = n19095 ^ n11459 ^ n10716 ;
  assign n19089 = n16653 ^ n13134 ^ n1238 ;
  assign n19090 = n19089 ^ n11177 ^ n961 ;
  assign n19091 = n14993 | n19090 ;
  assign n19092 = n19091 ^ n10910 ^ 1'b0 ;
  assign n19093 = n19092 ^ n15251 ^ n1694 ;
  assign n19094 = n19093 ^ n8639 ^ n2553 ;
  assign n19097 = n19096 ^ n19094 ^ 1'b0 ;
  assign n19098 = n16084 ^ n1781 ^ n655 ;
  assign n19099 = ( ~n922 & n9190 ) | ( ~n922 & n15363 ) | ( n9190 & n15363 ) ;
  assign n19100 = n13256 ^ n12884 ^ 1'b0 ;
  assign n19101 = ( n3707 & ~n11195 ) | ( n3707 & n14318 ) | ( ~n11195 & n14318 ) ;
  assign n19102 = ( n1357 & n1888 ) | ( n1357 & n2671 ) | ( n1888 & n2671 ) ;
  assign n19103 = n19102 ^ n11012 ^ n1198 ;
  assign n19104 = n6016 ^ n4386 ^ n3287 ;
  assign n19105 = ( n10132 & ~n19103 ) | ( n10132 & n19104 ) | ( ~n19103 & n19104 ) ;
  assign n19106 = ( n4283 & ~n10059 ) | ( n4283 & n17973 ) | ( ~n10059 & n17973 ) ;
  assign n19107 = ( n1819 & n19105 ) | ( n1819 & ~n19106 ) | ( n19105 & ~n19106 ) ;
  assign n19108 = n12368 ^ n10485 ^ n4590 ;
  assign n19109 = n11249 ^ n8472 ^ n3435 ;
  assign n19110 = n19109 ^ n16504 ^ n5479 ;
  assign n19111 = n19110 ^ n18825 ^ n7266 ;
  assign n19112 = ( n8272 & ~n13073 ) | ( n8272 & n19111 ) | ( ~n13073 & n19111 ) ;
  assign n19113 = n5363 ^ n4022 ^ n2536 ;
  assign n19114 = ( n797 & n7461 ) | ( n797 & ~n19113 ) | ( n7461 & ~n19113 ) ;
  assign n19115 = ~n486 & n2103 ;
  assign n19116 = ( n3677 & n4437 ) | ( n3677 & n19115 ) | ( n4437 & n19115 ) ;
  assign n19117 = ( n4704 & n10012 ) | ( n4704 & n11768 ) | ( n10012 & n11768 ) ;
  assign n19118 = n4561 | n19117 ;
  assign n19119 = n9508 | n19118 ;
  assign n19120 = n11954 ^ n5550 ^ 1'b0 ;
  assign n19121 = n19119 & n19120 ;
  assign n19122 = ( n19114 & n19116 ) | ( n19114 & n19121 ) | ( n19116 & n19121 ) ;
  assign n19123 = ( n865 & n3132 ) | ( n865 & ~n7313 ) | ( n3132 & ~n7313 ) ;
  assign n19124 = n5270 & ~n19123 ;
  assign n19125 = n19124 ^ n12533 ^ n3207 ;
  assign n19126 = n7818 ^ n7470 ^ n5803 ;
  assign n19127 = n19126 ^ n13631 ^ n7043 ;
  assign n19128 = n19127 ^ n18260 ^ n15144 ;
  assign n19129 = ( n3794 & n7183 ) | ( n3794 & n9679 ) | ( n7183 & n9679 ) ;
  assign n19130 = n12093 & n18612 ;
  assign n19131 = n10187 & ~n10563 ;
  assign n19132 = ~n13552 & n19131 ;
  assign n19133 = ( n648 & n1242 ) | ( n648 & n9613 ) | ( n1242 & n9613 ) ;
  assign n19134 = n19133 ^ n8201 ^ n1506 ;
  assign n19135 = n16967 ^ n14653 ^ n7722 ;
  assign n19136 = n19135 ^ n17005 ^ n7909 ;
  assign n19143 = ( n2903 & n8355 ) | ( n2903 & n14045 ) | ( n8355 & n14045 ) ;
  assign n19144 = n4812 & n19143 ;
  assign n19137 = ( n2159 & ~n2431 ) | ( n2159 & n3878 ) | ( ~n2431 & n3878 ) ;
  assign n19138 = ( n1511 & n7744 ) | ( n1511 & n11347 ) | ( n7744 & n11347 ) ;
  assign n19139 = ( n3945 & ~n7202 ) | ( n3945 & n19138 ) | ( ~n7202 & n19138 ) ;
  assign n19140 = ( n10261 & n10943 ) | ( n10261 & n19139 ) | ( n10943 & n19139 ) ;
  assign n19141 = ( n6591 & n7079 ) | ( n6591 & n19140 ) | ( n7079 & n19140 ) ;
  assign n19142 = ( n7174 & n19137 ) | ( n7174 & ~n19141 ) | ( n19137 & ~n19141 ) ;
  assign n19145 = n19144 ^ n19142 ^ n8034 ;
  assign n19146 = n16363 ^ n14439 ^ n8038 ;
  assign n19147 = n15192 ^ n11438 ^ n10792 ;
  assign n19148 = ( n282 & ~n3145 ) | ( n282 & n9079 ) | ( ~n3145 & n9079 ) ;
  assign n19150 = n6039 ^ n4861 ^ n4612 ;
  assign n19149 = n1634 & ~n9464 ;
  assign n19151 = n19150 ^ n19149 ^ n9340 ;
  assign n19152 = ( ~n5697 & n7419 ) | ( ~n5697 & n11139 ) | ( n7419 & n11139 ) ;
  assign n19153 = n10955 & n19152 ;
  assign n19154 = n19153 ^ n8671 ^ 1'b0 ;
  assign n19155 = n19154 ^ n6504 ^ n2457 ;
  assign n19156 = n13184 ^ n12136 ^ n2821 ;
  assign n19157 = ( ~n11513 & n19155 ) | ( ~n11513 & n19156 ) | ( n19155 & n19156 ) ;
  assign n19164 = n2791 ^ n2659 ^ n671 ;
  assign n19165 = n19164 ^ n7100 ^ n2735 ;
  assign n19161 = ( ~n977 & n1556 ) | ( ~n977 & n2642 ) | ( n1556 & n2642 ) ;
  assign n19162 = n19161 ^ n8010 ^ n3883 ;
  assign n19160 = ~n12348 & n16015 ;
  assign n19163 = n19162 ^ n19160 ^ n7757 ;
  assign n19166 = n19165 ^ n19163 ^ n2977 ;
  assign n19158 = n10484 ^ n920 ^ x93 ;
  assign n19159 = ( n2480 & n10568 ) | ( n2480 & ~n19158 ) | ( n10568 & ~n19158 ) ;
  assign n19167 = n19166 ^ n19159 ^ n12425 ;
  assign n19168 = n3928 | n5559 ;
  assign n19169 = n19168 ^ n12872 ^ n6484 ;
  assign n19170 = n7648 ^ n6473 ^ n6089 ;
  assign n19171 = n19170 ^ n1741 ^ 1'b0 ;
  assign n19172 = n19169 & n19171 ;
  assign n19173 = ( n9005 & ~n12077 ) | ( n9005 & n16385 ) | ( ~n12077 & n16385 ) ;
  assign n19178 = ( n6429 & ~n7141 ) | ( n6429 & n7813 ) | ( ~n7141 & n7813 ) ;
  assign n19174 = n17223 ^ n15115 ^ n882 ;
  assign n19175 = ( n5482 & n12416 ) | ( n5482 & ~n14682 ) | ( n12416 & ~n14682 ) ;
  assign n19176 = n19175 ^ n17339 ^ n4594 ;
  assign n19177 = ( n12525 & ~n19174 ) | ( n12525 & n19176 ) | ( ~n19174 & n19176 ) ;
  assign n19179 = n19178 ^ n19177 ^ n12565 ;
  assign n19180 = n14600 ^ n6120 ^ n4395 ;
  assign n19181 = ( n3897 & n12594 ) | ( n3897 & n19180 ) | ( n12594 & n19180 ) ;
  assign n19187 = n6493 ^ n926 ^ 1'b0 ;
  assign n19182 = n2013 & ~n7738 ;
  assign n19183 = n19182 ^ n2305 ^ 1'b0 ;
  assign n19184 = n19183 ^ n8251 ^ n2209 ;
  assign n19185 = n6386 | n19184 ;
  assign n19186 = ( n2606 & n16054 ) | ( n2606 & n19185 ) | ( n16054 & n19185 ) ;
  assign n19188 = n19187 ^ n19186 ^ n12855 ;
  assign n19189 = n1033 ^ n360 ^ x112 ;
  assign n19190 = n19189 ^ n15880 ^ n2431 ;
  assign n19191 = ( n12225 & ~n12868 ) | ( n12225 & n15422 ) | ( ~n12868 & n15422 ) ;
  assign n19192 = ( n5143 & ~n12057 ) | ( n5143 & n12100 ) | ( ~n12057 & n12100 ) ;
  assign n19193 = n8380 & ~n8932 ;
  assign n19194 = ~n6568 & n19193 ;
  assign n19196 = ( n4429 & ~n5235 ) | ( n4429 & n7679 ) | ( ~n5235 & n7679 ) ;
  assign n19197 = ( n221 & n9842 ) | ( n221 & n19196 ) | ( n9842 & n19196 ) ;
  assign n19198 = ( n871 & n3056 ) | ( n871 & ~n19197 ) | ( n3056 & ~n19197 ) ;
  assign n19195 = n6880 & n10982 ;
  assign n19199 = n19198 ^ n19195 ^ n8005 ;
  assign n19200 = n7257 | n19199 ;
  assign n19201 = ( n2085 & n2159 ) | ( n2085 & ~n10393 ) | ( n2159 & ~n10393 ) ;
  assign n19202 = ( n14725 & ~n16557 ) | ( n14725 & n19201 ) | ( ~n16557 & n19201 ) ;
  assign n19203 = ( ~n6952 & n8953 ) | ( ~n6952 & n19202 ) | ( n8953 & n19202 ) ;
  assign n19204 = n13266 ^ n5066 ^ n1429 ;
  assign n19205 = n19204 ^ n11060 ^ n1842 ;
  assign n19206 = n12660 ^ n7429 ^ n5433 ;
  assign n19207 = n19206 ^ n15622 ^ n11842 ;
  assign n19208 = n16360 ^ n6602 ^ n4419 ;
  assign n19209 = ( n854 & n2960 ) | ( n854 & ~n19208 ) | ( n2960 & ~n19208 ) ;
  assign n19210 = ~n1901 & n2404 ;
  assign n19211 = n19210 ^ n1114 ^ 1'b0 ;
  assign n19212 = n11556 ^ n8003 ^ 1'b0 ;
  assign n19213 = ( ~n1785 & n5638 ) | ( ~n1785 & n19212 ) | ( n5638 & n19212 ) ;
  assign n19214 = n19213 ^ n16535 ^ n11060 ;
  assign n19215 = n17237 ^ n16260 ^ n3715 ;
  assign n19216 = ( n1197 & n14017 ) | ( n1197 & ~n19215 ) | ( n14017 & ~n19215 ) ;
  assign n19217 = n19216 ^ n14581 ^ n4572 ;
  assign n19218 = ( n7481 & n16658 ) | ( n7481 & n19217 ) | ( n16658 & n19217 ) ;
  assign n19220 = n2632 | n5270 ;
  assign n19221 = n1849 | n19220 ;
  assign n19219 = n10951 ^ n10302 ^ n2493 ;
  assign n19222 = n19221 ^ n19219 ^ n4419 ;
  assign n19223 = ~n2592 & n15224 ;
  assign n19224 = ( n154 & n4191 ) | ( n154 & n4482 ) | ( n4191 & n4482 ) ;
  assign n19225 = ( n9628 & n19223 ) | ( n9628 & ~n19224 ) | ( n19223 & ~n19224 ) ;
  assign n19226 = n19225 ^ n12043 ^ n4183 ;
  assign n19227 = ( n2712 & n11673 ) | ( n2712 & n19226 ) | ( n11673 & n19226 ) ;
  assign n19228 = n13906 ^ n11166 ^ n1963 ;
  assign n19229 = n19228 ^ n18357 ^ 1'b0 ;
  assign n19233 = n11362 ^ n6476 ^ n3669 ;
  assign n19230 = n8719 ^ n3479 ^ 1'b0 ;
  assign n19231 = ~n16939 & n19230 ;
  assign n19232 = n19231 ^ n16478 ^ n8435 ;
  assign n19234 = n19233 ^ n19232 ^ n9237 ;
  assign n19236 = ( n742 & n9182 ) | ( n742 & n11284 ) | ( n9182 & n11284 ) ;
  assign n19237 = ( n8528 & n14727 ) | ( n8528 & n19236 ) | ( n14727 & n19236 ) ;
  assign n19235 = n6548 ^ n5548 ^ 1'b0 ;
  assign n19238 = n19237 ^ n19235 ^ n164 ;
  assign n19239 = ( n8943 & ~n13745 ) | ( n8943 & n17795 ) | ( ~n13745 & n17795 ) ;
  assign n19240 = n19239 ^ n10674 ^ n8196 ;
  assign n19241 = n10168 ^ n10077 ^ n474 ;
  assign n19242 = n19241 ^ n6201 ^ n2348 ;
  assign n19243 = n9229 ^ n4958 ^ n3519 ;
  assign n19247 = ( n5822 & ~n8850 ) | ( n5822 & n9437 ) | ( ~n8850 & n9437 ) ;
  assign n19244 = n7576 ^ n2514 ^ 1'b0 ;
  assign n19245 = ( n2876 & n6770 ) | ( n2876 & n19244 ) | ( n6770 & n19244 ) ;
  assign n19246 = n19245 ^ n11466 ^ 1'b0 ;
  assign n19248 = n19247 ^ n19246 ^ n4772 ;
  assign n19251 = ( n8194 & n13074 ) | ( n8194 & ~n13130 ) | ( n13074 & ~n13130 ) ;
  assign n19249 = n18611 ^ n16432 ^ n10239 ;
  assign n19250 = ~n13679 & n19249 ;
  assign n19252 = n19251 ^ n19250 ^ n18157 ;
  assign n19253 = n11061 ^ n9808 ^ n2511 ;
  assign n19254 = n19253 ^ n17181 ^ n9687 ;
  assign n19255 = n15892 ^ n508 ^ 1'b0 ;
  assign n19256 = n5228 ^ n5209 ^ n924 ;
  assign n19257 = n17507 ^ n12969 ^ n10307 ;
  assign n19258 = n19257 ^ n5560 ^ n1562 ;
  assign n19259 = n6932 ^ n5012 ^ 1'b0 ;
  assign n19260 = n2684 & ~n19259 ;
  assign n19261 = n19260 ^ n17371 ^ n3180 ;
  assign n19262 = n19261 ^ n5298 ^ n5249 ;
  assign n19263 = ( n15555 & n16503 ) | ( n15555 & n19262 ) | ( n16503 & n19262 ) ;
  assign n19264 = n5986 ^ n1892 ^ n339 ;
  assign n19277 = ~n4668 & n14493 ;
  assign n19274 = ( n716 & n4751 ) | ( n716 & ~n12252 ) | ( n4751 & ~n12252 ) ;
  assign n19275 = n19274 ^ n17433 ^ n6981 ;
  assign n19276 = n19275 ^ n14751 ^ n9816 ;
  assign n19269 = n536 & n5508 ;
  assign n19270 = n19269 ^ n5682 ^ n526 ;
  assign n19271 = n19270 ^ n5377 ^ n738 ;
  assign n19266 = ( n4275 & n5420 ) | ( n4275 & n15672 ) | ( n5420 & n15672 ) ;
  assign n19265 = n5330 & n6954 ;
  assign n19267 = n19266 ^ n19265 ^ n9957 ;
  assign n19268 = ( n10290 & n14807 ) | ( n10290 & n19267 ) | ( n14807 & n19267 ) ;
  assign n19272 = n19271 ^ n19268 ^ n3627 ;
  assign n19273 = n19272 ^ n13256 ^ n3499 ;
  assign n19278 = n19277 ^ n19276 ^ n19273 ;
  assign n19279 = ( n232 & n10713 ) | ( n232 & ~n11734 ) | ( n10713 & ~n11734 ) ;
  assign n19280 = ( n10143 & n13171 ) | ( n10143 & n13243 ) | ( n13171 & n13243 ) ;
  assign n19284 = n3951 & n16247 ;
  assign n19281 = n6070 & ~n7767 ;
  assign n19282 = n19281 ^ n3400 ^ 1'b0 ;
  assign n19283 = n19282 ^ n6764 ^ n3997 ;
  assign n19285 = n19284 ^ n19283 ^ x82 ;
  assign n19288 = n2769 ^ n2381 ^ n1313 ;
  assign n19289 = n19288 ^ n11233 ^ n411 ;
  assign n19286 = n9464 | n12013 ;
  assign n19287 = ( n15705 & n17589 ) | ( n15705 & ~n19286 ) | ( n17589 & ~n19286 ) ;
  assign n19290 = n19289 ^ n19287 ^ x25 ;
  assign n19291 = n19290 ^ n7505 ^ n6255 ;
  assign n19292 = ( n1940 & ~n12945 ) | ( n1940 & n13326 ) | ( ~n12945 & n13326 ) ;
  assign n19293 = ( x99 & n1767 ) | ( x99 & ~n6696 ) | ( n1767 & ~n6696 ) ;
  assign n19294 = ~n4896 & n5629 ;
  assign n19295 = n19294 ^ n2064 ^ 1'b0 ;
  assign n19296 = ( ~n8642 & n11792 ) | ( ~n8642 & n18453 ) | ( n11792 & n18453 ) ;
  assign n19297 = ( n4809 & ~n19295 ) | ( n4809 & n19296 ) | ( ~n19295 & n19296 ) ;
  assign n19298 = ( n7244 & ~n19293 ) | ( n7244 & n19297 ) | ( ~n19293 & n19297 ) ;
  assign n19299 = ( n384 & ~n2597 ) | ( n384 & n7413 ) | ( ~n2597 & n7413 ) ;
  assign n19300 = ( n3823 & n14231 ) | ( n3823 & ~n19299 ) | ( n14231 & ~n19299 ) ;
  assign n19301 = n19300 ^ n10419 ^ n1369 ;
  assign n19302 = n19301 ^ n11311 ^ n949 ;
  assign n19303 = ( n1467 & ~n7366 ) | ( n1467 & n13418 ) | ( ~n7366 & n13418 ) ;
  assign n19304 = ( n4011 & n7266 ) | ( n4011 & n14061 ) | ( n7266 & n14061 ) ;
  assign n19305 = n7394 ^ n5081 ^ n1203 ;
  assign n19306 = ( n12123 & n13695 ) | ( n12123 & ~n19305 ) | ( n13695 & ~n19305 ) ;
  assign n19307 = ( ~n19303 & n19304 ) | ( ~n19303 & n19306 ) | ( n19304 & n19306 ) ;
  assign n19308 = ( n2083 & n5450 ) | ( n2083 & ~n7324 ) | ( n5450 & ~n7324 ) ;
  assign n19309 = n19308 ^ n11786 ^ n11478 ;
  assign n19310 = n15472 ^ n8598 ^ n7320 ;
  assign n19311 = n2410 & ~n8247 ;
  assign n19312 = ~n19310 & n19311 ;
  assign n19313 = n15752 ^ n7631 ^ n7516 ;
  assign n19314 = ~n2941 & n4108 ;
  assign n19315 = n19314 ^ n7129 ^ 1'b0 ;
  assign n19316 = n19315 ^ n11795 ^ 1'b0 ;
  assign n19317 = n19313 & n19316 ;
  assign n19325 = ~n2704 & n5446 ;
  assign n19326 = n2406 & n19325 ;
  assign n19323 = n11839 ^ n4776 ^ n1383 ;
  assign n19324 = n19323 ^ n8360 ^ n206 ;
  assign n19318 = ( n1899 & n1913 ) | ( n1899 & ~n8798 ) | ( n1913 & ~n8798 ) ;
  assign n19319 = ( n3983 & n15836 ) | ( n3983 & n19318 ) | ( n15836 & n19318 ) ;
  assign n19320 = n19319 ^ n1331 ^ 1'b0 ;
  assign n19321 = n6154 | n19320 ;
  assign n19322 = n19321 ^ n11356 ^ n519 ;
  assign n19327 = n19326 ^ n19324 ^ n19322 ;
  assign n19328 = n14357 ^ n4205 ^ n708 ;
  assign n19329 = ( n6594 & ~n18802 ) | ( n6594 & n19328 ) | ( ~n18802 & n19328 ) ;
  assign n19330 = n13909 ^ n9950 ^ 1'b0 ;
  assign n19331 = n19329 & ~n19330 ;
  assign n19332 = n19331 ^ n6600 ^ 1'b0 ;
  assign n19333 = n8043 ^ n2032 ^ 1'b0 ;
  assign n19334 = n16825 & ~n19333 ;
  assign n19335 = ( n10384 & ~n13527 ) | ( n10384 & n19334 ) | ( ~n13527 & n19334 ) ;
  assign n19340 = ( n1399 & ~n4463 ) | ( n1399 & n11570 ) | ( ~n4463 & n11570 ) ;
  assign n19336 = ( ~n297 & n4549 ) | ( ~n297 & n5213 ) | ( n4549 & n5213 ) ;
  assign n19337 = n19336 ^ n2942 ^ x117 ;
  assign n19338 = n19337 ^ n10515 ^ 1'b0 ;
  assign n19339 = n5516 & ~n19338 ;
  assign n19341 = n19340 ^ n19339 ^ n5302 ;
  assign n19342 = n16299 ^ n14347 ^ n3794 ;
  assign n19343 = ( ~n3678 & n17061 ) | ( ~n3678 & n17075 ) | ( n17061 & n17075 ) ;
  assign n19344 = ( ~n2012 & n3364 ) | ( ~n2012 & n19343 ) | ( n3364 & n19343 ) ;
  assign n19345 = ( n3983 & ~n8395 ) | ( n3983 & n11426 ) | ( ~n8395 & n11426 ) ;
  assign n19346 = ( ~n9056 & n9124 ) | ( ~n9056 & n19345 ) | ( n9124 & n19345 ) ;
  assign n19347 = n19346 ^ n9748 ^ n6444 ;
  assign n19350 = n13806 & ~n15404 ;
  assign n19351 = ( n187 & n196 ) | ( n187 & ~n11161 ) | ( n196 & ~n11161 ) ;
  assign n19352 = n3566 & n19351 ;
  assign n19353 = n19352 ^ n5249 ^ 1'b0 ;
  assign n19354 = ( n8644 & n19350 ) | ( n8644 & ~n19353 ) | ( n19350 & ~n19353 ) ;
  assign n19348 = n8361 ^ n854 ^ n345 ;
  assign n19349 = n19348 ^ n17784 ^ n404 ;
  assign n19355 = n19354 ^ n19349 ^ n774 ;
  assign n19372 = n13073 ^ n3594 ^ n448 ;
  assign n19369 = ( n3286 & n4349 ) | ( n3286 & ~n18118 ) | ( n4349 & ~n18118 ) ;
  assign n19370 = n19369 ^ n2943 ^ n1771 ;
  assign n19362 = n9212 ^ n6858 ^ n4808 ;
  assign n19363 = n1626 & n2564 ;
  assign n19364 = ~x84 & n19363 ;
  assign n19365 = ( ~n3716 & n3956 ) | ( ~n3716 & n19364 ) | ( n3956 & n19364 ) ;
  assign n19366 = n2516 ^ n1443 ^ n722 ;
  assign n19367 = ( n779 & n7054 ) | ( n779 & n19366 ) | ( n7054 & n19366 ) ;
  assign n19368 = ( ~n19362 & n19365 ) | ( ~n19362 & n19367 ) | ( n19365 & n19367 ) ;
  assign n19371 = n19370 ^ n19368 ^ n3280 ;
  assign n19358 = ( n591 & n5643 ) | ( n591 & ~n6235 ) | ( n5643 & ~n6235 ) ;
  assign n19359 = n1670 & ~n8294 ;
  assign n19360 = ~n19358 & n19359 ;
  assign n19356 = n15484 ^ n3573 ^ n1889 ;
  assign n19357 = ~n1964 & n19356 ;
  assign n19361 = n19360 ^ n19357 ^ 1'b0 ;
  assign n19373 = n19372 ^ n19371 ^ n19361 ;
  assign n19374 = n15597 ^ n9024 ^ n4252 ;
  assign n19375 = n16355 & ~n19374 ;
  assign n19376 = n19375 ^ n11415 ^ n1393 ;
  assign n19377 = n7153 & ~n19376 ;
  assign n19378 = n9995 ^ n6835 ^ n4446 ;
  assign n19379 = ( n3394 & ~n9209 ) | ( n3394 & n13861 ) | ( ~n9209 & n13861 ) ;
  assign n19380 = n19379 ^ n11765 ^ n6120 ;
  assign n19381 = n17784 ^ n8925 ^ 1'b0 ;
  assign n19382 = ( n13184 & n14716 ) | ( n13184 & n19381 ) | ( n14716 & n19381 ) ;
  assign n19383 = n1374 & n18906 ;
  assign n19384 = ( n1388 & n3753 ) | ( n1388 & ~n13468 ) | ( n3753 & ~n13468 ) ;
  assign n19385 = n12890 ^ n11839 ^ 1'b0 ;
  assign n19386 = n19384 & ~n19385 ;
  assign n19387 = n19386 ^ n16244 ^ n15208 ;
  assign n19388 = n12232 ^ n736 ^ n654 ;
  assign n19389 = n19388 ^ n15579 ^ n10544 ;
  assign n19390 = n18876 ^ n14954 ^ n13352 ;
  assign n19391 = ( n4513 & n11491 ) | ( n4513 & ~n13173 ) | ( n11491 & ~n13173 ) ;
  assign n19392 = n19391 ^ n15092 ^ n12290 ;
  assign n19396 = n16475 ^ n12969 ^ n3266 ;
  assign n19393 = n7330 ^ n6894 ^ 1'b0 ;
  assign n19394 = n7995 & n19393 ;
  assign n19395 = n14719 & n19394 ;
  assign n19397 = n19396 ^ n19395 ^ 1'b0 ;
  assign n19398 = ( n1566 & ~n9469 ) | ( n1566 & n17582 ) | ( ~n9469 & n17582 ) ;
  assign n19399 = n19398 ^ n10381 ^ 1'b0 ;
  assign n19400 = n19399 ^ n13631 ^ n11708 ;
  assign n19401 = n16286 | n17886 ;
  assign n19402 = ( ~n959 & n3033 ) | ( ~n959 & n7624 ) | ( n3033 & n7624 ) ;
  assign n19403 = n11069 ^ n9776 ^ n218 ;
  assign n19404 = ( n1853 & n18469 ) | ( n1853 & n19403 ) | ( n18469 & n19403 ) ;
  assign n19405 = n6900 & n13776 ;
  assign n19406 = ~n8612 & n19405 ;
  assign n19407 = n7707 ^ n2079 ^ n1260 ;
  assign n19408 = ~n19406 & n19407 ;
  assign n19410 = n8979 ^ n6189 ^ n2511 ;
  assign n19411 = ~n8948 & n19410 ;
  assign n19409 = ( n206 & n5866 ) | ( n206 & ~n9105 ) | ( n5866 & ~n9105 ) ;
  assign n19412 = n19411 ^ n19409 ^ n2473 ;
  assign n19413 = ( n2589 & ~n2977 ) | ( n2589 & n12448 ) | ( ~n2977 & n12448 ) ;
  assign n19414 = ( ~n3360 & n7232 ) | ( ~n3360 & n7760 ) | ( n7232 & n7760 ) ;
  assign n19415 = ( x43 & n19413 ) | ( x43 & ~n19414 ) | ( n19413 & ~n19414 ) ;
  assign n19424 = ( n3466 & n4400 ) | ( n3466 & n17504 ) | ( n4400 & n17504 ) ;
  assign n19425 = ( n9341 & n13803 ) | ( n9341 & ~n19424 ) | ( n13803 & ~n19424 ) ;
  assign n19426 = ( n1357 & n1454 ) | ( n1357 & ~n19425 ) | ( n1454 & ~n19425 ) ;
  assign n19416 = ( ~n1473 & n2928 ) | ( ~n1473 & n9327 ) | ( n2928 & n9327 ) ;
  assign n19417 = n19416 ^ n4436 ^ n2167 ;
  assign n19419 = ( n2923 & n4519 ) | ( n2923 & ~n8661 ) | ( n4519 & ~n8661 ) ;
  assign n19418 = n12433 ^ n11185 ^ n5308 ;
  assign n19420 = n19419 ^ n19418 ^ n2613 ;
  assign n19421 = ( ~n1945 & n19417 ) | ( ~n1945 & n19420 ) | ( n19417 & n19420 ) ;
  assign n19422 = n19421 ^ n19277 ^ n8470 ;
  assign n19423 = n19422 ^ n16898 ^ n8963 ;
  assign n19427 = n19426 ^ n19423 ^ n18686 ;
  assign n19428 = n10425 ^ n6157 ^ n2195 ;
  assign n19429 = n13331 ^ n8959 ^ n545 ;
  assign n19430 = n19429 ^ n14488 ^ n9181 ;
  assign n19431 = ( n11733 & n19428 ) | ( n11733 & ~n19430 ) | ( n19428 & ~n19430 ) ;
  assign n19432 = ( ~n10919 & n13178 ) | ( ~n10919 & n19431 ) | ( n13178 & n19431 ) ;
  assign n19435 = ( n4708 & ~n7876 ) | ( n4708 & n9658 ) | ( ~n7876 & n9658 ) ;
  assign n19434 = ( n200 & n2110 ) | ( n200 & ~n16727 ) | ( n2110 & ~n16727 ) ;
  assign n19436 = n19435 ^ n19434 ^ n772 ;
  assign n19433 = ~n3072 & n18250 ;
  assign n19437 = n19436 ^ n19433 ^ 1'b0 ;
  assign n19438 = ( n2291 & n12130 ) | ( n2291 & ~n17290 ) | ( n12130 & ~n17290 ) ;
  assign n19439 = n16068 ^ n9275 ^ 1'b0 ;
  assign n19440 = ( n1566 & n2450 ) | ( n1566 & n3484 ) | ( n2450 & n3484 ) ;
  assign n19441 = n19440 ^ n12715 ^ n3136 ;
  assign n19442 = ( n193 & n12260 ) | ( n193 & n19441 ) | ( n12260 & n19441 ) ;
  assign n19445 = ( n1023 & n5019 ) | ( n1023 & ~n9735 ) | ( n5019 & ~n9735 ) ;
  assign n19446 = n19445 ^ n2810 ^ n2204 ;
  assign n19444 = n18438 ^ n11571 ^ n2609 ;
  assign n19443 = ( n5535 & n13335 ) | ( n5535 & ~n14368 ) | ( n13335 & ~n14368 ) ;
  assign n19447 = n19446 ^ n19444 ^ n19443 ;
  assign n19448 = n19442 & ~n19447 ;
  assign n19451 = n12047 ^ n1858 ^ 1'b0 ;
  assign n19452 = n628 & ~n19451 ;
  assign n19449 = ( n494 & n3294 ) | ( n494 & ~n10598 ) | ( n3294 & ~n10598 ) ;
  assign n19450 = n1476 & n19449 ;
  assign n19453 = n19452 ^ n19450 ^ n7418 ;
  assign n19454 = n6976 ^ n2870 ^ x106 ;
  assign n19455 = ( n4607 & n14830 ) | ( n4607 & n19454 ) | ( n14830 & n19454 ) ;
  assign n19456 = n19455 ^ n13079 ^ n10995 ;
  assign n19457 = ( n2065 & n3465 ) | ( n2065 & ~n17210 ) | ( n3465 & ~n17210 ) ;
  assign n19458 = ( n8050 & ~n13776 ) | ( n8050 & n19457 ) | ( ~n13776 & n19457 ) ;
  assign n19459 = ( n1455 & n3603 ) | ( n1455 & n19016 ) | ( n3603 & n19016 ) ;
  assign n19460 = ( x20 & n14348 ) | ( x20 & n19459 ) | ( n14348 & n19459 ) ;
  assign n19461 = n19460 ^ n16248 ^ n571 ;
  assign n19462 = n19461 ^ n7771 ^ n623 ;
  assign n19463 = ( n10749 & ~n15670 ) | ( n10749 & n19462 ) | ( ~n15670 & n19462 ) ;
  assign n19464 = n3170 & ~n7724 ;
  assign n19465 = n19464 ^ n15184 ^ 1'b0 ;
  assign n19466 = ( n2524 & n9197 ) | ( n2524 & ~n19465 ) | ( n9197 & ~n19465 ) ;
  assign n19469 = n10491 ^ n10464 ^ n4744 ;
  assign n19470 = n19469 ^ n17019 ^ 1'b0 ;
  assign n19467 = n7199 & ~n14543 ;
  assign n19468 = n19467 ^ n14810 ^ 1'b0 ;
  assign n19471 = n19470 ^ n19468 ^ n9513 ;
  assign n19477 = ( ~n7489 & n8492 ) | ( ~n7489 & n14104 ) | ( n8492 & n14104 ) ;
  assign n19472 = n6086 & ~n9477 ;
  assign n19473 = n19472 ^ n10179 ^ 1'b0 ;
  assign n19474 = ( n196 & ~n2784 ) | ( n196 & n5991 ) | ( ~n2784 & n5991 ) ;
  assign n19475 = n19474 ^ n18000 ^ n8384 ;
  assign n19476 = ( n10820 & ~n19473 ) | ( n10820 & n19475 ) | ( ~n19473 & n19475 ) ;
  assign n19478 = n19477 ^ n19476 ^ n9267 ;
  assign n19479 = ( n5449 & n7708 ) | ( n5449 & ~n11230 ) | ( n7708 & ~n11230 ) ;
  assign n19483 = ( n7571 & n18245 ) | ( n7571 & n18537 ) | ( n18245 & n18537 ) ;
  assign n19480 = x2 & n4876 ;
  assign n19481 = n19480 ^ n4799 ^ 1'b0 ;
  assign n19482 = ( ~n4045 & n9356 ) | ( ~n4045 & n19481 ) | ( n9356 & n19481 ) ;
  assign n19484 = n19483 ^ n19482 ^ n18578 ;
  assign n19485 = n12686 ^ n8454 ^ n4650 ;
  assign n19486 = n19485 ^ n14404 ^ n6845 ;
  assign n19487 = n18139 ^ n2077 ^ 1'b0 ;
  assign n19489 = n5428 ^ n1932 ^ 1'b0 ;
  assign n19488 = n19315 ^ n9400 ^ n3914 ;
  assign n19490 = n19489 ^ n19488 ^ 1'b0 ;
  assign n19491 = n10357 ^ n9837 ^ n6878 ;
  assign n19492 = ( n5127 & ~n6130 ) | ( n5127 & n7164 ) | ( ~n6130 & n7164 ) ;
  assign n19493 = n19492 ^ n4632 ^ 1'b0 ;
  assign n19494 = ~n19491 & n19493 ;
  assign n19495 = ( x48 & n5575 ) | ( x48 & n11253 ) | ( n5575 & n11253 ) ;
  assign n19496 = n19495 ^ n1663 ^ n564 ;
  assign n19497 = n5154 ^ n4207 ^ n178 ;
  assign n19498 = n19497 ^ n3953 ^ n3476 ;
  assign n19499 = n19498 ^ n16779 ^ n5353 ;
  assign n19501 = n1285 | n3506 ;
  assign n19502 = n19501 ^ n10925 ^ 1'b0 ;
  assign n19500 = ( ~n1985 & n2269 ) | ( ~n1985 & n6808 ) | ( n2269 & n6808 ) ;
  assign n19503 = n19502 ^ n19500 ^ n11891 ;
  assign n19511 = ( ~n7847 & n8595 ) | ( ~n7847 & n9554 ) | ( n8595 & n9554 ) ;
  assign n19512 = n19511 ^ n17560 ^ 1'b0 ;
  assign n19513 = ( n2991 & n10894 ) | ( n2991 & n12533 ) | ( n10894 & n12533 ) ;
  assign n19514 = n19512 & n19513 ;
  assign n19515 = n19514 ^ n4788 ^ 1'b0 ;
  assign n19504 = ( n1611 & n2432 ) | ( n1611 & n6709 ) | ( n2432 & n6709 ) ;
  assign n19506 = ~n6459 & n7733 ;
  assign n19507 = n19506 ^ n7665 ^ 1'b0 ;
  assign n19505 = n3806 ^ n3514 ^ 1'b0 ;
  assign n19508 = n19507 ^ n19505 ^ n4126 ;
  assign n19509 = ( ~n2619 & n5669 ) | ( ~n2619 & n19508 ) | ( n5669 & n19508 ) ;
  assign n19510 = ( n13978 & ~n19504 ) | ( n13978 & n19509 ) | ( ~n19504 & n19509 ) ;
  assign n19516 = n19515 ^ n19510 ^ n6884 ;
  assign n19517 = ( n1825 & ~n10461 ) | ( n1825 & n18507 ) | ( ~n10461 & n18507 ) ;
  assign n19518 = n19517 ^ n12024 ^ n7230 ;
  assign n19519 = n17637 ^ n5319 ^ n895 ;
  assign n19520 = n19519 ^ n16558 ^ n8375 ;
  assign n19521 = n19520 ^ n19216 ^ n17554 ;
  assign n19524 = ( n3340 & n6592 ) | ( n3340 & n9811 ) | ( n6592 & n9811 ) ;
  assign n19522 = n6098 & n11185 ;
  assign n19523 = n19522 ^ n17681 ^ 1'b0 ;
  assign n19525 = n19524 ^ n19523 ^ n7666 ;
  assign n19526 = n5763 & n7618 ;
  assign n19527 = ( n5880 & n10121 ) | ( n5880 & ~n19526 ) | ( n10121 & ~n19526 ) ;
  assign n19528 = ( n421 & n2861 ) | ( n421 & ~n19527 ) | ( n2861 & ~n19527 ) ;
  assign n19529 = n17574 ^ n17145 ^ n401 ;
  assign n19534 = n9721 & ~n13028 ;
  assign n19531 = n13517 ^ n13447 ^ 1'b0 ;
  assign n19532 = n8965 & n19531 ;
  assign n19530 = n1112 & n9487 ;
  assign n19533 = n19532 ^ n19530 ^ 1'b0 ;
  assign n19535 = n19534 ^ n19533 ^ n16327 ;
  assign n19536 = n19052 ^ n5947 ^ 1'b0 ;
  assign n19537 = n5756 ^ n4441 ^ 1'b0 ;
  assign n19538 = n4778 & ~n19537 ;
  assign n19539 = n11615 ^ n9972 ^ n1198 ;
  assign n19540 = n15424 ^ n12309 ^ n10636 ;
  assign n19541 = n5278 & n19540 ;
  assign n19542 = n19541 ^ n12116 ^ 1'b0 ;
  assign n19543 = ( n4669 & n9717 ) | ( n4669 & ~n19542 ) | ( n9717 & ~n19542 ) ;
  assign n19546 = n14684 ^ n9212 ^ n7320 ;
  assign n19544 = n17706 ^ n10942 ^ n4539 ;
  assign n19545 = n6364 & n19544 ;
  assign n19547 = n19546 ^ n19545 ^ 1'b0 ;
  assign n19548 = ~n3417 & n12402 ;
  assign n19549 = n19548 ^ n15383 ^ 1'b0 ;
  assign n19550 = n19549 ^ n17986 ^ n5673 ;
  assign n19551 = ( ~n5619 & n8528 ) | ( ~n5619 & n17875 ) | ( n8528 & n17875 ) ;
  assign n19552 = ( x37 & n19550 ) | ( x37 & ~n19551 ) | ( n19550 & ~n19551 ) ;
  assign n19553 = ( n7185 & n15672 ) | ( n7185 & ~n16040 ) | ( n15672 & ~n16040 ) ;
  assign n19554 = n13759 ^ n9371 ^ n3398 ;
  assign n19555 = n19369 ^ n16634 ^ x31 ;
  assign n19556 = ( n11869 & n19554 ) | ( n11869 & ~n19555 ) | ( n19554 & ~n19555 ) ;
  assign n19557 = ( n3302 & n5322 ) | ( n3302 & n6527 ) | ( n5322 & n6527 ) ;
  assign n19558 = ( ~n197 & n1977 ) | ( ~n197 & n19557 ) | ( n1977 & n19557 ) ;
  assign n19559 = ( x86 & n2667 ) | ( x86 & ~n5488 ) | ( n2667 & ~n5488 ) ;
  assign n19560 = n4318 & n19559 ;
  assign n19563 = ( n6733 & n16351 ) | ( n6733 & n18753 ) | ( n16351 & n18753 ) ;
  assign n19561 = ( ~n1118 & n2208 ) | ( ~n1118 & n3933 ) | ( n2208 & n3933 ) ;
  assign n19562 = ~n6910 & n19561 ;
  assign n19564 = n19563 ^ n19562 ^ 1'b0 ;
  assign n19567 = n7765 ^ n3121 ^ 1'b0 ;
  assign n19568 = n4443 | n19567 ;
  assign n19565 = ( n439 & ~n3156 ) | ( n439 & n5486 ) | ( ~n3156 & n5486 ) ;
  assign n19566 = n19565 ^ n711 ^ 1'b0 ;
  assign n19569 = n19568 ^ n19566 ^ n9998 ;
  assign n19570 = n19569 ^ n17532 ^ n743 ;
  assign n19571 = n9686 & ~n12096 ;
  assign n19572 = n19571 ^ n2415 ^ 1'b0 ;
  assign n19573 = ( x51 & n7527 ) | ( x51 & n19572 ) | ( n7527 & n19572 ) ;
  assign n19574 = ( ~n5761 & n7626 ) | ( ~n5761 & n13473 ) | ( n7626 & n13473 ) ;
  assign n19575 = ( ~n13866 & n16072 ) | ( ~n13866 & n17462 ) | ( n16072 & n17462 ) ;
  assign n19576 = n17245 ^ n16275 ^ n16172 ;
  assign n19577 = n19576 ^ n13400 ^ n10001 ;
  assign n19578 = ( ~n18663 & n19575 ) | ( ~n18663 & n19577 ) | ( n19575 & n19577 ) ;
  assign n19582 = n13282 ^ n12770 ^ n6839 ;
  assign n19579 = ( n2094 & n3471 ) | ( n2094 & ~n6285 ) | ( n3471 & ~n6285 ) ;
  assign n19580 = ( n931 & n12014 ) | ( n931 & n19579 ) | ( n12014 & n19579 ) ;
  assign n19581 = n4712 & ~n19580 ;
  assign n19583 = n19582 ^ n19581 ^ 1'b0 ;
  assign n19588 = n18499 ^ n3349 ^ 1'b0 ;
  assign n19585 = ( n3428 & n3983 ) | ( n3428 & n10330 ) | ( n3983 & n10330 ) ;
  assign n19586 = ( ~n9484 & n15719 ) | ( ~n9484 & n19585 ) | ( n15719 & n19585 ) ;
  assign n19584 = n4263 & n5036 ;
  assign n19587 = n19586 ^ n19584 ^ 1'b0 ;
  assign n19589 = n19588 ^ n19587 ^ n14250 ;
  assign n19590 = n19527 ^ n13581 ^ n6752 ;
  assign n19591 = n19590 ^ n9124 ^ n5214 ;
  assign n19592 = n10165 ^ n6666 ^ n4796 ;
  assign n19593 = ( n1486 & ~n3421 ) | ( n1486 & n16895 ) | ( ~n3421 & n16895 ) ;
  assign n19594 = n19593 ^ n3630 ^ n2243 ;
  assign n19595 = n19594 ^ n5881 ^ n4896 ;
  assign n19596 = n5954 | n6566 ;
  assign n19597 = n15683 ^ n11986 ^ n8374 ;
  assign n19598 = ( n919 & n1293 ) | ( n919 & ~n5385 ) | ( n1293 & ~n5385 ) ;
  assign n19599 = n7568 & n19598 ;
  assign n19600 = ~n19597 & n19599 ;
  assign n19601 = ( n1527 & n8250 ) | ( n1527 & n17020 ) | ( n8250 & n17020 ) ;
  assign n19602 = n19601 ^ n14958 ^ n5591 ;
  assign n19603 = n12171 ^ n4840 ^ n2889 ;
  assign n19604 = ( n3555 & n11439 ) | ( n3555 & n19603 ) | ( n11439 & n19603 ) ;
  assign n19605 = n12186 ^ n9374 ^ n5024 ;
  assign n19606 = ( ~n1162 & n5355 ) | ( ~n1162 & n7130 ) | ( n5355 & n7130 ) ;
  assign n19607 = n1077 | n17339 ;
  assign n19608 = n19606 & ~n19607 ;
  assign n19609 = ( n740 & ~n5482 ) | ( n740 & n19608 ) | ( ~n5482 & n19608 ) ;
  assign n19610 = n13352 | n17356 ;
  assign n19611 = n1661 | n19610 ;
  assign n19612 = n19611 ^ n11671 ^ n2266 ;
  assign n19613 = ~n5887 & n12548 ;
  assign n19614 = ( ~n6991 & n16416 ) | ( ~n6991 & n19613 ) | ( n16416 & n19613 ) ;
  assign n19615 = ( ~n2100 & n7621 ) | ( ~n2100 & n11363 ) | ( n7621 & n11363 ) ;
  assign n19616 = n9834 ^ n486 ^ 1'b0 ;
  assign n19617 = n19615 | n19616 ;
  assign n19618 = ( n2784 & n4192 ) | ( n2784 & ~n19617 ) | ( n4192 & ~n19617 ) ;
  assign n19619 = n18951 ^ n17485 ^ 1'b0 ;
  assign n19620 = ( ~n9061 & n9395 ) | ( ~n9061 & n9682 ) | ( n9395 & n9682 ) ;
  assign n19621 = ( n4443 & n9172 ) | ( n4443 & ~n14942 ) | ( n9172 & ~n14942 ) ;
  assign n19622 = n19620 & ~n19621 ;
  assign n19623 = n10061 ^ n8129 ^ n4027 ;
  assign n19624 = n19623 ^ n7883 ^ 1'b0 ;
  assign n19625 = n19624 ^ n18453 ^ n17113 ;
  assign n19626 = n17826 ^ n4146 ^ n775 ;
  assign n19627 = ( n8640 & n15399 ) | ( n8640 & ~n19626 ) | ( n15399 & ~n19626 ) ;
  assign n19631 = ( n1904 & n10658 ) | ( n1904 & n17527 ) | ( n10658 & n17527 ) ;
  assign n19630 = n3237 & ~n4240 ;
  assign n19632 = n19631 ^ n19630 ^ 1'b0 ;
  assign n19628 = ( n5116 & n10178 ) | ( n5116 & ~n10505 ) | ( n10178 & ~n10505 ) ;
  assign n19629 = n19628 ^ n12832 ^ n6891 ;
  assign n19633 = n19632 ^ n19629 ^ n19457 ;
  assign n19634 = n1166 & ~n9469 ;
  assign n19635 = ~n13695 & n19634 ;
  assign n19636 = ( n3850 & ~n8889 ) | ( n3850 & n15062 ) | ( ~n8889 & n15062 ) ;
  assign n19637 = n17576 ^ n8897 ^ n7287 ;
  assign n19638 = ~n2071 & n19637 ;
  assign n19639 = ~n19636 & n19638 ;
  assign n19640 = ( n276 & ~n8857 ) | ( n276 & n10818 ) | ( ~n8857 & n10818 ) ;
  assign n19641 = ( ~n5853 & n9225 ) | ( ~n5853 & n19640 ) | ( n9225 & n19640 ) ;
  assign n19642 = n527 | n19641 ;
  assign n19643 = ~n3591 & n12766 ;
  assign n19644 = ( n15404 & ~n16536 ) | ( n15404 & n19643 ) | ( ~n16536 & n19643 ) ;
  assign n19645 = n3404 & ~n11972 ;
  assign n19646 = n12482 ^ n1074 ^ 1'b0 ;
  assign n19647 = ( ~n9766 & n19645 ) | ( ~n9766 & n19646 ) | ( n19645 & n19646 ) ;
  assign n19648 = ( n2662 & n7210 ) | ( n2662 & n12433 ) | ( n7210 & n12433 ) ;
  assign n19649 = n19648 ^ n14076 ^ n10951 ;
  assign n19650 = n9555 ^ n6883 ^ n4166 ;
  assign n19651 = ( n3779 & n10765 ) | ( n3779 & ~n17635 ) | ( n10765 & ~n17635 ) ;
  assign n19652 = ( n10292 & n12926 ) | ( n10292 & ~n19651 ) | ( n12926 & ~n19651 ) ;
  assign n19653 = n8849 ^ n6210 ^ n469 ;
  assign n19654 = n19653 ^ n6174 ^ n3145 ;
  assign n19655 = ( n646 & ~n649 ) | ( n646 & n659 ) | ( ~n649 & n659 ) ;
  assign n19656 = ( n3011 & n4138 ) | ( n3011 & ~n19655 ) | ( n4138 & ~n19655 ) ;
  assign n19657 = n19656 ^ n10923 ^ n801 ;
  assign n19658 = ( ~n854 & n1651 ) | ( ~n854 & n19585 ) | ( n1651 & n19585 ) ;
  assign n19659 = ( n1405 & n4479 ) | ( n1405 & ~n19658 ) | ( n4479 & ~n19658 ) ;
  assign n19660 = ( ~n14797 & n14904 ) | ( ~n14797 & n19659 ) | ( n14904 & n19659 ) ;
  assign n19661 = n19660 ^ n14338 ^ n5019 ;
  assign n19662 = n7651 ^ n6152 ^ n2918 ;
  assign n19663 = ( n6362 & n9742 ) | ( n6362 & ~n19662 ) | ( n9742 & ~n19662 ) ;
  assign n19664 = ~n1982 & n3117 ;
  assign n19665 = n5119 & n19664 ;
  assign n19666 = ( n4370 & n10714 ) | ( n4370 & n19036 ) | ( n10714 & n19036 ) ;
  assign n19667 = ( ~n1606 & n5332 ) | ( ~n1606 & n19631 ) | ( n5332 & n19631 ) ;
  assign n19668 = ( n10879 & ~n19666 ) | ( n10879 & n19667 ) | ( ~n19666 & n19667 ) ;
  assign n19669 = ~n19665 & n19668 ;
  assign n19673 = ( n1844 & n7462 ) | ( n1844 & n10845 ) | ( n7462 & n10845 ) ;
  assign n19674 = n19673 ^ n1141 ^ 1'b0 ;
  assign n19675 = ( n6985 & ~n7122 ) | ( n6985 & n19674 ) | ( ~n7122 & n19674 ) ;
  assign n19671 = n15348 ^ n7158 ^ n2758 ;
  assign n19670 = n838 & n877 ;
  assign n19672 = n19671 ^ n19670 ^ n3976 ;
  assign n19676 = n19675 ^ n19672 ^ n6476 ;
  assign n19677 = n11235 ^ n7243 ^ n2814 ;
  assign n19678 = n13253 ^ n10385 ^ 1'b0 ;
  assign n19679 = n1708 | n19678 ;
  assign n19680 = n19679 ^ n17242 ^ 1'b0 ;
  assign n19681 = ( n391 & ~n8942 ) | ( n391 & n10691 ) | ( ~n8942 & n10691 ) ;
  assign n19682 = ( n3202 & ~n4237 ) | ( n3202 & n19681 ) | ( ~n4237 & n19681 ) ;
  assign n19685 = ( ~n1316 & n3839 ) | ( ~n1316 & n8162 ) | ( n3839 & n8162 ) ;
  assign n19686 = n688 & n7403 ;
  assign n19687 = n19686 ^ n8286 ^ n1084 ;
  assign n19688 = ( n6823 & ~n19685 ) | ( n6823 & n19687 ) | ( ~n19685 & n19687 ) ;
  assign n19689 = n8513 ^ n3977 ^ 1'b0 ;
  assign n19690 = n19688 & n19689 ;
  assign n19683 = ( n249 & n5504 ) | ( n249 & n9480 ) | ( n5504 & n9480 ) ;
  assign n19684 = ( ~n6312 & n6849 ) | ( ~n6312 & n19683 ) | ( n6849 & n19683 ) ;
  assign n19691 = n19690 ^ n19684 ^ n8704 ;
  assign n19693 = ( ~n1531 & n3259 ) | ( ~n1531 & n11933 ) | ( n3259 & n11933 ) ;
  assign n19692 = n17063 ^ n16553 ^ 1'b0 ;
  assign n19694 = n19693 ^ n19692 ^ n14205 ;
  assign n19695 = ~n7729 & n16587 ;
  assign n19696 = n19695 ^ n18600 ^ n1717 ;
  assign n19697 = ( n2811 & n3971 ) | ( n2811 & ~n8212 ) | ( n3971 & ~n8212 ) ;
  assign n19699 = ( ~n1392 & n5537 ) | ( ~n1392 & n10779 ) | ( n5537 & n10779 ) ;
  assign n19698 = ~n4574 & n6840 ;
  assign n19700 = n19699 ^ n19698 ^ n1931 ;
  assign n19701 = n13030 ^ n5408 ^ 1'b0 ;
  assign n19702 = ~n466 & n19701 ;
  assign n19703 = ~n14748 & n19702 ;
  assign n19704 = n14499 ^ n11146 ^ n7406 ;
  assign n19705 = n8534 ^ n4940 ^ n3725 ;
  assign n19706 = ( n7136 & n10228 ) | ( n7136 & n12549 ) | ( n10228 & n12549 ) ;
  assign n19707 = ( n4081 & n8051 ) | ( n4081 & n10085 ) | ( n8051 & n10085 ) ;
  assign n19708 = ~n3889 & n7173 ;
  assign n19709 = n19708 ^ n5863 ^ 1'b0 ;
  assign n19710 = n18431 | n19709 ;
  assign n19711 = n19710 ^ n11774 ^ n10620 ;
  assign n19712 = n12234 | n14090 ;
  assign n19713 = n3832 ^ n3691 ^ 1'b0 ;
  assign n19714 = ( n605 & ~n3154 ) | ( n605 & n19713 ) | ( ~n3154 & n19713 ) ;
  assign n19715 = n4795 ^ x118 ^ 1'b0 ;
  assign n19716 = n19714 & ~n19715 ;
  assign n19717 = ( ~n2010 & n19712 ) | ( ~n2010 & n19716 ) | ( n19712 & n19716 ) ;
  assign n19718 = n10571 ^ n4627 ^ x0 ;
  assign n19719 = ( n2119 & n3667 ) | ( n2119 & n4838 ) | ( n3667 & n4838 ) ;
  assign n19720 = ( n232 & ~n12146 ) | ( n232 & n19719 ) | ( ~n12146 & n19719 ) ;
  assign n19721 = n12190 ^ n6725 ^ n5014 ;
  assign n19722 = ( ~n1057 & n15737 ) | ( ~n1057 & n19721 ) | ( n15737 & n19721 ) ;
  assign n19723 = n19722 ^ n5174 ^ 1'b0 ;
  assign n19724 = n19723 ^ n3433 ^ n2426 ;
  assign n19725 = ( n346 & ~n2411 ) | ( n346 & n3635 ) | ( ~n2411 & n3635 ) ;
  assign n19726 = n19725 ^ n9795 ^ n3474 ;
  assign n19727 = n3609 ^ n3041 ^ n167 ;
  assign n19728 = ( n2309 & n10219 ) | ( n2309 & ~n11688 ) | ( n10219 & ~n11688 ) ;
  assign n19729 = ( ~n6273 & n19727 ) | ( ~n6273 & n19728 ) | ( n19727 & n19728 ) ;
  assign n19730 = ( n3396 & n19726 ) | ( n3396 & n19729 ) | ( n19726 & n19729 ) ;
  assign n19731 = ( n139 & n4390 ) | ( n139 & ~n7042 ) | ( n4390 & ~n7042 ) ;
  assign n19732 = ( ~n8465 & n11937 ) | ( ~n8465 & n16132 ) | ( n11937 & n16132 ) ;
  assign n19733 = ( n4303 & n6330 ) | ( n4303 & ~n13413 ) | ( n6330 & ~n13413 ) ;
  assign n19734 = ( n17489 & n19732 ) | ( n17489 & n19733 ) | ( n19732 & n19733 ) ;
  assign n19735 = ( ~n5754 & n13544 ) | ( ~n5754 & n19734 ) | ( n13544 & n19734 ) ;
  assign n19736 = ( ~n5755 & n19731 ) | ( ~n5755 & n19735 ) | ( n19731 & n19735 ) ;
  assign n19737 = n4790 ^ x126 ^ 1'b0 ;
  assign n19738 = ( n2014 & n8605 ) | ( n2014 & n19737 ) | ( n8605 & n19737 ) ;
  assign n19739 = ( n1084 & n3453 ) | ( n1084 & n9343 ) | ( n3453 & n9343 ) ;
  assign n19746 = n761 & n5609 ;
  assign n19747 = ~n13715 & n19746 ;
  assign n19745 = ( n10011 & ~n10291 ) | ( n10011 & n10523 ) | ( ~n10291 & n10523 ) ;
  assign n19740 = ( n5367 & n5755 ) | ( n5367 & ~n6070 ) | ( n5755 & ~n6070 ) ;
  assign n19741 = ~n7531 & n19740 ;
  assign n19742 = ~n4395 & n19741 ;
  assign n19743 = ( n4810 & n17049 ) | ( n4810 & n19742 ) | ( n17049 & n19742 ) ;
  assign n19744 = ( ~n746 & n7292 ) | ( ~n746 & n19743 ) | ( n7292 & n19743 ) ;
  assign n19748 = n19747 ^ n19745 ^ n19744 ;
  assign n19749 = n18511 ^ n16870 ^ 1'b0 ;
  assign n19750 = n9917 & ~n19749 ;
  assign n19751 = n19750 ^ n19274 ^ n1100 ;
  assign n19753 = ( n3908 & n7499 ) | ( n3908 & ~n7837 ) | ( n7499 & ~n7837 ) ;
  assign n19754 = n19753 ^ n13282 ^ n2068 ;
  assign n19752 = n1329 & ~n9257 ;
  assign n19755 = n19754 ^ n19752 ^ n4874 ;
  assign n19756 = n19755 ^ n9549 ^ n9497 ;
  assign n19762 = n12061 ^ n6171 ^ n4392 ;
  assign n19757 = n11008 ^ n9899 ^ n1440 ;
  assign n19758 = n5429 & n8946 ;
  assign n19759 = n19758 ^ n4237 ^ 1'b0 ;
  assign n19760 = ( ~n9003 & n10449 ) | ( ~n9003 & n19759 ) | ( n10449 & n19759 ) ;
  assign n19761 = ( n2203 & n19757 ) | ( n2203 & n19760 ) | ( n19757 & n19760 ) ;
  assign n19763 = n19762 ^ n19761 ^ n13976 ;
  assign n19765 = ( n6239 & n8644 ) | ( n6239 & n17681 ) | ( n8644 & n17681 ) ;
  assign n19764 = n12084 ^ n5978 ^ n1739 ;
  assign n19766 = n19765 ^ n19764 ^ n10877 ;
  assign n19767 = ( ~n8450 & n9616 ) | ( ~n8450 & n19766 ) | ( n9616 & n19766 ) ;
  assign n19768 = ( n293 & n9147 ) | ( n293 & n19199 ) | ( n9147 & n19199 ) ;
  assign n19769 = n2813 & ~n8738 ;
  assign n19770 = n19769 ^ n11146 ^ 1'b0 ;
  assign n19771 = n4105 & ~n19770 ;
  assign n19772 = n6449 ^ n1599 ^ 1'b0 ;
  assign n19773 = n19772 ^ n11624 ^ n6782 ;
  assign n19774 = n19773 ^ n7068 ^ n3814 ;
  assign n19775 = ( n8840 & n16644 ) | ( n8840 & n19774 ) | ( n16644 & n19774 ) ;
  assign n19776 = n19775 ^ n7390 ^ n215 ;
  assign n19777 = ~n16669 & n19776 ;
  assign n19778 = n19777 ^ n7372 ^ 1'b0 ;
  assign n19779 = ( n772 & ~n873 ) | ( n772 & n6799 ) | ( ~n873 & n6799 ) ;
  assign n19781 = ~n5488 & n7050 ;
  assign n19782 = n19781 ^ n3891 ^ 1'b0 ;
  assign n19783 = ( n424 & n5140 ) | ( n424 & n19782 ) | ( n5140 & n19782 ) ;
  assign n19780 = ( ~n1814 & n2444 ) | ( ~n1814 & n3515 ) | ( n2444 & n3515 ) ;
  assign n19784 = n19783 ^ n19780 ^ n10669 ;
  assign n19785 = n2774 | n19784 ;
  assign n19786 = ( n4658 & n7717 ) | ( n4658 & ~n19785 ) | ( n7717 & ~n19785 ) ;
  assign n19787 = n10783 ^ n6583 ^ n767 ;
  assign n19788 = ( n5961 & n19504 ) | ( n5961 & ~n19787 ) | ( n19504 & ~n19787 ) ;
  assign n19789 = ( ~n14072 & n19786 ) | ( ~n14072 & n19788 ) | ( n19786 & n19788 ) ;
  assign n19790 = ( n974 & ~n3199 ) | ( n974 & n6011 ) | ( ~n3199 & n6011 ) ;
  assign n19791 = ( n1354 & n1792 ) | ( n1354 & n3706 ) | ( n1792 & n3706 ) ;
  assign n19792 = n19790 | n19791 ;
  assign n19793 = n19792 ^ n11297 ^ 1'b0 ;
  assign n19794 = n19793 ^ n14668 ^ n13423 ;
  assign n19795 = n11333 ^ n8646 ^ n2120 ;
  assign n19796 = ( n9383 & n19794 ) | ( n9383 & ~n19795 ) | ( n19794 & ~n19795 ) ;
  assign n19797 = n19796 ^ n12108 ^ n11480 ;
  assign n19798 = ( n5895 & n6125 ) | ( n5895 & ~n10236 ) | ( n6125 & ~n10236 ) ;
  assign n19799 = n7989 ^ n4085 ^ 1'b0 ;
  assign n19800 = n5775 | n19799 ;
  assign n19801 = n19800 ^ n176 ^ 1'b0 ;
  assign n19802 = n15870 ^ n4588 ^ n4188 ;
  assign n19803 = n19802 ^ n9721 ^ n1496 ;
  assign n19804 = ( n19798 & n19801 ) | ( n19798 & n19803 ) | ( n19801 & n19803 ) ;
  assign n19806 = n16775 ^ n13855 ^ n10268 ;
  assign n19805 = n10636 | n12206 ;
  assign n19807 = n19806 ^ n19805 ^ 1'b0 ;
  assign n19808 = ( n4168 & n18938 ) | ( n4168 & n19807 ) | ( n18938 & n19807 ) ;
  assign n19810 = ( n3064 & n3999 ) | ( n3064 & n14603 ) | ( n3999 & n14603 ) ;
  assign n19809 = ( n6199 & ~n7966 ) | ( n6199 & n9785 ) | ( ~n7966 & n9785 ) ;
  assign n19811 = n19810 ^ n19809 ^ n11254 ;
  assign n19812 = n13324 ^ n5992 ^ n4023 ;
  assign n19813 = ( n9313 & n9504 ) | ( n9313 & ~n19812 ) | ( n9504 & ~n19812 ) ;
  assign n19816 = ( n4394 & n6629 ) | ( n4394 & n8657 ) | ( n6629 & n8657 ) ;
  assign n19814 = ( ~n6696 & n10520 ) | ( ~n6696 & n17645 ) | ( n10520 & n17645 ) ;
  assign n19815 = n19814 ^ n17772 ^ n11375 ;
  assign n19817 = n19816 ^ n19815 ^ n14796 ;
  assign n19818 = ( ~n5515 & n9538 ) | ( ~n5515 & n18176 ) | ( n9538 & n18176 ) ;
  assign n19819 = n17203 ^ n1583 ^ 1'b0 ;
  assign n19820 = n19818 | n19819 ;
  assign n19821 = n19820 ^ n15432 ^ 1'b0 ;
  assign n19822 = ( n1833 & n10545 ) | ( n1833 & n14973 ) | ( n10545 & n14973 ) ;
  assign n19823 = ~n5987 & n16025 ;
  assign n19824 = n19823 ^ n7499 ^ 1'b0 ;
  assign n19825 = n18835 ^ n328 ^ 1'b0 ;
  assign n19826 = n19825 ^ n6493 ^ n1561 ;
  assign n19827 = ( n2018 & ~n4140 ) | ( n2018 & n19826 ) | ( ~n4140 & n19826 ) ;
  assign n19828 = ( n1514 & ~n4623 ) | ( n1514 & n5139 ) | ( ~n4623 & n5139 ) ;
  assign n19829 = x65 & n5233 ;
  assign n19830 = n19829 ^ n8865 ^ n4319 ;
  assign n19831 = n19830 ^ n10190 ^ n1965 ;
  assign n19832 = ( n2303 & n13561 ) | ( n2303 & ~n15093 ) | ( n13561 & ~n15093 ) ;
  assign n19833 = n19832 ^ n15558 ^ n11816 ;
  assign n19834 = n2862 & ~n19833 ;
  assign n19837 = n13654 ^ n9431 ^ n2878 ;
  assign n19835 = n5926 ^ n908 ^ n477 ;
  assign n19836 = ( ~n2133 & n15583 ) | ( ~n2133 & n19835 ) | ( n15583 & n19835 ) ;
  assign n19838 = n19837 ^ n19836 ^ n15255 ;
  assign n19839 = n16844 ^ n8713 ^ 1'b0 ;
  assign n19840 = ( n17696 & ~n19838 ) | ( n17696 & n19839 ) | ( ~n19838 & n19839 ) ;
  assign n19841 = ( n10786 & n15652 ) | ( n10786 & n18928 ) | ( n15652 & n18928 ) ;
  assign n19842 = n16375 ^ n4064 ^ n1714 ;
  assign n19843 = n924 ^ n797 ^ n775 ;
  assign n19844 = n6559 & n19843 ;
  assign n19845 = n19844 ^ n15347 ^ n8229 ;
  assign n19846 = n18062 ^ n15426 ^ n811 ;
  assign n19847 = n14772 ^ n4394 ^ n4177 ;
  assign n19848 = n19847 ^ n14151 ^ n1463 ;
  assign n19849 = ( ~n3922 & n8758 ) | ( ~n3922 & n12956 ) | ( n8758 & n12956 ) ;
  assign n19850 = n3104 ^ n1348 ^ 1'b0 ;
  assign n19851 = n19850 ^ n7008 ^ n1590 ;
  assign n19852 = ( n11500 & n18940 ) | ( n11500 & n19851 ) | ( n18940 & n19851 ) ;
  assign n19853 = ( n530 & n2920 ) | ( n530 & ~n12660 ) | ( n2920 & ~n12660 ) ;
  assign n19854 = n19853 ^ n6845 ^ n6398 ;
  assign n19855 = n13904 ^ n7860 ^ n2820 ;
  assign n19856 = n19855 ^ n12177 ^ n3445 ;
  assign n19857 = ( n3561 & n19854 ) | ( n3561 & n19856 ) | ( n19854 & n19856 ) ;
  assign n19858 = ( n1579 & n4358 ) | ( n1579 & ~n19058 ) | ( n4358 & ~n19058 ) ;
  assign n19859 = ( n1904 & n7186 ) | ( n1904 & n13512 ) | ( n7186 & n13512 ) ;
  assign n19860 = n19859 ^ n15866 ^ n15221 ;
  assign n19861 = ( n3383 & n6645 ) | ( n3383 & n12968 ) | ( n6645 & n12968 ) ;
  assign n19862 = n19502 ^ n16351 ^ n8412 ;
  assign n19863 = ( n863 & ~n3953 ) | ( n863 & n5700 ) | ( ~n3953 & n5700 ) ;
  assign n19864 = n19863 ^ n14418 ^ n11522 ;
  assign n19865 = ( n3920 & n3999 ) | ( n3920 & n7309 ) | ( n3999 & n7309 ) ;
  assign n19866 = ( n7780 & ~n15417 ) | ( n7780 & n19865 ) | ( ~n15417 & n19865 ) ;
  assign n19867 = n15794 ^ n3406 ^ n1933 ;
  assign n19870 = n7302 ^ n3242 ^ n192 ;
  assign n19868 = ( n6283 & n8603 ) | ( n6283 & ~n9396 ) | ( n8603 & ~n9396 ) ;
  assign n19869 = n19868 ^ n13568 ^ n4201 ;
  assign n19871 = n19870 ^ n19869 ^ n6853 ;
  assign n19872 = ~n4406 & n16232 ;
  assign n19874 = ( ~n6390 & n10491 ) | ( ~n6390 & n15192 ) | ( n10491 & n15192 ) ;
  assign n19875 = n19874 ^ n4225 ^ 1'b0 ;
  assign n19876 = n4750 | n19875 ;
  assign n19873 = ( ~n3117 & n10073 ) | ( ~n3117 & n13856 ) | ( n10073 & n13856 ) ;
  assign n19877 = n19876 ^ n19873 ^ n3993 ;
  assign n19879 = ( n2360 & ~n6493 ) | ( n2360 & n18698 ) | ( ~n6493 & n18698 ) ;
  assign n19878 = ~n833 & n9058 ;
  assign n19880 = n19879 ^ n19878 ^ 1'b0 ;
  assign n19881 = ( ~n1634 & n3427 ) | ( ~n1634 & n12008 ) | ( n3427 & n12008 ) ;
  assign n19882 = n10442 ^ n9995 ^ n2359 ;
  assign n19883 = ( ~n257 & n455 ) | ( ~n257 & n19882 ) | ( n455 & n19882 ) ;
  assign n19884 = n8164 ^ n7940 ^ n5012 ;
  assign n19885 = n19884 ^ n6893 ^ n4945 ;
  assign n19886 = n3594 & n6848 ;
  assign n19887 = ~n6653 & n19886 ;
  assign n19888 = n19441 ^ n15926 ^ n702 ;
  assign n19889 = n19888 ^ n10841 ^ n8939 ;
  assign n19890 = ( n8760 & ~n19887 ) | ( n8760 & n19889 ) | ( ~n19887 & n19889 ) ;
  assign n19891 = ( ~n5843 & n8899 ) | ( ~n5843 & n19890 ) | ( n8899 & n19890 ) ;
  assign n19892 = ( n10765 & n19885 ) | ( n10765 & ~n19891 ) | ( n19885 & ~n19891 ) ;
  assign n19893 = n15033 ^ n4039 ^ n1017 ;
  assign n19894 = ~n9698 & n15682 ;
  assign n19895 = n1447 & n19894 ;
  assign n19896 = ( x36 & n13985 ) | ( x36 & n19895 ) | ( n13985 & n19895 ) ;
  assign n19897 = ( n10005 & n19893 ) | ( n10005 & ~n19896 ) | ( n19893 & ~n19896 ) ;
  assign n19898 = ( n3962 & n6666 ) | ( n3962 & n17977 ) | ( n6666 & n17977 ) ;
  assign n19899 = ( x8 & ~n379 ) | ( x8 & n2638 ) | ( ~n379 & n2638 ) ;
  assign n19900 = ( ~n6407 & n6581 ) | ( ~n6407 & n19899 ) | ( n6581 & n19899 ) ;
  assign n19901 = n19900 ^ n930 ^ x42 ;
  assign n19902 = n8017 ^ n6445 ^ 1'b0 ;
  assign n19903 = n1647 & ~n19902 ;
  assign n19904 = ( ~n4124 & n10224 ) | ( ~n4124 & n19903 ) | ( n10224 & n19903 ) ;
  assign n19905 = n17153 ^ n8028 ^ n1280 ;
  assign n19906 = ( n3300 & n5742 ) | ( n3300 & ~n18533 ) | ( n5742 & ~n18533 ) ;
  assign n19907 = n19906 ^ n12841 ^ n252 ;
  assign n19908 = ( n2727 & n11998 ) | ( n2727 & ~n14844 ) | ( n11998 & ~n14844 ) ;
  assign n19909 = n19908 ^ n14468 ^ 1'b0 ;
  assign n19910 = ( n6383 & ~n13244 ) | ( n6383 & n19909 ) | ( ~n13244 & n19909 ) ;
  assign n19911 = ~n4688 & n14161 ;
  assign n19912 = ~n6369 & n19911 ;
  assign n19913 = ( n1158 & n4044 ) | ( n1158 & n6091 ) | ( n4044 & n6091 ) ;
  assign n19914 = n19913 ^ n4996 ^ n3999 ;
  assign n19915 = ~n12572 & n19914 ;
  assign n19916 = ( n4191 & n19912 ) | ( n4191 & ~n19915 ) | ( n19912 & ~n19915 ) ;
  assign n19917 = ( n3128 & ~n4097 ) | ( n3128 & n14936 ) | ( ~n4097 & n14936 ) ;
  assign n19918 = ~n1103 & n19917 ;
  assign n19925 = ( ~n6287 & n10105 ) | ( ~n6287 & n12385 ) | ( n10105 & n12385 ) ;
  assign n19919 = ( n1887 & n9795 ) | ( n1887 & n16855 ) | ( n9795 & n16855 ) ;
  assign n19920 = n13175 ^ n7059 ^ n2255 ;
  assign n19921 = ( x65 & n19919 ) | ( x65 & n19920 ) | ( n19919 & n19920 ) ;
  assign n19922 = ( n2303 & n2798 ) | ( n2303 & n6808 ) | ( n2798 & n6808 ) ;
  assign n19923 = ( n10836 & ~n15940 ) | ( n10836 & n19922 ) | ( ~n15940 & n19922 ) ;
  assign n19924 = ( n17321 & n19921 ) | ( n17321 & n19923 ) | ( n19921 & n19923 ) ;
  assign n19926 = n19925 ^ n19924 ^ n5531 ;
  assign n19927 = n19926 ^ n5126 ^ x121 ;
  assign n19928 = ~n781 & n8838 ;
  assign n19929 = ~n2696 & n19928 ;
  assign n19930 = ( ~n1660 & n9570 ) | ( ~n1660 & n19929 ) | ( n9570 & n19929 ) ;
  assign n19931 = n18295 ^ n7171 ^ 1'b0 ;
  assign n19932 = n19931 ^ n6802 ^ n625 ;
  assign n19933 = n10702 ^ n2765 ^ n1208 ;
  assign n19934 = ( n2305 & ~n12356 ) | ( n2305 & n13384 ) | ( ~n12356 & n13384 ) ;
  assign n19935 = ( n3754 & ~n14448 ) | ( n3754 & n19934 ) | ( ~n14448 & n19934 ) ;
  assign n19936 = ( ~n3447 & n5537 ) | ( ~n3447 & n8438 ) | ( n5537 & n8438 ) ;
  assign n19937 = n19936 ^ n11950 ^ n1010 ;
  assign n19938 = n19937 ^ n17206 ^ n499 ;
  assign n19939 = ( n11185 & n19935 ) | ( n11185 & n19938 ) | ( n19935 & n19938 ) ;
  assign n19940 = ( n4438 & n11666 ) | ( n4438 & n19221 ) | ( n11666 & n19221 ) ;
  assign n19941 = ( n4139 & n19939 ) | ( n4139 & ~n19940 ) | ( n19939 & ~n19940 ) ;
  assign n19942 = ( ~n4869 & n6031 ) | ( ~n4869 & n8943 ) | ( n6031 & n8943 ) ;
  assign n19943 = ( ~n4168 & n4936 ) | ( ~n4168 & n13404 ) | ( n4936 & n13404 ) ;
  assign n19944 = ( n2515 & ~n8613 ) | ( n2515 & n10728 ) | ( ~n8613 & n10728 ) ;
  assign n19945 = n12905 ^ n11194 ^ 1'b0 ;
  assign n19946 = n19944 | n19945 ;
  assign n19947 = ( n11854 & n18913 ) | ( n11854 & ~n19946 ) | ( n18913 & ~n19946 ) ;
  assign n19948 = n19947 ^ n11168 ^ n7384 ;
  assign n19949 = n19948 ^ n12500 ^ n9854 ;
  assign n19950 = n13297 ^ n6506 ^ n1077 ;
  assign n19951 = n13450 & n16569 ;
  assign n19952 = ~n18356 & n19951 ;
  assign n19953 = n19952 ^ n15344 ^ 1'b0 ;
  assign n19954 = ( n4635 & n4902 ) | ( n4635 & n7282 ) | ( n4902 & n7282 ) ;
  assign n19955 = n2645 ^ n2063 ^ n1563 ;
  assign n19956 = n14995 ^ n8222 ^ n3563 ;
  assign n19957 = ( n14083 & n19955 ) | ( n14083 & ~n19956 ) | ( n19955 & ~n19956 ) ;
  assign n19958 = ( n1447 & ~n8060 ) | ( n1447 & n14072 ) | ( ~n8060 & n14072 ) ;
  assign n19959 = n8640 ^ n4559 ^ n370 ;
  assign n19960 = n5429 & n19959 ;
  assign n19961 = ~n19958 & n19960 ;
  assign n19962 = n14506 ^ n2928 ^ 1'b0 ;
  assign n19967 = n12734 ^ n4038 ^ 1'b0 ;
  assign n19968 = ~n3008 & n19967 ;
  assign n19965 = n3120 ^ n1444 ^ n601 ;
  assign n19964 = ( n566 & n2342 ) | ( n566 & n13566 ) | ( n2342 & n13566 ) ;
  assign n19963 = ( n7698 & n8010 ) | ( n7698 & n9193 ) | ( n8010 & n9193 ) ;
  assign n19966 = n19965 ^ n19964 ^ n19963 ;
  assign n19969 = n19968 ^ n19966 ^ n6008 ;
  assign n19970 = n19969 ^ n17067 ^ n13037 ;
  assign n19971 = ( n1297 & n7877 ) | ( n1297 & ~n9236 ) | ( n7877 & ~n9236 ) ;
  assign n19972 = n4686 & ~n7536 ;
  assign n19973 = ~n3485 & n8221 ;
  assign n19974 = ~n4351 & n19973 ;
  assign n19975 = n6140 & n8135 ;
  assign n19976 = n1482 & n19975 ;
  assign n19977 = ( n1995 & ~n5933 ) | ( n1995 & n13534 ) | ( ~n5933 & n13534 ) ;
  assign n19978 = n9947 ^ n8297 ^ n6620 ;
  assign n19979 = ( n1811 & n3510 ) | ( n1811 & n19978 ) | ( n3510 & n19978 ) ;
  assign n19980 = n13340 ^ n5655 ^ n4658 ;
  assign n19981 = n19980 ^ n8018 ^ n7166 ;
  assign n19982 = n1739 | n3391 ;
  assign n19983 = ( ~n389 & n5433 ) | ( ~n389 & n18762 ) | ( n5433 & n18762 ) ;
  assign n19984 = ( n1311 & n14069 ) | ( n1311 & n16866 ) | ( n14069 & n16866 ) ;
  assign n19985 = n10904 & ~n12015 ;
  assign n19986 = n19985 ^ n3036 ^ 1'b0 ;
  assign n19987 = n2648 & n17463 ;
  assign n19988 = n19986 & n19987 ;
  assign n19989 = ( ~n5476 & n5480 ) | ( ~n5476 & n19588 ) | ( n5480 & n19588 ) ;
  assign n19990 = ( n4811 & n18563 ) | ( n4811 & ~n19989 ) | ( n18563 & ~n19989 ) ;
  assign n19991 = ( n2183 & n5228 ) | ( n2183 & ~n19990 ) | ( n5228 & ~n19990 ) ;
  assign n19992 = n14195 ^ n7238 ^ 1'b0 ;
  assign n19993 = ~n15807 & n19992 ;
  assign n19994 = n5860 & n19993 ;
  assign n19995 = ~n19991 & n19994 ;
  assign n19996 = ( n5476 & n13981 ) | ( n5476 & ~n14795 ) | ( n13981 & ~n14795 ) ;
  assign n19997 = n15229 ^ n5298 ^ 1'b0 ;
  assign n19998 = ( ~n3902 & n19996 ) | ( ~n3902 & n19997 ) | ( n19996 & n19997 ) ;
  assign n19999 = ( x10 & ~n3433 ) | ( x10 & n19449 ) | ( ~n3433 & n19449 ) ;
  assign n20000 = ( n888 & n8838 ) | ( n888 & n9552 ) | ( n8838 & n9552 ) ;
  assign n20001 = n10073 ^ n8991 ^ n8364 ;
  assign n20002 = ( ~n14215 & n14550 ) | ( ~n14215 & n20001 ) | ( n14550 & n20001 ) ;
  assign n20003 = ( x29 & n298 ) | ( x29 & ~n2277 ) | ( n298 & ~n2277 ) ;
  assign n20004 = n20003 ^ n8304 ^ 1'b0 ;
  assign n20005 = n20004 ^ n7183 ^ n1308 ;
  assign n20006 = ( ~n17583 & n20002 ) | ( ~n17583 & n20005 ) | ( n20002 & n20005 ) ;
  assign n20007 = n12600 ^ n7529 ^ n7255 ;
  assign n20008 = n20007 ^ n13782 ^ n12072 ;
  assign n20010 = n14379 ^ n4205 ^ n1535 ;
  assign n20009 = ( n5106 & n7029 ) | ( n5106 & n14499 ) | ( n7029 & n14499 ) ;
  assign n20011 = n20010 ^ n20009 ^ 1'b0 ;
  assign n20012 = n15709 & ~n20011 ;
  assign n20013 = n7593 & n16929 ;
  assign n20014 = n10988 & n20013 ;
  assign n20016 = ~n10865 & n11159 ;
  assign n20015 = ~n1663 & n13363 ;
  assign n20017 = n20016 ^ n20015 ^ n9101 ;
  assign n20021 = n1392 & n9391 ;
  assign n20022 = n1830 & n20021 ;
  assign n20023 = ( n13529 & n15705 ) | ( n13529 & ~n20022 ) | ( n15705 & ~n20022 ) ;
  assign n20018 = n12226 ^ n2431 ^ n1395 ;
  assign n20019 = ( ~n3183 & n4153 ) | ( ~n3183 & n20018 ) | ( n4153 & n20018 ) ;
  assign n20020 = n20019 ^ n11908 ^ 1'b0 ;
  assign n20024 = n20023 ^ n20020 ^ 1'b0 ;
  assign n20026 = n3699 | n3807 ;
  assign n20027 = n369 & ~n20026 ;
  assign n20025 = n15776 ^ n1775 ^ n1162 ;
  assign n20028 = n20027 ^ n20025 ^ n12327 ;
  assign n20029 = ( n1705 & ~n8602 ) | ( n1705 & n20028 ) | ( ~n8602 & n20028 ) ;
  assign n20030 = ( n967 & n4581 ) | ( n967 & ~n13193 ) | ( n4581 & ~n13193 ) ;
  assign n20031 = ( n923 & n19540 ) | ( n923 & n20030 ) | ( n19540 & n20030 ) ;
  assign n20032 = ( x63 & n2489 ) | ( x63 & ~n2636 ) | ( n2489 & ~n2636 ) ;
  assign n20033 = n20032 ^ n16462 ^ 1'b0 ;
  assign n20034 = n20033 ^ n13736 ^ n9619 ;
  assign n20035 = ( n6115 & ~n9836 ) | ( n6115 & n20034 ) | ( ~n9836 & n20034 ) ;
  assign n20036 = n16851 ^ n16086 ^ n12421 ;
  assign n20037 = n20036 ^ n15048 ^ n12546 ;
  assign n20045 = n13271 ^ n5462 ^ n2874 ;
  assign n20042 = ~n8943 & n17762 ;
  assign n20043 = ~n2717 & n20042 ;
  assign n20044 = ( ~n7661 & n12758 ) | ( ~n7661 & n20043 ) | ( n12758 & n20043 ) ;
  assign n20038 = n15879 ^ n620 ^ n453 ;
  assign n20039 = n8940 & n18177 ;
  assign n20040 = n20038 & ~n20039 ;
  assign n20041 = ( n904 & n6405 ) | ( n904 & n20040 ) | ( n6405 & n20040 ) ;
  assign n20046 = n20045 ^ n20044 ^ n20041 ;
  assign n20047 = ( n6534 & ~n8801 ) | ( n6534 & n12001 ) | ( ~n8801 & n12001 ) ;
  assign n20048 = ( ~n5895 & n16162 ) | ( ~n5895 & n20047 ) | ( n16162 & n20047 ) ;
  assign n20049 = ( ~n8106 & n11036 ) | ( ~n8106 & n20048 ) | ( n11036 & n20048 ) ;
  assign n20050 = ( ~n5666 & n17717 ) | ( ~n5666 & n20049 ) | ( n17717 & n20049 ) ;
  assign n20051 = n16721 ^ n12126 ^ n2182 ;
  assign n20052 = ( ~n341 & n1383 ) | ( ~n341 & n20051 ) | ( n1383 & n20051 ) ;
  assign n20053 = ( x48 & n8496 ) | ( x48 & n11292 ) | ( n8496 & n11292 ) ;
  assign n20054 = n1802 & n20053 ;
  assign n20055 = n6504 & n20054 ;
  assign n20056 = n9161 ^ n9013 ^ 1'b0 ;
  assign n20057 = n170 & ~n9095 ;
  assign n20058 = ~n516 & n20057 ;
  assign n20059 = ( n3079 & n3231 ) | ( n3079 & n20058 ) | ( n3231 & n20058 ) ;
  assign n20060 = n20059 ^ n17211 ^ n15493 ;
  assign n20061 = ( n4079 & n5977 ) | ( n4079 & n8520 ) | ( n5977 & n8520 ) ;
  assign n20062 = n20061 ^ n17047 ^ n2383 ;
  assign n20063 = n20062 ^ n4637 ^ n4429 ;
  assign n20064 = n5365 ^ n374 ^ n202 ;
  assign n20065 = ( n7925 & n13936 ) | ( n7925 & ~n20064 ) | ( n13936 & ~n20064 ) ;
  assign n20066 = ( n1933 & n2862 ) | ( n1933 & ~n19481 ) | ( n2862 & ~n19481 ) ;
  assign n20067 = n20066 ^ n16988 ^ n679 ;
  assign n20068 = n20067 ^ n3945 ^ 1'b0 ;
  assign n20069 = ( n4413 & ~n9209 ) | ( n4413 & n20068 ) | ( ~n9209 & n20068 ) ;
  assign n20070 = ( n11258 & n13878 ) | ( n11258 & n20069 ) | ( n13878 & n20069 ) ;
  assign n20071 = ( n3931 & n10353 ) | ( n3931 & n14157 ) | ( n10353 & n14157 ) ;
  assign n20072 = ( n8418 & ~n16529 ) | ( n8418 & n19271 ) | ( ~n16529 & n19271 ) ;
  assign n20073 = x97 | n20072 ;
  assign n20074 = ( n1179 & n3447 ) | ( n1179 & ~n16863 ) | ( n3447 & ~n16863 ) ;
  assign n20075 = n18480 ^ n10263 ^ n9957 ;
  assign n20076 = ( n2388 & n18467 ) | ( n2388 & n20075 ) | ( n18467 & n20075 ) ;
  assign n20078 = ( ~n963 & n3767 ) | ( ~n963 & n6329 ) | ( n3767 & n6329 ) ;
  assign n20079 = ( ~n3101 & n17337 ) | ( ~n3101 & n20078 ) | ( n17337 & n20078 ) ;
  assign n20077 = n1102 | n11323 ;
  assign n20080 = n20079 ^ n20077 ^ 1'b0 ;
  assign n20081 = n4060 ^ n2730 ^ n1354 ;
  assign n20082 = n20081 ^ n18473 ^ n10586 ;
  assign n20083 = n20082 ^ n11339 ^ n8254 ;
  assign n20084 = ( ~n1239 & n2240 ) | ( ~n1239 & n10180 ) | ( n2240 & n10180 ) ;
  assign n20085 = ( n2976 & n14733 ) | ( n2976 & n19449 ) | ( n14733 & n19449 ) ;
  assign n20086 = ( n739 & n10934 ) | ( n739 & n16722 ) | ( n10934 & n16722 ) ;
  assign n20087 = ( n20084 & n20085 ) | ( n20084 & n20086 ) | ( n20085 & n20086 ) ;
  assign n20088 = ( n4414 & ~n8591 ) | ( n4414 & n8776 ) | ( ~n8591 & n8776 ) ;
  assign n20089 = ( n9903 & ~n10529 ) | ( n9903 & n20088 ) | ( ~n10529 & n20088 ) ;
  assign n20090 = n20089 ^ n16263 ^ n1365 ;
  assign n20091 = n11804 ^ n10623 ^ n4679 ;
  assign n20092 = n20091 ^ n5284 ^ n1935 ;
  assign n20093 = n7500 ^ n6278 ^ n354 ;
  assign n20094 = n15477 ^ n11048 ^ n2701 ;
  assign n20095 = n17450 ^ n9970 ^ n7877 ;
  assign n20096 = n5013 & ~n20095 ;
  assign n20097 = n20096 ^ n5277 ^ 1'b0 ;
  assign n20098 = n11584 ^ n7469 ^ 1'b0 ;
  assign n20099 = n12211 & n20098 ;
  assign n20100 = n6112 ^ n2664 ^ n1991 ;
  assign n20108 = ( n1141 & ~n5776 ) | ( n1141 & n10388 ) | ( ~n5776 & n10388 ) ;
  assign n20105 = ( n3334 & ~n7478 ) | ( n3334 & n9671 ) | ( ~n7478 & n9671 ) ;
  assign n20106 = ( n4931 & n5614 ) | ( n4931 & ~n20105 ) | ( n5614 & ~n20105 ) ;
  assign n20102 = ( ~n2642 & n3771 ) | ( ~n2642 & n6544 ) | ( n3771 & n6544 ) ;
  assign n20103 = ( n1971 & n9836 ) | ( n1971 & n20102 ) | ( n9836 & n20102 ) ;
  assign n20101 = n2788 | n8041 ;
  assign n20104 = n20103 ^ n20101 ^ 1'b0 ;
  assign n20107 = n20106 ^ n20104 ^ n5904 ;
  assign n20109 = n20108 ^ n20107 ^ n994 ;
  assign n20110 = n15268 ^ n14205 ^ n5492 ;
  assign n20111 = n387 | n4350 ;
  assign n20112 = n5898 ^ n3940 ^ n2447 ;
  assign n20113 = ( n3795 & n3889 ) | ( n3795 & ~n7148 ) | ( n3889 & ~n7148 ) ;
  assign n20114 = ( n3094 & ~n6922 ) | ( n3094 & n20113 ) | ( ~n6922 & n20113 ) ;
  assign n20115 = n20112 | n20114 ;
  assign n20116 = n20115 ^ n12569 ^ n3491 ;
  assign n20117 = n6797 & n10072 ;
  assign n20118 = n14567 & n20117 ;
  assign n20119 = n8781 & ~n15263 ;
  assign n20120 = n11377 & n20119 ;
  assign n20121 = n6658 | n20120 ;
  assign n20122 = n9244 ^ n6215 ^ n4029 ;
  assign n20123 = ( n2624 & ~n11038 ) | ( n2624 & n19163 ) | ( ~n11038 & n19163 ) ;
  assign n20124 = ( n5923 & n8728 ) | ( n5923 & n10714 ) | ( n8728 & n10714 ) ;
  assign n20125 = n20124 ^ n7030 ^ 1'b0 ;
  assign n20126 = n20125 ^ n16781 ^ n15266 ;
  assign n20127 = n7093 & n17540 ;
  assign n20128 = ( n6259 & ~n12864 ) | ( n6259 & n20127 ) | ( ~n12864 & n20127 ) ;
  assign n20129 = n11783 & n12177 ;
  assign n20130 = n18910 ^ n4241 ^ 1'b0 ;
  assign n20131 = n20130 ^ n6520 ^ 1'b0 ;
  assign n20132 = n18227 & ~n20131 ;
  assign n20133 = n20132 ^ n7853 ^ n746 ;
  assign n20134 = ( n3013 & n4461 ) | ( n3013 & ~n18622 ) | ( n4461 & ~n18622 ) ;
  assign n20137 = n6501 ^ n3042 ^ 1'b0 ;
  assign n20138 = n12513 & ~n20137 ;
  assign n20139 = n20138 ^ n6424 ^ 1'b0 ;
  assign n20135 = ( n3365 & ~n3456 ) | ( n3365 & n5484 ) | ( ~n3456 & n5484 ) ;
  assign n20136 = n20135 ^ n8280 ^ n1887 ;
  assign n20140 = n20139 ^ n20136 ^ n15919 ;
  assign n20141 = n19923 ^ n15684 ^ n8644 ;
  assign n20142 = n5368 & ~n19241 ;
  assign n20143 = ( n7365 & ~n7563 ) | ( n7365 & n7759 ) | ( ~n7563 & n7759 ) ;
  assign n20144 = n17271 ^ n14896 ^ n12386 ;
  assign n20145 = n13235 ^ n7583 ^ 1'b0 ;
  assign n20146 = n5897 | n14996 ;
  assign n20147 = n20146 ^ n6966 ^ 1'b0 ;
  assign n20148 = ( n1191 & ~n20145 ) | ( n1191 & n20147 ) | ( ~n20145 & n20147 ) ;
  assign n20149 = ( n4551 & ~n8803 ) | ( n4551 & n20148 ) | ( ~n8803 & n20148 ) ;
  assign n20150 = ( ~n12489 & n14295 ) | ( ~n12489 & n15033 ) | ( n14295 & n15033 ) ;
  assign n20151 = n752 & n14638 ;
  assign n20152 = ( n7880 & ~n10349 ) | ( n7880 & n20151 ) | ( ~n10349 & n20151 ) ;
  assign n20153 = n15208 | n20152 ;
  assign n20154 = ( ~n19497 & n20150 ) | ( ~n19497 & n20153 ) | ( n20150 & n20153 ) ;
  assign n20155 = ( n1251 & n9706 ) | ( n1251 & ~n13583 ) | ( n9706 & ~n13583 ) ;
  assign n20156 = n9801 ^ n8469 ^ n4546 ;
  assign n20157 = ( ~n6562 & n8446 ) | ( ~n6562 & n20156 ) | ( n8446 & n20156 ) ;
  assign n20158 = ( ~n8317 & n9121 ) | ( ~n8317 & n20157 ) | ( n9121 & n20157 ) ;
  assign n20159 = n1942 | n16904 ;
  assign n20160 = ( n6612 & n17330 ) | ( n6612 & n20159 ) | ( n17330 & n20159 ) ;
  assign n20161 = n20158 & ~n20160 ;
  assign n20162 = n15997 ^ n11645 ^ n1580 ;
  assign n20163 = ( n421 & ~n5970 ) | ( n421 & n11971 ) | ( ~n5970 & n11971 ) ;
  assign n20164 = n20163 ^ n11082 ^ n8352 ;
  assign n20165 = ( n10457 & ~n20162 ) | ( n10457 & n20164 ) | ( ~n20162 & n20164 ) ;
  assign n20166 = n5245 ^ n4577 ^ n1260 ;
  assign n20167 = n20166 ^ n12981 ^ n7502 ;
  assign n20168 = n20167 ^ n10150 ^ 1'b0 ;
  assign n20169 = n5937 & ~n20168 ;
  assign n20170 = ( n4319 & n15426 ) | ( n4319 & n20169 ) | ( n15426 & n20169 ) ;
  assign n20171 = n11225 & n15672 ;
  assign n20172 = n20171 ^ n3517 ^ n363 ;
  assign n20173 = n14071 ^ n3274 ^ n1637 ;
  assign n20174 = n8518 ^ n8139 ^ n5487 ;
  assign n20175 = n14790 ^ n10125 ^ n1246 ;
  assign n20178 = n5084 ^ n2149 ^ n340 ;
  assign n20179 = ( n5780 & ~n8325 ) | ( n5780 & n20178 ) | ( ~n8325 & n20178 ) ;
  assign n20176 = n2010 | n3973 ;
  assign n20177 = n20176 ^ n17732 ^ 1'b0 ;
  assign n20180 = n20179 ^ n20177 ^ n19884 ;
  assign n20181 = n2632 | n10102 ;
  assign n20182 = n7357 & ~n20181 ;
  assign n20183 = n11027 ^ n6398 ^ n3847 ;
  assign n20184 = n20183 ^ n11259 ^ n1491 ;
  assign n20185 = ( ~n5719 & n10275 ) | ( ~n5719 & n11130 ) | ( n10275 & n11130 ) ;
  assign n20186 = ( ~n17443 & n18302 ) | ( ~n17443 & n20185 ) | ( n18302 & n20185 ) ;
  assign n20189 = n6179 ^ n2082 ^ 1'b0 ;
  assign n20187 = ( n209 & ~n2623 ) | ( n209 & n5709 ) | ( ~n2623 & n5709 ) ;
  assign n20188 = ~n16653 & n20187 ;
  assign n20190 = n20189 ^ n20188 ^ 1'b0 ;
  assign n20191 = ( n7574 & n12605 ) | ( n7574 & ~n20190 ) | ( n12605 & ~n20190 ) ;
  assign n20192 = ( ~n3684 & n19374 ) | ( ~n3684 & n20191 ) | ( n19374 & n20191 ) ;
  assign n20193 = n20192 ^ n19761 ^ n1585 ;
  assign n20194 = n4240 ^ n3884 ^ n1716 ;
  assign n20195 = n20194 ^ n11156 ^ n9706 ;
  assign n20196 = n9573 ^ n7080 ^ n5483 ;
  assign n20197 = n16783 ^ n8932 ^ x47 ;
  assign n20198 = ( n6489 & n11054 ) | ( n6489 & n20197 ) | ( n11054 & n20197 ) ;
  assign n20199 = ( n13650 & ~n20196 ) | ( n13650 & n20198 ) | ( ~n20196 & n20198 ) ;
  assign n20200 = n7538 ^ n4788 ^ 1'b0 ;
  assign n20201 = n9481 & n20200 ;
  assign n20202 = n20201 ^ n18191 ^ n13134 ;
  assign n20203 = n7563 ^ n3425 ^ 1'b0 ;
  assign n20204 = n3176 | n20203 ;
  assign n20208 = ( n2204 & n2753 ) | ( n2204 & ~n5704 ) | ( n2753 & ~n5704 ) ;
  assign n20207 = n19198 ^ n12440 ^ x75 ;
  assign n20205 = n9563 | n13283 ;
  assign n20206 = ( n11055 & n19399 ) | ( n11055 & n20205 ) | ( n19399 & n20205 ) ;
  assign n20209 = n20208 ^ n20207 ^ n20206 ;
  assign n20210 = ( n3199 & ~n14665 ) | ( n3199 & n20209 ) | ( ~n14665 & n20209 ) ;
  assign n20211 = n18729 & ~n20210 ;
  assign n20212 = n5109 ^ n2114 ^ n582 ;
  assign n20213 = ( n8816 & n14596 ) | ( n8816 & n16160 ) | ( n14596 & n16160 ) ;
  assign n20214 = ( ~n6487 & n7341 ) | ( ~n6487 & n20213 ) | ( n7341 & n20213 ) ;
  assign n20215 = ( n18736 & n20212 ) | ( n18736 & ~n20214 ) | ( n20212 & ~n20214 ) ;
  assign n20216 = ( n848 & n6727 ) | ( n848 & n10083 ) | ( n6727 & n10083 ) ;
  assign n20217 = n4713 ^ n3717 ^ 1'b0 ;
  assign n20218 = ( n3870 & ~n8151 ) | ( n3870 & n20217 ) | ( ~n8151 & n20217 ) ;
  assign n20219 = n20218 ^ n8707 ^ n4599 ;
  assign n20220 = ( ~n1438 & n2637 ) | ( ~n1438 & n20219 ) | ( n2637 & n20219 ) ;
  assign n20221 = ( n11235 & n20216 ) | ( n11235 & n20220 ) | ( n20216 & n20220 ) ;
  assign n20222 = ( ~n629 & n4359 ) | ( ~n629 & n9375 ) | ( n4359 & n9375 ) ;
  assign n20223 = ( n4504 & n7635 ) | ( n4504 & n17543 ) | ( n7635 & n17543 ) ;
  assign n20227 = ( x40 & n164 ) | ( x40 & n1097 ) | ( n164 & n1097 ) ;
  assign n20224 = n10175 ^ n9174 ^ n6480 ;
  assign n20225 = ( n4528 & ~n6489 ) | ( n4528 & n20224 ) | ( ~n6489 & n20224 ) ;
  assign n20226 = ( n6840 & n10042 ) | ( n6840 & ~n20225 ) | ( n10042 & ~n20225 ) ;
  assign n20228 = n20227 ^ n20226 ^ n18280 ;
  assign n20230 = n3749 ^ n2051 ^ 1'b0 ;
  assign n20231 = n363 | n20230 ;
  assign n20232 = ( n1451 & n11494 ) | ( n1451 & n20231 ) | ( n11494 & n20231 ) ;
  assign n20229 = ( ~n12163 & n13111 ) | ( ~n12163 & n16133 ) | ( n13111 & n16133 ) ;
  assign n20233 = n20232 ^ n20229 ^ n17871 ;
  assign n20234 = n20233 ^ n14503 ^ n3287 ;
  assign n20235 = ( n1233 & n4569 ) | ( n1233 & ~n8750 ) | ( n4569 & ~n8750 ) ;
  assign n20236 = n10458 & n20235 ;
  assign n20237 = ~n20234 & n20236 ;
  assign n20238 = n7219 ^ n2383 ^ n1097 ;
  assign n20239 = n19843 ^ n7963 ^ x16 ;
  assign n20240 = n20239 ^ n7174 ^ n637 ;
  assign n20241 = ( ~n18503 & n20238 ) | ( ~n18503 & n20240 ) | ( n20238 & n20240 ) ;
  assign n20242 = ( ~n1046 & n1463 ) | ( ~n1046 & n2439 ) | ( n1463 & n2439 ) ;
  assign n20243 = ( n350 & n8852 ) | ( n350 & n10940 ) | ( n8852 & n10940 ) ;
  assign n20246 = ( ~n12184 & n12347 ) | ( ~n12184 & n18380 ) | ( n12347 & n18380 ) ;
  assign n20244 = ( ~n187 & n6120 ) | ( ~n187 & n17605 ) | ( n6120 & n17605 ) ;
  assign n20245 = ( n1404 & n4470 ) | ( n1404 & n20244 ) | ( n4470 & n20244 ) ;
  assign n20247 = n20246 ^ n20245 ^ n4602 ;
  assign n20248 = ( n3204 & n6299 ) | ( n3204 & n10010 ) | ( n6299 & n10010 ) ;
  assign n20249 = ( n2118 & n5823 ) | ( n2118 & n20248 ) | ( n5823 & n20248 ) ;
  assign n20250 = ( n523 & ~n3912 ) | ( n523 & n9922 ) | ( ~n3912 & n9922 ) ;
  assign n20251 = ( n1533 & n9329 ) | ( n1533 & n20250 ) | ( n9329 & n20250 ) ;
  assign n20252 = n2388 & ~n3395 ;
  assign n20253 = n20252 ^ n1391 ^ 1'b0 ;
  assign n20254 = n20253 ^ n8300 ^ n6702 ;
  assign n20255 = ( n190 & ~n14045 ) | ( n190 & n17112 ) | ( ~n14045 & n17112 ) ;
  assign n20256 = ( ~n20251 & n20254 ) | ( ~n20251 & n20255 ) | ( n20254 & n20255 ) ;
  assign n20257 = ~n13584 & n20256 ;
  assign n20258 = ( n4244 & n15024 ) | ( n4244 & ~n17061 ) | ( n15024 & ~n17061 ) ;
  assign n20259 = n2985 & ~n20258 ;
  assign n20260 = ( n1655 & n5362 ) | ( n1655 & n7893 ) | ( n5362 & n7893 ) ;
  assign n20261 = n12636 & n20260 ;
  assign n20262 = n20261 ^ n2678 ^ 1'b0 ;
  assign n20263 = ( ~n1241 & n7714 ) | ( ~n1241 & n20262 ) | ( n7714 & n20262 ) ;
  assign n20264 = n18002 ^ n13748 ^ n12908 ;
  assign n20265 = ( n7144 & ~n14071 ) | ( n7144 & n15952 ) | ( ~n14071 & n15952 ) ;
  assign n20266 = n20265 ^ n15069 ^ n6236 ;
  assign n20267 = ( n7474 & ~n12523 ) | ( n7474 & n20062 ) | ( ~n12523 & n20062 ) ;
  assign n20268 = n6433 & n12893 ;
  assign n20269 = n20268 ^ n13592 ^ 1'b0 ;
  assign n20270 = ~n6278 & n20269 ;
  assign n20271 = n5733 & ~n11981 ;
  assign n20277 = n9977 ^ n7550 ^ 1'b0 ;
  assign n20276 = ( n4233 & n8890 ) | ( n4233 & n9563 ) | ( n8890 & n9563 ) ;
  assign n20272 = ( ~n3796 & n6823 ) | ( ~n3796 & n11165 ) | ( n6823 & n11165 ) ;
  assign n20273 = ( n5591 & n12614 ) | ( n5591 & n20272 ) | ( n12614 & n20272 ) ;
  assign n20274 = ~n8508 & n14183 ;
  assign n20275 = ~n20273 & n20274 ;
  assign n20278 = n20277 ^ n20276 ^ n20275 ;
  assign n20279 = ( x118 & ~n3305 ) | ( x118 & n14523 ) | ( ~n3305 & n14523 ) ;
  assign n20280 = n20279 ^ n3488 ^ n1100 ;
  assign n20281 = n19870 ^ n15585 ^ n4555 ;
  assign n20282 = ( n8106 & n11035 ) | ( n8106 & ~n20281 ) | ( n11035 & ~n20281 ) ;
  assign n20285 = ( n3013 & n9836 ) | ( n3013 & ~n17542 ) | ( n9836 & ~n17542 ) ;
  assign n20284 = ( ~n2870 & n10585 ) | ( ~n2870 & n15103 ) | ( n10585 & n15103 ) ;
  assign n20283 = n14688 ^ n6029 ^ n4468 ;
  assign n20286 = n20285 ^ n20284 ^ n20283 ;
  assign n20287 = n16969 ^ n8165 ^ n423 ;
  assign n20289 = ( ~n4886 & n6008 ) | ( ~n4886 & n8528 ) | ( n6008 & n8528 ) ;
  assign n20288 = n11969 ^ n10046 ^ n7571 ;
  assign n20290 = n20289 ^ n20288 ^ 1'b0 ;
  assign n20296 = ( n5666 & n7388 ) | ( n5666 & n8425 ) | ( n7388 & n8425 ) ;
  assign n20293 = ~n6467 & n11895 ;
  assign n20294 = n3229 & n20293 ;
  assign n20295 = ( n2395 & n3987 ) | ( n2395 & ~n20294 ) | ( n3987 & ~n20294 ) ;
  assign n20291 = n9005 ^ n8259 ^ n3378 ;
  assign n20292 = n20291 ^ n17551 ^ n11277 ;
  assign n20297 = n20296 ^ n20295 ^ n20292 ;
  assign n20298 = ( n8821 & ~n11279 ) | ( n8821 & n15821 ) | ( ~n11279 & n15821 ) ;
  assign n20299 = n20298 ^ n16375 ^ n14194 ;
  assign n20300 = ~n280 & n17934 ;
  assign n20301 = n20300 ^ n15419 ^ 1'b0 ;
  assign n20302 = ( n8816 & n9479 ) | ( n8816 & n20301 ) | ( n9479 & n20301 ) ;
  assign n20303 = ( n1031 & n14103 ) | ( n1031 & n20302 ) | ( n14103 & n20302 ) ;
  assign n20304 = n6802 & ~n15864 ;
  assign n20305 = n20304 ^ n3510 ^ 1'b0 ;
  assign n20306 = ( n3940 & n9061 ) | ( n3940 & ~n16261 ) | ( n9061 & ~n16261 ) ;
  assign n20307 = ( n8612 & n13367 ) | ( n8612 & ~n20233 ) | ( n13367 & ~n20233 ) ;
  assign n20308 = ( n7321 & n20306 ) | ( n7321 & ~n20307 ) | ( n20306 & ~n20307 ) ;
  assign n20309 = ( n4708 & n20305 ) | ( n4708 & ~n20308 ) | ( n20305 & ~n20308 ) ;
  assign n20310 = ( ~n647 & n5417 ) | ( ~n647 & n7931 ) | ( n5417 & n7931 ) ;
  assign n20311 = n20310 ^ n14225 ^ n1954 ;
  assign n20312 = n15689 ^ n7792 ^ 1'b0 ;
  assign n20313 = n4460 & n20312 ;
  assign n20314 = ( n421 & n11733 ) | ( n421 & ~n20313 ) | ( n11733 & ~n20313 ) ;
  assign n20315 = n8895 ^ n8816 ^ n7537 ;
  assign n20316 = n129 & ~n3804 ;
  assign n20317 = n20315 & n20316 ;
  assign n20318 = n20317 ^ n9709 ^ n4096 ;
  assign n20319 = x81 & n13021 ;
  assign n20320 = n14273 & n20319 ;
  assign n20321 = n3588 | n10495 ;
  assign n20322 = ( ~n681 & n1809 ) | ( ~n681 & n19123 ) | ( n1809 & n19123 ) ;
  assign n20323 = n20322 ^ n17886 ^ n1645 ;
  assign n20324 = n3259 & ~n4158 ;
  assign n20325 = n12365 ^ n9053 ^ x78 ;
  assign n20326 = n9211 ^ n2749 ^ 1'b0 ;
  assign n20327 = n7557 & n20326 ;
  assign n20328 = n20327 ^ n10941 ^ n6796 ;
  assign n20329 = n20328 ^ n12241 ^ n12061 ;
  assign n20330 = ( ~n7668 & n15708 ) | ( ~n7668 & n18825 ) | ( n15708 & n18825 ) ;
  assign n20331 = ( ~n5700 & n11565 ) | ( ~n5700 & n20330 ) | ( n11565 & n20330 ) ;
  assign n20332 = n9431 ^ n8228 ^ n6677 ;
  assign n20333 = n13730 ^ n8828 ^ n2813 ;
  assign n20334 = n20333 ^ n16402 ^ n982 ;
  assign n20335 = ( ~n1917 & n5128 ) | ( ~n1917 & n20334 ) | ( n5128 & n20334 ) ;
  assign n20337 = ( ~n321 & n4347 ) | ( ~n321 & n6932 ) | ( n4347 & n6932 ) ;
  assign n20336 = n12170 | n16607 ;
  assign n20338 = n20337 ^ n20336 ^ n8398 ;
  assign n20339 = ( n4091 & n6238 ) | ( n4091 & n17565 ) | ( n6238 & n17565 ) ;
  assign n20340 = n18883 ^ n7942 ^ n3417 ;
  assign n20341 = ( ~n8719 & n9970 ) | ( ~n8719 & n20340 ) | ( n9970 & n20340 ) ;
  assign n20347 = ( ~n2149 & n6121 ) | ( ~n2149 & n10156 ) | ( n6121 & n10156 ) ;
  assign n20348 = ( n237 & n3356 ) | ( n237 & n20347 ) | ( n3356 & n20347 ) ;
  assign n20343 = ( ~x1 & n134 ) | ( ~x1 & n17243 ) | ( n134 & n17243 ) ;
  assign n20344 = ( n1896 & ~n5079 ) | ( n1896 & n20343 ) | ( ~n5079 & n20343 ) ;
  assign n20342 = ( n10074 & n10434 ) | ( n10074 & n11533 ) | ( n10434 & n11533 ) ;
  assign n20345 = n20344 ^ n20342 ^ n1074 ;
  assign n20346 = n19597 & n20345 ;
  assign n20349 = n20348 ^ n20346 ^ 1'b0 ;
  assign n20350 = n6086 ^ n4737 ^ n194 ;
  assign n20351 = n20350 ^ n12323 ^ n8233 ;
  assign n20352 = ( ~n229 & n1463 ) | ( ~n229 & n9042 ) | ( n1463 & n9042 ) ;
  assign n20353 = n10443 ^ n9549 ^ n492 ;
  assign n20354 = ( ~n12406 & n13406 ) | ( ~n12406 & n19685 ) | ( n13406 & n19685 ) ;
  assign n20355 = n20354 ^ n7284 ^ n3586 ;
  assign n20356 = ( n20352 & ~n20353 ) | ( n20352 & n20355 ) | ( ~n20353 & n20355 ) ;
  assign n20357 = ( n5611 & n7380 ) | ( n5611 & ~n7773 ) | ( n7380 & ~n7773 ) ;
  assign n20358 = ( n2665 & n10109 ) | ( n2665 & n20357 ) | ( n10109 & n20357 ) ;
  assign n20359 = n20358 ^ n12290 ^ n3175 ;
  assign n20360 = n20359 ^ n11063 ^ n1445 ;
  assign n20361 = n9185 & ~n19237 ;
  assign n20363 = ( n5036 & n6099 ) | ( n5036 & ~n18125 ) | ( n6099 & ~n18125 ) ;
  assign n20362 = n8582 ^ n914 ^ 1'b0 ;
  assign n20364 = n20363 ^ n20362 ^ n385 ;
  assign n20365 = n14954 ^ n5696 ^ n1052 ;
  assign n20366 = n6489 & n20365 ;
  assign n20367 = n10010 ^ n9905 ^ n6567 ;
  assign n20368 = n20367 ^ n12251 ^ n9424 ;
  assign n20369 = n18857 ^ n13928 ^ n10364 ;
  assign n20370 = ( n3424 & n4175 ) | ( n3424 & ~n13208 ) | ( n4175 & ~n13208 ) ;
  assign n20371 = ( n460 & ~n4530 ) | ( n460 & n13458 ) | ( ~n4530 & n13458 ) ;
  assign n20372 = n1707 & ~n3993 ;
  assign n20373 = ( n2291 & n12511 ) | ( n2291 & n20372 ) | ( n12511 & n20372 ) ;
  assign n20374 = ( n5396 & n11153 ) | ( n5396 & n20373 ) | ( n11153 & n20373 ) ;
  assign n20375 = n15077 ^ n3359 ^ 1'b0 ;
  assign n20376 = n3290 & ~n3643 ;
  assign n20377 = n16922 & n20376 ;
  assign n20384 = ~n2518 & n9745 ;
  assign n20385 = n20384 ^ n2997 ^ 1'b0 ;
  assign n20383 = n9866 ^ n7738 ^ n6704 ;
  assign n20386 = n20385 ^ n20383 ^ 1'b0 ;
  assign n20378 = n10266 ^ n4032 ^ 1'b0 ;
  assign n20379 = n16611 | n20378 ;
  assign n20380 = n20379 ^ n17284 ^ n7366 ;
  assign n20381 = n20380 ^ n4358 ^ n3571 ;
  assign n20382 = n5468 | n20381 ;
  assign n20387 = n20386 ^ n20382 ^ 1'b0 ;
  assign n20388 = n12267 ^ n6756 ^ n4622 ;
  assign n20389 = n14653 ^ n13217 ^ n12851 ;
  assign n20390 = n20389 ^ n15669 ^ n1827 ;
  assign n20391 = ( ~n4339 & n5637 ) | ( ~n4339 & n7725 ) | ( n5637 & n7725 ) ;
  assign n20392 = ( n1157 & n11058 ) | ( n1157 & ~n20391 ) | ( n11058 & ~n20391 ) ;
  assign n20393 = ( n7477 & n16431 ) | ( n7477 & n20392 ) | ( n16431 & n20392 ) ;
  assign n20394 = ( n20388 & n20390 ) | ( n20388 & n20393 ) | ( n20390 & n20393 ) ;
  assign n20395 = n17796 ^ n5092 ^ n4858 ;
  assign n20396 = n8687 ^ n5644 ^ n3124 ;
  assign n20397 = ( x39 & n7178 ) | ( x39 & n17291 ) | ( n7178 & n17291 ) ;
  assign n20398 = ( n18748 & n20396 ) | ( n18748 & ~n20397 ) | ( n20396 & ~n20397 ) ;
  assign n20399 = ( n4216 & n20395 ) | ( n4216 & n20398 ) | ( n20395 & n20398 ) ;
  assign n20400 = n19772 ^ n16732 ^ n13376 ;
  assign n20401 = ( n3289 & n8151 ) | ( n3289 & n20400 ) | ( n8151 & n20400 ) ;
  assign n20402 = ( n6242 & n18895 ) | ( n6242 & ~n20401 ) | ( n18895 & ~n20401 ) ;
  assign n20403 = ( n1434 & n11671 ) | ( n1434 & ~n20402 ) | ( n11671 & ~n20402 ) ;
  assign n20404 = ~n14692 & n18796 ;
  assign n20405 = ( n343 & n788 ) | ( n343 & ~n6042 ) | ( n788 & ~n6042 ) ;
  assign n20406 = ( ~n8040 & n9895 ) | ( ~n8040 & n12867 ) | ( n9895 & n12867 ) ;
  assign n20407 = ( n12812 & n20405 ) | ( n12812 & n20406 ) | ( n20405 & n20406 ) ;
  assign n20408 = n18249 ^ n15424 ^ n11548 ;
  assign n20409 = n9413 ^ n4566 ^ n4168 ;
  assign n20410 = n20409 ^ n5363 ^ 1'b0 ;
  assign n20411 = ( n5549 & n9058 ) | ( n5549 & n20410 ) | ( n9058 & n20410 ) ;
  assign n20412 = n12743 ^ n9991 ^ n2277 ;
  assign n20413 = n3594 ^ n2141 ^ 1'b0 ;
  assign n20414 = n20413 ^ n7037 ^ 1'b0 ;
  assign n20415 = n20412 & ~n20414 ;
  assign n20416 = ( n8023 & n9717 ) | ( n8023 & n20415 ) | ( n9717 & n20415 ) ;
  assign n20417 = n19740 ^ n15436 ^ 1'b0 ;
  assign n20418 = n7565 | n20417 ;
  assign n20419 = n20418 ^ n16849 ^ n6481 ;
  assign n20420 = ( n3429 & n4896 ) | ( n3429 & n20419 ) | ( n4896 & n20419 ) ;
  assign n20424 = n9096 ^ n8421 ^ 1'b0 ;
  assign n20425 = n7407 & ~n20424 ;
  assign n20421 = n9263 ^ n3904 ^ n2933 ;
  assign n20422 = ( n3971 & n10981 ) | ( n3971 & n20421 ) | ( n10981 & n20421 ) ;
  assign n20423 = n20422 ^ n19441 ^ n2174 ;
  assign n20426 = n20425 ^ n20423 ^ n9228 ;
  assign n20427 = ( x32 & n9675 ) | ( x32 & ~n20426 ) | ( n9675 & ~n20426 ) ;
  assign n20428 = ( n881 & n1187 ) | ( n881 & ~n9183 ) | ( n1187 & ~n9183 ) ;
  assign n20429 = ( ~n2426 & n13177 ) | ( ~n2426 & n20428 ) | ( n13177 & n20428 ) ;
  assign n20430 = n15853 ^ n4172 ^ n2420 ;
  assign n20431 = n6077 ^ n1366 ^ n827 ;
  assign n20432 = n20431 ^ n10371 ^ n8848 ;
  assign n20433 = n4022 & ~n20432 ;
  assign n20434 = n20433 ^ n1879 ^ 1'b0 ;
  assign n20435 = ( n3554 & n5816 ) | ( n3554 & n5922 ) | ( n5816 & n5922 ) ;
  assign n20436 = ( n5575 & ~n12511 ) | ( n5575 & n20435 ) | ( ~n12511 & n20435 ) ;
  assign n20437 = n20436 ^ n9938 ^ n1013 ;
  assign n20438 = ( n5262 & n9780 ) | ( n5262 & ~n13531 ) | ( n9780 & ~n13531 ) ;
  assign n20439 = ( n2645 & n10546 ) | ( n2645 & n14688 ) | ( n10546 & n14688 ) ;
  assign n20440 = ( n433 & n20438 ) | ( n433 & ~n20439 ) | ( n20438 & ~n20439 ) ;
  assign n20441 = ( n1456 & n7578 ) | ( n1456 & n9933 ) | ( n7578 & n9933 ) ;
  assign n20442 = ( n12191 & n14969 ) | ( n12191 & n20441 ) | ( n14969 & n20441 ) ;
  assign n20443 = n4206 ^ n2428 ^ n417 ;
  assign n20444 = ( ~n6255 & n11035 ) | ( ~n6255 & n20443 ) | ( n11035 & n20443 ) ;
  assign n20445 = ( ~n11467 & n20442 ) | ( ~n11467 & n20444 ) | ( n20442 & n20444 ) ;
  assign n20446 = ( n9178 & ~n17502 ) | ( n9178 & n18828 ) | ( ~n17502 & n18828 ) ;
  assign n20447 = n9184 ^ n273 ^ 1'b0 ;
  assign n20448 = ( n6741 & ~n11446 ) | ( n6741 & n20447 ) | ( ~n11446 & n20447 ) ;
  assign n20449 = n11805 ^ n2659 ^ 1'b0 ;
  assign n20450 = n20449 ^ n3190 ^ n2778 ;
  assign n20453 = n5169 ^ n4862 ^ n3416 ;
  assign n20451 = n9386 ^ n1906 ^ 1'b0 ;
  assign n20452 = n20451 ^ n6267 ^ n3102 ;
  assign n20454 = n20453 ^ n20452 ^ n14632 ;
  assign n20455 = n8383 ^ n5544 ^ n2618 ;
  assign n20456 = ( n4334 & ~n12462 ) | ( n4334 & n18936 ) | ( ~n12462 & n18936 ) ;
  assign n20457 = n20456 ^ n6444 ^ 1'b0 ;
  assign n20458 = n5158 ^ n4249 ^ n2921 ;
  assign n20459 = ( ~n20455 & n20457 ) | ( ~n20455 & n20458 ) | ( n20457 & n20458 ) ;
  assign n20460 = n14335 ^ n4440 ^ n4145 ;
  assign n20461 = ( n8548 & ~n15559 ) | ( n8548 & n20460 ) | ( ~n15559 & n20460 ) ;
  assign n20462 = n18971 ^ n13432 ^ n3810 ;
  assign n20463 = n18014 & n18296 ;
  assign n20464 = ~n20462 & n20463 ;
  assign n20469 = n1497 & n14765 ;
  assign n20470 = n20469 ^ n19481 ^ 1'b0 ;
  assign n20468 = n11546 ^ n8815 ^ 1'b0 ;
  assign n20465 = n16475 ^ n4364 ^ n1878 ;
  assign n20466 = ( x39 & n12569 ) | ( x39 & ~n20465 ) | ( n12569 & ~n20465 ) ;
  assign n20467 = n16458 & n20466 ;
  assign n20471 = n20470 ^ n20468 ^ n20467 ;
  assign n20472 = ( n2478 & n15022 ) | ( n2478 & ~n17928 ) | ( n15022 & ~n17928 ) ;
  assign n20473 = n20010 ^ n16561 ^ n2140 ;
  assign n20474 = n540 & ~n3260 ;
  assign n20475 = n20474 ^ n10003 ^ 1'b0 ;
  assign n20476 = n6282 & ~n18100 ;
  assign n20477 = n20476 ^ n1865 ^ 1'b0 ;
  assign n20478 = ( ~n4755 & n9127 ) | ( ~n4755 & n20477 ) | ( n9127 & n20477 ) ;
  assign n20479 = n20475 | n20478 ;
  assign n20480 = n9225 ^ n8355 ^ n3604 ;
  assign n20481 = n16557 ^ n15621 ^ n6220 ;
  assign n20482 = n12267 ^ n6450 ^ 1'b0 ;
  assign n20483 = n20482 ^ n4120 ^ 1'b0 ;
  assign n20484 = ( ~n1972 & n10639 ) | ( ~n1972 & n20483 ) | ( n10639 & n20483 ) ;
  assign n20485 = ( n5065 & ~n9357 ) | ( n5065 & n11529 ) | ( ~n9357 & n11529 ) ;
  assign n20486 = n20485 ^ n9575 ^ 1'b0 ;
  assign n20487 = n20484 | n20486 ;
  assign n20488 = ( n1898 & n4550 ) | ( n1898 & ~n12466 ) | ( n4550 & ~n12466 ) ;
  assign n20492 = ( n2481 & n9324 ) | ( n2481 & ~n13297 ) | ( n9324 & ~n13297 ) ;
  assign n20489 = n17574 ^ n5899 ^ n4415 ;
  assign n20490 = ~n9748 & n20489 ;
  assign n20491 = n13173 & n20490 ;
  assign n20493 = n20492 ^ n20491 ^ n331 ;
  assign n20494 = n5303 ^ n2812 ^ n2335 ;
  assign n20495 = n20494 ^ n11880 ^ n11249 ;
  assign n20497 = ( ~n1530 & n11691 ) | ( ~n1530 & n16980 ) | ( n11691 & n16980 ) ;
  assign n20496 = n18850 ^ n15128 ^ n6962 ;
  assign n20498 = n20497 ^ n20496 ^ n4963 ;
  assign n20499 = ( n12108 & n20495 ) | ( n12108 & n20498 ) | ( n20495 & n20498 ) ;
  assign n20500 = ( n7302 & ~n12757 ) | ( n7302 & n20499 ) | ( ~n12757 & n20499 ) ;
  assign n20501 = n963 & ~n8383 ;
  assign n20502 = ( n536 & n6457 ) | ( n536 & n20501 ) | ( n6457 & n20501 ) ;
  assign n20503 = n7805 ^ n6884 ^ n555 ;
  assign n20504 = ( n10921 & ~n12683 ) | ( n10921 & n20503 ) | ( ~n12683 & n20503 ) ;
  assign n20505 = ( ~n2276 & n18882 ) | ( ~n2276 & n20504 ) | ( n18882 & n20504 ) ;
  assign n20506 = n11520 ^ n11498 ^ n7431 ;
  assign n20507 = n13263 ^ n10505 ^ n7909 ;
  assign n20508 = ~n1856 & n8944 ;
  assign n20509 = n20508 ^ n11992 ^ n8331 ;
  assign n20510 = n16833 ^ n12918 ^ n3640 ;
  assign n20511 = n18970 ^ n3029 ^ 1'b0 ;
  assign n20513 = n5114 & ~n10076 ;
  assign n20512 = n1707 ^ n945 ^ n556 ;
  assign n20514 = n20513 ^ n20512 ^ n14191 ;
  assign n20515 = ( n2695 & ~n5904 ) | ( n2695 & n19844 ) | ( ~n5904 & n19844 ) ;
  assign n20516 = ( n2041 & n2066 ) | ( n2041 & ~n10516 ) | ( n2066 & ~n10516 ) ;
  assign n20517 = n20516 ^ n10950 ^ n9269 ;
  assign n20518 = n20517 ^ n14122 ^ n1199 ;
  assign n20519 = ( ~n20514 & n20515 ) | ( ~n20514 & n20518 ) | ( n20515 & n20518 ) ;
  assign n20520 = ( n4417 & n12708 ) | ( n4417 & n15625 ) | ( n12708 & n15625 ) ;
  assign n20521 = ( ~n1137 & n9610 ) | ( ~n1137 & n20520 ) | ( n9610 & n20520 ) ;
  assign n20522 = n12281 & n12285 ;
  assign n20523 = ~n3444 & n20522 ;
  assign n20524 = ( n9806 & ~n16824 ) | ( n9806 & n19489 ) | ( ~n16824 & n19489 ) ;
  assign n20525 = ( n7739 & ~n12229 ) | ( n7739 & n20524 ) | ( ~n12229 & n20524 ) ;
  assign n20526 = ( n12660 & n20523 ) | ( n12660 & ~n20525 ) | ( n20523 & ~n20525 ) ;
  assign n20527 = n20526 ^ n9762 ^ n867 ;
  assign n20528 = n7084 & n9623 ;
  assign n20529 = ~n10814 & n20528 ;
  assign n20530 = n20529 ^ n17507 ^ n4895 ;
  assign n20531 = n8250 ^ n8243 ^ n4083 ;
  assign n20532 = ( n15518 & n20089 ) | ( n15518 & n20531 ) | ( n20089 & n20531 ) ;
  assign n20533 = ( n10298 & n13133 ) | ( n10298 & ~n20532 ) | ( n13133 & ~n20532 ) ;
  assign n20534 = ( n2562 & n5656 ) | ( n2562 & ~n7574 ) | ( n5656 & ~n7574 ) ;
  assign n20535 = ( n200 & n16451 ) | ( n200 & ~n19336 ) | ( n16451 & ~n19336 ) ;
  assign n20536 = ~n20534 & n20535 ;
  assign n20537 = n20536 ^ n216 ^ 1'b0 ;
  assign n20538 = n19816 ^ n5127 ^ 1'b0 ;
  assign n20539 = ( ~n564 & n1352 ) | ( ~n564 & n20538 ) | ( n1352 & n20538 ) ;
  assign n20540 = ( ~n8932 & n9240 ) | ( ~n8932 & n9379 ) | ( n9240 & n9379 ) ;
  assign n20541 = n20540 ^ n18927 ^ n15682 ;
  assign n20542 = n6360 & n20541 ;
  assign n20543 = n2671 ^ n2309 ^ 1'b0 ;
  assign n20544 = n20542 | n20543 ;
  assign n20545 = n20544 ^ n15374 ^ n12498 ;
  assign n20546 = ( ~x65 & n5847 ) | ( ~x65 & n9502 ) | ( n5847 & n9502 ) ;
  assign n20547 = n4157 & ~n5528 ;
  assign n20548 = n7378 & n20547 ;
  assign n20549 = n20548 ^ n12941 ^ n2122 ;
  assign n20550 = n12671 ^ n2298 ^ 1'b0 ;
  assign n20551 = ( ~n2784 & n8750 ) | ( ~n2784 & n18091 ) | ( n8750 & n18091 ) ;
  assign n20554 = n17587 ^ x87 ^ 1'b0 ;
  assign n20552 = ( n9091 & n15445 ) | ( n9091 & n19062 ) | ( n15445 & n19062 ) ;
  assign n20553 = ( n4605 & n19117 ) | ( n4605 & n20552 ) | ( n19117 & n20552 ) ;
  assign n20555 = n20554 ^ n20553 ^ n17213 ;
  assign n20556 = n5692 & n17163 ;
  assign n20557 = ~n9701 & n20556 ;
  assign n20558 = n3083 ^ n1665 ^ 1'b0 ;
  assign n20559 = n7106 & n20558 ;
  assign n20560 = n20559 ^ n4326 ^ n1260 ;
  assign n20561 = n20560 ^ n6894 ^ n4612 ;
  assign n20562 = n20561 ^ n17627 ^ n9551 ;
  assign n20566 = n10375 ^ n5637 ^ n317 ;
  assign n20563 = n368 & ~n9748 ;
  assign n20564 = n20563 ^ n10578 ^ n8432 ;
  assign n20565 = ( n7804 & ~n8791 ) | ( n7804 & n20564 ) | ( ~n8791 & n20564 ) ;
  assign n20567 = n20566 ^ n20565 ^ n523 ;
  assign n20568 = n18155 ^ n3183 ^ 1'b0 ;
  assign n20569 = ( n10988 & ~n18786 ) | ( n10988 & n20568 ) | ( ~n18786 & n20568 ) ;
  assign n20570 = ( ~n1079 & n2616 ) | ( ~n1079 & n6807 ) | ( n2616 & n6807 ) ;
  assign n20571 = ( n7505 & ~n10576 ) | ( n7505 & n20570 ) | ( ~n10576 & n20570 ) ;
  assign n20572 = n20571 ^ n19628 ^ n7880 ;
  assign n20573 = n8753 ^ n8640 ^ n1655 ;
  assign n20574 = ( n3689 & ~n7431 ) | ( n3689 & n20573 ) | ( ~n7431 & n20573 ) ;
  assign n20575 = ( n10836 & n10951 ) | ( n10836 & n11209 ) | ( n10951 & n11209 ) ;
  assign n20576 = ( n2975 & n7183 ) | ( n2975 & n12952 ) | ( n7183 & n12952 ) ;
  assign n20577 = n20576 ^ n17047 ^ n4028 ;
  assign n20578 = ( n1328 & n8107 ) | ( n1328 & n20577 ) | ( n8107 & n20577 ) ;
  assign n20579 = n16392 & ~n20578 ;
  assign n20580 = n20575 & n20579 ;
  assign n20581 = n657 & n5677 ;
  assign n20582 = ~n11153 & n20581 ;
  assign n20583 = n883 & n6309 ;
  assign n20584 = ~n8091 & n20583 ;
  assign n20585 = ( n10070 & ~n12630 ) | ( n10070 & n20584 ) | ( ~n12630 & n20584 ) ;
  assign n20586 = ( ~n19324 & n20582 ) | ( ~n19324 & n20585 ) | ( n20582 & n20585 ) ;
  assign n20587 = n1827 & n2814 ;
  assign n20588 = n19853 ^ n11409 ^ n7474 ;
  assign n20589 = ( n15602 & n20587 ) | ( n15602 & ~n20588 ) | ( n20587 & ~n20588 ) ;
  assign n20590 = ( n11035 & n18017 ) | ( n11035 & n18960 ) | ( n18017 & n18960 ) ;
  assign n20591 = n14965 ^ n6922 ^ n4369 ;
  assign n20592 = ( ~n5335 & n11693 ) | ( ~n5335 & n13846 ) | ( n11693 & n13846 ) ;
  assign n20593 = ( n15596 & ~n20591 ) | ( n15596 & n20592 ) | ( ~n20591 & n20592 ) ;
  assign n20594 = ( n10761 & ~n14676 ) | ( n10761 & n14990 ) | ( ~n14676 & n14990 ) ;
  assign n20595 = n14692 ^ n982 ^ 1'b0 ;
  assign n20596 = n20595 ^ n13037 ^ n9612 ;
  assign n20597 = n8298 ^ n7228 ^ n2227 ;
  assign n20603 = ( n3009 & n8716 ) | ( n3009 & ~n9294 ) | ( n8716 & ~n9294 ) ;
  assign n20600 = ( n2735 & n11138 ) | ( n2735 & n18256 ) | ( n11138 & n18256 ) ;
  assign n20601 = n20600 ^ n5498 ^ 1'b0 ;
  assign n20602 = n3614 & n20601 ;
  assign n20598 = n1897 & n7276 ;
  assign n20599 = n20598 ^ n8759 ^ 1'b0 ;
  assign n20604 = n20603 ^ n20602 ^ n20599 ;
  assign n20605 = ( ~n11741 & n14396 ) | ( ~n11741 & n20604 ) | ( n14396 & n20604 ) ;
  assign n20606 = n20605 ^ n5253 ^ 1'b0 ;
  assign n20607 = n20597 & n20606 ;
  assign n20608 = ( n1045 & n5278 ) | ( n1045 & n11362 ) | ( n5278 & n11362 ) ;
  assign n20609 = n20608 ^ n18372 ^ n9683 ;
  assign n20610 = n20609 ^ n1880 ^ 1'b0 ;
  assign n20611 = n1794 & n4434 ;
  assign n20612 = n20611 ^ n16485 ^ n9704 ;
  assign n20613 = ( n1485 & ~n10482 ) | ( n1485 & n20612 ) | ( ~n10482 & n20612 ) ;
  assign n20614 = ~n12275 & n17820 ;
  assign n20615 = n20614 ^ n3253 ^ n1150 ;
  assign n20616 = ( n477 & n1907 ) | ( n477 & n20615 ) | ( n1907 & n20615 ) ;
  assign n20617 = ( ~n5815 & n18193 ) | ( ~n5815 & n20616 ) | ( n18193 & n20616 ) ;
  assign n20618 = ( n3084 & n6217 ) | ( n3084 & ~n14797 ) | ( n6217 & ~n14797 ) ;
  assign n20619 = ( n4233 & n11351 ) | ( n4233 & n20618 ) | ( n11351 & n20618 ) ;
  assign n20621 = ( n6270 & ~n8587 ) | ( n6270 & n15779 ) | ( ~n8587 & n15779 ) ;
  assign n20622 = n18210 ^ n3135 ^ 1'b0 ;
  assign n20623 = n20621 & n20622 ;
  assign n20620 = ~n7508 & n14506 ;
  assign n20624 = n20623 ^ n20620 ^ n486 ;
  assign n20625 = ( n6606 & ~n8715 ) | ( n6606 & n9413 ) | ( ~n8715 & n9413 ) ;
  assign n20626 = n8807 ^ n3593 ^ n3070 ;
  assign n20627 = n14619 ^ n7249 ^ n6075 ;
  assign n20628 = n20627 ^ n12343 ^ n8939 ;
  assign n20629 = n8809 ^ n7138 ^ n4896 ;
  assign n20630 = n20629 ^ n15633 ^ n7156 ;
  assign n20631 = ( n7587 & n9656 ) | ( n7587 & n9872 ) | ( n9656 & n9872 ) ;
  assign n20632 = n20631 ^ n19241 ^ n1543 ;
  assign n20633 = n20632 ^ n17031 ^ n7604 ;
  assign n20634 = n19681 ^ n8203 ^ n736 ;
  assign n20635 = n14847 ^ n2151 ^ n1391 ;
  assign n20636 = n14660 ^ n4953 ^ n227 ;
  assign n20637 = ( n5129 & n20635 ) | ( n5129 & n20636 ) | ( n20635 & n20636 ) ;
  assign n20638 = n14046 ^ n8103 ^ n1707 ;
  assign n20639 = n20638 ^ n12213 ^ n11195 ;
  assign n20640 = n18790 ^ n18352 ^ n11868 ;
  assign n20641 = ( n2139 & n20639 ) | ( n2139 & ~n20640 ) | ( n20639 & ~n20640 ) ;
  assign n20642 = ( n3670 & n7794 ) | ( n3670 & ~n13579 ) | ( n7794 & ~n13579 ) ;
  assign n20643 = ( n2996 & ~n3729 ) | ( n2996 & n20642 ) | ( ~n3729 & n20642 ) ;
  assign n20644 = n20643 ^ n11003 ^ n8230 ;
  assign n20645 = n6627 ^ n6085 ^ n1595 ;
  assign n20646 = ( n3244 & ~n8788 ) | ( n3244 & n20645 ) | ( ~n8788 & n20645 ) ;
  assign n20647 = ( n3760 & n10088 ) | ( n3760 & ~n10465 ) | ( n10088 & ~n10465 ) ;
  assign n20648 = n7552 & ~n20647 ;
  assign n20649 = ( n825 & ~n18620 ) | ( n825 & n20648 ) | ( ~n18620 & n20648 ) ;
  assign n20650 = n16770 ^ n13157 ^ 1'b0 ;
  assign n20651 = n20650 ^ n2268 ^ 1'b0 ;
  assign n20652 = n20649 & n20651 ;
  assign n20653 = ( n9050 & n20646 ) | ( n9050 & ~n20652 ) | ( n20646 & ~n20652 ) ;
  assign n20654 = n2062 & n4571 ;
  assign n20655 = n20654 ^ n266 ^ 1'b0 ;
  assign n20656 = ( ~n2331 & n6962 ) | ( ~n2331 & n20655 ) | ( n6962 & n20655 ) ;
  assign n20657 = ( n6199 & n9894 ) | ( n6199 & n20656 ) | ( n9894 & n20656 ) ;
  assign n20658 = ( n633 & ~n17912 ) | ( n633 & n20657 ) | ( ~n17912 & n20657 ) ;
  assign n20659 = n2592 & ~n14263 ;
  assign n20660 = n20659 ^ n3678 ^ 1'b0 ;
  assign n20661 = n20660 ^ n12890 ^ n7513 ;
  assign n20662 = n17242 ^ n13695 ^ n1686 ;
  assign n20663 = n20662 ^ n16103 ^ n15802 ;
  assign n20664 = n16969 ^ n1138 ^ 1'b0 ;
  assign n20665 = n4966 & ~n20664 ;
  assign n20666 = ( n8944 & n20663 ) | ( n8944 & n20665 ) | ( n20663 & n20665 ) ;
  assign n20667 = n4759 ^ n1671 ^ n1424 ;
  assign n20668 = ( n2120 & n18612 ) | ( n2120 & ~n20667 ) | ( n18612 & ~n20667 ) ;
  assign n20669 = n7746 & n20668 ;
  assign n20670 = ( ~x78 & n7218 ) | ( ~x78 & n17102 ) | ( n7218 & n17102 ) ;
  assign n20671 = n20670 ^ n19268 ^ x50 ;
  assign n20672 = n15897 ^ n14964 ^ 1'b0 ;
  assign n20673 = n16184 & n20672 ;
  assign n20675 = n13297 ^ n12100 ^ n8482 ;
  assign n20676 = n20675 ^ n19695 ^ n307 ;
  assign n20674 = n7192 ^ n4291 ^ n612 ;
  assign n20677 = n20676 ^ n20674 ^ n150 ;
  assign n20678 = n15157 ^ n10386 ^ 1'b0 ;
  assign n20679 = n20678 ^ n11494 ^ n8281 ;
  assign n20681 = n1387 & ~n9713 ;
  assign n20680 = n5375 | n13638 ;
  assign n20682 = n20681 ^ n20680 ^ n5210 ;
  assign n20683 = n9920 ^ n1505 ^ 1'b0 ;
  assign n20684 = n20683 ^ n8598 ^ n975 ;
  assign n20685 = ( n5750 & n7603 ) | ( n5750 & ~n9423 ) | ( n7603 & ~n9423 ) ;
  assign n20686 = n18016 ^ n11077 ^ n9109 ;
  assign n20691 = n1264 & n6897 ;
  assign n20692 = n20691 ^ n8086 ^ 1'b0 ;
  assign n20693 = n20692 ^ n16693 ^ n10423 ;
  assign n20687 = n9419 ^ n8384 ^ n701 ;
  assign n20688 = ( n17915 & n19765 ) | ( n17915 & n20687 ) | ( n19765 & n20687 ) ;
  assign n20689 = n7139 & ~n20688 ;
  assign n20690 = n20689 ^ n18491 ^ n18191 ;
  assign n20694 = n20693 ^ n20690 ^ n1245 ;
  assign n20695 = n20694 ^ n11543 ^ n3572 ;
  assign n20696 = n14801 ^ n9364 ^ n933 ;
  assign n20697 = ( n4487 & ~n7302 ) | ( n4487 & n12132 ) | ( ~n7302 & n12132 ) ;
  assign n20698 = n20697 ^ n12172 ^ n7285 ;
  assign n20699 = ( n6624 & ~n7048 ) | ( n6624 & n10053 ) | ( ~n7048 & n10053 ) ;
  assign n20700 = n20699 ^ n18533 ^ n4864 ;
  assign n20701 = n10516 ^ n8392 ^ n7570 ;
  assign n20702 = n2295 ^ n2116 ^ 1'b0 ;
  assign n20703 = n20701 | n20702 ;
  assign n20704 = ( n769 & ~n20700 ) | ( n769 & n20703 ) | ( ~n20700 & n20703 ) ;
  assign n20708 = n18597 ^ n5959 ^ 1'b0 ;
  assign n20707 = ( n958 & ~n3889 ) | ( n958 & n7636 ) | ( ~n3889 & n7636 ) ;
  assign n20705 = n6831 & ~n8788 ;
  assign n20706 = n6694 & n20705 ;
  assign n20709 = n20708 ^ n20707 ^ n20706 ;
  assign n20710 = n20709 ^ n19142 ^ n6798 ;
  assign n20716 = ( n1004 & n1795 ) | ( n1004 & ~n6333 ) | ( n1795 & ~n6333 ) ;
  assign n20714 = ( ~n6137 & n9193 ) | ( ~n6137 & n12017 ) | ( n9193 & n12017 ) ;
  assign n20715 = ( ~n7596 & n16273 ) | ( ~n7596 & n20714 ) | ( n16273 & n20714 ) ;
  assign n20712 = ( n15845 & ~n17028 ) | ( n15845 & n20038 ) | ( ~n17028 & n20038 ) ;
  assign n20711 = n16730 ^ n4770 ^ n2970 ;
  assign n20713 = n20712 ^ n20711 ^ n10180 ;
  assign n20717 = n20716 ^ n20715 ^ n20713 ;
  assign n20718 = n10728 ^ n9915 ^ n388 ;
  assign n20719 = ( n2735 & n4183 ) | ( n2735 & n20718 ) | ( n4183 & n20718 ) ;
  assign n20720 = n11970 ^ n7999 ^ n5776 ;
  assign n20721 = n20719 & ~n20720 ;
  assign n20728 = n7030 ^ n6588 ^ n191 ;
  assign n20727 = ( x19 & n1497 ) | ( x19 & n16494 ) | ( n1497 & n16494 ) ;
  assign n20729 = n20728 ^ n20727 ^ n6960 ;
  assign n20730 = n20729 ^ n17988 ^ 1'b0 ;
  assign n20723 = n7001 ^ n2504 ^ n1775 ;
  assign n20724 = ~n2470 & n20723 ;
  assign n20725 = ( n1020 & n2751 ) | ( n1020 & n20724 ) | ( n2751 & n20724 ) ;
  assign n20722 = n19515 ^ n11039 ^ n3866 ;
  assign n20726 = n20725 ^ n20722 ^ n11691 ;
  assign n20731 = n20730 ^ n20726 ^ n14049 ;
  assign n20732 = ( ~n2903 & n4388 ) | ( ~n2903 & n14314 ) | ( n4388 & n14314 ) ;
  assign n20733 = n3721 | n20732 ;
  assign n20734 = n20733 ^ n9741 ^ 1'b0 ;
  assign n20735 = n20313 ^ n18737 ^ 1'b0 ;
  assign n20736 = n13583 & ~n20735 ;
  assign n20739 = n20112 ^ n9651 ^ 1'b0 ;
  assign n20737 = n13133 ^ n9500 ^ n2528 ;
  assign n20738 = n20737 ^ n9431 ^ 1'b0 ;
  assign n20740 = n20739 ^ n20738 ^ n13731 ;
  assign n20741 = ( n10334 & ~n10474 ) | ( n10334 & n11739 ) | ( ~n10474 & n11739 ) ;
  assign n20742 = n20741 ^ n530 ^ 1'b0 ;
  assign n20743 = n19606 ^ n13504 ^ 1'b0 ;
  assign n20744 = n11057 & ~n20743 ;
  assign n20745 = n20744 ^ n12195 ^ n1509 ;
  assign n20746 = n519 & n2935 ;
  assign n20747 = n20746 ^ n12267 ^ n9008 ;
  assign n20752 = n6104 ^ n3789 ^ n530 ;
  assign n20748 = ( n2303 & n7040 ) | ( n2303 & n12317 ) | ( n7040 & n12317 ) ;
  assign n20749 = n20748 ^ n13534 ^ 1'b0 ;
  assign n20750 = n5669 & ~n20749 ;
  assign n20751 = n20750 ^ x88 ^ 1'b0 ;
  assign n20753 = n20752 ^ n20751 ^ n1003 ;
  assign n20754 = n4539 & n8677 ;
  assign n20755 = n19391 ^ n8260 ^ n2527 ;
  assign n20756 = ( n809 & n20754 ) | ( n809 & n20755 ) | ( n20754 & n20755 ) ;
  assign n20757 = n16163 ^ n16103 ^ n7737 ;
  assign n20758 = n9447 ^ n3453 ^ n2575 ;
  assign n20759 = ( n5446 & ~n14655 ) | ( n5446 & n20758 ) | ( ~n14655 & n20758 ) ;
  assign n20760 = ( x61 & ~n7837 ) | ( x61 & n11270 ) | ( ~n7837 & n11270 ) ;
  assign n20761 = n19594 ^ n249 ^ 1'b0 ;
  assign n20762 = n2806 | n20761 ;
  assign n20763 = ( ~n6447 & n20760 ) | ( ~n6447 & n20762 ) | ( n20760 & n20762 ) ;
  assign n20764 = ( ~n576 & n3274 ) | ( ~n576 & n7046 ) | ( n3274 & n7046 ) ;
  assign n20765 = n17496 ^ n11018 ^ n5380 ;
  assign n20766 = ( ~n15041 & n20764 ) | ( ~n15041 & n20765 ) | ( n20764 & n20765 ) ;
  assign n20767 = n11003 ^ n1434 ^ 1'b0 ;
  assign n20768 = n1977 | n20767 ;
  assign n20769 = ~n2421 & n20768 ;
  assign n20770 = ( n6749 & n10061 ) | ( n6749 & ~n11521 ) | ( n10061 & ~n11521 ) ;
  assign n20771 = n20770 ^ n18602 ^ 1'b0 ;
  assign n20772 = n9619 & n16194 ;
  assign n20773 = n13146 ^ n4663 ^ 1'b0 ;
  assign n20774 = n11080 ^ n3051 ^ 1'b0 ;
  assign n20775 = n20774 ^ n15247 ^ n13119 ;
  assign n20776 = ( n800 & ~n3203 ) | ( n800 & n7839 ) | ( ~n3203 & n7839 ) ;
  assign n20777 = n20776 ^ n13004 ^ n1769 ;
  assign n20778 = ( n777 & n1576 ) | ( n777 & n14956 ) | ( n1576 & n14956 ) ;
  assign n20779 = n20778 ^ n8635 ^ x38 ;
  assign n20780 = n2699 & n7254 ;
  assign n20781 = n20780 ^ n3173 ^ 1'b0 ;
  assign n20782 = n20781 ^ n5608 ^ n3851 ;
  assign n20783 = n20782 ^ n8764 ^ 1'b0 ;
  assign n20784 = ~n11964 & n20783 ;
  assign n20785 = n17337 ^ n7458 ^ 1'b0 ;
  assign n20786 = ( ~n15804 & n18718 ) | ( ~n15804 & n20785 ) | ( n18718 & n20785 ) ;
  assign n20787 = n12533 & ~n15004 ;
  assign n20788 = ( n8956 & n19340 ) | ( n8956 & ~n20787 ) | ( n19340 & ~n20787 ) ;
  assign n20789 = ( n3179 & n9820 ) | ( n3179 & ~n12825 ) | ( n9820 & ~n12825 ) ;
  assign n20790 = n20789 ^ n13097 ^ n7508 ;
  assign n20791 = ~n4760 & n8645 ;
  assign n20792 = n3434 | n5239 ;
  assign n20793 = n20792 ^ n13261 ^ 1'b0 ;
  assign n20795 = n11376 ^ n3789 ^ n1158 ;
  assign n20794 = n13377 ^ n5597 ^ n163 ;
  assign n20796 = n20795 ^ n20794 ^ n18023 ;
  assign n20797 = n139 & n15429 ;
  assign n20798 = ( ~x123 & n9900 ) | ( ~x123 & n20797 ) | ( n9900 & n20797 ) ;
  assign n20799 = x83 & ~n20456 ;
  assign n20800 = ~n12687 & n20799 ;
  assign n20801 = ( n6294 & ~n20798 ) | ( n6294 & n20800 ) | ( ~n20798 & n20800 ) ;
  assign n20802 = n14778 ^ n207 ^ 1'b0 ;
  assign n20803 = n19340 & ~n20802 ;
  assign n20804 = ( ~n1363 & n2536 ) | ( ~n1363 & n4809 ) | ( n2536 & n4809 ) ;
  assign n20805 = n20804 ^ n9097 ^ n3305 ;
  assign n20806 = n3085 ^ n3074 ^ n1837 ;
  assign n20807 = n20806 ^ n17275 ^ n6729 ;
  assign n20808 = ( n15066 & ~n16078 ) | ( n15066 & n20807 ) | ( ~n16078 & n20807 ) ;
  assign n20809 = n20805 | n20808 ;
  assign n20810 = n8715 | n20809 ;
  assign n20811 = n15853 ^ n11227 ^ n1357 ;
  assign n20812 = ( ~n1933 & n13681 ) | ( ~n1933 & n14564 ) | ( n13681 & n14564 ) ;
  assign n20813 = ( n5382 & ~n7191 ) | ( n5382 & n20812 ) | ( ~n7191 & n20812 ) ;
  assign n20814 = n11063 ^ n7105 ^ n1957 ;
  assign n20815 = ( n9452 & n14000 ) | ( n9452 & ~n20814 ) | ( n14000 & ~n20814 ) ;
  assign n20816 = n10065 ^ n8991 ^ 1'b0 ;
  assign n20817 = ( n2504 & n3995 ) | ( n2504 & ~n20816 ) | ( n3995 & ~n20816 ) ;
  assign n20818 = n20817 ^ n13534 ^ n1878 ;
  assign n20819 = n3199 | n3397 ;
  assign n20820 = n20819 ^ n12855 ^ n436 ;
  assign n20821 = n20820 ^ n15993 ^ n3517 ;
  assign n20822 = n20821 ^ n8657 ^ n6850 ;
  assign n20823 = ( ~n4737 & n14025 ) | ( ~n4737 & n16049 ) | ( n14025 & n16049 ) ;
  assign n20824 = n20823 ^ n9183 ^ 1'b0 ;
  assign n20825 = ( n3360 & n7351 ) | ( n3360 & n9128 ) | ( n7351 & n9128 ) ;
  assign n20826 = n20825 ^ n19095 ^ n13428 ;
  assign n20827 = ( ~n8691 & n15879 ) | ( ~n8691 & n17988 ) | ( n15879 & n17988 ) ;
  assign n20828 = n2668 ^ n951 ^ 1'b0 ;
  assign n20829 = n545 & n20828 ;
  assign n20830 = ( n927 & n15897 ) | ( n927 & ~n20829 ) | ( n15897 & ~n20829 ) ;
  assign n20831 = n10071 ^ n9425 ^ 1'b0 ;
  assign n20832 = ( n669 & n3033 ) | ( n669 & n5754 ) | ( n3033 & n5754 ) ;
  assign n20833 = ( ~n2375 & n15858 ) | ( ~n2375 & n17494 ) | ( n15858 & n17494 ) ;
  assign n20834 = ( n2281 & ~n14417 ) | ( n2281 & n20833 ) | ( ~n14417 & n20833 ) ;
  assign n20835 = ( ~n5743 & n10880 ) | ( ~n5743 & n20834 ) | ( n10880 & n20834 ) ;
  assign n20836 = n17621 ^ n14853 ^ n12448 ;
  assign n20838 = ( n161 & n2637 ) | ( n161 & n11217 ) | ( n2637 & n11217 ) ;
  assign n20837 = ( n2556 & n10210 ) | ( n2556 & n19338 ) | ( n10210 & n19338 ) ;
  assign n20839 = n20838 ^ n20837 ^ n15229 ;
  assign n20840 = ( n4112 & n12365 ) | ( n4112 & n20839 ) | ( n12365 & n20839 ) ;
  assign n20841 = n6336 ^ n273 ^ 1'b0 ;
  assign n20842 = n11858 & n20841 ;
  assign n20843 = ( n9146 & ~n12926 ) | ( n9146 & n20842 ) | ( ~n12926 & n20842 ) ;
  assign n20844 = ( n9997 & n15515 ) | ( n9997 & ~n16248 ) | ( n15515 & ~n16248 ) ;
  assign n20845 = ( n7915 & ~n10353 ) | ( n7915 & n20844 ) | ( ~n10353 & n20844 ) ;
  assign n20846 = n3712 & n12784 ;
  assign n20847 = n5795 & n20846 ;
  assign n20848 = ( n4843 & ~n8031 ) | ( n4843 & n12205 ) | ( ~n8031 & n12205 ) ;
  assign n20849 = n2412 & n20848 ;
  assign n20850 = ~n1170 & n20849 ;
  assign n20851 = ( n4686 & n6864 ) | ( n4686 & ~n7352 ) | ( n6864 & ~n7352 ) ;
  assign n20852 = n20851 ^ n5974 ^ n2537 ;
  assign n20853 = n12228 ^ n9729 ^ n1030 ;
  assign n20854 = n20853 ^ n3678 ^ n1385 ;
  assign n20855 = ( n390 & n1930 ) | ( n390 & ~n8686 ) | ( n1930 & ~n8686 ) ;
  assign n20856 = n20855 ^ n15145 ^ n13018 ;
  assign n20857 = n4289 & n17701 ;
  assign n20858 = n11925 & n20857 ;
  assign n20859 = n20858 ^ n18507 ^ n9283 ;
  assign n20860 = ( n6515 & n12889 ) | ( n6515 & n20859 ) | ( n12889 & n20859 ) ;
  assign n20865 = n14499 ^ n6922 ^ n2999 ;
  assign n20863 = n19764 ^ n12511 ^ n3091 ;
  assign n20861 = ( ~n2431 & n4335 ) | ( ~n2431 & n4937 ) | ( n4335 & n4937 ) ;
  assign n20862 = ( n4188 & ~n7040 ) | ( n4188 & n20861 ) | ( ~n7040 & n20861 ) ;
  assign n20864 = n20863 ^ n20862 ^ n10397 ;
  assign n20866 = n20865 ^ n20864 ^ n16508 ;
  assign n20867 = ( n2888 & ~n14187 ) | ( n2888 & n16515 ) | ( ~n14187 & n16515 ) ;
  assign n20868 = ( n3104 & n9588 ) | ( n3104 & n19899 ) | ( n9588 & n19899 ) ;
  assign n20869 = n20868 ^ n15099 ^ n6487 ;
  assign n20870 = n20869 ^ n1598 ^ 1'b0 ;
  assign n20872 = ( n3990 & ~n5743 ) | ( n3990 & n11926 ) | ( ~n5743 & n11926 ) ;
  assign n20871 = n3575 | n4457 ;
  assign n20873 = n20872 ^ n20871 ^ 1'b0 ;
  assign n20874 = n20873 ^ n6805 ^ n5515 ;
  assign n20875 = ( ~n448 & n5966 ) | ( ~n448 & n11412 ) | ( n5966 & n11412 ) ;
  assign n20881 = n14278 ^ n10842 ^ n8987 ;
  assign n20882 = n11029 & n20881 ;
  assign n20879 = n14843 ^ n13454 ^ n12475 ;
  assign n20880 = ( n5919 & n12447 ) | ( n5919 & n20879 ) | ( n12447 & n20879 ) ;
  assign n20877 = n18032 ^ n2795 ^ n2642 ;
  assign n20876 = n13350 ^ n7529 ^ n1667 ;
  assign n20878 = n20877 ^ n20876 ^ 1'b0 ;
  assign n20883 = n20882 ^ n20880 ^ n20878 ;
  assign n20884 = ( n1109 & ~n3346 ) | ( n1109 & n3869 ) | ( ~n3346 & n3869 ) ;
  assign n20885 = n20884 ^ n9551 ^ n5937 ;
  assign n20886 = ( ~n950 & n3764 ) | ( ~n950 & n14578 ) | ( n3764 & n14578 ) ;
  assign n20887 = ( n6591 & n7139 ) | ( n6591 & n13836 ) | ( n7139 & n13836 ) ;
  assign n20888 = ( n8648 & n15551 ) | ( n8648 & ~n20887 ) | ( n15551 & ~n20887 ) ;
  assign n20889 = ( n6462 & n20886 ) | ( n6462 & n20888 ) | ( n20886 & n20888 ) ;
  assign n20890 = ( n5870 & n20885 ) | ( n5870 & ~n20889 ) | ( n20885 & ~n20889 ) ;
  assign n20891 = n951 & n20890 ;
  assign n20892 = ( n6268 & ~n7738 ) | ( n6268 & n13090 ) | ( ~n7738 & n13090 ) ;
  assign n20893 = n20727 ^ n13918 ^ 1'b0 ;
  assign n20894 = n10299 ^ n7879 ^ 1'b0 ;
  assign n20895 = n14552 | n20894 ;
  assign n20897 = ( n517 & n5091 ) | ( n517 & n9611 ) | ( n5091 & n9611 ) ;
  assign n20896 = n18868 ^ n9480 ^ n8514 ;
  assign n20898 = n20897 ^ n20896 ^ 1'b0 ;
  assign n20899 = ( ~n3596 & n4790 ) | ( ~n3596 & n9376 ) | ( n4790 & n9376 ) ;
  assign n20900 = n10926 ^ n5386 ^ n1147 ;
  assign n20901 = ~x68 & n15073 ;
  assign n20902 = ( ~n379 & n8735 ) | ( ~n379 & n14651 ) | ( n8735 & n14651 ) ;
  assign n20903 = ( ~n5320 & n20901 ) | ( ~n5320 & n20902 ) | ( n20901 & n20902 ) ;
  assign n20904 = n20419 ^ n18017 ^ n13238 ;
  assign n20905 = ( n6008 & n12270 ) | ( n6008 & n20396 ) | ( n12270 & n20396 ) ;
  assign n20906 = n17086 ^ n15265 ^ n9512 ;
  assign n20907 = n18171 ^ n7640 ^ n5039 ;
  assign n20913 = ~n4674 & n5782 ;
  assign n20914 = n20913 ^ n16618 ^ 1'b0 ;
  assign n20911 = ( n459 & ~n4275 ) | ( n459 & n17183 ) | ( ~n4275 & n17183 ) ;
  assign n20912 = ( n421 & n8224 ) | ( n421 & n20911 ) | ( n8224 & n20911 ) ;
  assign n20908 = n19838 ^ n3179 ^ 1'b0 ;
  assign n20909 = n18005 & ~n20908 ;
  assign n20910 = n20909 ^ n10419 ^ n4536 ;
  assign n20915 = n20914 ^ n20912 ^ n20910 ;
  assign n20920 = n20514 ^ n10681 ^ n5470 ;
  assign n20916 = n5120 ^ n4165 ^ n4014 ;
  assign n20917 = n20916 ^ n8850 ^ n2156 ;
  assign n20918 = ( n12328 & n15905 ) | ( n12328 & ~n20797 ) | ( n15905 & ~n20797 ) ;
  assign n20919 = ( n18553 & n20917 ) | ( n18553 & n20918 ) | ( n20917 & n20918 ) ;
  assign n20921 = n20920 ^ n20919 ^ n19391 ;
  assign n20922 = n19675 ^ n2110 ^ n942 ;
  assign n20923 = ( ~n2887 & n3031 ) | ( ~n2887 & n6842 ) | ( n3031 & n6842 ) ;
  assign n20924 = n20923 ^ n20053 ^ n14884 ;
  assign n20925 = ( n10455 & n16650 ) | ( n10455 & ~n20924 ) | ( n16650 & ~n20924 ) ;
  assign n20926 = n11771 ^ n9729 ^ n4595 ;
  assign n20927 = ( ~n2748 & n20265 ) | ( ~n2748 & n20926 ) | ( n20265 & n20926 ) ;
  assign n20928 = n14318 | n20927 ;
  assign n20931 = n977 & n3834 ;
  assign n20932 = ~n3360 & n20931 ;
  assign n20930 = n5256 & n6626 ;
  assign n20929 = ( n4626 & n18531 ) | ( n4626 & ~n20023 ) | ( n18531 & ~n20023 ) ;
  assign n20933 = n20932 ^ n20930 ^ n20929 ;
  assign n20934 = n9204 | n11548 ;
  assign n20935 = ( n3539 & ~n3580 ) | ( n3539 & n4281 ) | ( ~n3580 & n4281 ) ;
  assign n20936 = n3266 & n20935 ;
  assign n20937 = n9972 & n20936 ;
  assign n20938 = n12343 ^ n3315 ^ 1'b0 ;
  assign n20939 = n20166 ^ n11829 ^ n7467 ;
  assign n20940 = n20939 ^ n5891 ^ n1817 ;
  assign n20941 = n11376 ^ n10986 ^ 1'b0 ;
  assign n20942 = n19253 | n20941 ;
  assign n20943 = ( n12955 & n17214 ) | ( n12955 & n20942 ) | ( n17214 & n20942 ) ;
  assign n20944 = n18198 ^ n9954 ^ n9595 ;
  assign n20945 = n2286 & n3999 ;
  assign n20946 = n2266 ^ n2221 ^ n1667 ;
  assign n20947 = ( n16829 & n20945 ) | ( n16829 & n20946 ) | ( n20945 & n20946 ) ;
  assign n20948 = n20947 ^ n8938 ^ n419 ;
  assign n20949 = n20948 ^ n14730 ^ n10598 ;
  assign n20950 = ( n1343 & n1666 ) | ( n1343 & n3154 ) | ( n1666 & n3154 ) ;
  assign n20951 = n20950 ^ n5290 ^ n4188 ;
  assign n20952 = ( n1373 & n2347 ) | ( n1373 & ~n5601 ) | ( n2347 & ~n5601 ) ;
  assign n20953 = n20952 ^ n2039 ^ n1684 ;
  assign n20954 = ( n13932 & n20951 ) | ( n13932 & ~n20953 ) | ( n20951 & ~n20953 ) ;
  assign n20955 = ( n1264 & n2286 ) | ( n1264 & n7908 ) | ( n2286 & n7908 ) ;
  assign n20956 = n20955 ^ n9483 ^ n4557 ;
  assign n20957 = ( ~n1642 & n1932 ) | ( ~n1642 & n3356 ) | ( n1932 & n3356 ) ;
  assign n20958 = ( n5459 & n8579 ) | ( n5459 & n20957 ) | ( n8579 & n20957 ) ;
  assign n20959 = ( n11057 & n20956 ) | ( n11057 & ~n20958 ) | ( n20956 & ~n20958 ) ;
  assign n20960 = ( ~n7539 & n13936 ) | ( ~n7539 & n18835 ) | ( n13936 & n18835 ) ;
  assign n20961 = ~n7079 & n20960 ;
  assign n20962 = n1454 & n16348 ;
  assign n20963 = n20962 ^ n9874 ^ 1'b0 ;
  assign n20964 = ( n4717 & ~n20449 ) | ( n4717 & n20963 ) | ( ~n20449 & n20963 ) ;
  assign n20965 = ( n3068 & n17311 ) | ( n3068 & n20964 ) | ( n17311 & n20964 ) ;
  assign n20966 = ( n2410 & n2716 ) | ( n2410 & n11362 ) | ( n2716 & n11362 ) ;
  assign n20967 = n11246 ^ n10258 ^ 1'b0 ;
  assign n20968 = ~n3565 & n20967 ;
  assign n20969 = n15631 ^ n11569 ^ n10003 ;
  assign n20970 = n20969 ^ n15602 ^ n10011 ;
  assign n20971 = ( n3427 & n17470 ) | ( n3427 & n20970 ) | ( n17470 & n20970 ) ;
  assign n20972 = ( n3220 & ~n6409 ) | ( n3220 & n20971 ) | ( ~n6409 & n20971 ) ;
  assign n20973 = ( n5805 & n11502 ) | ( n5805 & ~n17252 ) | ( n11502 & ~n17252 ) ;
  assign n20974 = n12735 ^ n3834 ^ n496 ;
  assign n20975 = ( ~n7441 & n7776 ) | ( ~n7441 & n16079 ) | ( n7776 & n16079 ) ;
  assign n20976 = ( ~n2008 & n19116 ) | ( ~n2008 & n20881 ) | ( n19116 & n20881 ) ;
  assign n20977 = n11385 & n20066 ;
  assign n20978 = n12290 ^ n11704 ^ 1'b0 ;
  assign n20979 = n13230 & n18147 ;
  assign n20980 = ~n4544 & n20979 ;
  assign n20981 = ~n2693 & n6188 ;
  assign n20982 = n7346 & n20981 ;
  assign n20983 = n20982 ^ n14450 ^ n2881 ;
  assign n20984 = n3469 & n20983 ;
  assign n20985 = n20984 ^ n11951 ^ 1'b0 ;
  assign n20987 = n7787 ^ n6011 ^ n4372 ;
  assign n20986 = ( n2530 & n20066 ) | ( n2530 & n20540 ) | ( n20066 & n20540 ) ;
  assign n20988 = n20987 ^ n20986 ^ n15807 ;
  assign n20989 = n20988 ^ n7308 ^ n3648 ;
  assign n20990 = n2175 ^ n2021 ^ n453 ;
  assign n20991 = n10989 | n20990 ;
  assign n20992 = n20989 | n20991 ;
  assign n20993 = n17985 ^ n7380 ^ n535 ;
  assign n20994 = ( n6311 & n14226 ) | ( n6311 & ~n14572 ) | ( n14226 & ~n14572 ) ;
  assign n20995 = ( n4018 & n7767 ) | ( n4018 & n12847 ) | ( n7767 & n12847 ) ;
  assign n20996 = n8209 ^ n5904 ^ n5572 ;
  assign n20997 = ( n14061 & n15257 ) | ( n14061 & n17195 ) | ( n15257 & n17195 ) ;
  assign n20998 = n2404 ^ n1053 ^ 1'b0 ;
  assign n20999 = n4842 & ~n20998 ;
  assign n21000 = n20999 ^ n12637 ^ x81 ;
  assign n21001 = ( x48 & n20997 ) | ( x48 & ~n21000 ) | ( n20997 & ~n21000 ) ;
  assign n21002 = n19665 ^ n13384 ^ n213 ;
  assign n21003 = n21002 ^ n19566 ^ n16544 ;
  assign n21004 = n11372 ^ n2450 ^ n1300 ;
  assign n21005 = n21004 ^ n18819 ^ n4180 ;
  assign n21009 = n17266 ^ n15434 ^ n3254 ;
  assign n21006 = ( n537 & n1027 ) | ( n537 & ~n1360 ) | ( n1027 & ~n1360 ) ;
  assign n21007 = n10675 ^ n4881 ^ 1'b0 ;
  assign n21008 = n21006 | n21007 ;
  assign n21010 = n21009 ^ n21008 ^ n4155 ;
  assign n21011 = n16732 ^ n16273 ^ n1425 ;
  assign n21012 = n21011 ^ n18203 ^ n13715 ;
  assign n21013 = ~n1086 & n8524 ;
  assign n21014 = ~n14158 & n21013 ;
  assign n21016 = n1163 & n12241 ;
  assign n21017 = n21016 ^ n4112 ^ 1'b0 ;
  assign n21015 = n15165 ^ n432 ^ 1'b0 ;
  assign n21018 = n21017 ^ n21015 ^ n20150 ;
  assign n21019 = n20824 | n21018 ;
  assign n21020 = n21019 ^ n5187 ^ 1'b0 ;
  assign n21021 = ( ~n6955 & n11688 ) | ( ~n6955 & n14489 ) | ( n11688 & n14489 ) ;
  assign n21022 = ~n323 & n9107 ;
  assign n21023 = n10745 ^ n10620 ^ n4253 ;
  assign n21024 = ( n17108 & n21022 ) | ( n17108 & n21023 ) | ( n21022 & n21023 ) ;
  assign n21025 = ( ~n17622 & n21021 ) | ( ~n17622 & n21024 ) | ( n21021 & n21024 ) ;
  assign n21026 = ( n9250 & ~n10265 ) | ( n9250 & n21025 ) | ( ~n10265 & n21025 ) ;
  assign n21027 = ( n380 & n1525 ) | ( n380 & ~n12956 ) | ( n1525 & ~n12956 ) ;
  assign n21028 = ( ~n5622 & n5660 ) | ( ~n5622 & n6466 ) | ( n5660 & n6466 ) ;
  assign n21029 = n17871 ^ n14945 ^ n4510 ;
  assign n21030 = ( n17037 & ~n19611 ) | ( n17037 & n21029 ) | ( ~n19611 & n21029 ) ;
  assign n21031 = n20534 ^ n14416 ^ n7141 ;
  assign n21032 = n7039 ^ n1110 ^ 1'b0 ;
  assign n21033 = n14629 | n21032 ;
  assign n21034 = ( ~n539 & n557 ) | ( ~n539 & n2531 ) | ( n557 & n2531 ) ;
  assign n21035 = n21034 ^ n8491 ^ 1'b0 ;
  assign n21036 = n4067 | n21035 ;
  assign n21037 = ( n4572 & ~n4690 ) | ( n4572 & n21036 ) | ( ~n4690 & n21036 ) ;
  assign n21038 = n13138 ^ n631 ^ 1'b0 ;
  assign n21039 = n21037 & n21038 ;
  assign n21040 = ~n2062 & n21039 ;
  assign n21041 = n17703 ^ n15549 ^ n4944 ;
  assign n21042 = n21041 ^ n18720 ^ n11431 ;
  assign n21043 = ( n518 & n9819 ) | ( n518 & ~n16091 ) | ( n9819 & ~n16091 ) ;
  assign n21044 = n7423 | n21043 ;
  assign n21045 = ( ~n1119 & n8100 ) | ( ~n1119 & n11570 ) | ( n8100 & n11570 ) ;
  assign n21046 = n21045 ^ n14996 ^ 1'b0 ;
  assign n21047 = ( n17543 & ~n20084 ) | ( n17543 & n21046 ) | ( ~n20084 & n21046 ) ;
  assign n21051 = n279 & ~n959 ;
  assign n21052 = n21051 ^ n5980 ^ 1'b0 ;
  assign n21049 = n7879 ^ n1588 ^ 1'b0 ;
  assign n21050 = n21049 ^ n1659 ^ n409 ;
  assign n21048 = ( ~n8259 & n12294 ) | ( ~n8259 & n14976 ) | ( n12294 & n14976 ) ;
  assign n21053 = n21052 ^ n21050 ^ n21048 ;
  assign n21055 = n13581 ^ n3424 ^ n1443 ;
  assign n21054 = ( n3776 & ~n4675 ) | ( n3776 & n17984 ) | ( ~n4675 & n17984 ) ;
  assign n21056 = n21055 ^ n21054 ^ n8681 ;
  assign n21057 = n4810 & n10916 ;
  assign n21058 = n21057 ^ n6333 ^ 1'b0 ;
  assign n21059 = n4182 & ~n7153 ;
  assign n21060 = n12114 & n21059 ;
  assign n21062 = n11473 ^ n9995 ^ n2008 ;
  assign n21063 = ( n1933 & ~n17871 ) | ( n1933 & n21062 ) | ( ~n17871 & n21062 ) ;
  assign n21061 = ~n9341 & n14204 ;
  assign n21064 = n21063 ^ n21061 ^ n1259 ;
  assign n21067 = ( n228 & ~n6544 ) | ( n228 & n10314 ) | ( ~n6544 & n10314 ) ;
  assign n21065 = n6395 ^ n3823 ^ n2846 ;
  assign n21066 = ( n6901 & n8567 ) | ( n6901 & n21065 ) | ( n8567 & n21065 ) ;
  assign n21068 = n21067 ^ n21066 ^ n15703 ;
  assign n21069 = ( n3406 & n20970 ) | ( n3406 & ~n21068 ) | ( n20970 & ~n21068 ) ;
  assign n21074 = n3371 ^ n2092 ^ n732 ;
  assign n21075 = n21074 ^ n8788 ^ x3 ;
  assign n21076 = n14083 ^ n6782 ^ 1'b0 ;
  assign n21077 = ( n10552 & n21075 ) | ( n10552 & n21076 ) | ( n21075 & n21076 ) ;
  assign n21070 = n14559 ^ n2763 ^ n1815 ;
  assign n21071 = n21070 ^ n9260 ^ n4365 ;
  assign n21072 = n15440 & n21071 ;
  assign n21073 = n21072 ^ n6589 ^ 1'b0 ;
  assign n21078 = n21077 ^ n21073 ^ n3851 ;
  assign n21079 = n21078 ^ n12128 ^ n1611 ;
  assign n21082 = n19289 ^ n13668 ^ n5997 ;
  assign n21083 = n21082 ^ n12685 ^ n6541 ;
  assign n21080 = n10932 ^ n955 ^ 1'b0 ;
  assign n21081 = ~n16568 & n21080 ;
  assign n21084 = n21083 ^ n21081 ^ n3327 ;
  assign n21085 = ( n5741 & n9538 ) | ( n5741 & ~n10112 ) | ( n9538 & ~n10112 ) ;
  assign n21086 = ( ~n3908 & n12152 ) | ( ~n3908 & n21085 ) | ( n12152 & n21085 ) ;
  assign n21088 = ( n157 & n8122 ) | ( n157 & n17000 ) | ( n8122 & n17000 ) ;
  assign n21089 = n21088 ^ n11264 ^ 1'b0 ;
  assign n21087 = ( n9453 & n15722 ) | ( n9453 & n16531 ) | ( n15722 & n16531 ) ;
  assign n21090 = n21089 ^ n21087 ^ n10958 ;
  assign n21091 = ( n139 & n8119 ) | ( n139 & ~n8904 ) | ( n8119 & ~n8904 ) ;
  assign n21092 = n21091 ^ n18130 ^ n12048 ;
  assign n21093 = ( ~n3349 & n3907 ) | ( ~n3349 & n21092 ) | ( n3907 & n21092 ) ;
  assign n21094 = n14608 | n15514 ;
  assign n21096 = ( n242 & n2168 ) | ( n242 & ~n2179 ) | ( n2168 & ~n2179 ) ;
  assign n21095 = ( n1503 & n2914 ) | ( n1503 & ~n3596 ) | ( n2914 & ~n3596 ) ;
  assign n21097 = n21096 ^ n21095 ^ n6492 ;
  assign n21098 = n19667 ^ n5718 ^ n172 ;
  assign n21099 = n21098 ^ n14530 ^ n11499 ;
  assign n21100 = ( ~n11350 & n11451 ) | ( ~n11350 & n20268 ) | ( n11451 & n20268 ) ;
  assign n21101 = ( n8189 & ~n14512 ) | ( n8189 & n16422 ) | ( ~n14512 & n16422 ) ;
  assign n21102 = n7438 & ~n12200 ;
  assign n21103 = n21102 ^ n7807 ^ 1'b0 ;
  assign n21104 = ~n7287 & n8691 ;
  assign n21105 = n8268 ^ n1384 ^ 1'b0 ;
  assign n21106 = ( ~n2733 & n12764 ) | ( ~n2733 & n19303 ) | ( n12764 & n19303 ) ;
  assign n21107 = n21106 ^ n12818 ^ n2748 ;
  assign n21108 = ~n4129 & n6276 ;
  assign n21109 = n21108 ^ n7792 ^ 1'b0 ;
  assign n21110 = n11343 ^ n2710 ^ n396 ;
  assign n21111 = n21110 ^ n6310 ^ 1'b0 ;
  assign n21112 = ~n21109 & n21111 ;
  assign n21113 = ( n10471 & n14885 ) | ( n10471 & ~n21112 ) | ( n14885 & ~n21112 ) ;
  assign n21114 = n18749 ^ n18640 ^ n16541 ;
  assign n21116 = ( ~n3109 & n6180 ) | ( ~n3109 & n9183 ) | ( n6180 & n9183 ) ;
  assign n21115 = ( n3704 & n9246 ) | ( n3704 & ~n17067 ) | ( n9246 & ~n17067 ) ;
  assign n21117 = n21116 ^ n21115 ^ n17096 ;
  assign n21118 = ( x17 & n13055 ) | ( x17 & ~n21117 ) | ( n13055 & ~n21117 ) ;
  assign n21120 = ( ~n2371 & n2673 ) | ( ~n2371 & n2763 ) | ( n2673 & n2763 ) ;
  assign n21119 = n715 & n16121 ;
  assign n21121 = n21120 ^ n21119 ^ 1'b0 ;
  assign n21122 = ( n4537 & ~n7971 ) | ( n4537 & n10842 ) | ( ~n7971 & n10842 ) ;
  assign n21123 = ( n2697 & n3090 ) | ( n2697 & ~n16777 ) | ( n3090 & ~n16777 ) ;
  assign n21124 = ( n8006 & n16814 ) | ( n8006 & ~n21123 ) | ( n16814 & ~n21123 ) ;
  assign n21125 = n21124 ^ n9617 ^ n2428 ;
  assign n21126 = n15477 ^ n10852 ^ n6928 ;
  assign n21127 = ( n6847 & ~n11672 ) | ( n6847 & n21126 ) | ( ~n11672 & n21126 ) ;
  assign n21128 = ( ~n2353 & n9493 ) | ( ~n2353 & n21127 ) | ( n9493 & n21127 ) ;
  assign n21129 = n21128 ^ n18656 ^ n11067 ;
  assign n21130 = n1636 & n3598 ;
  assign n21131 = n21130 ^ n8842 ^ 1'b0 ;
  assign n21132 = n21131 ^ n12070 ^ n7487 ;
  assign n21133 = ( n3849 & ~n14422 ) | ( n3849 & n17954 ) | ( ~n14422 & n17954 ) ;
  assign n21134 = ( n7683 & n10079 ) | ( n7683 & n20135 ) | ( n10079 & n20135 ) ;
  assign n21135 = n19284 ^ n10365 ^ n1557 ;
  assign n21136 = n3575 & n16753 ;
  assign n21137 = n15823 ^ n10979 ^ n398 ;
  assign n21138 = n11161 ^ n6086 ^ n5061 ;
  assign n21139 = n20736 ^ n19119 ^ n5566 ;
  assign n21140 = n10691 ^ n6946 ^ n5754 ;
  assign n21141 = n7199 ^ n7004 ^ 1'b0 ;
  assign n21142 = ~n2958 & n21141 ;
  assign n21143 = n10472 ^ n6040 ^ n2767 ;
  assign n21144 = ( n5351 & n11786 ) | ( n5351 & n21143 ) | ( n11786 & n21143 ) ;
  assign n21145 = n6455 | n20132 ;
  assign n21146 = n6955 ^ n1543 ^ n721 ;
  assign n21147 = n21146 ^ n12576 ^ n9121 ;
  assign n21148 = n17320 ^ n9288 ^ n2514 ;
  assign n21149 = n16898 ^ n6109 ^ n5136 ;
  assign n21150 = ( n21147 & n21148 ) | ( n21147 & ~n21149 ) | ( n21148 & ~n21149 ) ;
  assign n21151 = ( n938 & n5668 ) | ( n938 & ~n8254 ) | ( n5668 & ~n8254 ) ;
  assign n21152 = n10520 ^ n7130 ^ n5803 ;
  assign n21153 = n5719 & ~n21152 ;
  assign n21154 = n9247 ^ n8337 ^ n2481 ;
  assign n21155 = n21154 ^ n13274 ^ n10449 ;
  assign n21156 = n20917 ^ n2864 ^ n1090 ;
  assign n21157 = ~n858 & n5410 ;
  assign n21158 = ( n5357 & ~n21156 ) | ( n5357 & n21157 ) | ( ~n21156 & n21157 ) ;
  assign n21159 = ( n2243 & ~n17724 ) | ( n2243 & n21158 ) | ( ~n17724 & n21158 ) ;
  assign n21160 = ( n14785 & n17682 ) | ( n14785 & n19812 ) | ( n17682 & n19812 ) ;
  assign n21161 = n330 & n14592 ;
  assign n21162 = n21161 ^ n9538 ^ 1'b0 ;
  assign n21163 = ~n19812 & n21162 ;
  assign n21164 = n21163 ^ n5252 ^ 1'b0 ;
  assign n21165 = ( n2549 & n18589 ) | ( n2549 & n21164 ) | ( n18589 & n21164 ) ;
  assign n21166 = ( n12048 & ~n20608 ) | ( n12048 & n21165 ) | ( ~n20608 & n21165 ) ;
  assign n21167 = n3697 ^ n3473 ^ n552 ;
  assign n21168 = n16561 & n21167 ;
  assign n21169 = n21168 ^ n11590 ^ n151 ;
  assign n21170 = ( n4487 & n4750 ) | ( n4487 & ~n6077 ) | ( n4750 & ~n6077 ) ;
  assign n21171 = n7054 | n21170 ;
  assign n21172 = n14026 & ~n21171 ;
  assign n21173 = n21172 ^ n4333 ^ 1'b0 ;
  assign n21174 = ~n18089 & n21173 ;
  assign n21175 = n19637 ^ n3954 ^ n3308 ;
  assign n21176 = n9065 & ~n21175 ;
  assign n21177 = ( n1514 & n2417 ) | ( n1514 & n2697 ) | ( n2417 & n2697 ) ;
  assign n21178 = ( ~n10463 & n14953 ) | ( ~n10463 & n21177 ) | ( n14953 & n21177 ) ;
  assign n21179 = ( n1520 & n3059 ) | ( n1520 & ~n6804 ) | ( n3059 & ~n6804 ) ;
  assign n21180 = ( n17642 & ~n18117 ) | ( n17642 & n21179 ) | ( ~n18117 & n21179 ) ;
  assign n21181 = ( n3365 & n13581 ) | ( n3365 & ~n19903 ) | ( n13581 & ~n19903 ) ;
  assign n21186 = n7922 & ~n10332 ;
  assign n21182 = ( n830 & n7096 ) | ( n830 & n7692 ) | ( n7096 & n7692 ) ;
  assign n21183 = ( ~n4904 & n13078 ) | ( ~n4904 & n21182 ) | ( n13078 & n21182 ) ;
  assign n21184 = ~n10631 & n21183 ;
  assign n21185 = n21184 ^ n13559 ^ 1'b0 ;
  assign n21187 = n21186 ^ n21185 ^ n19890 ;
  assign n21188 = ( n565 & ~n2663 ) | ( n565 & n8628 ) | ( ~n2663 & n8628 ) ;
  assign n21189 = n21188 ^ n10099 ^ n3538 ;
  assign n21190 = n1311 & ~n4124 ;
  assign n21191 = ~n5025 & n20988 ;
  assign n21192 = n21190 & n21191 ;
  assign n21193 = n13376 ^ n8107 ^ n1090 ;
  assign n21194 = ( n1774 & n6809 ) | ( n1774 & n20272 ) | ( n6809 & n20272 ) ;
  assign n21195 = ( n10688 & n21193 ) | ( n10688 & n21194 ) | ( n21193 & n21194 ) ;
  assign n21196 = n17759 ^ n2339 ^ 1'b0 ;
  assign n21197 = n15664 | n21196 ;
  assign n21198 = ( n7727 & ~n20217 ) | ( n7727 & n21197 ) | ( ~n20217 & n21197 ) ;
  assign n21201 = n14806 ^ n4758 ^ n633 ;
  assign n21200 = ( n3188 & n9602 ) | ( n3188 & ~n10539 ) | ( n9602 & ~n10539 ) ;
  assign n21199 = ( ~n8411 & n12760 ) | ( ~n8411 & n19588 ) | ( n12760 & n19588 ) ;
  assign n21202 = n21201 ^ n21200 ^ n21199 ;
  assign n21203 = n21202 ^ n20187 ^ n8917 ;
  assign n21208 = ( n189 & n5834 ) | ( n189 & n7208 ) | ( n5834 & n7208 ) ;
  assign n21204 = n2134 & ~n13406 ;
  assign n21205 = n21204 ^ n4814 ^ 1'b0 ;
  assign n21206 = ( n4796 & n9978 ) | ( n4796 & n13582 ) | ( n9978 & n13582 ) ;
  assign n21207 = ( n9552 & n21205 ) | ( n9552 & ~n21206 ) | ( n21205 & ~n21206 ) ;
  assign n21209 = n21208 ^ n21207 ^ n6037 ;
  assign n21210 = n21209 ^ n18292 ^ n8480 ;
  assign n21211 = ~n5581 & n13770 ;
  assign n21212 = ( n13320 & n21210 ) | ( n13320 & ~n21211 ) | ( n21210 & ~n21211 ) ;
  assign n21213 = n19103 ^ n12413 ^ n1653 ;
  assign n21214 = x70 & n8432 ;
  assign n21215 = ~n21213 & n21214 ;
  assign n21216 = n21215 ^ n5865 ^ n452 ;
  assign n21217 = n21216 ^ n15399 ^ n4614 ;
  assign n21218 = ( n4505 & ~n6857 ) | ( n4505 & n19922 ) | ( ~n6857 & n19922 ) ;
  assign n21219 = n14670 ^ n12308 ^ n3431 ;
  assign n21220 = ( n10861 & ~n21218 ) | ( n10861 & n21219 ) | ( ~n21218 & n21219 ) ;
  assign n21221 = n184 | n5147 ;
  assign n21222 = n18576 ^ n12449 ^ n11081 ;
  assign n21223 = n21221 & n21222 ;
  assign n21224 = ( n2158 & ~n11906 ) | ( n2158 & n13141 ) | ( ~n11906 & n13141 ) ;
  assign n21225 = ( n2121 & ~n13091 ) | ( n2121 & n21224 ) | ( ~n13091 & n21224 ) ;
  assign n21226 = ( ~n5622 & n9249 ) | ( ~n5622 & n21225 ) | ( n9249 & n21225 ) ;
  assign n21227 = n8550 ^ n3127 ^ 1'b0 ;
  assign n21228 = n21227 ^ n6596 ^ n6534 ;
  assign n21229 = ( n12780 & n14037 ) | ( n12780 & ~n21228 ) | ( n14037 & ~n21228 ) ;
  assign n21230 = n21229 ^ n1597 ^ n1466 ;
  assign n21231 = ( n524 & n1379 ) | ( n524 & n14421 ) | ( n1379 & n14421 ) ;
  assign n21232 = n21231 ^ n12890 ^ n2240 ;
  assign n21233 = n21232 ^ n16483 ^ n5062 ;
  assign n21234 = ( n3222 & n10828 ) | ( n3222 & ~n14022 ) | ( n10828 & ~n14022 ) ;
  assign n21235 = n19920 ^ n1992 ^ 1'b0 ;
  assign n21236 = n8863 & n21235 ;
  assign n21237 = ( n3412 & ~n12983 ) | ( n3412 & n14844 ) | ( ~n12983 & n14844 ) ;
  assign n21238 = n21237 ^ n19447 ^ n3268 ;
  assign n21239 = n16147 ^ n10725 ^ n4133 ;
  assign n21240 = ( n4090 & n14715 ) | ( n4090 & n21239 ) | ( n14715 & n21239 ) ;
  assign n21241 = ( ~n764 & n779 ) | ( ~n764 & n5303 ) | ( n779 & n5303 ) ;
  assign n21242 = n21241 ^ n15832 ^ n2314 ;
  assign n21243 = ( n2887 & n11156 ) | ( n2887 & ~n13107 ) | ( n11156 & ~n13107 ) ;
  assign n21244 = n9590 ^ n5889 ^ 1'b0 ;
  assign n21245 = n21244 ^ n15857 ^ 1'b0 ;
  assign n21246 = ~n6551 & n21245 ;
  assign n21247 = n21246 ^ n14097 ^ n2309 ;
  assign n21248 = ( ~n4148 & n7971 ) | ( ~n4148 & n21110 ) | ( n7971 & n21110 ) ;
  assign n21249 = ( n2570 & n3583 ) | ( n2570 & n21248 ) | ( n3583 & n21248 ) ;
  assign n21250 = n21249 ^ n15189 ^ n13529 ;
  assign n21251 = n10680 ^ n8513 ^ 1'b0 ;
  assign n21252 = n19386 & n21251 ;
  assign n21253 = n11500 ^ n4939 ^ n1636 ;
  assign n21254 = n19326 ^ n2590 ^ 1'b0 ;
  assign n21255 = n8490 | n21254 ;
  assign n21259 = ( n1202 & n5108 ) | ( n1202 & n6727 ) | ( n5108 & n6727 ) ;
  assign n21256 = ( ~n6794 & n9561 ) | ( ~n6794 & n11339 ) | ( n9561 & n11339 ) ;
  assign n21257 = ~n12347 & n20781 ;
  assign n21258 = n21256 & n21257 ;
  assign n21260 = n21259 ^ n21258 ^ n2801 ;
  assign n21261 = ( n6260 & ~n21255 ) | ( n6260 & n21260 ) | ( ~n21255 & n21260 ) ;
  assign n21262 = ( n3752 & n21253 ) | ( n3752 & n21261 ) | ( n21253 & n21261 ) ;
  assign n21263 = n16243 ^ n11120 ^ 1'b0 ;
  assign n21264 = ~n8445 & n21263 ;
  assign n21265 = n21262 | n21264 ;
  assign n21266 = ( ~n20350 & n21252 ) | ( ~n20350 & n21265 ) | ( n21252 & n21265 ) ;
  assign n21267 = ~n5304 & n12562 ;
  assign n21273 = n11806 ^ n5286 ^ n3206 ;
  assign n21274 = n21273 ^ n8021 ^ n7812 ;
  assign n21268 = ( n3878 & n4596 ) | ( n3878 & n6094 ) | ( n4596 & n6094 ) ;
  assign n21269 = ~n1172 & n11975 ;
  assign n21270 = n21268 | n21269 ;
  assign n21271 = n21270 ^ n14413 ^ 1'b0 ;
  assign n21272 = ( n9310 & n11891 ) | ( n9310 & n21271 ) | ( n11891 & n21271 ) ;
  assign n21275 = n21274 ^ n21272 ^ n17556 ;
  assign n21276 = ~n670 & n4378 ;
  assign n21277 = n21276 ^ n4846 ^ 1'b0 ;
  assign n21278 = ( n4319 & n15115 ) | ( n4319 & ~n16938 ) | ( n15115 & ~n16938 ) ;
  assign n21279 = n19033 ^ n9731 ^ n6665 ;
  assign n21280 = ( ~n12409 & n19425 ) | ( ~n12409 & n21279 ) | ( n19425 & n21279 ) ;
  assign n21281 = ( n8939 & n20443 ) | ( n8939 & n21280 ) | ( n20443 & n21280 ) ;
  assign n21282 = n2686 & ~n3740 ;
  assign n21283 = ( n2952 & n4121 ) | ( n2952 & ~n21282 ) | ( n4121 & ~n21282 ) ;
  assign n21284 = ( n1085 & n8815 ) | ( n1085 & n15623 ) | ( n8815 & n15623 ) ;
  assign n21285 = ( n1580 & n6527 ) | ( n1580 & n21284 ) | ( n6527 & n21284 ) ;
  assign n21286 = n14212 ^ n14000 ^ n2454 ;
  assign n21287 = ( n1105 & n1551 ) | ( n1105 & n1855 ) | ( n1551 & n1855 ) ;
  assign n21288 = n21287 ^ n4271 ^ n698 ;
  assign n21289 = n21288 ^ n1696 ^ 1'b0 ;
  assign n21290 = n17208 & n21289 ;
  assign n21291 = ( n5218 & ~n7541 ) | ( n5218 & n8243 ) | ( ~n7541 & n8243 ) ;
  assign n21292 = n20715 ^ n15808 ^ n4493 ;
  assign n21293 = ( n433 & n21291 ) | ( n433 & n21292 ) | ( n21291 & n21292 ) ;
  assign n21294 = n4996 ^ n1141 ^ n352 ;
  assign n21295 = ( n3020 & n11287 ) | ( n3020 & n21149 ) | ( n11287 & n21149 ) ;
  assign n21298 = n7170 ^ n2556 ^ n662 ;
  assign n21299 = n21298 ^ n12572 ^ 1'b0 ;
  assign n21296 = ( n1488 & n6555 ) | ( n1488 & ~n9607 ) | ( n6555 & ~n9607 ) ;
  assign n21297 = ( n11684 & n18735 ) | ( n11684 & ~n21296 ) | ( n18735 & ~n21296 ) ;
  assign n21300 = n21299 ^ n21297 ^ n824 ;
  assign n21301 = ( n3802 & n11041 ) | ( n3802 & n14855 ) | ( n11041 & n14855 ) ;
  assign n21302 = n19199 ^ n18011 ^ n2382 ;
  assign n21303 = n9136 ^ n8530 ^ n5042 ;
  assign n21304 = n6582 ^ n2794 ^ 1'b0 ;
  assign n21305 = ~n21303 & n21304 ;
  assign n21306 = n18287 ^ n4039 ^ 1'b0 ;
  assign n21307 = n10171 & ~n21306 ;
  assign n21308 = n21307 ^ n19549 ^ 1'b0 ;
  assign n21309 = ( n3552 & ~n3780 ) | ( n3552 & n3898 ) | ( ~n3780 & n3898 ) ;
  assign n21310 = n21309 ^ n18910 ^ n12493 ;
  assign n21311 = ( ~n1167 & n8887 ) | ( ~n1167 & n21310 ) | ( n8887 & n21310 ) ;
  assign n21317 = n18304 ^ n12615 ^ n2340 ;
  assign n21313 = n5105 ^ n2039 ^ 1'b0 ;
  assign n21314 = ~n4829 & n21313 ;
  assign n21315 = ( n3382 & n4979 ) | ( n3382 & ~n5074 ) | ( n4979 & ~n5074 ) ;
  assign n21316 = ( n18620 & n21314 ) | ( n18620 & ~n21315 ) | ( n21314 & ~n21315 ) ;
  assign n21312 = ( n2503 & n5881 ) | ( n2503 & ~n7011 ) | ( n5881 & ~n7011 ) ;
  assign n21318 = n21317 ^ n21316 ^ n21312 ;
  assign n21320 = n19315 ^ n15994 ^ n7693 ;
  assign n21319 = n10673 ^ n9542 ^ n1840 ;
  assign n21321 = n21320 ^ n21319 ^ n17458 ;
  assign n21322 = n3520 | n7472 ;
  assign n21323 = n16065 | n21322 ;
  assign n21324 = n9373 ^ n4979 ^ n2661 ;
  assign n21325 = ( n15459 & ~n21323 ) | ( n15459 & n21324 ) | ( ~n21323 & n21324 ) ;
  assign n21326 = n7499 ^ n3085 ^ n2839 ;
  assign n21327 = n21326 ^ n5079 ^ n3338 ;
  assign n21328 = n21327 ^ n19812 ^ n18352 ;
  assign n21329 = n21328 ^ n9184 ^ n5651 ;
  assign n21330 = n20932 ^ n7768 ^ 1'b0 ;
  assign n21331 = ~n1105 & n21330 ;
  assign n21332 = n17155 ^ n12385 ^ n9930 ;
  assign n21333 = n9056 & ~n21332 ;
  assign n21334 = n18180 ^ n6833 ^ n326 ;
  assign n21335 = ( ~n20986 & n21333 ) | ( ~n20986 & n21334 ) | ( n21333 & n21334 ) ;
  assign n21336 = ( n1971 & n2902 ) | ( n1971 & ~n5588 ) | ( n2902 & ~n5588 ) ;
  assign n21337 = ( ~n1620 & n1898 ) | ( ~n1620 & n3428 ) | ( n1898 & n3428 ) ;
  assign n21338 = ( n638 & ~n2956 ) | ( n638 & n21337 ) | ( ~n2956 & n21337 ) ;
  assign n21339 = ( ~n7595 & n7929 ) | ( ~n7595 & n21338 ) | ( n7929 & n21338 ) ;
  assign n21340 = ( n2208 & ~n6864 ) | ( n2208 & n10463 ) | ( ~n6864 & n10463 ) ;
  assign n21341 = ( n610 & n11191 ) | ( n610 & n21340 ) | ( n11191 & n21340 ) ;
  assign n21342 = n9816 | n21341 ;
  assign n21343 = n21342 ^ n7519 ^ 1'b0 ;
  assign n21344 = ( n6467 & n21339 ) | ( n6467 & ~n21343 ) | ( n21339 & ~n21343 ) ;
  assign n21345 = n3398 & ~n3410 ;
  assign n21346 = n4067 & n21345 ;
  assign n21347 = ( ~n242 & n2637 ) | ( ~n242 & n4188 ) | ( n2637 & n4188 ) ;
  assign n21348 = ( n11422 & n15872 ) | ( n11422 & ~n21347 ) | ( n15872 & ~n21347 ) ;
  assign n21349 = ( ~n5155 & n21346 ) | ( ~n5155 & n21348 ) | ( n21346 & n21348 ) ;
  assign n21350 = n21349 ^ n20752 ^ n5194 ;
  assign n21352 = ( n4066 & n8057 ) | ( n4066 & n13437 ) | ( n8057 & n13437 ) ;
  assign n21351 = n15980 ^ n11166 ^ n7472 ;
  assign n21353 = n21352 ^ n21351 ^ n16676 ;
  assign n21354 = ( ~n8939 & n10878 ) | ( ~n8939 & n11472 ) | ( n10878 & n11472 ) ;
  assign n21355 = n14143 & n21354 ;
  assign n21356 = n21355 ^ n6436 ^ 1'b0 ;
  assign n21357 = ( n5448 & ~n15689 ) | ( n5448 & n21356 ) | ( ~n15689 & n21356 ) ;
  assign n21358 = ( n345 & n7475 ) | ( n345 & n7647 ) | ( n7475 & n7647 ) ;
  assign n21359 = ( x48 & n11229 ) | ( x48 & n21358 ) | ( n11229 & n21358 ) ;
  assign n21360 = n1879 & ~n10773 ;
  assign n21361 = n7757 & n21360 ;
  assign n21362 = ( n475 & n5515 ) | ( n475 & n21361 ) | ( n5515 & n21361 ) ;
  assign n21363 = ( x39 & n5282 ) | ( x39 & n21362 ) | ( n5282 & n21362 ) ;
  assign n21364 = n21363 ^ n5846 ^ n5380 ;
  assign n21365 = ( n5843 & n19225 ) | ( n5843 & n21364 ) | ( n19225 & n21364 ) ;
  assign n21366 = ( n1968 & ~n10703 ) | ( n1968 & n19337 ) | ( ~n10703 & n19337 ) ;
  assign n21367 = n16181 ^ n8951 ^ n1137 ;
  assign n21368 = ( x81 & n5014 ) | ( x81 & ~n7848 ) | ( n5014 & ~n7848 ) ;
  assign n21369 = n21368 ^ n10321 ^ n8864 ;
  assign n21370 = ( ~n7893 & n21367 ) | ( ~n7893 & n21369 ) | ( n21367 & n21369 ) ;
  assign n21372 = n5198 ^ n2500 ^ n400 ;
  assign n21371 = n13468 ^ n11736 ^ n8187 ;
  assign n21373 = n21372 ^ n21371 ^ n5483 ;
  assign n21374 = n17649 & ~n21373 ;
  assign n21375 = ( n5746 & n15084 ) | ( n5746 & ~n21374 ) | ( n15084 & ~n21374 ) ;
  assign n21376 = ( n3908 & ~n4650 ) | ( n3908 & n12992 ) | ( ~n4650 & n12992 ) ;
  assign n21377 = ( ~n9185 & n9464 ) | ( ~n9185 & n21376 ) | ( n9464 & n21376 ) ;
  assign n21378 = n15263 ^ n5594 ^ 1'b0 ;
  assign n21379 = n21378 ^ n19344 ^ n7116 ;
  assign n21381 = ( n1281 & n2486 ) | ( n1281 & n6887 ) | ( n2486 & n6887 ) ;
  assign n21380 = n20930 ^ n11933 ^ n10193 ;
  assign n21382 = n21381 ^ n21380 ^ n5315 ;
  assign n21383 = ( n2407 & n15188 ) | ( n2407 & n21382 ) | ( n15188 & n21382 ) ;
  assign n21384 = n12338 & n13330 ;
  assign n21385 = n21384 ^ n8717 ^ 1'b0 ;
  assign n21391 = n10544 ^ n6362 ^ n2340 ;
  assign n21392 = n15057 ^ n11060 ^ n1896 ;
  assign n21393 = ( n6516 & n21391 ) | ( n6516 & n21392 ) | ( n21391 & n21392 ) ;
  assign n21387 = n9392 ^ n3014 ^ n2793 ;
  assign n21388 = ( n2456 & ~n12505 ) | ( n2456 & n21387 ) | ( ~n12505 & n21387 ) ;
  assign n21389 = n14472 ^ n7737 ^ x93 ;
  assign n21390 = n21388 | n21389 ;
  assign n21386 = n6447 ^ n2184 ^ n1351 ;
  assign n21394 = n21393 ^ n21390 ^ n21386 ;
  assign n21395 = n9347 ^ n7051 ^ 1'b0 ;
  assign n21396 = n21395 ^ n5831 ^ n4062 ;
  assign n21397 = n13551 & ~n21396 ;
  assign n21398 = n1968 ^ n1503 ^ n1084 ;
  assign n21399 = ( n2589 & n17770 ) | ( n2589 & ~n21398 ) | ( n17770 & ~n21398 ) ;
  assign n21400 = n6790 ^ n3706 ^ 1'b0 ;
  assign n21401 = ~n11948 & n21400 ;
  assign n21402 = n21401 ^ n17229 ^ n13552 ;
  assign n21403 = ( n1813 & n9372 ) | ( n1813 & ~n13124 ) | ( n9372 & ~n13124 ) ;
  assign n21404 = n14406 & n21403 ;
  assign n21405 = n2953 & n21404 ;
  assign n21406 = n16118 ^ n11995 ^ 1'b0 ;
  assign n21407 = n21405 | n21406 ;
  assign n21408 = n21407 ^ n5498 ^ 1'b0 ;
  assign n21409 = n21408 ^ n15039 ^ n5475 ;
  assign n21410 = ~n5078 & n21409 ;
  assign n21411 = n20125 ^ n12531 ^ n5538 ;
  assign n21412 = ( ~n8530 & n10117 ) | ( ~n8530 & n21411 ) | ( n10117 & n21411 ) ;
  assign n21413 = n9760 ^ n9240 ^ n6504 ;
  assign n21414 = n1134 & ~n5559 ;
  assign n21415 = n21414 ^ n746 ^ 1'b0 ;
  assign n21416 = n21415 ^ n13688 ^ 1'b0 ;
  assign n21417 = ( n906 & n2757 ) | ( n906 & ~n10395 ) | ( n2757 & ~n10395 ) ;
  assign n21418 = ( n2466 & n3241 ) | ( n2466 & ~n21417 ) | ( n3241 & ~n21417 ) ;
  assign n21419 = ( ~n10871 & n12549 ) | ( ~n10871 & n16825 ) | ( n12549 & n16825 ) ;
  assign n21420 = n6055 ^ n5172 ^ 1'b0 ;
  assign n21421 = n21420 ^ n20531 ^ n11288 ;
  assign n21422 = ( n305 & n2570 ) | ( n305 & n8233 ) | ( n2570 & n8233 ) ;
  assign n21423 = n21422 ^ n5499 ^ 1'b0 ;
  assign n21424 = ( ~n5299 & n13830 ) | ( ~n5299 & n21423 ) | ( n13830 & n21423 ) ;
  assign n21425 = n21424 ^ n19774 ^ n10962 ;
  assign n21426 = ( ~n9633 & n9642 ) | ( ~n9633 & n11523 ) | ( n9642 & n11523 ) ;
  assign n21427 = ( n19504 & ~n21425 ) | ( n19504 & n21426 ) | ( ~n21425 & n21426 ) ;
  assign n21428 = n20040 ^ n2281 ^ n192 ;
  assign n21429 = ( n8596 & ~n14356 ) | ( n8596 & n21428 ) | ( ~n14356 & n21428 ) ;
  assign n21430 = ( n549 & ~n8438 ) | ( n549 & n9313 ) | ( ~n8438 & n9313 ) ;
  assign n21431 = n21430 ^ n15751 ^ n4767 ;
  assign n21432 = ( n9650 & ~n18176 ) | ( n9650 & n21431 ) | ( ~n18176 & n21431 ) ;
  assign n21433 = n21432 ^ n13096 ^ 1'b0 ;
  assign n21435 = n16327 ^ n129 ^ 1'b0 ;
  assign n21436 = n8526 & n21435 ;
  assign n21434 = ~n9351 & n18985 ;
  assign n21437 = n21436 ^ n21434 ^ 1'b0 ;
  assign n21438 = n14535 & ~n21437 ;
  assign n21439 = n8962 & n21438 ;
  assign n21440 = ( n814 & ~n1075 ) | ( n814 & n14280 ) | ( ~n1075 & n14280 ) ;
  assign n21441 = ( n5026 & n17736 ) | ( n5026 & ~n21440 ) | ( n17736 & ~n21440 ) ;
  assign n21442 = ( n4585 & ~n5027 ) | ( n4585 & n5991 ) | ( ~n5027 & n5991 ) ;
  assign n21443 = ( n1939 & n21228 ) | ( n1939 & ~n21442 ) | ( n21228 & ~n21442 ) ;
  assign n21444 = n8450 & ~n15020 ;
  assign n21446 = n9997 ^ n5659 ^ n2810 ;
  assign n21445 = ( n8525 & ~n10643 ) | ( n8525 & n17210 ) | ( ~n10643 & n17210 ) ;
  assign n21447 = n21446 ^ n21445 ^ n19931 ;
  assign n21448 = n21447 ^ n8684 ^ n6598 ;
  assign n21449 = n21082 ^ n12072 ^ 1'b0 ;
  assign n21450 = n18825 ^ n6896 ^ n6436 ;
  assign n21451 = n21450 ^ n6431 ^ n2877 ;
  assign n21452 = n21451 ^ n10833 ^ 1'b0 ;
  assign n21453 = ~n11503 & n21452 ;
  assign n21458 = n3577 ^ n2492 ^ n1808 ;
  assign n21455 = n16084 ^ n6458 ^ n6364 ;
  assign n21456 = ~n14682 & n21455 ;
  assign n21457 = n568 & n21456 ;
  assign n21454 = n9786 ^ n4046 ^ n3008 ;
  assign n21459 = n21458 ^ n21457 ^ n21454 ;
  assign n21462 = n15821 ^ n15272 ^ n12529 ;
  assign n21460 = n8917 ^ n1094 ^ n481 ;
  assign n21461 = n21460 ^ n9886 ^ n798 ;
  assign n21463 = n21462 ^ n21461 ^ n239 ;
  assign n21464 = ( n3043 & n5745 ) | ( n3043 & n7618 ) | ( n5745 & n7618 ) ;
  assign n21465 = ( ~n469 & n20882 ) | ( ~n469 & n21464 ) | ( n20882 & n21464 ) ;
  assign n21466 = ( ~n6143 & n18190 ) | ( ~n6143 & n21000 ) | ( n18190 & n21000 ) ;
  assign n21467 = n11950 ^ n8706 ^ n4247 ;
  assign n21468 = n6771 | n13910 ;
  assign n21469 = n16071 | n21468 ;
  assign n21470 = ( n1686 & ~n9861 ) | ( n1686 & n11061 ) | ( ~n9861 & n11061 ) ;
  assign n21471 = ( n4344 & n14778 ) | ( n4344 & n21470 ) | ( n14778 & n21470 ) ;
  assign n21472 = ~n361 & n814 ;
  assign n21473 = ( n3229 & n13441 ) | ( n3229 & ~n20701 ) | ( n13441 & ~n20701 ) ;
  assign n21474 = ( n549 & n2324 ) | ( n549 & ~n9533 ) | ( n2324 & ~n9533 ) ;
  assign n21475 = ( n910 & n11797 ) | ( n910 & ~n21474 ) | ( n11797 & ~n21474 ) ;
  assign n21476 = ( n7815 & ~n8489 ) | ( n7815 & n21475 ) | ( ~n8489 & n21475 ) ;
  assign n21477 = n21476 ^ n16568 ^ 1'b0 ;
  assign n21478 = n21477 ^ x92 ^ 1'b0 ;
  assign n21479 = n21473 & n21478 ;
  assign n21480 = ( ~n5811 & n11537 ) | ( ~n5811 & n13051 ) | ( n11537 & n13051 ) ;
  assign n21481 = n21480 ^ n18461 ^ n17757 ;
  assign n21482 = ( n21472 & n21479 ) | ( n21472 & ~n21481 ) | ( n21479 & ~n21481 ) ;
  assign n21483 = ( n1960 & n11810 ) | ( n1960 & n15587 ) | ( n11810 & n15587 ) ;
  assign n21484 = ( ~n3525 & n20226 ) | ( ~n3525 & n21483 ) | ( n20226 & n21483 ) ;
  assign n21485 = ( n8062 & ~n21482 ) | ( n8062 & n21484 ) | ( ~n21482 & n21484 ) ;
  assign n21486 = n11064 ^ n2754 ^ n2232 ;
  assign n21487 = ( ~n1385 & n4906 ) | ( ~n1385 & n6122 ) | ( n4906 & n6122 ) ;
  assign n21488 = ( ~n8129 & n21486 ) | ( ~n8129 & n21487 ) | ( n21486 & n21487 ) ;
  assign n21489 = n9953 ^ n9732 ^ n4388 ;
  assign n21490 = ( n1062 & n19144 ) | ( n1062 & n21489 ) | ( n19144 & n21489 ) ;
  assign n21491 = ( n5046 & n12336 ) | ( n5046 & ~n16547 ) | ( n12336 & ~n16547 ) ;
  assign n21492 = n21491 ^ n10624 ^ n2677 ;
  assign n21493 = n21492 ^ n10142 ^ n2539 ;
  assign n21494 = n3563 | n10115 ;
  assign n21495 = n21493 & ~n21494 ;
  assign n21496 = n20169 ^ n12270 ^ n10382 ;
  assign n21497 = n15228 ^ n9695 ^ n5059 ;
  assign n21498 = n21497 ^ n12947 ^ n7965 ;
  assign n21503 = n16228 ^ n6307 ^ 1'b0 ;
  assign n21499 = n4483 ^ n937 ^ x67 ;
  assign n21500 = n9547 ^ n7175 ^ n5054 ;
  assign n21501 = ( n6974 & n21499 ) | ( n6974 & n21500 ) | ( n21499 & n21500 ) ;
  assign n21502 = ( n12260 & ~n19435 ) | ( n12260 & n21501 ) | ( ~n19435 & n21501 ) ;
  assign n21504 = n21503 ^ n21502 ^ n6169 ;
  assign n21505 = ( n2073 & n5610 ) | ( n2073 & n6435 ) | ( n5610 & n6435 ) ;
  assign n21506 = ~n7563 & n16937 ;
  assign n21507 = n13065 & n21506 ;
  assign n21508 = ( x4 & n8062 ) | ( x4 & n16549 ) | ( n8062 & n16549 ) ;
  assign n21509 = ~n21507 & n21508 ;
  assign n21510 = n21505 | n21509 ;
  assign n21511 = ( n2717 & ~n3037 ) | ( n2717 & n19262 ) | ( ~n3037 & n19262 ) ;
  assign n21512 = n1884 ^ n683 ^ 1'b0 ;
  assign n21513 = n9777 & n21512 ;
  assign n21514 = ( n3184 & n5168 ) | ( n3184 & n21513 ) | ( n5168 & n21513 ) ;
  assign n21515 = ( ~n5611 & n17357 ) | ( ~n5611 & n21514 ) | ( n17357 & n21514 ) ;
  assign n21517 = n3051 | n6640 ;
  assign n21518 = n21517 ^ n1369 ^ 1'b0 ;
  assign n21516 = ( n3191 & n7707 ) | ( n3191 & n10348 ) | ( n7707 & n10348 ) ;
  assign n21519 = n21518 ^ n21516 ^ n3168 ;
  assign n21520 = ( ~n4100 & n17454 ) | ( ~n4100 & n21519 ) | ( n17454 & n21519 ) ;
  assign n21521 = ( n2309 & ~n2787 ) | ( n2309 & n21348 ) | ( ~n2787 & n21348 ) ;
  assign n21522 = n16351 ^ n8469 ^ n3120 ;
  assign n21523 = n21522 ^ n5061 ^ 1'b0 ;
  assign n21524 = n18476 ^ n5917 ^ n5364 ;
  assign n21525 = ( ~n7101 & n8614 ) | ( ~n7101 & n21524 ) | ( n8614 & n21524 ) ;
  assign n21526 = n21525 ^ n17284 ^ n582 ;
  assign n21527 = n17581 ^ n16215 ^ n410 ;
  assign n21528 = ( n14469 & ~n21526 ) | ( n14469 & n21527 ) | ( ~n21526 & n21527 ) ;
  assign n21529 = n12195 & ~n16264 ;
  assign n21530 = n9164 ^ n3102 ^ 1'b0 ;
  assign n21531 = n16949 & ~n21530 ;
  assign n21534 = n15274 ^ n7531 ^ n3082 ;
  assign n21533 = n11885 & n15254 ;
  assign n21535 = n21534 ^ n21533 ^ n4608 ;
  assign n21536 = ( n8562 & ~n14676 ) | ( n8562 & n21535 ) | ( ~n14676 & n21535 ) ;
  assign n21532 = n12828 ^ n3028 ^ x12 ;
  assign n21537 = n21536 ^ n21532 ^ n7132 ;
  assign n21538 = ( n3614 & ~n9329 ) | ( n3614 & n11798 ) | ( ~n9329 & n11798 ) ;
  assign n21539 = n12541 ^ n9570 ^ n9524 ;
  assign n21540 = n8089 ^ n2387 ^ 1'b0 ;
  assign n21541 = ( ~n2821 & n4483 ) | ( ~n2821 & n21540 ) | ( n4483 & n21540 ) ;
  assign n21542 = ( n21538 & ~n21539 ) | ( n21538 & n21541 ) | ( ~n21539 & n21541 ) ;
  assign n21543 = n7042 ^ n1202 ^ 1'b0 ;
  assign n21544 = ( n5622 & n19835 ) | ( n5622 & n21543 ) | ( n19835 & n21543 ) ;
  assign n21545 = ( ~n5622 & n11064 ) | ( ~n5622 & n21544 ) | ( n11064 & n21544 ) ;
  assign n21546 = n9178 ^ n4970 ^ n2973 ;
  assign n21547 = ( n19095 & ~n21545 ) | ( n19095 & n21546 ) | ( ~n21545 & n21546 ) ;
  assign n21549 = n12018 ^ n9614 ^ n834 ;
  assign n21548 = ( n3406 & ~n5799 ) | ( n3406 & n8006 ) | ( ~n5799 & n8006 ) ;
  assign n21550 = n21549 ^ n21548 ^ 1'b0 ;
  assign n21551 = n2400 & ~n21550 ;
  assign n21552 = ( n2436 & n4932 ) | ( n2436 & ~n8679 ) | ( n4932 & ~n8679 ) ;
  assign n21553 = n714 | n11798 ;
  assign n21554 = n21553 ^ n7230 ^ 1'b0 ;
  assign n21555 = n11272 ^ n3535 ^ n907 ;
  assign n21556 = n21555 ^ n5418 ^ n3944 ;
  assign n21557 = ( n19876 & n21554 ) | ( n19876 & n21556 ) | ( n21554 & n21556 ) ;
  assign n21558 = n21557 ^ n6343 ^ 1'b0 ;
  assign n21559 = ( n10386 & n21552 ) | ( n10386 & n21558 ) | ( n21552 & n21558 ) ;
  assign n21560 = n14931 ^ n11288 ^ n8773 ;
  assign n21561 = n21560 ^ n15331 ^ n6687 ;
  assign n21562 = ( n4742 & ~n14389 ) | ( n4742 & n21561 ) | ( ~n14389 & n21561 ) ;
  assign n21563 = n6445 ^ n6157 ^ n1956 ;
  assign n21564 = ( n637 & ~n14772 ) | ( n637 & n21563 ) | ( ~n14772 & n21563 ) ;
  assign n21565 = n5402 ^ n3826 ^ n1995 ;
  assign n21566 = ( n1610 & n16222 ) | ( n1610 & n21565 ) | ( n16222 & n21565 ) ;
  assign n21567 = n21287 ^ n12178 ^ n2674 ;
  assign n21568 = ( ~n1335 & n19915 ) | ( ~n1335 & n21567 ) | ( n19915 & n21567 ) ;
  assign n21569 = n21256 ^ n20289 ^ n1249 ;
  assign n21570 = n14791 ^ n8667 ^ n502 ;
  assign n21571 = n21570 ^ n12804 ^ n9533 ;
  assign n21572 = n21571 ^ n17062 ^ n9080 ;
  assign n21573 = n14174 ^ n3857 ^ 1'b0 ;
  assign n21574 = n12030 ^ n9520 ^ n1306 ;
  assign n21575 = n21574 ^ n2419 ^ 1'b0 ;
  assign n21577 = ( n543 & n793 ) | ( n543 & n17321 ) | ( n793 & n17321 ) ;
  assign n21576 = n1517 | n5872 ;
  assign n21578 = n21577 ^ n21576 ^ 1'b0 ;
  assign n21579 = ( ~n21573 & n21575 ) | ( ~n21573 & n21578 ) | ( n21575 & n21578 ) ;
  assign n21580 = ( ~n611 & n4335 ) | ( ~n611 & n5782 ) | ( n4335 & n5782 ) ;
  assign n21581 = n10893 | n21580 ;
  assign n21582 = n21581 ^ n16596 ^ 1'b0 ;
  assign n21583 = n21582 ^ n20848 ^ n8109 ;
  assign n21584 = n16103 ^ n10774 ^ n9715 ;
  assign n21587 = n11835 ^ n431 ^ 1'b0 ;
  assign n21588 = ~n6057 & n21587 ;
  assign n21589 = n21588 ^ n20151 ^ 1'b0 ;
  assign n21590 = ~n4628 & n21589 ;
  assign n21586 = n13927 ^ n198 ^ 1'b0 ;
  assign n21585 = ( n6182 & ~n10979 ) | ( n6182 & n13998 ) | ( ~n10979 & n13998 ) ;
  assign n21591 = n21590 ^ n21586 ^ n21585 ;
  assign n21592 = ( n172 & ~n536 ) | ( n172 & n7847 ) | ( ~n536 & n7847 ) ;
  assign n21593 = ( ~n11307 & n17637 ) | ( ~n11307 & n21592 ) | ( n17637 & n21592 ) ;
  assign n21594 = ( n3609 & ~n5211 ) | ( n3609 & n11760 ) | ( ~n5211 & n11760 ) ;
  assign n21595 = ( ~n10710 & n10883 ) | ( ~n10710 & n21594 ) | ( n10883 & n21594 ) ;
  assign n21596 = n15193 ^ n8670 ^ 1'b0 ;
  assign n21597 = n9731 & n21596 ;
  assign n21598 = ( n1587 & n4846 ) | ( n1587 & ~n12448 ) | ( n4846 & ~n12448 ) ;
  assign n21599 = n21597 & n21598 ;
  assign n21601 = ( ~n9178 & n9493 ) | ( ~n9178 & n15130 ) | ( n9493 & n15130 ) ;
  assign n21602 = ( n6668 & n11202 ) | ( n6668 & ~n21601 ) | ( n11202 & ~n21601 ) ;
  assign n21600 = ( n8493 & n18171 ) | ( n8493 & n20627 ) | ( n18171 & n20627 ) ;
  assign n21603 = n21602 ^ n21600 ^ n12421 ;
  assign n21604 = n14889 ^ n12411 ^ n7228 ;
  assign n21605 = ( n6536 & n8438 ) | ( n6536 & n13099 ) | ( n8438 & n13099 ) ;
  assign n21606 = n20353 ^ n8153 ^ n4969 ;
  assign n21607 = ( ~n7529 & n11741 ) | ( ~n7529 & n14976 ) | ( n11741 & n14976 ) ;
  assign n21608 = ( n13652 & n21606 ) | ( n13652 & n21607 ) | ( n21606 & n21607 ) ;
  assign n21609 = n3412 & n6941 ;
  assign n21610 = n21609 ^ n13619 ^ n9343 ;
  assign n21611 = n9604 ^ n3954 ^ n1372 ;
  assign n21612 = ( n8720 & n14637 ) | ( n8720 & n21611 ) | ( n14637 & n21611 ) ;
  assign n21613 = n14604 ^ n8074 ^ n7988 ;
  assign n21615 = n17020 ^ n242 ^ x117 ;
  assign n21614 = ( ~n4055 & n7496 ) | ( ~n4055 & n14073 ) | ( n7496 & n14073 ) ;
  assign n21616 = n21615 ^ n21614 ^ 1'b0 ;
  assign n21617 = n9714 & ~n20431 ;
  assign n21618 = n21617 ^ n11371 ^ 1'b0 ;
  assign n21619 = n19300 ^ n12967 ^ n9284 ;
  assign n21620 = ( n2504 & ~n4327 ) | ( n2504 & n9435 ) | ( ~n4327 & n9435 ) ;
  assign n21621 = n16713 ^ n4546 ^ n2047 ;
  assign n21622 = n21621 ^ n10893 ^ n8862 ;
  assign n21623 = ( n2706 & n14983 ) | ( n2706 & ~n21622 ) | ( n14983 & ~n21622 ) ;
  assign n21624 = n13116 ^ n13106 ^ 1'b0 ;
  assign n21625 = ( n585 & n1434 ) | ( n585 & n3970 ) | ( n1434 & n3970 ) ;
  assign n21626 = n21625 ^ n16371 ^ n2513 ;
  assign n21627 = n14983 ^ n14134 ^ n2120 ;
  assign n21628 = ( n4231 & n8528 ) | ( n4231 & ~n9759 ) | ( n8528 & ~n9759 ) ;
  assign n21629 = n16730 ^ n15203 ^ n10184 ;
  assign n21630 = ( n3270 & n3729 ) | ( n3270 & ~n17055 ) | ( n3729 & ~n17055 ) ;
  assign n21631 = ( n4144 & ~n7262 ) | ( n4144 & n21630 ) | ( ~n7262 & n21630 ) ;
  assign n21632 = ( n11948 & ~n21629 ) | ( n11948 & n21631 ) | ( ~n21629 & n21631 ) ;
  assign n21633 = ( n10175 & n12652 ) | ( n10175 & ~n19737 ) | ( n12652 & ~n19737 ) ;
  assign n21634 = n14840 ^ n9400 ^ n8605 ;
  assign n21635 = ( n9383 & n17579 ) | ( n9383 & n21634 ) | ( n17579 & n21634 ) ;
  assign n21636 = n13951 | n16031 ;
  assign n21637 = ~n6850 & n21636 ;
  assign n21638 = ~n12898 & n14564 ;
  assign n21639 = n21638 ^ n7237 ^ 1'b0 ;
  assign n21640 = n13793 ^ n10393 ^ n4983 ;
  assign n21641 = n21640 ^ n12812 ^ n10945 ;
  assign n21642 = ( ~n18539 & n19851 ) | ( ~n18539 & n21641 ) | ( n19851 & n21641 ) ;
  assign n21643 = n13852 ^ n3591 ^ n3310 ;
  assign n21644 = ( n4057 & ~n4146 ) | ( n4057 & n12610 ) | ( ~n4146 & n12610 ) ;
  assign n21645 = ( n6928 & ~n7710 ) | ( n6928 & n15793 ) | ( ~n7710 & n15793 ) ;
  assign n21646 = n7377 & ~n10186 ;
  assign n21647 = ( n12915 & n17658 ) | ( n12915 & ~n21646 ) | ( n17658 & ~n21646 ) ;
  assign n21648 = n11495 ^ n4594 ^ x61 ;
  assign n21649 = n21648 ^ n13319 ^ n5690 ;
  assign n21650 = n5985 ^ n144 ^ 1'b0 ;
  assign n21651 = n21649 & n21650 ;
  assign n21652 = n6135 ^ n3691 ^ n270 ;
  assign n21653 = ( n7445 & n11147 ) | ( n7445 & n21652 ) | ( n11147 & n21652 ) ;
  assign n21654 = n21653 ^ n18297 ^ n9854 ;
  assign n21656 = ( n1095 & n3625 ) | ( n1095 & n11135 ) | ( n3625 & n11135 ) ;
  assign n21655 = n13919 ^ n9696 ^ n7834 ;
  assign n21657 = n21656 ^ n21655 ^ n10767 ;
  assign n21658 = n13423 ^ n11552 ^ n6686 ;
  assign n21659 = ( ~n13450 & n15398 ) | ( ~n13450 & n21658 ) | ( n15398 & n21658 ) ;
  assign n21660 = n19319 & ~n21659 ;
  assign n21665 = ( ~n1521 & n3403 ) | ( ~n1521 & n12634 ) | ( n3403 & n12634 ) ;
  assign n21662 = ( n2046 & n12032 ) | ( n2046 & n18481 ) | ( n12032 & n18481 ) ;
  assign n21661 = n12244 & n17653 ;
  assign n21663 = n21662 ^ n21661 ^ 1'b0 ;
  assign n21664 = n21663 ^ n7739 ^ n6687 ;
  assign n21666 = n21665 ^ n21664 ^ n271 ;
  assign n21667 = n15887 | n21417 ;
  assign n21668 = n19296 ^ n14368 ^ n10014 ;
  assign n21669 = n21668 ^ n12177 ^ n12001 ;
  assign n21670 = n12767 ^ n3814 ^ 1'b0 ;
  assign n21671 = n19708 ^ n14819 ^ n12850 ;
  assign n21672 = n21671 ^ n14149 ^ n1571 ;
  assign n21673 = n14833 ^ n3924 ^ n3786 ;
  assign n21674 = ( n7134 & n13478 ) | ( n7134 & n21673 ) | ( n13478 & n21673 ) ;
  assign n21675 = ( n4706 & n17620 ) | ( n4706 & n21674 ) | ( n17620 & n21674 ) ;
  assign n21676 = n11478 ^ n6957 ^ n5869 ;
  assign n21677 = n1148 | n12132 ;
  assign n21678 = ( n6819 & ~n7079 ) | ( n6819 & n21677 ) | ( ~n7079 & n21677 ) ;
  assign n21679 = n20400 ^ n15596 ^ n1576 ;
  assign n21680 = n16066 & n21679 ;
  assign n21681 = n21680 ^ n15972 ^ n10404 ;
  assign n21682 = n21082 ^ n19765 ^ n11385 ;
  assign n21683 = ( n678 & n10636 ) | ( n678 & n21682 ) | ( n10636 & n21682 ) ;
  assign n21684 = ( n815 & ~n6642 ) | ( n815 & n6792 ) | ( ~n6642 & n6792 ) ;
  assign n21685 = ~n12858 & n18221 ;
  assign n21686 = n2781 & ~n18266 ;
  assign n21687 = ~n19409 & n21686 ;
  assign n21688 = n15827 ^ n12087 ^ n5080 ;
  assign n21689 = n17564 ^ n4250 ^ n822 ;
  assign n21690 = ( n6555 & ~n20022 ) | ( n6555 & n21689 ) | ( ~n20022 & n21689 ) ;
  assign n21691 = ( n1211 & ~n7832 ) | ( n1211 & n11450 ) | ( ~n7832 & n11450 ) ;
  assign n21692 = ( ~n2181 & n5986 ) | ( ~n2181 & n14190 ) | ( n5986 & n14190 ) ;
  assign n21693 = n10588 & ~n17555 ;
  assign n21694 = n6315 & n21693 ;
  assign n21695 = n16260 ^ n5893 ^ 1'b0 ;
  assign n21696 = ( n7660 & n11057 ) | ( n7660 & n15500 ) | ( n11057 & n15500 ) ;
  assign n21697 = ( ~n4772 & n21695 ) | ( ~n4772 & n21696 ) | ( n21695 & n21696 ) ;
  assign n21698 = n16967 ^ n14391 ^ n10345 ;
  assign n21699 = ( n20848 & ~n21477 ) | ( n20848 & n21698 ) | ( ~n21477 & n21698 ) ;
  assign n21700 = ( n8411 & n12913 ) | ( n8411 & n21699 ) | ( n12913 & n21699 ) ;
  assign n21701 = ( ~n2012 & n3743 ) | ( ~n2012 & n6653 ) | ( n3743 & n6653 ) ;
  assign n21702 = ( n5200 & n9795 ) | ( n5200 & ~n11537 ) | ( n9795 & ~n11537 ) ;
  assign n21703 = ( n462 & n9016 ) | ( n462 & n21702 ) | ( n9016 & n21702 ) ;
  assign n21704 = n21703 ^ n14110 ^ n1647 ;
  assign n21705 = n21701 & ~n21704 ;
  assign n21706 = n21705 ^ n18646 ^ n224 ;
  assign n21707 = n6004 ^ n3733 ^ n1785 ;
  assign n21708 = n21707 ^ n10632 ^ n961 ;
  assign n21709 = ( ~n7362 & n12188 ) | ( ~n7362 & n21708 ) | ( n12188 & n21708 ) ;
  assign n21710 = ( n382 & n1820 ) | ( n382 & ~n7071 ) | ( n1820 & ~n7071 ) ;
  assign n21711 = n21710 ^ n3127 ^ 1'b0 ;
  assign n21712 = n17915 ^ n12417 ^ n183 ;
  assign n21713 = ( n5091 & n21711 ) | ( n5091 & n21712 ) | ( n21711 & n21712 ) ;
  assign n21714 = n18530 ^ n2781 ^ n1650 ;
  assign n21717 = n7579 ^ n3969 ^ n1963 ;
  assign n21715 = n6622 ^ n5231 ^ 1'b0 ;
  assign n21716 = ( n13953 & ~n18556 ) | ( n13953 & n21715 ) | ( ~n18556 & n21715 ) ;
  assign n21718 = n21717 ^ n21716 ^ n1069 ;
  assign n21722 = n11442 ^ n8681 ^ n4727 ;
  assign n21719 = ( n4091 & n4334 ) | ( n4091 & n15206 ) | ( n4334 & n15206 ) ;
  assign n21720 = n21719 ^ n3628 ^ n660 ;
  assign n21721 = n21720 ^ n20162 ^ n14237 ;
  assign n21723 = n21722 ^ n21721 ^ n18873 ;
  assign n21724 = ( n410 & ~n4565 ) | ( n410 & n14314 ) | ( ~n4565 & n14314 ) ;
  assign n21725 = n21724 ^ n17869 ^ n7652 ;
  assign n21727 = ( n5062 & ~n8371 ) | ( n5062 & n17436 ) | ( ~n8371 & n17436 ) ;
  assign n21728 = n21727 ^ n2854 ^ n2701 ;
  assign n21726 = n21679 ^ n16056 ^ n12391 ;
  assign n21729 = n21728 ^ n21726 ^ n15544 ;
  assign n21730 = n7990 & n19033 ;
  assign n21731 = ~n283 & n21730 ;
  assign n21732 = n21731 ^ n18543 ^ n13177 ;
  assign n21733 = n13879 ^ n3548 ^ 1'b0 ;
  assign n21734 = ( n1480 & ~n13802 ) | ( n1480 & n21733 ) | ( ~n13802 & n21733 ) ;
  assign n21735 = n4565 ^ n1783 ^ 1'b0 ;
  assign n21736 = n6717 | n21735 ;
  assign n21737 = n21736 ^ n9467 ^ n3066 ;
  assign n21740 = ~n3392 & n7706 ;
  assign n21738 = n12789 & ~n21168 ;
  assign n21739 = n21738 ^ n6166 ^ 1'b0 ;
  assign n21741 = n21740 ^ n21739 ^ n7254 ;
  assign n21744 = ( n7827 & n11357 ) | ( n7827 & ~n19299 ) | ( n11357 & ~n19299 ) ;
  assign n21742 = ~n5442 & n13804 ;
  assign n21743 = ~n6243 & n21742 ;
  assign n21745 = n21744 ^ n21743 ^ n17519 ;
  assign n21746 = n11746 ^ n8107 ^ n6986 ;
  assign n21747 = n21746 ^ n7539 ^ n1598 ;
  assign n21748 = ~n8696 & n9127 ;
  assign n21749 = n8003 & n21748 ;
  assign n21750 = ( n13722 & n17188 ) | ( n13722 & n21749 ) | ( n17188 & n21749 ) ;
  assign n21751 = n14133 ^ n9956 ^ n312 ;
  assign n21752 = n1020 & n4676 ;
  assign n21753 = ( ~n2652 & n4234 ) | ( ~n2652 & n13404 ) | ( n4234 & n13404 ) ;
  assign n21754 = ( n16102 & n21752 ) | ( n16102 & ~n21753 ) | ( n21752 & ~n21753 ) ;
  assign n21755 = n21754 ^ n4344 ^ n375 ;
  assign n21756 = ( ~n2175 & n4130 ) | ( ~n2175 & n12294 ) | ( n4130 & n12294 ) ;
  assign n21757 = n21756 ^ n20475 ^ n18379 ;
  assign n21765 = ( n7725 & n8619 ) | ( n7725 & n16526 ) | ( n8619 & n16526 ) ;
  assign n21764 = ( n390 & n4036 ) | ( n390 & n17583 ) | ( n4036 & n17583 ) ;
  assign n21766 = n21765 ^ n21764 ^ n9555 ;
  assign n21763 = n5903 ^ n5625 ^ n2101 ;
  assign n21758 = n3107 ^ n2784 ^ n2682 ;
  assign n21759 = n21758 ^ n1431 ^ 1'b0 ;
  assign n21760 = ( ~n856 & n4122 ) | ( ~n856 & n21759 ) | ( n4122 & n21759 ) ;
  assign n21761 = n21760 ^ n16597 ^ n1049 ;
  assign n21762 = n21761 ^ n17977 ^ n10580 ;
  assign n21767 = n21766 ^ n21763 ^ n21762 ;
  assign n21768 = ( n9941 & n13578 ) | ( n9941 & n17956 ) | ( n13578 & n17956 ) ;
  assign n21769 = n21768 ^ n12846 ^ n6895 ;
  assign n21770 = ( ~n919 & n2402 ) | ( ~n919 & n21749 ) | ( n2402 & n21749 ) ;
  assign n21771 = ( x122 & n20183 ) | ( x122 & n21770 ) | ( n20183 & n21770 ) ;
  assign n21772 = n349 | n21771 ;
  assign n21773 = n21769 | n21772 ;
  assign n21774 = ( n9146 & n9193 ) | ( n9146 & ~n17663 ) | ( n9193 & ~n17663 ) ;
  assign n21775 = ( n11386 & n16371 ) | ( n11386 & ~n21774 ) | ( n16371 & ~n21774 ) ;
  assign n21776 = n21775 ^ n12645 ^ n7773 ;
  assign n21777 = n21776 ^ n21560 ^ n8372 ;
  assign n21778 = n14977 ^ n4593 ^ n2352 ;
  assign n21779 = ( n563 & n10659 ) | ( n563 & n21070 ) | ( n10659 & n21070 ) ;
  assign n21780 = n12816 ^ n11797 ^ n5074 ;
  assign n21781 = n16753 ^ n8854 ^ 1'b0 ;
  assign n21782 = ( n19160 & n21780 ) | ( n19160 & ~n21781 ) | ( n21780 & ~n21781 ) ;
  assign n21783 = ( n3965 & n5239 ) | ( n3965 & n21782 ) | ( n5239 & n21782 ) ;
  assign n21784 = ( n256 & n3141 ) | ( n256 & n9642 ) | ( n3141 & n9642 ) ;
  assign n21785 = n21784 ^ n11285 ^ n1620 ;
  assign n21786 = n21785 ^ n10357 ^ n9482 ;
  assign n21787 = n10635 ^ n4198 ^ n1703 ;
  assign n21788 = n15484 | n21787 ;
  assign n21789 = n21788 ^ n18413 ^ n4674 ;
  assign n21790 = n19199 & ~n21789 ;
  assign n21791 = ~n8106 & n21790 ;
  assign n21792 = n21791 ^ n17958 ^ 1'b0 ;
  assign n21793 = ( n5378 & n8716 ) | ( n5378 & n21792 ) | ( n8716 & n21792 ) ;
  assign n21794 = ( n4325 & ~n21786 ) | ( n4325 & n21793 ) | ( ~n21786 & n21793 ) ;
  assign n21795 = n5167 ^ n1867 ^ n285 ;
  assign n21796 = ( ~n6982 & n12071 ) | ( ~n6982 & n21795 ) | ( n12071 & n21795 ) ;
  assign n21797 = n5748 ^ n4982 ^ n1729 ;
  assign n21798 = n21797 ^ n9575 ^ n2977 ;
  assign n21799 = ( ~n3750 & n19255 ) | ( ~n3750 & n21798 ) | ( n19255 & n21798 ) ;
  assign n21800 = n12900 & ~n20885 ;
  assign n21801 = n13901 ^ n9217 ^ n4420 ;
  assign n21802 = ( n3150 & n5256 ) | ( n3150 & n7313 ) | ( n5256 & n7313 ) ;
  assign n21803 = n21802 ^ n8938 ^ n3583 ;
  assign n21804 = n21110 ^ n5066 ^ 1'b0 ;
  assign n21805 = ~n3667 & n21804 ;
  assign n21806 = ( ~n5942 & n21803 ) | ( ~n5942 & n21805 ) | ( n21803 & n21805 ) ;
  assign n21807 = ( ~n5508 & n15987 ) | ( ~n5508 & n21806 ) | ( n15987 & n21806 ) ;
  assign n21808 = ( n5066 & ~n13483 ) | ( n5066 & n21807 ) | ( ~n13483 & n21807 ) ;
  assign n21810 = n18237 ^ n13597 ^ n9514 ;
  assign n21809 = ( n645 & n10988 ) | ( n645 & ~n15248 ) | ( n10988 & ~n15248 ) ;
  assign n21811 = n21810 ^ n21809 ^ n1934 ;
  assign n21812 = n20956 ^ n19533 ^ n10724 ;
  assign n21813 = n13965 | n21812 ;
  assign n21814 = n21813 ^ n5746 ^ 1'b0 ;
  assign n21815 = ( ~n6751 & n7504 ) | ( ~n6751 & n21442 ) | ( n7504 & n21442 ) ;
  assign n21816 = n11235 ^ n2758 ^ 1'b0 ;
  assign n21817 = ( ~n1858 & n16988 ) | ( ~n1858 & n20197 ) | ( n16988 & n20197 ) ;
  assign n21818 = ( ~n3171 & n21816 ) | ( ~n3171 & n21817 ) | ( n21816 & n21817 ) ;
  assign n21819 = n15296 ^ n1957 ^ 1'b0 ;
  assign n21820 = n20688 ^ n7276 ^ n4793 ;
  assign n21821 = ( ~n19532 & n21819 ) | ( ~n19532 & n21820 ) | ( n21819 & n21820 ) ;
  assign n21822 = ( ~n14593 & n20674 ) | ( ~n14593 & n21821 ) | ( n20674 & n21821 ) ;
  assign n21823 = n14076 ^ n10105 ^ n1592 ;
  assign n21824 = n14803 ^ n12082 ^ n10519 ;
  assign n21825 = ( n5103 & n9159 ) | ( n5103 & ~n14136 ) | ( n9159 & ~n14136 ) ;
  assign n21826 = ( n8966 & ~n9721 ) | ( n8966 & n21825 ) | ( ~n9721 & n21825 ) ;
  assign n21827 = n15720 ^ n5231 ^ n3517 ;
  assign n21828 = n2656 | n21827 ;
  assign n21829 = n21828 ^ n692 ^ 1'b0 ;
  assign n21830 = n17407 ^ n7932 ^ n471 ;
  assign n21831 = n19237 ^ n8859 ^ 1'b0 ;
  assign n21832 = ( ~n2536 & n12316 ) | ( ~n2536 & n16758 ) | ( n12316 & n16758 ) ;
  assign n21833 = ( ~n16079 & n21831 ) | ( ~n16079 & n21832 ) | ( n21831 & n21832 ) ;
  assign n21834 = n21830 | n21833 ;
  assign n21835 = n8370 | n8736 ;
  assign n21836 = n21835 ^ n3983 ^ 1'b0 ;
  assign n21837 = n3541 ^ n3226 ^ n2122 ;
  assign n21838 = ( ~n812 & n3424 ) | ( ~n812 & n21837 ) | ( n3424 & n21837 ) ;
  assign n21839 = ( n6998 & n21836 ) | ( n6998 & n21838 ) | ( n21836 & n21838 ) ;
  assign n21840 = ~n2101 & n5291 ;
  assign n21841 = ( n1324 & n5863 ) | ( n1324 & n21840 ) | ( n5863 & n21840 ) ;
  assign n21842 = n21841 ^ n9872 ^ n9013 ;
  assign n21844 = n15226 ^ n10937 ^ n10276 ;
  assign n21845 = ( n2248 & ~n5015 ) | ( n2248 & n21844 ) | ( ~n5015 & n21844 ) ;
  assign n21843 = ( n1711 & ~n6301 ) | ( n1711 & n14286 ) | ( ~n6301 & n14286 ) ;
  assign n21846 = n21845 ^ n21843 ^ n21535 ;
  assign n21847 = ( ~n3235 & n13579 ) | ( ~n3235 & n21846 ) | ( n13579 & n21846 ) ;
  assign n21848 = n9937 ^ n2123 ^ 1'b0 ;
  assign n21849 = ( n3496 & n17214 ) | ( n3496 & n21848 ) | ( n17214 & n21848 ) ;
  assign n21850 = ~n8386 & n18942 ;
  assign n21851 = ~n21849 & n21850 ;
  assign n21852 = n21851 ^ n17357 ^ n3343 ;
  assign n21856 = n9708 ^ n3726 ^ n1729 ;
  assign n21853 = ~n5966 & n6775 ;
  assign n21854 = n14048 ^ n8715 ^ n6014 ;
  assign n21855 = ( n15345 & n21853 ) | ( n15345 & ~n21854 ) | ( n21853 & ~n21854 ) ;
  assign n21857 = n21856 ^ n21855 ^ x34 ;
  assign n21858 = ( n4680 & n10668 ) | ( n4680 & ~n17667 ) | ( n10668 & ~n17667 ) ;
  assign n21859 = n14528 ^ n13189 ^ n4836 ;
  assign n21860 = n19300 ^ n15233 ^ n1822 ;
  assign n21864 = ( n826 & n1836 ) | ( n826 & n10257 ) | ( n1836 & n10257 ) ;
  assign n21862 = ( n5369 & n6237 ) | ( n5369 & ~n13745 ) | ( n6237 & ~n13745 ) ;
  assign n21863 = n21862 ^ n20358 ^ n3521 ;
  assign n21861 = ( n8164 & n18994 ) | ( n8164 & ~n20061 ) | ( n18994 & ~n20061 ) ;
  assign n21865 = n21864 ^ n21863 ^ n21861 ;
  assign n21866 = n9584 ^ n5192 ^ 1'b0 ;
  assign n21867 = ( n1234 & n9684 ) | ( n1234 & ~n13935 ) | ( n9684 & ~n13935 ) ;
  assign n21868 = ( n2287 & n8820 ) | ( n2287 & n13770 ) | ( n8820 & n13770 ) ;
  assign n21869 = n8142 ^ n5549 ^ n1405 ;
  assign n21870 = ( n2471 & n6163 ) | ( n2471 & ~n14776 ) | ( n6163 & ~n14776 ) ;
  assign n21871 = ( n2038 & n9277 ) | ( n2038 & ~n21870 ) | ( n9277 & ~n21870 ) ;
  assign n21872 = n21871 ^ n5043 ^ 1'b0 ;
  assign n21873 = ~n12316 & n18673 ;
  assign n21874 = ( n3264 & ~n4126 ) | ( n3264 & n18164 ) | ( ~n4126 & n18164 ) ;
  assign n21875 = ( n1395 & n7851 ) | ( n1395 & ~n9607 ) | ( n7851 & ~n9607 ) ;
  assign n21876 = n21875 ^ n10729 ^ n5442 ;
  assign n21878 = ( n5463 & n12695 ) | ( n5463 & n13037 ) | ( n12695 & n13037 ) ;
  assign n21877 = ( ~n800 & n6229 ) | ( ~n800 & n13694 ) | ( n6229 & n13694 ) ;
  assign n21879 = n21878 ^ n21877 ^ n164 ;
  assign n21880 = n4895 ^ n4570 ^ n1585 ;
  assign n21881 = ~n8967 & n10306 ;
  assign n21882 = n21881 ^ n5472 ^ 1'b0 ;
  assign n21883 = ( n12442 & n13162 ) | ( n12442 & ~n21882 ) | ( n13162 & ~n21882 ) ;
  assign n21884 = n14915 & n16355 ;
  assign n21885 = n21884 ^ n8713 ^ n7038 ;
  assign n21886 = n15349 ^ n5101 ^ 1'b0 ;
  assign n21887 = n2957 & ~n21886 ;
  assign n21888 = n19184 ^ n14624 ^ n8059 ;
  assign n21889 = n8948 & ~n21888 ;
  assign n21890 = n2196 & n21889 ;
  assign n21891 = ~n9143 & n18743 ;
  assign n21892 = n21891 ^ n21809 ^ n20104 ;
  assign n21893 = ( n8486 & ~n10439 ) | ( n8486 & n14842 ) | ( ~n10439 & n14842 ) ;
  assign n21894 = ( n7372 & ~n7622 ) | ( n7372 & n19111 ) | ( ~n7622 & n19111 ) ;
  assign n21895 = n21894 ^ n10765 ^ n8191 ;
  assign n21896 = ~n21893 & n21895 ;
  assign n21900 = n19505 ^ n10783 ^ 1'b0 ;
  assign n21901 = ~n17112 & n21900 ;
  assign n21897 = ~n3885 & n16871 ;
  assign n21898 = ~n17502 & n21897 ;
  assign n21899 = n21898 ^ n15103 ^ n7484 ;
  assign n21902 = n21901 ^ n21899 ^ n13246 ;
  assign n21903 = n15331 & n20838 ;
  assign n21904 = ~n10134 & n21903 ;
  assign n21905 = n21904 ^ n18559 ^ n6351 ;
  assign n21906 = ( ~n234 & n10052 ) | ( ~n234 & n16597 ) | ( n10052 & n16597 ) ;
  assign n21907 = n19367 ^ n7465 ^ n201 ;
  assign n21908 = n3844 ^ n2542 ^ 1'b0 ;
  assign n21909 = n21908 ^ n8778 ^ n3835 ;
  assign n21910 = n3199 & n3626 ;
  assign n21911 = ~n21909 & n21910 ;
  assign n21912 = n21911 ^ n14708 ^ 1'b0 ;
  assign n21913 = ~n21907 & n21912 ;
  assign n21914 = n7233 ^ n3709 ^ 1'b0 ;
  assign n21915 = n7662 ^ n5902 ^ 1'b0 ;
  assign n21916 = n16845 | n21915 ;
  assign n21917 = ( ~n3128 & n12624 ) | ( ~n3128 & n21916 ) | ( n12624 & n21916 ) ;
  assign n21918 = ( n15718 & ~n21914 ) | ( n15718 & n21917 ) | ( ~n21914 & n21917 ) ;
  assign n21919 = ~n5204 & n9366 ;
  assign n21920 = n21919 ^ n11271 ^ 1'b0 ;
  assign n21921 = n12246 ^ n4578 ^ n3287 ;
  assign n21922 = n5838 | n5990 ;
  assign n21923 = n21922 ^ n3893 ^ n3034 ;
  assign n21928 = ( n5592 & ~n7143 ) | ( n5592 & n13918 ) | ( ~n7143 & n13918 ) ;
  assign n21924 = n7656 | n19052 ;
  assign n21925 = n9854 | n21924 ;
  assign n21926 = ( n3892 & ~n7276 ) | ( n3892 & n21925 ) | ( ~n7276 & n21925 ) ;
  assign n21927 = n21926 ^ n15801 ^ n13643 ;
  assign n21929 = n21928 ^ n21927 ^ n19668 ;
  assign n21930 = ( n14097 & n21923 ) | ( n14097 & n21929 ) | ( n21923 & n21929 ) ;
  assign n21931 = n18538 ^ n11734 ^ 1'b0 ;
  assign n21932 = n19755 ^ n19265 ^ n3430 ;
  assign n21933 = n8242 ^ n4770 ^ 1'b0 ;
  assign n21934 = n14476 & ~n21933 ;
  assign n21935 = ( n9267 & ~n18414 ) | ( n9267 & n21934 ) | ( ~n18414 & n21934 ) ;
  assign n21936 = ( ~n6894 & n10282 ) | ( ~n6894 & n21935 ) | ( n10282 & n21935 ) ;
  assign n21937 = n463 & ~n1299 ;
  assign n21938 = n21937 ^ n10580 ^ 1'b0 ;
  assign n21939 = n5634 ^ n1048 ^ 1'b0 ;
  assign n21940 = ~n10120 & n21939 ;
  assign n21941 = n21940 ^ n14368 ^ n3291 ;
  assign n21942 = n13077 ^ n12232 ^ n2848 ;
  assign n21943 = ( n2642 & ~n10282 ) | ( n2642 & n17760 ) | ( ~n10282 & n17760 ) ;
  assign n21944 = ~n4180 & n12539 ;
  assign n21945 = n21944 ^ n6715 ^ 1'b0 ;
  assign n21946 = ( n14655 & n21358 ) | ( n14655 & n21945 ) | ( n21358 & n21945 ) ;
  assign n21950 = n8352 ^ n6672 ^ n1169 ;
  assign n21951 = ( ~n6754 & n11154 ) | ( ~n6754 & n21950 ) | ( n11154 & n21950 ) ;
  assign n21952 = n21951 ^ n2814 ^ n2491 ;
  assign n21948 = ( n2012 & n3234 ) | ( n2012 & ~n5225 ) | ( n3234 & ~n5225 ) ;
  assign n21947 = n2114 ^ n2090 ^ n1876 ;
  assign n21949 = n21948 ^ n21947 ^ n1447 ;
  assign n21953 = n21952 ^ n21949 ^ n19955 ;
  assign n21956 = n19315 ^ n493 ^ 1'b0 ;
  assign n21957 = ~n7611 & n16040 ;
  assign n21958 = n21957 ^ n1762 ^ 1'b0 ;
  assign n21959 = ( ~n15325 & n21956 ) | ( ~n15325 & n21958 ) | ( n21956 & n21958 ) ;
  assign n21954 = ~n1172 & n13551 ;
  assign n21955 = ~n21856 & n21954 ;
  assign n21960 = n21959 ^ n21955 ^ n2335 ;
  assign n21961 = n16804 ^ n15090 ^ 1'b0 ;
  assign n21962 = ( n11672 & n21960 ) | ( n11672 & ~n21961 ) | ( n21960 & ~n21961 ) ;
  assign n21965 = ( ~n1446 & n11460 ) | ( ~n1446 & n17548 ) | ( n11460 & n17548 ) ;
  assign n21966 = n21965 ^ n1551 ^ 1'b0 ;
  assign n21963 = ( ~n2472 & n3115 ) | ( ~n2472 & n11540 ) | ( n3115 & n11540 ) ;
  assign n21964 = n3980 | n21963 ;
  assign n21967 = n21966 ^ n21964 ^ 1'b0 ;
  assign n21968 = n4007 ^ n1181 ^ n1076 ;
  assign n21969 = n21968 ^ n11035 ^ n7283 ;
  assign n21970 = n21834 ^ n16923 ^ 1'b0 ;
  assign n21971 = n21969 | n21970 ;
  assign n21972 = ( n4519 & ~n10578 ) | ( n4519 & n12627 ) | ( ~n10578 & n12627 ) ;
  assign n21973 = n668 & ~n2514 ;
  assign n21974 = n21973 ^ n7379 ^ n6740 ;
  assign n21975 = n21974 ^ n1130 ^ x93 ;
  assign n21978 = ( n1304 & n6562 ) | ( n1304 & ~n15982 ) | ( n6562 & ~n15982 ) ;
  assign n21979 = n4262 & n21978 ;
  assign n21980 = n21979 ^ n3616 ^ 1'b0 ;
  assign n21976 = n18410 ^ n16952 ^ 1'b0 ;
  assign n21977 = n6413 & ~n21976 ;
  assign n21981 = n21980 ^ n21977 ^ n15770 ;
  assign n21982 = n17433 ^ n4683 ^ n1260 ;
  assign n21983 = n21982 ^ n16228 ^ 1'b0 ;
  assign n21984 = n16987 ^ n16073 ^ n5774 ;
  assign n21985 = ( n10384 & ~n16684 ) | ( n10384 & n21984 ) | ( ~n16684 & n21984 ) ;
  assign n21986 = n12071 ^ n4182 ^ 1'b0 ;
  assign n21987 = n21985 & ~n21986 ;
  assign n21988 = ( n10741 & ~n20917 ) | ( n10741 & n21987 ) | ( ~n20917 & n21987 ) ;
  assign n21989 = n21988 ^ n16518 ^ n7381 ;
  assign n21990 = ( n6733 & n13194 ) | ( n6733 & ~n15187 ) | ( n13194 & ~n15187 ) ;
  assign n21991 = n18395 ^ n13498 ^ n8065 ;
  assign n21992 = n3503 & ~n4279 ;
  assign n21993 = ( n3613 & ~n21991 ) | ( n3613 & n21992 ) | ( ~n21991 & n21992 ) ;
  assign n21994 = n19637 ^ n17622 ^ 1'b0 ;
  assign n21995 = n4539 ^ n3158 ^ n2833 ;
  assign n21996 = n6502 ^ n2880 ^ x56 ;
  assign n21997 = n17190 ^ n9175 ^ n3109 ;
  assign n21998 = n528 & n9342 ;
  assign n21999 = ( n2147 & n16008 ) | ( n2147 & ~n21998 ) | ( n16008 & ~n21998 ) ;
  assign n22000 = ( n11191 & ~n13002 ) | ( n11191 & n19613 ) | ( ~n13002 & n19613 ) ;
  assign n22005 = ( n1671 & n1679 ) | ( n1671 & ~n2960 ) | ( n1679 & ~n2960 ) ;
  assign n22006 = ( ~n709 & n10566 ) | ( ~n709 & n22005 ) | ( n10566 & n22005 ) ;
  assign n22001 = n3019 & ~n16717 ;
  assign n22002 = n18124 & n22001 ;
  assign n22003 = ( n960 & n10395 ) | ( n960 & ~n22002 ) | ( n10395 & ~n22002 ) ;
  assign n22004 = ( n2864 & n5546 ) | ( n2864 & ~n22003 ) | ( n5546 & ~n22003 ) ;
  assign n22007 = n22006 ^ n22004 ^ n7884 ;
  assign n22008 = n15274 ^ n7120 ^ n3391 ;
  assign n22010 = n14389 ^ n13724 ^ n1232 ;
  assign n22009 = n14072 ^ n1617 ^ n1368 ;
  assign n22011 = n22010 ^ n22009 ^ n6832 ;
  assign n22012 = n543 & ~n22011 ;
  assign n22014 = ( n14041 & n17738 ) | ( n14041 & n21518 ) | ( n17738 & n21518 ) ;
  assign n22013 = ( n2349 & n5306 ) | ( n2349 & n5419 ) | ( n5306 & n5419 ) ;
  assign n22015 = n22014 ^ n22013 ^ n17500 ;
  assign n22016 = ( ~n169 & n536 ) | ( ~n169 & n11798 ) | ( n536 & n11798 ) ;
  assign n22017 = ( n1653 & ~n9559 ) | ( n1653 & n22016 ) | ( ~n9559 & n22016 ) ;
  assign n22018 = n19024 ^ n9967 ^ 1'b0 ;
  assign n22019 = ( n19406 & n22017 ) | ( n19406 & n22018 ) | ( n22017 & n22018 ) ;
  assign n22020 = n14753 ^ n13491 ^ n11754 ;
  assign n22021 = ( ~n923 & n14217 ) | ( ~n923 & n21324 ) | ( n14217 & n21324 ) ;
  assign n22022 = ( n7187 & ~n9571 ) | ( n7187 & n15585 ) | ( ~n9571 & n15585 ) ;
  assign n22023 = ( n1467 & n12876 ) | ( n1467 & n12995 ) | ( n12876 & n12995 ) ;
  assign n22024 = ( n11852 & ~n22022 ) | ( n11852 & n22023 ) | ( ~n22022 & n22023 ) ;
  assign n22025 = ( n8479 & n17997 ) | ( n8479 & n22024 ) | ( n17997 & n22024 ) ;
  assign n22026 = n10539 ^ n7216 ^ 1'b0 ;
  assign n22027 = n22026 ^ n21509 ^ n15597 ;
  assign n22028 = ( ~n11286 & n12102 ) | ( ~n11286 & n17682 ) | ( n12102 & n17682 ) ;
  assign n22029 = n15466 ^ n8528 ^ n3199 ;
  assign n22031 = n984 & n7072 ;
  assign n22032 = n11085 & n22031 ;
  assign n22030 = n12229 ^ n4644 ^ n971 ;
  assign n22033 = n22032 ^ n22030 ^ n21386 ;
  assign n22034 = n22033 ^ n18728 ^ n3479 ;
  assign n22035 = ( n4591 & ~n14301 ) | ( n4591 & n16550 ) | ( ~n14301 & n16550 ) ;
  assign n22036 = ( n1717 & n19037 ) | ( n1717 & ~n22035 ) | ( n19037 & ~n22035 ) ;
  assign n22037 = ( n9362 & ~n12570 ) | ( n9362 & n18898 ) | ( ~n12570 & n18898 ) ;
  assign n22038 = n22037 ^ n21831 ^ 1'b0 ;
  assign n22039 = ( n1795 & n4596 ) | ( n1795 & ~n5559 ) | ( n4596 & ~n5559 ) ;
  assign n22040 = n1637 ^ n253 ^ 1'b0 ;
  assign n22041 = n1891 & ~n22040 ;
  assign n22042 = ( n7309 & n14964 ) | ( n7309 & ~n22041 ) | ( n14964 & ~n22041 ) ;
  assign n22043 = ( n1445 & ~n13194 ) | ( n1445 & n22042 ) | ( ~n13194 & n22042 ) ;
  assign n22044 = n22043 ^ n7490 ^ n6860 ;
  assign n22045 = n13301 ^ n12294 ^ n2444 ;
  assign n22046 = n8142 | n14600 ;
  assign n22047 = n22046 ^ n1601 ^ 1'b0 ;
  assign n22048 = n726 | n22047 ;
  assign n22049 = ( n9528 & n9860 ) | ( n9528 & ~n13208 ) | ( n9860 & ~n13208 ) ;
  assign n22050 = n22049 ^ n15455 ^ 1'b0 ;
  assign n22051 = n22048 & n22050 ;
  assign n22053 = n8271 ^ n5639 ^ n1497 ;
  assign n22054 = ( n788 & ~n17748 ) | ( n788 & n22053 ) | ( ~n17748 & n22053 ) ;
  assign n22052 = ~n1537 & n12668 ;
  assign n22055 = n22054 ^ n22052 ^ n12146 ;
  assign n22056 = n6868 ^ n936 ^ n315 ;
  assign n22057 = n4820 | n7897 ;
  assign n22058 = n12376 ^ n10187 ^ n3055 ;
  assign n22059 = n10419 ^ n9543 ^ n3517 ;
  assign n22060 = n22059 ^ n4902 ^ n1172 ;
  assign n22061 = ( n5108 & n12965 ) | ( n5108 & ~n22060 ) | ( n12965 & ~n22060 ) ;
  assign n22062 = n3800 & n18508 ;
  assign n22063 = n22062 ^ n3145 ^ 1'b0 ;
  assign n22064 = ( ~n2870 & n14764 ) | ( ~n2870 & n22063 ) | ( n14764 & n22063 ) ;
  assign n22065 = n22061 | n22064 ;
  assign n22066 = n22065 ^ n310 ^ 1'b0 ;
  assign n22067 = n10879 ^ n1708 ^ n1257 ;
  assign n22068 = n9628 ^ n8269 ^ n3831 ;
  assign n22069 = ( n7394 & n15352 ) | ( n7394 & ~n22068 ) | ( n15352 & ~n22068 ) ;
  assign n22070 = n22069 ^ n3064 ^ 1'b0 ;
  assign n22071 = n22070 ^ n18537 ^ n341 ;
  assign n22072 = ( n20276 & n22067 ) | ( n20276 & n22071 ) | ( n22067 & n22071 ) ;
  assign n22073 = ( n22058 & n22066 ) | ( n22058 & ~n22072 ) | ( n22066 & ~n22072 ) ;
  assign n22074 = ~n3687 & n4183 ;
  assign n22075 = n22074 ^ n16166 ^ 1'b0 ;
  assign n22076 = n20246 ^ n15548 ^ 1'b0 ;
  assign n22077 = ( n2934 & ~n19701 ) | ( n2934 & n21431 ) | ( ~n19701 & n21431 ) ;
  assign n22078 = n10704 ^ n5843 ^ n716 ;
  assign n22079 = n22078 ^ n17554 ^ n957 ;
  assign n22080 = ( n2024 & ~n8073 ) | ( n2024 & n10650 ) | ( ~n8073 & n10650 ) ;
  assign n22081 = n10472 ^ n5260 ^ n3016 ;
  assign n22082 = n22081 ^ n8794 ^ n5900 ;
  assign n22083 = ( n3781 & ~n4822 ) | ( n3781 & n15555 ) | ( ~n4822 & n15555 ) ;
  assign n22084 = ( n15092 & n22082 ) | ( n15092 & n22083 ) | ( n22082 & n22083 ) ;
  assign n22085 = n7164 & ~n12264 ;
  assign n22086 = n22085 ^ n1182 ^ 1'b0 ;
  assign n22087 = n22086 ^ n14863 ^ n7407 ;
  assign n22088 = ( n2167 & n8178 ) | ( n2167 & ~n22087 ) | ( n8178 & ~n22087 ) ;
  assign n22089 = n7009 & n22088 ;
  assign n22090 = n22089 ^ n1921 ^ 1'b0 ;
  assign n22091 = ( n8226 & ~n8820 ) | ( n8226 & n15752 ) | ( ~n8820 & n15752 ) ;
  assign n22092 = ( n5275 & n9939 ) | ( n5275 & n19266 ) | ( n9939 & n19266 ) ;
  assign n22093 = n10053 ^ x82 ^ 1'b0 ;
  assign n22094 = n22093 ^ n8716 ^ n6491 ;
  assign n22095 = ( n16962 & n20496 ) | ( n16962 & n22094 ) | ( n20496 & n22094 ) ;
  assign n22096 = n13701 ^ n10905 ^ n4398 ;
  assign n22097 = n22096 ^ n20909 ^ 1'b0 ;
  assign n22098 = n9960 ^ n8742 ^ 1'b0 ;
  assign n22099 = n14416 ^ n8666 ^ n3681 ;
  assign n22100 = ( n877 & n5063 ) | ( n877 & n22099 ) | ( n5063 & n22099 ) ;
  assign n22101 = ~n13986 & n22100 ;
  assign n22102 = ~n17410 & n22101 ;
  assign n22108 = n19170 ^ n16853 ^ 1'b0 ;
  assign n22109 = n5338 & ~n22108 ;
  assign n22110 = n22109 ^ n12072 ^ 1'b0 ;
  assign n22107 = ( ~n410 & n4052 ) | ( ~n410 & n13649 ) | ( n4052 & n13649 ) ;
  assign n22103 = n3962 ^ n2360 ^ 1'b0 ;
  assign n22104 = ~n2785 & n22103 ;
  assign n22105 = ~n9279 & n22104 ;
  assign n22106 = n10623 & n22105 ;
  assign n22111 = n22110 ^ n22107 ^ n22106 ;
  assign n22112 = n7693 ^ n7414 ^ n4694 ;
  assign n22113 = ( n4838 & n5032 ) | ( n4838 & n11391 ) | ( n5032 & n11391 ) ;
  assign n22114 = ( n3310 & n14862 ) | ( n3310 & ~n22113 ) | ( n14862 & ~n22113 ) ;
  assign n22115 = n560 | n4158 ;
  assign n22116 = n22115 ^ n4660 ^ 1'b0 ;
  assign n22117 = n16669 ^ n8153 ^ 1'b0 ;
  assign n22118 = n16355 | n22117 ;
  assign n22119 = ( ~n3993 & n22116 ) | ( ~n3993 & n22118 ) | ( n22116 & n22118 ) ;
  assign n22120 = n13520 ^ n5625 ^ n4744 ;
  assign n22121 = n11184 & n16705 ;
  assign n22122 = n22121 ^ n12962 ^ n9628 ;
  assign n22123 = n19346 ^ n13652 ^ 1'b0 ;
  assign n22124 = ~n968 & n22123 ;
  assign n22125 = ( n5248 & n21312 ) | ( n5248 & ~n22124 ) | ( n21312 & ~n22124 ) ;
  assign n22126 = ( n2651 & ~n13737 ) | ( n2651 & n20212 ) | ( ~n13737 & n20212 ) ;
  assign n22127 = ( n812 & ~n9347 ) | ( n812 & n22126 ) | ( ~n9347 & n22126 ) ;
  assign n22128 = ( n2478 & ~n7805 ) | ( n2478 & n10186 ) | ( ~n7805 & n10186 ) ;
  assign n22129 = n22128 ^ n15478 ^ n12097 ;
  assign n22130 = n9114 & ~n13965 ;
  assign n22131 = n22130 ^ n335 ^ 1'b0 ;
  assign n22132 = ( ~n5838 & n14198 ) | ( ~n5838 & n22131 ) | ( n14198 & n22131 ) ;
  assign n22133 = n7107 ^ n5015 ^ n4099 ;
  assign n22134 = n12235 ^ n8998 ^ n8381 ;
  assign n22135 = n12840 ^ n5977 ^ n3064 ;
  assign n22136 = n7963 ^ n4071 ^ n1574 ;
  assign n22137 = ( ~n309 & n5044 ) | ( ~n309 & n22136 ) | ( n5044 & n22136 ) ;
  assign n22138 = ( ~n4550 & n18625 ) | ( ~n4550 & n20058 ) | ( n18625 & n20058 ) ;
  assign n22139 = ( ~n10416 & n11472 ) | ( ~n10416 & n17155 ) | ( n11472 & n17155 ) ;
  assign n22140 = ( ~n11507 & n18423 ) | ( ~n11507 & n22139 ) | ( n18423 & n22139 ) ;
  assign n22141 = n22140 ^ n16396 ^ n10962 ;
  assign n22142 = ( n22137 & ~n22138 ) | ( n22137 & n22141 ) | ( ~n22138 & n22141 ) ;
  assign n22143 = n19731 ^ n12231 ^ n11297 ;
  assign n22145 = n4612 ^ n2815 ^ n2760 ;
  assign n22146 = n22145 ^ n5042 ^ n340 ;
  assign n22144 = n10823 ^ n6579 ^ n5893 ;
  assign n22147 = n22146 ^ n22144 ^ 1'b0 ;
  assign n22148 = n14034 & ~n22147 ;
  assign n22149 = ( n9059 & n22143 ) | ( n9059 & n22148 ) | ( n22143 & n22148 ) ;
  assign n22150 = n7356 ^ n6677 ^ n4750 ;
  assign n22151 = n7879 ^ n5436 ^ 1'b0 ;
  assign n22152 = n22151 ^ n9329 ^ n4259 ;
  assign n22153 = ( n4739 & ~n22150 ) | ( n4739 & n22152 ) | ( ~n22150 & n22152 ) ;
  assign n22154 = n11456 ^ n8114 ^ n7722 ;
  assign n22155 = ( ~n4150 & n8629 ) | ( ~n4150 & n10148 ) | ( n8629 & n10148 ) ;
  assign n22156 = n2293 & n3833 ;
  assign n22157 = n9142 & n22156 ;
  assign n22158 = n22157 ^ n5949 ^ n5359 ;
  assign n22159 = ( n9704 & n22155 ) | ( n9704 & ~n22158 ) | ( n22155 & ~n22158 ) ;
  assign n22160 = ~n22154 & n22159 ;
  assign n22161 = n7417 & n22160 ;
  assign n22162 = n14494 ^ n3152 ^ 1'b0 ;
  assign n22163 = n239 & n22162 ;
  assign n22164 = ( ~n6448 & n6853 ) | ( ~n6448 & n11118 ) | ( n6853 & n11118 ) ;
  assign n22165 = ( n4465 & ~n5921 ) | ( n4465 & n22164 ) | ( ~n5921 & n22164 ) ;
  assign n22166 = ( n7985 & n10738 ) | ( n7985 & n22165 ) | ( n10738 & n22165 ) ;
  assign n22167 = ( n716 & n3170 ) | ( n716 & n6442 ) | ( n3170 & n6442 ) ;
  assign n22168 = ~n6093 & n22167 ;
  assign n22169 = n2609 & n6098 ;
  assign n22170 = ( n3565 & n7377 ) | ( n3565 & n22169 ) | ( n7377 & n22169 ) ;
  assign n22171 = n17392 ^ n12502 ^ n11963 ;
  assign n22172 = ( ~n2165 & n22170 ) | ( ~n2165 & n22171 ) | ( n22170 & n22171 ) ;
  assign n22173 = n20650 ^ n14828 ^ n8525 ;
  assign n22174 = ( n4230 & n5516 ) | ( n4230 & ~n10807 ) | ( n5516 & ~n10807 ) ;
  assign n22175 = n22174 ^ n1584 ^ x109 ;
  assign n22177 = n15840 ^ n8590 ^ 1'b0 ;
  assign n22178 = n3105 | n22177 ;
  assign n22179 = n12759 ^ n5235 ^ n4004 ;
  assign n22180 = ( ~n12403 & n14715 ) | ( ~n12403 & n22179 ) | ( n14715 & n22179 ) ;
  assign n22181 = ~n22178 & n22180 ;
  assign n22182 = ~n2463 & n22181 ;
  assign n22176 = n14446 ^ n3578 ^ n3222 ;
  assign n22183 = n22182 ^ n22176 ^ n454 ;
  assign n22184 = ( n2217 & n16079 ) | ( n2217 & n16829 ) | ( n16079 & n16829 ) ;
  assign n22185 = ( n3777 & n4048 ) | ( n3777 & n22184 ) | ( n4048 & n22184 ) ;
  assign n22186 = ( n1863 & n22183 ) | ( n1863 & ~n22185 ) | ( n22183 & ~n22185 ) ;
  assign n22187 = ( n278 & n1246 ) | ( n278 & n14660 ) | ( n1246 & n14660 ) ;
  assign n22190 = n4491 | n5382 ;
  assign n22189 = n13164 ^ n12039 ^ n11761 ;
  assign n22188 = n9878 ^ n3016 ^ n683 ;
  assign n22191 = n22190 ^ n22189 ^ n22188 ;
  assign n22192 = ( n132 & ~n4934 ) | ( n132 & n5705 ) | ( ~n4934 & n5705 ) ;
  assign n22193 = n16454 ^ n16144 ^ n11737 ;
  assign n22194 = n22193 ^ n523 ^ 1'b0 ;
  assign n22195 = ~n22192 & n22194 ;
  assign n22196 = ( n10481 & n13231 ) | ( n10481 & ~n19758 ) | ( n13231 & ~n19758 ) ;
  assign n22197 = ( n456 & ~n8462 ) | ( n456 & n22196 ) | ( ~n8462 & n22196 ) ;
  assign n22198 = ( n9568 & n22195 ) | ( n9568 & n22197 ) | ( n22195 & n22197 ) ;
  assign n22199 = ( n8611 & n17550 ) | ( n8611 & n18367 ) | ( n17550 & n18367 ) ;
  assign n22200 = n21560 ^ n3163 ^ 1'b0 ;
  assign n22201 = ( n2892 & n12703 ) | ( n2892 & ~n22179 ) | ( n12703 & ~n22179 ) ;
  assign n22202 = n22201 ^ n20952 ^ n17214 ;
  assign n22203 = n9299 ^ n8530 ^ 1'b0 ;
  assign n22204 = n3692 & n22203 ;
  assign n22205 = n18096 ^ n4843 ^ n1478 ;
  assign n22206 = ( n624 & ~n7288 ) | ( n624 & n10127 ) | ( ~n7288 & n10127 ) ;
  assign n22207 = n5424 ^ n2100 ^ 1'b0 ;
  assign n22208 = ( n16402 & n22206 ) | ( n16402 & n22207 ) | ( n22206 & n22207 ) ;
  assign n22209 = n22208 ^ n21447 ^ n15061 ;
  assign n22210 = n22064 ^ n18812 ^ n2052 ;
  assign n22211 = ( ~n13985 & n18378 ) | ( ~n13985 & n22210 ) | ( n18378 & n22210 ) ;
  assign n22212 = ~n281 & n22211 ;
  assign n22213 = n14614 ^ n10235 ^ n9302 ;
  assign n22217 = n5049 ^ n704 ^ 1'b0 ;
  assign n22218 = n22217 ^ n4482 ^ n1635 ;
  assign n22214 = ( n3277 & ~n3795 ) | ( n3277 & n19293 ) | ( ~n3795 & n19293 ) ;
  assign n22215 = ( n8764 & n20025 ) | ( n8764 & n22214 ) | ( n20025 & n22214 ) ;
  assign n22216 = ( n8205 & n15909 ) | ( n8205 & n22215 ) | ( n15909 & n22215 ) ;
  assign n22219 = n22218 ^ n22216 ^ n10571 ;
  assign n22220 = n22219 ^ n5960 ^ 1'b0 ;
  assign n22221 = ~n8625 & n22220 ;
  assign n22222 = n10744 & n22221 ;
  assign n22223 = ( n14592 & ~n22213 ) | ( n14592 & n22222 ) | ( ~n22213 & n22222 ) ;
  assign n22224 = ( n3123 & n9180 ) | ( n3123 & ~n14002 ) | ( n9180 & ~n14002 ) ;
  assign n22225 = n22224 ^ n18115 ^ n16326 ;
  assign n22226 = n581 | n3914 ;
  assign n22227 = n22226 ^ n5551 ^ 1'b0 ;
  assign n22228 = ( n2461 & n16618 ) | ( n2461 & ~n22227 ) | ( n16618 & ~n22227 ) ;
  assign n22229 = n22228 ^ n4047 ^ n1633 ;
  assign n22230 = n1315 & n19877 ;
  assign n22231 = ( ~n6309 & n7460 ) | ( ~n6309 & n18250 ) | ( n7460 & n18250 ) ;
  assign n22232 = n3181 ^ n992 ^ 1'b0 ;
  assign n22233 = n11835 | n22232 ;
  assign n22234 = ( n534 & n18781 ) | ( n534 & ~n22233 ) | ( n18781 & ~n22233 ) ;
  assign n22235 = n14900 ^ n12063 ^ 1'b0 ;
  assign n22236 = ~n5971 & n18979 ;
  assign n22237 = ( ~n2449 & n16677 ) | ( ~n2449 & n22236 ) | ( n16677 & n22236 ) ;
  assign n22239 = ( n6267 & ~n6970 ) | ( n6267 & n7109 ) | ( ~n6970 & n7109 ) ;
  assign n22240 = ( ~n9268 & n20635 ) | ( ~n9268 & n22239 ) | ( n20635 & n22239 ) ;
  assign n22238 = ( n4553 & n8777 ) | ( n4553 & n16470 ) | ( n8777 & n16470 ) ;
  assign n22241 = n22240 ^ n22238 ^ n21782 ;
  assign n22242 = ( n1735 & n2156 ) | ( n1735 & ~n22241 ) | ( n2156 & ~n22241 ) ;
  assign n22243 = n4896 ^ n4761 ^ n3343 ;
  assign n22244 = n19446 ^ n702 ^ 1'b0 ;
  assign n22245 = n17966 & n22244 ;
  assign n22246 = n20573 ^ n13967 ^ n1997 ;
  assign n22247 = n22043 ^ n13677 ^ n10085 ;
  assign n22250 = n9843 ^ n7076 ^ n3358 ;
  assign n22251 = ( n440 & n13882 ) | ( n440 & ~n22250 ) | ( n13882 & ~n22250 ) ;
  assign n22248 = n1097 & ~n8234 ;
  assign n22249 = n22248 ^ n16901 ^ 1'b0 ;
  assign n22252 = n22251 ^ n22249 ^ n16612 ;
  assign n22253 = n21715 ^ n2481 ^ n1531 ;
  assign n22254 = ( n11786 & n19865 ) | ( n11786 & n22253 ) | ( n19865 & n22253 ) ;
  assign n22255 = n13703 ^ n10016 ^ n8718 ;
  assign n22256 = n811 & n6625 ;
  assign n22257 = n22256 ^ n5204 ^ n1531 ;
  assign n22258 = ( n2297 & n3523 ) | ( n2297 & n3792 ) | ( n3523 & n3792 ) ;
  assign n22259 = n10151 & n17775 ;
  assign n22260 = ( ~n8302 & n22258 ) | ( ~n8302 & n22259 ) | ( n22258 & n22259 ) ;
  assign n22262 = n10622 ^ n5474 ^ 1'b0 ;
  assign n22263 = ( n3453 & n10720 ) | ( n3453 & n22262 ) | ( n10720 & n22262 ) ;
  assign n22261 = n856 & n3774 ;
  assign n22264 = n22263 ^ n22261 ^ 1'b0 ;
  assign n22265 = n12451 ^ n684 ^ 1'b0 ;
  assign n22266 = n22265 ^ n19844 ^ n5829 ;
  assign n22267 = n15659 ^ n6094 ^ 1'b0 ;
  assign n22268 = ( ~n1176 & n3713 ) | ( ~n1176 & n5316 ) | ( n3713 & n5316 ) ;
  assign n22269 = n2388 & n22268 ;
  assign n22270 = ~n22267 & n22269 ;
  assign n22271 = n20689 ^ n12561 ^ n5646 ;
  assign n22272 = ( n4725 & n9356 ) | ( n4725 & n22271 ) | ( n9356 & n22271 ) ;
  assign n22273 = ( n16582 & ~n22270 ) | ( n16582 & n22272 ) | ( ~n22270 & n22272 ) ;
  assign n22274 = n9595 ^ n2151 ^ n713 ;
  assign n22275 = n22274 ^ n2953 ^ 1'b0 ;
  assign n22276 = ( ~n5899 & n12054 ) | ( ~n5899 & n12139 ) | ( n12054 & n12139 ) ;
  assign n22277 = ( n3320 & n4380 ) | ( n3320 & n7619 ) | ( n4380 & n7619 ) ;
  assign n22278 = ( n15559 & ~n22276 ) | ( n15559 & n22277 ) | ( ~n22276 & n22277 ) ;
  assign n22279 = n13827 ^ n2797 ^ 1'b0 ;
  assign n22280 = ~n22278 & n22279 ;
  assign n22281 = ( n12480 & n21197 ) | ( n12480 & n22280 ) | ( n21197 & n22280 ) ;
  assign n22282 = ~n471 & n20706 ;
  assign n22283 = n22282 ^ n4955 ^ n2128 ;
  assign n22284 = ( n3217 & ~n10566 ) | ( n3217 & n22283 ) | ( ~n10566 & n22283 ) ;
  assign n22285 = ( n8535 & n14029 ) | ( n8535 & ~n20343 ) | ( n14029 & ~n20343 ) ;
  assign n22286 = n22285 ^ n15245 ^ n12102 ;
  assign n22287 = n14270 ^ n12177 ^ n7798 ;
  assign n22288 = n5274 | n22287 ;
  assign n22289 = n885 & n2755 ;
  assign n22290 = n22289 ^ n3234 ^ 1'b0 ;
  assign n22291 = n22290 ^ n13688 ^ n9124 ;
  assign n22292 = ( n2837 & n4104 ) | ( n2837 & n5713 ) | ( n4104 & n5713 ) ;
  assign n22293 = n13511 ^ n2774 ^ 1'b0 ;
  assign n22294 = n22293 ^ n7357 ^ 1'b0 ;
  assign n22295 = n16605 ^ n1472 ^ n452 ;
  assign n22296 = n7349 | n15997 ;
  assign n22297 = n22296 ^ n5508 ^ 1'b0 ;
  assign n22298 = n22297 ^ n11208 ^ n5875 ;
  assign n22299 = n3868 & ~n14899 ;
  assign n22300 = ( n6308 & n6333 ) | ( n6308 & ~n21968 ) | ( n6333 & ~n21968 ) ;
  assign n22301 = n22300 ^ n6014 ^ n671 ;
  assign n22302 = ( n11869 & n12607 ) | ( n11869 & ~n14684 ) | ( n12607 & ~n14684 ) ;
  assign n22303 = n12855 ^ n9000 ^ n603 ;
  assign n22304 = ( n6126 & ~n8310 ) | ( n6126 & n11636 ) | ( ~n8310 & n11636 ) ;
  assign n22305 = n15064 ^ n12124 ^ n7412 ;
  assign n22306 = n22305 ^ n6022 ^ n1705 ;
  assign n22307 = n16467 ^ n11923 ^ x34 ;
  assign n22308 = n3708 ^ n248 ^ 1'b0 ;
  assign n22309 = n22308 ^ n12687 ^ n8496 ;
  assign n22310 = n5187 & ~n9349 ;
  assign n22312 = n9065 ^ n8610 ^ n1739 ;
  assign n22311 = n14275 ^ n7341 ^ n4067 ;
  assign n22313 = n22312 ^ n22311 ^ n13523 ;
  assign n22314 = ~n2485 & n7278 ;
  assign n22315 = n8639 ^ n8197 ^ 1'b0 ;
  assign n22316 = n22315 ^ n11308 ^ n9736 ;
  assign n22317 = n22316 ^ n11448 ^ n3676 ;
  assign n22318 = n19398 ^ n10836 ^ n7027 ;
  assign n22320 = n11563 ^ n10943 ^ n1545 ;
  assign n22319 = ( n2594 & ~n3571 ) | ( n2594 & n6955 ) | ( ~n3571 & n6955 ) ;
  assign n22321 = n22320 ^ n22319 ^ n11519 ;
  assign n22322 = n21486 ^ n7468 ^ n3305 ;
  assign n22323 = n22322 ^ n8687 ^ n1300 ;
  assign n22324 = n7274 | n9053 ;
  assign n22325 = n12241 | n22324 ;
  assign n22326 = ( ~n2740 & n7080 ) | ( ~n2740 & n10645 ) | ( n7080 & n10645 ) ;
  assign n22327 = ( ~n4002 & n9450 ) | ( ~n4002 & n21698 ) | ( n9450 & n21698 ) ;
  assign n22328 = n4065 ^ n430 ^ x118 ;
  assign n22330 = ( n3060 & ~n6843 ) | ( n3060 & n20897 ) | ( ~n6843 & n20897 ) ;
  assign n22329 = ( n4707 & n10102 ) | ( n4707 & n13775 ) | ( n10102 & n13775 ) ;
  assign n22331 = n22330 ^ n22329 ^ n1401 ;
  assign n22332 = n20151 ^ n4930 ^ n193 ;
  assign n22333 = n7062 | n22332 ;
  assign n22335 = n14340 ^ n13367 ^ n10246 ;
  assign n22334 = ( n2462 & ~n7283 ) | ( n2462 & n11447 ) | ( ~n7283 & n11447 ) ;
  assign n22336 = n22335 ^ n22334 ^ n5758 ;
  assign n22337 = ( n4907 & n10234 ) | ( n4907 & ~n16887 ) | ( n10234 & ~n16887 ) ;
  assign n22338 = n3035 | n7656 ;
  assign n22339 = n14810 | n22338 ;
  assign n22340 = n6611 & n15192 ;
  assign n22341 = ~n10612 & n22340 ;
  assign n22342 = ( n3997 & n6384 ) | ( n3997 & n19161 ) | ( n6384 & n19161 ) ;
  assign n22346 = ( n1441 & n10390 ) | ( n1441 & n11880 ) | ( n10390 & n11880 ) ;
  assign n22347 = ( n5109 & n14216 ) | ( n5109 & ~n22346 ) | ( n14216 & ~n22346 ) ;
  assign n22343 = ( n2260 & ~n12709 ) | ( n2260 & n17739 ) | ( ~n12709 & n17739 ) ;
  assign n22344 = ( ~n855 & n2935 ) | ( ~n855 & n22343 ) | ( n2935 & n22343 ) ;
  assign n22345 = n22344 ^ n12343 ^ n4576 ;
  assign n22348 = n22347 ^ n22345 ^ 1'b0 ;
  assign n22349 = ( ~n11270 & n22342 ) | ( ~n11270 & n22348 ) | ( n22342 & n22348 ) ;
  assign n22350 = ( ~n1848 & n2952 ) | ( ~n1848 & n22349 ) | ( n2952 & n22349 ) ;
  assign n22351 = ( n639 & n20885 ) | ( n639 & ~n22350 ) | ( n20885 & ~n22350 ) ;
  assign n22352 = ( n7783 & n8052 ) | ( n7783 & n9953 ) | ( n8052 & n9953 ) ;
  assign n22353 = n22352 ^ n9911 ^ n6623 ;
  assign n22354 = ( n1860 & n9265 ) | ( n1860 & ~n22353 ) | ( n9265 & ~n22353 ) ;
  assign n22355 = ( ~n1485 & n8729 ) | ( ~n1485 & n22354 ) | ( n8729 & n22354 ) ;
  assign n22356 = ( x7 & n14960 ) | ( x7 & n22355 ) | ( n14960 & n22355 ) ;
  assign n22357 = ( n6863 & n19621 ) | ( n6863 & ~n22272 ) | ( n19621 & ~n22272 ) ;
  assign n22362 = n14920 ^ n4349 ^ n527 ;
  assign n22358 = ( n7539 & n9566 ) | ( n7539 & ~n13883 ) | ( n9566 & ~n13883 ) ;
  assign n22359 = ( ~n9451 & n11891 ) | ( ~n9451 & n22358 ) | ( n11891 & n22358 ) ;
  assign n22360 = n13314 & ~n22359 ;
  assign n22361 = n22360 ^ n15701 ^ n14284 ;
  assign n22363 = n22362 ^ n22361 ^ 1'b0 ;
  assign n22364 = n20781 ^ n20358 ^ n19713 ;
  assign n22365 = ( n403 & n472 ) | ( n403 & ~n20061 ) | ( n472 & ~n20061 ) ;
  assign n22366 = ( n6899 & n11799 ) | ( n6899 & n22365 ) | ( n11799 & n22365 ) ;
  assign n22367 = ~n22364 & n22366 ;
  assign n22370 = ( n2316 & n7829 ) | ( n2316 & n13585 ) | ( n7829 & n13585 ) ;
  assign n22368 = n874 & ~n7016 ;
  assign n22369 = ~n6738 & n22368 ;
  assign n22371 = n22370 ^ n22369 ^ 1'b0 ;
  assign n22372 = ~n452 & n22371 ;
  assign n22373 = n17132 ^ n9264 ^ n3665 ;
  assign n22374 = ~n18588 & n22373 ;
  assign n22375 = n20982 ^ n17607 ^ 1'b0 ;
  assign n22376 = ( x68 & n17235 ) | ( x68 & ~n22375 ) | ( n17235 & ~n22375 ) ;
  assign n22377 = n12799 ^ n9217 ^ 1'b0 ;
  assign n22378 = n22376 & ~n22377 ;
  assign n22379 = n20971 ^ n14889 ^ n1457 ;
  assign n22380 = ( n4472 & ~n22378 ) | ( n4472 & n22379 ) | ( ~n22378 & n22379 ) ;
  assign n22381 = n1038 ^ n253 ^ x93 ;
  assign n22382 = n22381 ^ n2929 ^ 1'b0 ;
  assign n22383 = n7665 ^ n457 ^ 1'b0 ;
  assign n22384 = n11413 ^ n10971 ^ n9506 ;
  assign n22385 = n2245 & n22384 ;
  assign n22386 = ( n15921 & n22383 ) | ( n15921 & ~n22385 ) | ( n22383 & ~n22385 ) ;
  assign n22387 = ( ~n12247 & n22382 ) | ( ~n12247 & n22386 ) | ( n22382 & n22386 ) ;
  assign n22388 = ( n1400 & ~n9125 ) | ( n1400 & n16147 ) | ( ~n9125 & n16147 ) ;
  assign n22389 = n15063 ^ n4457 ^ n799 ;
  assign n22390 = n20053 ^ n4944 ^ 1'b0 ;
  assign n22391 = n14402 ^ n3681 ^ 1'b0 ;
  assign n22392 = ~n18107 & n22391 ;
  assign n22393 = n21925 ^ n11799 ^ n10660 ;
  assign n22394 = n1882 & n3497 ;
  assign n22395 = n22394 ^ n6188 ^ n418 ;
  assign n22396 = n22395 ^ n10232 ^ n9417 ;
  assign n22397 = n14653 ^ n3374 ^ n1102 ;
  assign n22398 = n18826 ^ n1889 ^ n997 ;
  assign n22399 = n22398 ^ n6234 ^ n2569 ;
  assign n22400 = ( n1826 & n3466 ) | ( n1826 & n22399 ) | ( n3466 & n22399 ) ;
  assign n22401 = n8956 ^ n3834 ^ 1'b0 ;
  assign n22402 = n4110 & ~n22401 ;
  assign n22403 = n22402 ^ n7951 ^ n2980 ;
  assign n22404 = ( n22397 & n22400 ) | ( n22397 & ~n22403 ) | ( n22400 & ~n22403 ) ;
  assign n22405 = ( x48 & n1310 ) | ( x48 & n2581 ) | ( n1310 & n2581 ) ;
  assign n22406 = ( n1932 & n7488 ) | ( n1932 & ~n22405 ) | ( n7488 & ~n22405 ) ;
  assign n22407 = ( n3702 & n17505 ) | ( n3702 & n21586 ) | ( n17505 & n21586 ) ;
  assign n22408 = n5295 | n20602 ;
  assign n22409 = n17679 ^ n10061 ^ 1'b0 ;
  assign n22410 = n22408 & ~n22409 ;
  assign n22411 = n22410 ^ n13643 ^ n9737 ;
  assign n22412 = n2206 | n7586 ;
  assign n22413 = n12755 ^ n10371 ^ n1603 ;
  assign n22414 = n22413 ^ n19559 ^ n3438 ;
  assign n22415 = n5019 ^ n2952 ^ 1'b0 ;
  assign n22416 = n22414 | n22415 ;
  assign n22417 = n20945 ^ n15884 ^ 1'b0 ;
  assign n22418 = ( ~n10495 & n15531 ) | ( ~n10495 & n21376 ) | ( n15531 & n21376 ) ;
  assign n22419 = ( n6364 & n6713 ) | ( n6364 & n22418 ) | ( n6713 & n22418 ) ;
  assign n22420 = ( n1921 & ~n11906 ) | ( n1921 & n15325 ) | ( ~n11906 & n15325 ) ;
  assign n22421 = n5284 & ~n5645 ;
  assign n22422 = n22421 ^ n20396 ^ n2332 ;
  assign n22423 = n22422 ^ n6265 ^ n4313 ;
  assign n22424 = ( n11720 & n22420 ) | ( n11720 & ~n22423 ) | ( n22420 & ~n22423 ) ;
  assign n22425 = n22424 ^ n20971 ^ n13692 ;
  assign n22426 = n9462 ^ n5825 ^ n4696 ;
  assign n22427 = ( n3466 & n6357 ) | ( n3466 & n22426 ) | ( n6357 & n22426 ) ;
  assign n22428 = ( ~n498 & n2250 ) | ( ~n498 & n2682 ) | ( n2250 & n2682 ) ;
  assign n22429 = ( ~n16257 & n22427 ) | ( ~n16257 & n22428 ) | ( n22427 & n22428 ) ;
  assign n22432 = n18683 ^ n963 ^ x21 ;
  assign n22430 = ( n943 & ~n4160 ) | ( n943 & n9591 ) | ( ~n4160 & n9591 ) ;
  assign n22431 = n11985 & ~n22430 ;
  assign n22433 = n22432 ^ n22431 ^ n15216 ;
  assign n22434 = n10204 | n10480 ;
  assign n22435 = n22434 ^ n20764 ^ n7351 ;
  assign n22436 = n20010 ^ n10619 ^ 1'b0 ;
  assign n22437 = n11227 ^ n5396 ^ n1086 ;
  assign n22438 = ( n12163 & n19620 ) | ( n12163 & ~n22437 ) | ( n19620 & ~n22437 ) ;
  assign n22439 = n22436 & n22438 ;
  assign n22440 = n16364 & n22439 ;
  assign n22441 = n17095 ^ n6605 ^ 1'b0 ;
  assign n22442 = n6588 | n22441 ;
  assign n22443 = n5591 | n6894 ;
  assign n22444 = n10995 | n22443 ;
  assign n22445 = n22444 ^ n13716 ^ n11259 ;
  assign n22447 = n8223 ^ n4609 ^ n2381 ;
  assign n22448 = n22447 ^ n7454 ^ n1309 ;
  assign n22446 = n22287 ^ n857 ^ 1'b0 ;
  assign n22449 = n22448 ^ n22446 ^ n20768 ;
  assign n22450 = ( ~n9399 & n13346 ) | ( ~n9399 & n13967 ) | ( n13346 & n13967 ) ;
  assign n22458 = n1799 & n3683 ;
  assign n22459 = n22458 ^ n6489 ^ 1'b0 ;
  assign n22460 = n22459 ^ n7686 ^ n917 ;
  assign n22461 = ( ~n4019 & n12292 ) | ( ~n4019 & n22460 ) | ( n12292 & n22460 ) ;
  assign n22451 = n2894 ^ n563 ^ 1'b0 ;
  assign n22452 = n894 | n11161 ;
  assign n22453 = n22452 ^ n1055 ^ 1'b0 ;
  assign n22454 = ( n11545 & n12042 ) | ( n11545 & n22453 ) | ( n12042 & n22453 ) ;
  assign n22455 = n22454 ^ n13014 ^ n9006 ;
  assign n22456 = n22455 ^ n3422 ^ 1'b0 ;
  assign n22457 = n22451 | n22456 ;
  assign n22462 = n22461 ^ n22457 ^ n6624 ;
  assign n22463 = ( ~n5101 & n7133 ) | ( ~n5101 & n19688 ) | ( n7133 & n19688 ) ;
  assign n22464 = ( n11407 & n17269 ) | ( n11407 & n22463 ) | ( n17269 & n22463 ) ;
  assign n22465 = n4812 | n22464 ;
  assign n22466 = ( n2989 & n5719 ) | ( n2989 & ~n17314 ) | ( n5719 & ~n17314 ) ;
  assign n22467 = ( n1043 & n13221 ) | ( n1043 & ~n14002 ) | ( n13221 & ~n14002 ) ;
  assign n22468 = ( ~n5467 & n22466 ) | ( ~n5467 & n22467 ) | ( n22466 & n22467 ) ;
  assign n22469 = ( ~n1787 & n6035 ) | ( ~n1787 & n20499 ) | ( n6035 & n20499 ) ;
  assign n22474 = ( ~n2604 & n3117 ) | ( ~n2604 & n20001 ) | ( n3117 & n20001 ) ;
  assign n22471 = ~n943 & n6153 ;
  assign n22472 = n22471 ^ n8691 ^ n2402 ;
  assign n22470 = n18210 ^ n9376 ^ n4403 ;
  assign n22473 = n22472 ^ n22470 ^ n7382 ;
  assign n22475 = n22474 ^ n22473 ^ n18145 ;
  assign n22476 = ( n8885 & ~n13499 ) | ( n8885 & n15060 ) | ( ~n13499 & n15060 ) ;
  assign n22477 = n705 & ~n1895 ;
  assign n22478 = n22477 ^ n1012 ^ 1'b0 ;
  assign n22479 = ( n1668 & ~n16222 ) | ( n1668 & n22478 ) | ( ~n16222 & n22478 ) ;
  assign n22480 = ~n4510 & n22479 ;
  assign n22481 = ( n8033 & n18125 ) | ( n8033 & n22480 ) | ( n18125 & n22480 ) ;
  assign n22482 = n17630 ^ n14908 ^ n14614 ;
  assign n22483 = n20701 ^ n12340 ^ n169 ;
  assign n22484 = n22145 ^ n15057 ^ 1'b0 ;
  assign n22485 = n22484 ^ n18243 ^ n13316 ;
  assign n22486 = n3030 ^ n882 ^ 1'b0 ;
  assign n22487 = n4561 | n22486 ;
  assign n22488 = ( n1663 & n7887 ) | ( n1663 & ~n16977 ) | ( n7887 & ~n16977 ) ;
  assign n22489 = n4384 ^ n3686 ^ n3063 ;
  assign n22490 = n22489 ^ n18282 ^ n17649 ;
  assign n22491 = ( ~n3338 & n8411 ) | ( ~n3338 & n16526 ) | ( n8411 & n16526 ) ;
  assign n22492 = n19168 & ~n22491 ;
  assign n22493 = ( n5793 & ~n6765 ) | ( n5793 & n19590 ) | ( ~n6765 & n19590 ) ;
  assign n22494 = ( n5425 & ~n8321 ) | ( n5425 & n22493 ) | ( ~n8321 & n22493 ) ;
  assign n22495 = ( n7412 & n11731 ) | ( n7412 & n15922 ) | ( n11731 & n15922 ) ;
  assign n22496 = n17314 ^ n15901 ^ 1'b0 ;
  assign n22497 = n22496 ^ n19874 ^ n8848 ;
  assign n22498 = n22497 ^ n12858 ^ 1'b0 ;
  assign n22499 = n13492 ^ n5228 ^ n4996 ;
  assign n22500 = n10750 ^ n2371 ^ 1'b0 ;
  assign n22501 = x18 & ~n22500 ;
  assign n22502 = n11595 ^ n9738 ^ 1'b0 ;
  assign n22503 = n3674 | n22502 ;
  assign n22504 = ( ~n3169 & n9400 ) | ( ~n3169 & n18625 ) | ( n9400 & n18625 ) ;
  assign n22505 = n22504 ^ n9429 ^ n3521 ;
  assign n22506 = n16671 ^ n3310 ^ n1747 ;
  assign n22507 = ( n5036 & n6166 ) | ( n5036 & ~n12903 ) | ( n6166 & ~n12903 ) ;
  assign n22508 = n19850 ^ n11308 ^ n5941 ;
  assign n22509 = ( ~n7937 & n9223 ) | ( ~n7937 & n22508 ) | ( n9223 & n22508 ) ;
  assign n22510 = n22507 & n22509 ;
  assign n22511 = ( n168 & ~n9962 ) | ( n168 & n12309 ) | ( ~n9962 & n12309 ) ;
  assign n22512 = ( n7803 & ~n17143 ) | ( n7803 & n22511 ) | ( ~n17143 & n22511 ) ;
  assign n22513 = n22512 ^ n17967 ^ 1'b0 ;
  assign n22514 = ( n4626 & n6832 ) | ( n4626 & ~n9485 ) | ( n6832 & ~n9485 ) ;
  assign n22515 = ( n5243 & n10600 ) | ( n5243 & n19492 ) | ( n10600 & n19492 ) ;
  assign n22516 = n12030 & n13642 ;
  assign n22517 = n22516 ^ n14351 ^ 1'b0 ;
  assign n22518 = n8316 & n22517 ;
  assign n22519 = ~n4945 & n22518 ;
  assign n22520 = ~n1916 & n9314 ;
  assign n22521 = n17266 ^ n3922 ^ 1'b0 ;
  assign n22522 = ~n22520 & n22521 ;
  assign n22523 = ( n3462 & n10946 ) | ( n3462 & ~n11842 ) | ( n10946 & ~n11842 ) ;
  assign n22524 = n22523 ^ n7265 ^ n3211 ;
  assign n22525 = ( n14488 & ~n17886 ) | ( n14488 & n22524 ) | ( ~n17886 & n22524 ) ;
  assign n22530 = ( ~n5882 & n15834 ) | ( ~n5882 & n17288 ) | ( n15834 & n17288 ) ;
  assign n22528 = ( ~n2391 & n7064 ) | ( ~n2391 & n12386 ) | ( n7064 & n12386 ) ;
  assign n22526 = ( ~n6042 & n7440 ) | ( ~n6042 & n14959 ) | ( n7440 & n14959 ) ;
  assign n22527 = n22526 ^ n7207 ^ n4776 ;
  assign n22529 = n22528 ^ n22527 ^ n18060 ;
  assign n22531 = n22530 ^ n22529 ^ n14564 ;
  assign n22532 = n19161 ^ n13251 ^ n11177 ;
  assign n22536 = n12553 ^ n4704 ^ n1286 ;
  assign n22533 = n11377 ^ n4071 ^ 1'b0 ;
  assign n22534 = ( n2710 & n3797 ) | ( n2710 & n22533 ) | ( n3797 & n22533 ) ;
  assign n22535 = n22534 ^ n8712 ^ n3784 ;
  assign n22537 = n22536 ^ n22535 ^ n12642 ;
  assign n22538 = n20501 ^ n8774 ^ n417 ;
  assign n22539 = ~n1730 & n22538 ;
  assign n22540 = n8378 & n22539 ;
  assign n22541 = n1659 & n5260 ;
  assign n22542 = n22541 ^ n224 ^ 1'b0 ;
  assign n22543 = ( n12279 & n17119 ) | ( n12279 & n22047 ) | ( n17119 & n22047 ) ;
  assign n22544 = ( n15477 & ~n16057 ) | ( n15477 & n20227 ) | ( ~n16057 & n20227 ) ;
  assign n22545 = n14097 ^ n8269 ^ n4018 ;
  assign n22546 = ~n7065 & n15979 ;
  assign n22547 = n22546 ^ n13943 ^ 1'b0 ;
  assign n22548 = ( n1926 & n22545 ) | ( n1926 & n22547 ) | ( n22545 & n22547 ) ;
  assign n22549 = ( n4028 & n20716 ) | ( n4028 & ~n22548 ) | ( n20716 & ~n22548 ) ;
  assign n22550 = n6960 ^ n4858 ^ n3672 ;
  assign n22551 = ( n7405 & n10175 ) | ( n7405 & ~n22550 ) | ( n10175 & ~n22550 ) ;
  assign n22552 = n14700 & n17202 ;
  assign n22553 = n22552 ^ n21156 ^ 1'b0 ;
  assign n22554 = ( n2977 & n6340 ) | ( n2977 & ~n12832 ) | ( n6340 & ~n12832 ) ;
  assign n22555 = ( ~n774 & n8565 ) | ( ~n774 & n13974 ) | ( n8565 & n13974 ) ;
  assign n22556 = n14861 ^ n510 ^ 1'b0 ;
  assign n22557 = n1801 & ~n5671 ;
  assign n22558 = ( ~n22555 & n22556 ) | ( ~n22555 & n22557 ) | ( n22556 & n22557 ) ;
  assign n22559 = ( n16376 & n20935 ) | ( n16376 & n22558 ) | ( n20935 & n22558 ) ;
  assign n22561 = n16591 ^ n6949 ^ n5846 ;
  assign n22560 = n8903 ^ n3939 ^ n1511 ;
  assign n22562 = n22561 ^ n22560 ^ n3453 ;
  assign n22563 = n22562 ^ n8716 ^ n4474 ;
  assign n22564 = n18958 ^ n10820 ^ n10274 ;
  assign n22565 = n22564 ^ n7406 ^ n6991 ;
  assign n22566 = n22565 ^ n21381 ^ n344 ;
  assign n22571 = n3807 ^ n528 ^ n477 ;
  assign n22572 = ( n6926 & n12474 ) | ( n6926 & ~n22571 ) | ( n12474 & ~n22571 ) ;
  assign n22573 = n22572 ^ n15031 ^ n5634 ;
  assign n22567 = n15283 ^ n8163 ^ n4372 ;
  assign n22568 = ( n7283 & n15672 ) | ( n7283 & n22567 ) | ( n15672 & n22567 ) ;
  assign n22569 = n14157 | n22568 ;
  assign n22570 = n3138 & ~n22569 ;
  assign n22574 = n22573 ^ n22570 ^ n18288 ;
  assign n22577 = ( ~n798 & n5879 ) | ( ~n798 & n6764 ) | ( n5879 & n6764 ) ;
  assign n22578 = ( n7116 & n17501 ) | ( n7116 & n22577 ) | ( n17501 & n22577 ) ;
  assign n22575 = n8020 ^ n1978 ^ n519 ;
  assign n22576 = ( n4085 & n14894 ) | ( n4085 & n22575 ) | ( n14894 & n22575 ) ;
  assign n22579 = n22578 ^ n22576 ^ n12088 ;
  assign n22580 = n5525 ^ n1909 ^ n1557 ;
  assign n22581 = ( ~n12232 & n20781 ) | ( ~n12232 & n22580 ) | ( n20781 & n22580 ) ;
  assign n22582 = n4648 & n14031 ;
  assign n22583 = n16660 & n22582 ;
  assign n22584 = ( ~n21088 & n22581 ) | ( ~n21088 & n22583 ) | ( n22581 & n22583 ) ;
  assign n22585 = n18739 ^ n13564 ^ n8567 ;
  assign n22586 = n10547 | n22585 ;
  assign n22587 = n22586 ^ n5683 ^ 1'b0 ;
  assign n22588 = n7230 & ~n17254 ;
  assign n22589 = n9163 ^ n3777 ^ 1'b0 ;
  assign n22590 = n12983 ^ n772 ^ 1'b0 ;
  assign n22591 = n9570 | n10449 ;
  assign n22592 = n226 | n22591 ;
  assign n22593 = ( n22589 & n22590 ) | ( n22589 & ~n22592 ) | ( n22590 & ~n22592 ) ;
  assign n22594 = n10395 ^ n5912 ^ 1'b0 ;
  assign n22595 = ( n8294 & n16154 ) | ( n8294 & n22594 ) | ( n16154 & n22594 ) ;
  assign n22596 = n8193 & ~n8736 ;
  assign n22597 = n22596 ^ n12685 ^ 1'b0 ;
  assign n22598 = ( ~n5540 & n8608 ) | ( ~n5540 & n8768 ) | ( n8608 & n8768 ) ;
  assign n22599 = n22598 ^ n10995 ^ n5944 ;
  assign n22600 = n22599 ^ n13266 ^ n10683 ;
  assign n22601 = ( n18182 & ~n22597 ) | ( n18182 & n22600 ) | ( ~n22597 & n22600 ) ;
  assign n22605 = ( n4266 & ~n4656 ) | ( n4266 & n16118 ) | ( ~n4656 & n16118 ) ;
  assign n22602 = ( n3409 & n5658 ) | ( n3409 & ~n7442 ) | ( n5658 & ~n7442 ) ;
  assign n22603 = ( n255 & n13432 ) | ( n255 & ~n22602 ) | ( n13432 & ~n22602 ) ;
  assign n22604 = n22603 ^ n19900 ^ n16684 ;
  assign n22606 = n22605 ^ n22604 ^ n1534 ;
  assign n22607 = n22463 ^ n9749 ^ n2705 ;
  assign n22610 = n3788 & n8015 ;
  assign n22611 = n22610 ^ n7713 ^ n1706 ;
  assign n22612 = n22611 ^ n18177 ^ n17302 ;
  assign n22608 = n11018 ^ n6145 ^ n2778 ;
  assign n22609 = ( ~n10371 & n15209 ) | ( ~n10371 & n22608 ) | ( n15209 & n22608 ) ;
  assign n22613 = n22612 ^ n22609 ^ n3145 ;
  assign n22614 = n22613 ^ n21500 ^ n9464 ;
  assign n22615 = n21958 ^ n12017 ^ n5066 ;
  assign n22616 = n467 & n6534 ;
  assign n22617 = n22616 ^ n17450 ^ 1'b0 ;
  assign n22618 = ( ~n2494 & n17883 ) | ( ~n2494 & n22617 ) | ( n17883 & n22617 ) ;
  assign n22625 = ( n3524 & ~n4232 ) | ( n3524 & n12665 ) | ( ~n4232 & n12665 ) ;
  assign n22626 = ( n5524 & n11716 ) | ( n5524 & n22625 ) | ( n11716 & n22625 ) ;
  assign n22624 = n4304 | n15648 ;
  assign n22627 = n22626 ^ n22624 ^ n5709 ;
  assign n22620 = n12281 ^ n10912 ^ n2314 ;
  assign n22619 = n8460 ^ n7260 ^ n681 ;
  assign n22621 = n22620 ^ n22619 ^ n9739 ;
  assign n22622 = ~n17062 & n22621 ;
  assign n22623 = ( n422 & ~n14966 ) | ( n422 & n22622 ) | ( ~n14966 & n22622 ) ;
  assign n22628 = n22627 ^ n22623 ^ n867 ;
  assign n22629 = n21074 ^ n7364 ^ 1'b0 ;
  assign n22630 = n2605 & n22629 ;
  assign n22631 = n2073 ^ n307 ^ 1'b0 ;
  assign n22632 = n794 & n4358 ;
  assign n22633 = ( n9390 & n22631 ) | ( n9390 & ~n22632 ) | ( n22631 & ~n22632 ) ;
  assign n22634 = ( n647 & n18203 ) | ( n647 & ~n22633 ) | ( n18203 & ~n22633 ) ;
  assign n22635 = ( ~n376 & n3420 ) | ( ~n376 & n4313 ) | ( n3420 & n4313 ) ;
  assign n22636 = n17461 ^ n13617 ^ n7162 ;
  assign n22637 = n22635 & n22636 ;
  assign n22638 = n12844 ^ n11754 ^ n7056 ;
  assign n22639 = ( ~n219 & n1523 ) | ( ~n219 & n19319 ) | ( n1523 & n19319 ) ;
  assign n22640 = ( n3745 & ~n11447 ) | ( n3745 & n18918 ) | ( ~n11447 & n18918 ) ;
  assign n22645 = n18620 ^ n1033 ^ 1'b0 ;
  assign n22641 = n15248 ^ n9170 ^ n5299 ;
  assign n22642 = n13621 ^ n7460 ^ n2215 ;
  assign n22643 = n22642 ^ n19959 ^ n19424 ;
  assign n22644 = ( n13279 & n22641 ) | ( n13279 & n22643 ) | ( n22641 & n22643 ) ;
  assign n22646 = n22645 ^ n22644 ^ 1'b0 ;
  assign n22647 = ( n8162 & ~n22640 ) | ( n8162 & n22646 ) | ( ~n22640 & n22646 ) ;
  assign n22648 = n3195 ^ n2847 ^ n2379 ;
  assign n22649 = n9215 ^ n7903 ^ n442 ;
  assign n22650 = ~n8339 & n18912 ;
  assign n22651 = ~n22649 & n22650 ;
  assign n22652 = n9435 ^ n2207 ^ n2012 ;
  assign n22653 = n7813 & ~n22652 ;
  assign n22654 = ( n1666 & n16596 ) | ( n1666 & ~n22653 ) | ( n16596 & ~n22653 ) ;
  assign n22655 = ( n5402 & n22611 ) | ( n5402 & n22654 ) | ( n22611 & n22654 ) ;
  assign n22656 = n22201 ^ n4473 ^ n2727 ;
  assign n22657 = n8804 ^ n4146 ^ 1'b0 ;
  assign n22658 = n12818 & n22657 ;
  assign n22659 = ( ~n12751 & n13077 ) | ( ~n12751 & n22658 ) | ( n13077 & n22658 ) ;
  assign n22660 = ( ~n3771 & n6733 ) | ( ~n3771 & n22659 ) | ( n6733 & n22659 ) ;
  assign n22661 = n2137 & ~n19086 ;
  assign n22662 = n22661 ^ n16124 ^ n2349 ;
  assign n22663 = ( n4492 & ~n5042 ) | ( n4492 & n9740 ) | ( ~n5042 & n9740 ) ;
  assign n22664 = n22663 ^ n12343 ^ n3855 ;
  assign n22665 = n10970 | n22664 ;
  assign n22666 = n4445 ^ n1061 ^ n474 ;
  assign n22669 = n5625 ^ n1837 ^ x105 ;
  assign n22667 = n11740 ^ n8770 ^ n8262 ;
  assign n22668 = n22667 ^ n10753 ^ n6947 ;
  assign n22670 = n22669 ^ n22668 ^ n962 ;
  assign n22671 = ( n11758 & n22666 ) | ( n11758 & ~n22670 ) | ( n22666 & ~n22670 ) ;
  assign n22672 = ( n2396 & n12615 ) | ( n2396 & n15082 ) | ( n12615 & n15082 ) ;
  assign n22673 = n18874 ^ n10611 ^ n521 ;
  assign n22674 = ~n4964 & n22673 ;
  assign n22675 = n14030 ^ n10678 ^ n4264 ;
  assign n22676 = n7360 & n8376 ;
  assign n22677 = n22676 ^ n20431 ^ n1103 ;
  assign n22678 = ( n5673 & n22675 ) | ( n5673 & ~n22677 ) | ( n22675 & ~n22677 ) ;
  assign n22679 = n14646 ^ n13355 ^ n8621 ;
  assign n22680 = n6568 & n16168 ;
  assign n22681 = ~n12363 & n22680 ;
  assign n22682 = ( n13860 & n22679 ) | ( n13860 & n22681 ) | ( n22679 & n22681 ) ;
  assign n22683 = ( n8740 & n13056 ) | ( n8740 & n22682 ) | ( n13056 & n22682 ) ;
  assign n22684 = n22683 ^ n12403 ^ n2378 ;
  assign n22685 = n13350 ^ n4468 ^ n2749 ;
  assign n22686 = ( n17793 & n18221 ) | ( n17793 & n22685 ) | ( n18221 & n22685 ) ;
  assign n22687 = ( n11955 & ~n20888 ) | ( n11955 & n22686 ) | ( ~n20888 & n22686 ) ;
  assign n22689 = n12669 ^ n510 ^ n502 ;
  assign n22688 = n14950 ^ n6607 ^ 1'b0 ;
  assign n22690 = n22689 ^ n22688 ^ n7495 ;
  assign n22691 = n22690 ^ n18388 ^ n8000 ;
  assign n22692 = n22691 ^ n18168 ^ n17213 ;
  assign n22693 = n2877 ^ n2630 ^ 1'b0 ;
  assign n22694 = n270 & n22693 ;
  assign n22695 = ( ~n5447 & n20033 ) | ( ~n5447 & n22694 ) | ( n20033 & n22694 ) ;
  assign n22697 = n1881 & ~n3429 ;
  assign n22698 = ( ~n7567 & n13294 ) | ( ~n7567 & n22697 ) | ( n13294 & n22697 ) ;
  assign n22696 = ( n11939 & n15257 ) | ( n11939 & n18429 ) | ( n15257 & n18429 ) ;
  assign n22699 = n22698 ^ n22696 ^ 1'b0 ;
  assign n22700 = n525 & ~n22699 ;
  assign n22701 = ( n3874 & ~n6283 ) | ( n3874 & n9726 ) | ( ~n6283 & n9726 ) ;
  assign n22702 = ( n13873 & n17604 ) | ( n13873 & ~n22701 ) | ( n17604 & ~n22701 ) ;
  assign n22704 = n9646 & n14160 ;
  assign n22703 = n20381 ^ n7661 ^ n3578 ;
  assign n22705 = n22704 ^ n22703 ^ n11500 ;
  assign n22706 = ( n6269 & n7730 ) | ( n6269 & n20185 ) | ( n7730 & n20185 ) ;
  assign n22707 = ( n394 & n8148 ) | ( n394 & ~n22706 ) | ( n8148 & ~n22706 ) ;
  assign n22708 = n22707 ^ n14754 ^ n14579 ;
  assign n22709 = n22708 ^ n11856 ^ n6926 ;
  assign n22710 = n2373 & n7562 ;
  assign n22711 = n22710 ^ n12582 ^ 1'b0 ;
  assign n22712 = ( n7237 & ~n8020 ) | ( n7237 & n22711 ) | ( ~n8020 & n22711 ) ;
  assign n22713 = n13617 ^ n5720 ^ n3251 ;
  assign n22714 = n22713 ^ n19732 ^ n1134 ;
  assign n22715 = ( n2007 & ~n5050 ) | ( n2007 & n7981 ) | ( ~n5050 & n7981 ) ;
  assign n22716 = n22715 ^ n8282 ^ 1'b0 ;
  assign n22717 = n7616 ^ n4044 ^ 1'b0 ;
  assign n22719 = n3827 & ~n4397 ;
  assign n22720 = ( n587 & n5067 ) | ( n587 & ~n22719 ) | ( n5067 & ~n22719 ) ;
  assign n22721 = ( n2680 & n12173 ) | ( n2680 & ~n22720 ) | ( n12173 & ~n22720 ) ;
  assign n22718 = n14467 ^ n12802 ^ n3558 ;
  assign n22722 = n22721 ^ n22718 ^ n2727 ;
  assign n22724 = n15357 ^ n3339 ^ n251 ;
  assign n22725 = n293 | n22724 ;
  assign n22726 = n22725 ^ n21109 ^ 1'b0 ;
  assign n22723 = n6876 | n12018 ;
  assign n22727 = n22726 ^ n22723 ^ n7859 ;
  assign n22733 = n3572 ^ n3519 ^ n559 ;
  assign n22728 = n11206 ^ n4335 ^ n1438 ;
  assign n22729 = ( n446 & n1859 ) | ( n446 & ~n22728 ) | ( n1859 & ~n22728 ) ;
  assign n22730 = ( n1741 & n13047 ) | ( n1741 & ~n19666 ) | ( n13047 & ~n19666 ) ;
  assign n22731 = n5439 & n22730 ;
  assign n22732 = n22729 & n22731 ;
  assign n22734 = n22733 ^ n22732 ^ n10127 ;
  assign n22735 = n9897 ^ n6821 ^ n4254 ;
  assign n22736 = n11684 ^ n11024 ^ n7233 ;
  assign n22737 = n16284 ^ n4554 ^ 1'b0 ;
  assign n22738 = n9200 & ~n22737 ;
  assign n22739 = ( ~n22735 & n22736 ) | ( ~n22735 & n22738 ) | ( n22736 & n22738 ) ;
  assign n22740 = n1173 & ~n9022 ;
  assign n22741 = n22740 ^ n5225 ^ 1'b0 ;
  assign n22742 = n22741 ^ n15986 ^ n1667 ;
  assign n22743 = n12768 ^ n5054 ^ 1'b0 ;
  assign n22744 = n12027 ^ n3280 ^ 1'b0 ;
  assign n22745 = ~n2339 & n22744 ;
  assign n22746 = n20603 ^ n4022 ^ n2281 ;
  assign n22747 = ( n2820 & n8575 ) | ( n2820 & n21067 ) | ( n8575 & n21067 ) ;
  assign n22748 = ( n2581 & ~n12815 ) | ( n2581 & n22747 ) | ( ~n12815 & n22747 ) ;
  assign n22749 = n22748 ^ n19249 ^ n475 ;
  assign n22750 = n10844 ^ n4138 ^ n3620 ;
  assign n22751 = ( n2547 & n14987 ) | ( n2547 & n22750 ) | ( n14987 & n22750 ) ;
  assign n22752 = ~n4683 & n13953 ;
  assign n22753 = ( ~n12086 & n13700 ) | ( ~n12086 & n22752 ) | ( n13700 & n22752 ) ;
  assign n22754 = n8162 ^ n2897 ^ n1558 ;
  assign n22760 = n6326 ^ n4414 ^ 1'b0 ;
  assign n22761 = ( n3843 & ~n11272 ) | ( n3843 & n22760 ) | ( ~n11272 & n22760 ) ;
  assign n22762 = n22761 ^ n9185 ^ n2357 ;
  assign n22755 = n2700 ^ n1878 ^ n1739 ;
  assign n22756 = ~n19922 & n22755 ;
  assign n22757 = ( ~n1606 & n10468 ) | ( ~n1606 & n22756 ) | ( n10468 & n22756 ) ;
  assign n22758 = n22757 ^ n4481 ^ 1'b0 ;
  assign n22759 = n22758 ^ n16021 ^ n2449 ;
  assign n22763 = n22762 ^ n22759 ^ n16689 ;
  assign n22764 = ( x123 & n1523 ) | ( x123 & n10741 ) | ( n1523 & n10741 ) ;
  assign n22765 = ( ~n2551 & n15283 ) | ( ~n2551 & n22764 ) | ( n15283 & n22764 ) ;
  assign n22766 = n17028 ^ n2511 ^ n1882 ;
  assign n22767 = ( n8825 & ~n16155 ) | ( n8825 & n22766 ) | ( ~n16155 & n22766 ) ;
  assign n22768 = n19919 ^ n19033 ^ n6137 ;
  assign n22769 = n7480 & ~n22768 ;
  assign n22770 = n22769 ^ n411 ^ 1'b0 ;
  assign n22771 = n17298 ^ n11992 ^ n6270 ;
  assign n22775 = ( n5340 & n5507 ) | ( n5340 & ~n10766 ) | ( n5507 & ~n10766 ) ;
  assign n22773 = n17463 ^ n1826 ^ 1'b0 ;
  assign n22772 = n20868 & n22082 ;
  assign n22774 = n22773 ^ n22772 ^ x68 ;
  assign n22776 = n22775 ^ n22774 ^ n22497 ;
  assign n22777 = n3694 ^ n867 ^ x30 ;
  assign n22778 = n9786 & n22777 ;
  assign n22779 = n16888 ^ n10745 ^ n3404 ;
  assign n22780 = n18352 ^ n9790 ^ n511 ;
  assign n22781 = n22780 ^ n18269 ^ 1'b0 ;
  assign n22782 = n10749 | n22781 ;
  assign n22783 = n12551 & ~n22782 ;
  assign n22784 = n22783 ^ n14162 ^ 1'b0 ;
  assign n22785 = ( n2255 & n2378 ) | ( n2255 & n19286 ) | ( n2378 & n19286 ) ;
  assign n22786 = n22785 ^ n17732 ^ n1797 ;
  assign n22787 = n2891 & n22786 ;
  assign n22788 = ( ~n8064 & n10897 ) | ( ~n8064 & n13071 ) | ( n10897 & n13071 ) ;
  assign n22789 = n14053 ^ n5463 ^ n4660 ;
  assign n22790 = ~n661 & n22789 ;
  assign n22791 = ~n14493 & n22790 ;
  assign n22792 = n22788 & n22791 ;
  assign n22793 = ~n1227 & n22170 ;
  assign n22794 = n7527 & ~n22782 ;
  assign n22795 = n22794 ^ n16352 ^ n5011 ;
  assign n22796 = n16393 ^ n7691 ^ n3612 ;
  assign n22797 = ( n6590 & n20069 ) | ( n6590 & n22796 ) | ( n20069 & n22796 ) ;
  assign n22798 = n14165 ^ n852 ^ x46 ;
  assign n22799 = ( n12429 & ~n18600 ) | ( n12429 & n22798 ) | ( ~n18600 & n22798 ) ;
  assign n22800 = ( n9685 & n13244 ) | ( n9685 & ~n22799 ) | ( n13244 & ~n22799 ) ;
  assign n22801 = ( n650 & n4011 ) | ( n650 & n9774 ) | ( n4011 & n9774 ) ;
  assign n22802 = n22801 ^ n10265 ^ n790 ;
  assign n22807 = n9001 ^ n4935 ^ n4862 ;
  assign n22808 = ( n3337 & n10600 ) | ( n3337 & ~n22807 ) | ( n10600 & ~n22807 ) ;
  assign n22809 = n22808 ^ n18645 ^ n9391 ;
  assign n22806 = n15839 ^ n3325 ^ n1335 ;
  assign n22803 = n9890 ^ n9312 ^ n5143 ;
  assign n22804 = ( n1570 & n10073 ) | ( n1570 & n21960 ) | ( n10073 & n21960 ) ;
  assign n22805 = ( n12584 & n22803 ) | ( n12584 & n22804 ) | ( n22803 & n22804 ) ;
  assign n22810 = n22809 ^ n22806 ^ n22805 ;
  assign n22811 = ( n2158 & ~n3371 ) | ( n2158 & n8696 ) | ( ~n3371 & n8696 ) ;
  assign n22812 = n22811 ^ n956 ^ 1'b0 ;
  assign n22813 = n22812 ^ n16215 ^ n1830 ;
  assign n22814 = n22813 ^ n9376 ^ n7345 ;
  assign n22815 = ( n15448 & ~n15636 ) | ( n15448 & n21045 ) | ( ~n15636 & n21045 ) ;
  assign n22816 = n22384 ^ n8685 ^ n363 ;
  assign n22817 = ( n2465 & ~n22815 ) | ( n2465 & n22816 ) | ( ~n22815 & n22816 ) ;
  assign n22818 = ( n3132 & ~n4372 ) | ( n3132 & n7144 ) | ( ~n4372 & n7144 ) ;
  assign n22819 = n22818 ^ n17676 ^ n10347 ;
  assign n22820 = n22819 ^ n8538 ^ n6399 ;
  assign n22821 = n22820 ^ n19602 ^ n2111 ;
  assign n22822 = n2050 & ~n9964 ;
  assign n22823 = n4007 | n9282 ;
  assign n22824 = n18152 | n22823 ;
  assign n22825 = n22824 ^ n9276 ^ 1'b0 ;
  assign n22826 = n8745 | n22825 ;
  assign n22827 = n22826 ^ n20754 ^ 1'b0 ;
  assign n22828 = ( n9284 & n22822 ) | ( n9284 & ~n22827 ) | ( n22822 & ~n22827 ) ;
  assign n22829 = ~n2601 & n8591 ;
  assign n22830 = n22829 ^ n1283 ^ n571 ;
  assign n22831 = n17541 ^ n8697 ^ n3959 ;
  assign n22832 = n22831 ^ n11986 ^ n11472 ;
  assign n22833 = n14902 ^ n9654 ^ n5570 ;
  assign n22834 = n13370 ^ n2400 ^ 1'b0 ;
  assign n22835 = n8706 | n22834 ;
  assign n22836 = n22835 ^ n18773 ^ n9506 ;
  assign n22837 = ( n539 & n16925 ) | ( n539 & n22836 ) | ( n16925 & n22836 ) ;
  assign n22838 = ( n11835 & ~n22833 ) | ( n11835 & n22837 ) | ( ~n22833 & n22837 ) ;
  assign n22839 = ( n1758 & n2766 ) | ( n1758 & n16801 ) | ( n2766 & n16801 ) ;
  assign n22840 = n7353 & ~n14931 ;
  assign n22841 = n22840 ^ n18615 ^ 1'b0 ;
  assign n22842 = ( n12251 & ~n22839 ) | ( n12251 & n22841 ) | ( ~n22839 & n22841 ) ;
  assign n22843 = ( n694 & n1840 ) | ( n694 & ~n20588 ) | ( n1840 & ~n20588 ) ;
  assign n22844 = n19925 ^ n14752 ^ n13987 ;
  assign n22845 = ( n463 & n2354 ) | ( n463 & n15894 ) | ( n2354 & n15894 ) ;
  assign n22846 = ( n22843 & ~n22844 ) | ( n22843 & n22845 ) | ( ~n22844 & n22845 ) ;
  assign n22848 = ( n3263 & ~n7923 ) | ( n3263 & n9745 ) | ( ~n7923 & n9745 ) ;
  assign n22847 = n2991 & ~n13986 ;
  assign n22849 = n22848 ^ n22847 ^ 1'b0 ;
  assign n22850 = n10580 ^ n5079 ^ n4172 ;
  assign n22851 = ~n22849 & n22850 ;
  assign n22852 = ~n4219 & n22851 ;
  assign n22853 = n21186 ^ n6242 ^ n2085 ;
  assign n22854 = ( n7202 & n11923 ) | ( n7202 & ~n18332 ) | ( n11923 & ~n18332 ) ;
  assign n22855 = ~n22853 & n22854 ;
  assign n22856 = ( ~n6473 & n8303 ) | ( ~n6473 & n12092 ) | ( n8303 & n12092 ) ;
  assign n22857 = n20306 ^ n12548 ^ x37 ;
  assign n22859 = ( n2254 & n11933 ) | ( n2254 & ~n15248 ) | ( n11933 & ~n15248 ) ;
  assign n22858 = n18274 ^ n1976 ^ n1707 ;
  assign n22860 = n22859 ^ n22858 ^ n2457 ;
  assign n22864 = ( n315 & ~n8530 ) | ( n315 & n13228 ) | ( ~n8530 & n13228 ) ;
  assign n22861 = n14033 ^ n8962 ^ n3548 ;
  assign n22862 = n22861 ^ n5096 ^ n2350 ;
  assign n22863 = n22862 ^ n1666 ^ 1'b0 ;
  assign n22865 = n22864 ^ n22863 ^ n13089 ;
  assign n22866 = n17077 ^ n14156 ^ n10104 ;
  assign n22867 = ( n3787 & ~n5528 ) | ( n3787 & n5749 ) | ( ~n5528 & n5749 ) ;
  assign n22868 = ~n17286 & n18774 ;
  assign n22869 = n22868 ^ n21663 ^ n9364 ;
  assign n22870 = ( ~n7858 & n22867 ) | ( ~n7858 & n22869 ) | ( n22867 & n22869 ) ;
  assign n22872 = n15125 ^ n9135 ^ n8607 ;
  assign n22873 = n22872 ^ n631 ^ n302 ;
  assign n22871 = n6982 ^ n5799 ^ n2679 ;
  assign n22874 = n22873 ^ n22871 ^ n5542 ;
  assign n22875 = n20053 ^ n6878 ^ n2851 ;
  assign n22876 = n22875 ^ n9076 ^ n6631 ;
  assign n22877 = n7626 & n10773 ;
  assign n22878 = n18436 ^ n10570 ^ x3 ;
  assign n22879 = n16842 ^ n6905 ^ n6057 ;
  assign n22880 = n11042 ^ n7706 ^ n3120 ;
  assign n22881 = n20240 ^ n9872 ^ n7434 ;
  assign n22882 = ( n9044 & n22880 ) | ( n9044 & ~n22881 ) | ( n22880 & ~n22881 ) ;
  assign n22883 = n9386 ^ n9004 ^ n6726 ;
  assign n22894 = n218 & n12984 ;
  assign n22895 = n22894 ^ n19667 ^ 1'b0 ;
  assign n22884 = n5137 ^ n2806 ^ n189 ;
  assign n22885 = ( n352 & n7715 ) | ( n352 & n22884 ) | ( n7715 & n22884 ) ;
  assign n22886 = n19366 ^ n4656 ^ n1785 ;
  assign n22887 = ~n8707 & n22886 ;
  assign n22888 = n22885 & n22887 ;
  assign n22889 = n10969 & ~n22888 ;
  assign n22890 = n8106 ^ n6992 ^ n3573 ;
  assign n22891 = n22890 ^ n10937 ^ n5234 ;
  assign n22892 = ( ~n7727 & n22889 ) | ( ~n7727 & n22891 ) | ( n22889 & n22891 ) ;
  assign n22893 = ( n1967 & ~n12246 ) | ( n1967 & n22892 ) | ( ~n12246 & n22892 ) ;
  assign n22896 = n22895 ^ n22893 ^ n5463 ;
  assign n22897 = ~n12125 & n21312 ;
  assign n22898 = n1099 & n22897 ;
  assign n22899 = n9551 ^ n4076 ^ n906 ;
  assign n22900 = n15231 | n15426 ;
  assign n22901 = ~n22899 & n22900 ;
  assign n22902 = n9977 ^ n5546 ^ n1148 ;
  assign n22903 = n22902 ^ n17986 ^ n7044 ;
  assign n22904 = ( n5708 & n18787 ) | ( n5708 & ~n22903 ) | ( n18787 & ~n22903 ) ;
  assign n22906 = n10434 ^ n5722 ^ n3471 ;
  assign n22907 = ( ~n7866 & n11308 ) | ( ~n7866 & n22906 ) | ( n11308 & n22906 ) ;
  assign n22905 = ( n13414 & n13909 ) | ( n13414 & ~n22144 ) | ( n13909 & ~n22144 ) ;
  assign n22908 = n22907 ^ n22905 ^ n15834 ;
  assign n22909 = n12680 ^ n10496 ^ n9754 ;
  assign n22910 = ( n15377 & n15747 ) | ( n15377 & n22909 ) | ( n15747 & n22909 ) ;
  assign n22911 = n7020 ^ n6539 ^ n1485 ;
  assign n22912 = n2928 & n6924 ;
  assign n22913 = ( n6344 & n22911 ) | ( n6344 & n22912 ) | ( n22911 & n22912 ) ;
  assign n22914 = ( n5500 & n9619 ) | ( n5500 & ~n13971 ) | ( n9619 & ~n13971 ) ;
  assign n22915 = ( n5757 & n22322 ) | ( n5757 & n22914 ) | ( n22322 & n22914 ) ;
  assign n22916 = n22915 ^ n13064 ^ n9054 ;
  assign n22917 = ~n2997 & n7164 ;
  assign n22918 = n22917 ^ n19737 ^ 1'b0 ;
  assign n22919 = ( n1248 & ~n11343 ) | ( n1248 & n22918 ) | ( ~n11343 & n22918 ) ;
  assign n22920 = ( ~n5223 & n7536 ) | ( ~n5223 & n14680 ) | ( n7536 & n14680 ) ;
  assign n22921 = n17635 | n20315 ;
  assign n22922 = n10521 & ~n22921 ;
  assign n22923 = ( ~n881 & n4853 ) | ( ~n881 & n22922 ) | ( n4853 & n22922 ) ;
  assign n22924 = ( n5903 & ~n9284 ) | ( n5903 & n9683 ) | ( ~n9284 & n9683 ) ;
  assign n22925 = ( n2624 & n8344 ) | ( n2624 & n22924 ) | ( n8344 & n22924 ) ;
  assign n22926 = n22925 ^ n12790 ^ n5985 ;
  assign n22927 = ( n12558 & n19879 ) | ( n12558 & n22893 ) | ( n19879 & n22893 ) ;
  assign n22928 = n13483 ^ n8666 ^ n7801 ;
  assign n22929 = ( ~n9693 & n17484 ) | ( ~n9693 & n22928 ) | ( n17484 & n22928 ) ;
  assign n22930 = n22929 ^ n19354 ^ n5667 ;
  assign n22934 = n10091 ^ n4582 ^ n2062 ;
  assign n22931 = n12199 ^ n6504 ^ n2438 ;
  assign n22932 = n22931 ^ n16091 ^ n15162 ;
  assign n22933 = ( ~n10860 & n13309 ) | ( ~n10860 & n22932 ) | ( n13309 & n22932 ) ;
  assign n22935 = n22934 ^ n22933 ^ n953 ;
  assign n22936 = n12054 ^ n7626 ^ n6602 ;
  assign n22937 = n20825 ^ n4962 ^ n1234 ;
  assign n22938 = n22035 ^ n21062 ^ n9720 ;
  assign n22939 = ( ~n4953 & n7050 ) | ( ~n4953 & n21825 ) | ( n7050 & n21825 ) ;
  assign n22940 = ( n3401 & ~n9534 ) | ( n3401 & n22939 ) | ( ~n9534 & n22939 ) ;
  assign n22941 = n14991 ^ n9020 ^ n1574 ;
  assign n22942 = ( n14668 & n14837 ) | ( n14668 & ~n22941 ) | ( n14837 & ~n22941 ) ;
  assign n22943 = n323 | n6045 ;
  assign n22944 = n3968 & ~n22943 ;
  assign n22945 = ( ~n5034 & n7383 ) | ( ~n5034 & n22944 ) | ( n7383 & n22944 ) ;
  assign n22946 = n22945 ^ n12396 ^ 1'b0 ;
  assign n22947 = ~n3666 & n12402 ;
  assign n22948 = n22947 ^ n14767 ^ 1'b0 ;
  assign n22949 = ( n2371 & ~n10513 ) | ( n2371 & n19231 ) | ( ~n10513 & n19231 ) ;
  assign n22950 = ( n1917 & ~n7723 ) | ( n1917 & n10797 ) | ( ~n7723 & n10797 ) ;
  assign n22952 = ( n4588 & n7813 ) | ( n4588 & ~n10002 ) | ( n7813 & ~n10002 ) ;
  assign n22951 = ( n3446 & n13526 ) | ( n3446 & n21526 ) | ( n13526 & n21526 ) ;
  assign n22953 = n22952 ^ n22951 ^ 1'b0 ;
  assign n22954 = ( ~n4556 & n5135 ) | ( ~n4556 & n11576 ) | ( n5135 & n11576 ) ;
  assign n22955 = ( n8177 & ~n9852 ) | ( n8177 & n16573 ) | ( ~n9852 & n16573 ) ;
  assign n22956 = n22955 ^ n10519 ^ n5603 ;
  assign n22957 = n1757 & n2336 ;
  assign n22958 = n8096 | n22957 ;
  assign n22959 = n8078 | n22958 ;
  assign n22960 = ( n1797 & n21862 ) | ( n1797 & n22959 ) | ( n21862 & n22959 ) ;
  assign n22961 = ( n22954 & n22956 ) | ( n22954 & ~n22960 ) | ( n22956 & ~n22960 ) ;
  assign n22962 = n18151 ^ n3548 ^ n1246 ;
  assign n22963 = ( n816 & n17207 ) | ( n816 & ~n22962 ) | ( n17207 & ~n22962 ) ;
  assign n22964 = n7709 & n22963 ;
  assign n22965 = n22964 ^ n18210 ^ 1'b0 ;
  assign n22966 = ( ~n5172 & n6257 ) | ( ~n5172 & n22965 ) | ( n6257 & n22965 ) ;
  assign n22967 = n21095 ^ n6951 ^ 1'b0 ;
  assign n22968 = n9036 & ~n22967 ;
  assign n22969 = n22968 ^ n19851 ^ n3008 ;
  assign n22970 = n17489 ^ n8584 ^ n4576 ;
  assign n22971 = n4506 & ~n22583 ;
  assign n22972 = n22971 ^ n2040 ^ 1'b0 ;
  assign n22973 = n7954 | n22453 ;
  assign n22974 = n12047 | n22973 ;
  assign n22975 = ( n11237 & n15701 ) | ( n11237 & n17940 ) | ( n15701 & n17940 ) ;
  assign n22976 = n18565 ^ n14828 ^ n390 ;
  assign n22977 = ( n3791 & ~n9965 ) | ( n3791 & n22190 ) | ( ~n9965 & n22190 ) ;
  assign n22978 = ( ~n16467 & n18572 ) | ( ~n16467 & n22915 ) | ( n18572 & n22915 ) ;
  assign n22979 = n463 & ~n13563 ;
  assign n22980 = n22979 ^ n10463 ^ 1'b0 ;
  assign n22981 = n14688 ^ n5467 ^ n3813 ;
  assign n22982 = n10755 ^ x73 ^ 1'b0 ;
  assign n22983 = n22982 ^ n20989 ^ n12802 ;
  assign n22984 = ( ~n14013 & n22981 ) | ( ~n14013 & n22983 ) | ( n22981 & n22983 ) ;
  assign n22985 = ( n9785 & n11347 ) | ( n9785 & ~n13482 ) | ( n11347 & ~n13482 ) ;
  assign n22986 = ( n4176 & ~n10778 ) | ( n4176 & n19546 ) | ( ~n10778 & n19546 ) ;
  assign n22987 = ( n11215 & n14716 ) | ( n11215 & n18248 ) | ( n14716 & n18248 ) ;
  assign n22988 = ( n17607 & n19708 ) | ( n17607 & n22987 ) | ( n19708 & n22987 ) ;
  assign n22989 = n22988 ^ n19321 ^ n18835 ;
  assign n22990 = ( n3715 & ~n9558 ) | ( n3715 & n10539 ) | ( ~n9558 & n10539 ) ;
  assign n22991 = n2150 & n12030 ;
  assign n22992 = n22991 ^ n1387 ^ 1'b0 ;
  assign n22996 = n15518 ^ n5350 ^ 1'b0 ;
  assign n22997 = n14029 & ~n22996 ;
  assign n22998 = n22997 ^ n1506 ^ 1'b0 ;
  assign n22999 = n22998 ^ n22611 ^ n1920 ;
  assign n22994 = ( n1978 & ~n8308 ) | ( n1978 & n11763 ) | ( ~n8308 & n11763 ) ;
  assign n22995 = ( n3669 & ~n6093 ) | ( n3669 & n22994 ) | ( ~n6093 & n22994 ) ;
  assign n22993 = ( n9105 & ~n12168 ) | ( n9105 & n18679 ) | ( ~n12168 & n18679 ) ;
  assign n23000 = n22999 ^ n22995 ^ n22993 ;
  assign n23001 = n9068 ^ n1294 ^ 1'b0 ;
  assign n23002 = n15297 ^ n9833 ^ n6675 ;
  assign n23004 = ( ~n2044 & n3051 ) | ( ~n2044 & n10659 ) | ( n3051 & n10659 ) ;
  assign n23003 = ( n7165 & ~n17454 ) | ( n7165 & n19253 ) | ( ~n17454 & n19253 ) ;
  assign n23005 = n23004 ^ n23003 ^ 1'b0 ;
  assign n23006 = ( ~n1883 & n23002 ) | ( ~n1883 & n23005 ) | ( n23002 & n23005 ) ;
  assign n23008 = ~n588 & n13928 ;
  assign n23007 = n16887 ^ n5223 ^ n3564 ;
  assign n23009 = n23008 ^ n23007 ^ n20383 ;
  assign n23012 = ( ~n1391 & n1452 ) | ( ~n1391 & n9857 ) | ( n1452 & n9857 ) ;
  assign n23010 = n3274 ^ n3122 ^ 1'b0 ;
  assign n23011 = ( ~n4066 & n7631 ) | ( ~n4066 & n23010 ) | ( n7631 & n23010 ) ;
  assign n23013 = n23012 ^ n23011 ^ 1'b0 ;
  assign n23014 = n893 | n23013 ;
  assign n23015 = n22366 ^ n12382 ^ 1'b0 ;
  assign n23016 = ~n13334 & n23015 ;
  assign n23017 = ( ~n825 & n2558 ) | ( ~n825 & n16811 ) | ( n2558 & n16811 ) ;
  assign n23018 = n16001 ^ n4863 ^ n3231 ;
  assign n23019 = n12528 ^ n11372 ^ n2179 ;
  assign n23020 = n12226 ^ n8591 ^ n4087 ;
  assign n23021 = ( n2183 & n12315 ) | ( n2183 & ~n23020 ) | ( n12315 & ~n23020 ) ;
  assign n23025 = ( x52 & ~n2843 ) | ( x52 & n12497 ) | ( ~n2843 & n12497 ) ;
  assign n23022 = n3437 ^ n370 ^ 1'b0 ;
  assign n23023 = n23022 ^ n7406 ^ n191 ;
  assign n23024 = n23023 ^ n16373 ^ n4067 ;
  assign n23026 = n23025 ^ n23024 ^ n13695 ;
  assign n23027 = n23026 ^ n16844 ^ n2196 ;
  assign n23028 = n20033 ^ n12115 ^ n6715 ;
  assign n23029 = n23028 ^ n15360 ^ n5403 ;
  assign n23030 = n23029 ^ n10374 ^ 1'b0 ;
  assign n23031 = ~n22179 & n23030 ;
  assign n23032 = ~n3502 & n9622 ;
  assign n23033 = n20713 ^ n13581 ^ n2065 ;
  assign n23034 = ( ~n782 & n2019 ) | ( ~n782 & n23033 ) | ( n2019 & n23033 ) ;
  assign n23035 = n1970 | n23034 ;
  assign n23036 = n19993 | n23035 ;
  assign n23037 = n12702 ^ n3257 ^ 1'b0 ;
  assign n23038 = ( n2787 & n7697 ) | ( n2787 & ~n23037 ) | ( n7697 & ~n23037 ) ;
  assign n23039 = ( n13060 & n16863 ) | ( n13060 & ~n23038 ) | ( n16863 & ~n23038 ) ;
  assign n23040 = n7411 & n23039 ;
  assign n23041 = ~n23036 & n23040 ;
  assign n23042 = ( n405 & n22410 ) | ( n405 & n23041 ) | ( n22410 & n23041 ) ;
  assign n23043 = n15666 ^ n9825 ^ n2843 ;
  assign n23044 = n23043 ^ n22764 ^ n7774 ;
  assign n23047 = ( n360 & ~n421 ) | ( n360 & n5827 ) | ( ~n421 & n5827 ) ;
  assign n23045 = ( n1395 & n3318 ) | ( n1395 & ~n7744 ) | ( n3318 & ~n7744 ) ;
  assign n23046 = ( n4336 & n16796 ) | ( n4336 & n23045 ) | ( n16796 & n23045 ) ;
  assign n23048 = n23047 ^ n23046 ^ n18478 ;
  assign n23049 = n23048 ^ n19386 ^ n6021 ;
  assign n23050 = ( n4512 & n10053 ) | ( n4512 & n20268 ) | ( n10053 & n20268 ) ;
  assign n23051 = n22495 ^ n9217 ^ 1'b0 ;
  assign n23052 = n17224 ^ n8106 ^ n1705 ;
  assign n23053 = n10738 ^ n8024 ^ 1'b0 ;
  assign n23056 = n12600 ^ n3084 ^ n2028 ;
  assign n23057 = ( ~n4687 & n19683 ) | ( ~n4687 & n23056 ) | ( n19683 & n23056 ) ;
  assign n23054 = n1151 & ~n18497 ;
  assign n23055 = n6642 & n23054 ;
  assign n23058 = n23057 ^ n23055 ^ n10746 ;
  assign n23059 = ( n4360 & ~n4392 ) | ( n4360 & n7055 ) | ( ~n4392 & n7055 ) ;
  assign n23060 = n23059 ^ n10750 ^ n6200 ;
  assign n23061 = ( n5098 & ~n12926 ) | ( n5098 & n23060 ) | ( ~n12926 & n23060 ) ;
  assign n23062 = ~n11936 & n15612 ;
  assign n23064 = n7278 ^ n2471 ^ n1784 ;
  assign n23065 = n23064 ^ n15979 ^ n2595 ;
  assign n23066 = ~n10143 & n23065 ;
  assign n23063 = ( ~n3635 & n11519 ) | ( ~n3635 & n22889 ) | ( n11519 & n22889 ) ;
  assign n23067 = n23066 ^ n23063 ^ n326 ;
  assign n23068 = n1417 | n20441 ;
  assign n23069 = n6094 ^ n1235 ^ 1'b0 ;
  assign n23070 = ~n16021 & n23069 ;
  assign n23071 = n23070 ^ n2963 ^ n595 ;
  assign n23072 = n3494 & ~n23071 ;
  assign n23073 = n23072 ^ n11761 ^ 1'b0 ;
  assign n23074 = ~n8303 & n9873 ;
  assign n23075 = n23074 ^ n4612 ^ 1'b0 ;
  assign n23076 = n23075 ^ n17576 ^ n14162 ;
  assign n23077 = n23076 ^ n22806 ^ n4846 ;
  assign n23078 = n23077 ^ n22853 ^ n164 ;
  assign n23079 = n23078 ^ n14828 ^ 1'b0 ;
  assign n23080 = n11441 & n23079 ;
  assign n23081 = n15610 ^ n12104 ^ n2969 ;
  assign n23082 = n6095 ^ n2187 ^ 1'b0 ;
  assign n23083 = n1752 & n23082 ;
  assign n23084 = n23083 ^ n17198 ^ n2782 ;
  assign n23085 = ( n18676 & n23081 ) | ( n18676 & n23084 ) | ( n23081 & n23084 ) ;
  assign n23086 = n23085 ^ n16745 ^ n15872 ;
  assign n23087 = n4322 ^ n3257 ^ n1257 ;
  assign n23088 = n23087 ^ n6095 ^ n5230 ;
  assign n23091 = n15733 ^ n14949 ^ n11083 ;
  assign n23089 = n7762 & n14469 ;
  assign n23090 = n23089 ^ n10016 ^ 1'b0 ;
  assign n23092 = n23091 ^ n23090 ^ n2107 ;
  assign n23093 = ( n1306 & ~n6357 ) | ( n1306 & n16148 ) | ( ~n6357 & n16148 ) ;
  assign n23095 = n18933 ^ n6193 ^ n3719 ;
  assign n23094 = n17698 & n18613 ;
  assign n23096 = n23095 ^ n23094 ^ n2784 ;
  assign n23097 = n10683 ^ n3107 ^ 1'b0 ;
  assign n23098 = ( n6230 & n18535 ) | ( n6230 & ~n23097 ) | ( n18535 & ~n23097 ) ;
  assign n23099 = ( n1529 & n7965 ) | ( n1529 & n10144 ) | ( n7965 & n10144 ) ;
  assign n23100 = n15248 ^ n10800 ^ n673 ;
  assign n23101 = n23100 ^ n14108 ^ n6449 ;
  assign n23102 = n23101 ^ n11249 ^ n2966 ;
  assign n23103 = n18667 ^ n13163 ^ n3556 ;
  assign n23105 = n3459 ^ n3049 ^ n2847 ;
  assign n23104 = n3827 & n16656 ;
  assign n23106 = n23105 ^ n23104 ^ 1'b0 ;
  assign n23107 = ( n6798 & ~n12356 ) | ( n6798 & n23106 ) | ( ~n12356 & n23106 ) ;
  assign n23113 = n22982 ^ n6072 ^ 1'b0 ;
  assign n23114 = n20706 | n23113 ;
  assign n23109 = n17794 ^ n3481 ^ 1'b0 ;
  assign n23110 = n1479 & ~n23109 ;
  assign n23111 = ( ~n1680 & n12013 ) | ( ~n1680 & n23110 ) | ( n12013 & n23110 ) ;
  assign n23108 = n12502 ^ n7945 ^ n2600 ;
  assign n23112 = n23111 ^ n23108 ^ n19817 ;
  assign n23115 = n23114 ^ n23112 ^ n8816 ;
  assign n23116 = ( ~x76 & n11618 ) | ( ~x76 & n16871 ) | ( n11618 & n16871 ) ;
  assign n23119 = ( n5774 & ~n8666 ) | ( n5774 & n12701 ) | ( ~n8666 & n12701 ) ;
  assign n23120 = n4770 ^ n767 ^ 1'b0 ;
  assign n23121 = n23119 & ~n23120 ;
  assign n23117 = n5564 | n11067 ;
  assign n23118 = n23117 ^ n18507 ^ 1'b0 ;
  assign n23122 = n23121 ^ n23118 ^ n7126 ;
  assign n23123 = n7605 | n19936 ;
  assign n23124 = n4160 | n23123 ;
  assign n23125 = ( n669 & n6891 ) | ( n669 & n15225 ) | ( n6891 & n15225 ) ;
  assign n23126 = ( n6703 & n12841 ) | ( n6703 & ~n17745 ) | ( n12841 & ~n17745 ) ;
  assign n23127 = ( n5840 & n7887 ) | ( n5840 & ~n11800 ) | ( n7887 & ~n11800 ) ;
  assign n23128 = ( ~n5059 & n9297 ) | ( ~n5059 & n16124 ) | ( n9297 & n16124 ) ;
  assign n23129 = ( n4533 & n7557 ) | ( n4533 & n23128 ) | ( n7557 & n23128 ) ;
  assign n23130 = n23129 ^ n15574 ^ n5519 ;
  assign n23131 = ( n3496 & n16552 ) | ( n3496 & n20383 ) | ( n16552 & n20383 ) ;
  assign n23132 = ( n14395 & n23130 ) | ( n14395 & n23131 ) | ( n23130 & n23131 ) ;
  assign n23133 = n17564 ^ n5604 ^ n3956 ;
  assign n23134 = n8499 ^ n3055 ^ n1248 ;
  assign n23135 = n23134 ^ n15549 ^ n6795 ;
  assign n23136 = n22594 ^ n13377 ^ n7612 ;
  assign n23137 = ~n3813 & n4839 ;
  assign n23138 = n23137 ^ n14063 ^ 1'b0 ;
  assign n23139 = ( n4904 & n15442 ) | ( n4904 & ~n18576 ) | ( n15442 & ~n18576 ) ;
  assign n23140 = ( n2356 & n4876 ) | ( n2356 & ~n13828 ) | ( n4876 & ~n13828 ) ;
  assign n23143 = ( n4934 & n6998 ) | ( n4934 & n11984 ) | ( n6998 & n11984 ) ;
  assign n23144 = n23143 ^ n15248 ^ n12367 ;
  assign n23145 = n23144 ^ n13060 ^ n4464 ;
  assign n23141 = ( n3362 & n3514 ) | ( n3362 & ~n19241 ) | ( n3514 & ~n19241 ) ;
  assign n23142 = n23141 ^ n13617 ^ n562 ;
  assign n23146 = n23145 ^ n23142 ^ n20587 ;
  assign n23147 = ~n7738 & n22093 ;
  assign n23148 = n23147 ^ n5846 ^ n4920 ;
  assign n23149 = n12110 ^ n5825 ^ n2023 ;
  assign n23150 = n4802 & ~n23149 ;
  assign n23151 = n23150 ^ n6606 ^ 1'b0 ;
  assign n23152 = ( n4346 & n10053 ) | ( n4346 & ~n23105 ) | ( n10053 & ~n23105 ) ;
  assign n23153 = n23152 ^ n4016 ^ 1'b0 ;
  assign n23154 = n7958 & ~n23153 ;
  assign n23155 = ~n3305 & n23154 ;
  assign n23156 = n14462 ^ n7780 ^ n6258 ;
  assign n23157 = ( n964 & ~n12400 ) | ( n964 & n19301 ) | ( ~n12400 & n19301 ) ;
  assign n23158 = n1562 & n8493 ;
  assign n23159 = ( n11936 & n16111 ) | ( n11936 & ~n23158 ) | ( n16111 & ~n23158 ) ;
  assign n23160 = n7540 ^ n1705 ^ 1'b0 ;
  assign n23161 = n23160 ^ n19398 ^ n4090 ;
  assign n23162 = ( n1671 & n7335 ) | ( n1671 & n23161 ) | ( n7335 & n23161 ) ;
  assign n23163 = ( n15862 & ~n18420 ) | ( n15862 & n19929 ) | ( ~n18420 & n19929 ) ;
  assign n23164 = n13891 ^ n8147 ^ 1'b0 ;
  assign n23165 = n15757 | n23164 ;
  assign n23166 = n5699 & ~n23165 ;
  assign n23167 = n23166 ^ n12000 ^ 1'b0 ;
  assign n23168 = ( n16906 & ~n22362 ) | ( n16906 & n22963 ) | ( ~n22362 & n22963 ) ;
  assign n23169 = ( n3401 & n5284 ) | ( n3401 & n10413 ) | ( n5284 & n10413 ) ;
  assign n23170 = n23169 ^ n19133 ^ n5535 ;
  assign n23171 = ( n1752 & ~n8159 ) | ( n1752 & n22169 ) | ( ~n8159 & n22169 ) ;
  assign n23172 = n23171 ^ n15987 ^ 1'b0 ;
  assign n23173 = n23172 ^ n23121 ^ n14656 ;
  assign n23174 = n3930 & ~n4852 ;
  assign n23175 = n23174 ^ n1201 ^ 1'b0 ;
  assign n23176 = ( ~n5061 & n12281 ) | ( ~n5061 & n13578 ) | ( n12281 & n13578 ) ;
  assign n23177 = ( n2216 & n23175 ) | ( n2216 & n23176 ) | ( n23175 & n23176 ) ;
  assign n23178 = n20520 ^ n2900 ^ n2756 ;
  assign n23179 = n6651 ^ n6165 ^ n4334 ;
  assign n23180 = ( n2558 & ~n5884 ) | ( n2558 & n7968 ) | ( ~n5884 & n7968 ) ;
  assign n23181 = n19159 ^ n15026 ^ n9301 ;
  assign n23182 = ( n289 & n473 ) | ( n289 & n11493 ) | ( n473 & n11493 ) ;
  assign n23183 = ( n5323 & n9185 ) | ( n5323 & ~n23182 ) | ( n9185 & ~n23182 ) ;
  assign n23184 = n20405 ^ n218 ^ 1'b0 ;
  assign n23185 = n23184 ^ n16426 ^ n1335 ;
  assign n23186 = n23185 ^ n13891 ^ 1'b0 ;
  assign n23187 = n17011 ^ n5454 ^ n1830 ;
  assign n23188 = n23187 ^ n14764 ^ 1'b0 ;
  assign n23189 = n1923 | n23188 ;
  assign n23190 = n23189 ^ n3400 ^ n2970 ;
  assign n23191 = n23190 ^ n18199 ^ n9905 ;
  assign n23193 = n14644 ^ n4658 ^ n3433 ;
  assign n23192 = n9404 ^ n8275 ^ n427 ;
  assign n23194 = n23193 ^ n23192 ^ n651 ;
  assign n23195 = ( ~n288 & n3192 ) | ( ~n288 & n3342 ) | ( n3192 & n3342 ) ;
  assign n23196 = n23195 ^ n11842 ^ n1459 ;
  assign n23197 = ( n7001 & ~n10923 ) | ( n7001 & n13149 ) | ( ~n10923 & n13149 ) ;
  assign n23198 = n1826 & ~n3414 ;
  assign n23199 = ~n23197 & n23198 ;
  assign n23200 = n7667 ^ n7278 ^ 1'b0 ;
  assign n23201 = n22035 ^ n18224 ^ 1'b0 ;
  assign n23202 = n14632 | n23201 ;
  assign n23203 = n23202 ^ n21197 ^ 1'b0 ;
  assign n23204 = n23200 & n23203 ;
  assign n23205 = n17463 & n23204 ;
  assign n23206 = n23205 ^ n328 ^ 1'b0 ;
  assign n23207 = n8887 & ~n10922 ;
  assign n23208 = ( n3912 & n18243 ) | ( n3912 & ~n23207 ) | ( n18243 & ~n23207 ) ;
  assign n23209 = n11639 ^ n11474 ^ n811 ;
  assign n23210 = ( n1354 & ~n5899 ) | ( n1354 & n23209 ) | ( ~n5899 & n23209 ) ;
  assign n23211 = ( n6669 & n21699 ) | ( n6669 & n23210 ) | ( n21699 & n23210 ) ;
  assign n23212 = n11433 ^ n9312 ^ n1995 ;
  assign n23213 = n19533 ^ n6109 ^ 1'b0 ;
  assign n23214 = n23213 ^ n17229 ^ n3590 ;
  assign n23215 = ( ~n988 & n23212 ) | ( ~n988 & n23214 ) | ( n23212 & n23214 ) ;
  assign n23216 = ( n1842 & ~n10053 ) | ( n1842 & n10556 ) | ( ~n10053 & n10556 ) ;
  assign n23217 = ( n2274 & ~n3340 ) | ( n2274 & n15276 ) | ( ~n3340 & n15276 ) ;
  assign n23218 = ( n2314 & ~n15317 ) | ( n2314 & n23217 ) | ( ~n15317 & n23217 ) ;
  assign n23219 = ( ~n7556 & n18802 ) | ( ~n7556 & n23218 ) | ( n18802 & n23218 ) ;
  assign n23220 = n3535 & n20938 ;
  assign n23221 = n23220 ^ n2157 ^ 1'b0 ;
  assign n23222 = n22428 ^ n21218 ^ n12231 ;
  assign n23223 = n21973 ^ n5379 ^ x22 ;
  assign n23224 = ( ~n14968 & n23222 ) | ( ~n14968 & n23223 ) | ( n23222 & n23223 ) ;
  assign n23225 = ( ~n424 & n3180 ) | ( ~n424 & n17151 ) | ( n3180 & n17151 ) ;
  assign n23226 = ( n1285 & ~n9054 ) | ( n1285 & n16818 ) | ( ~n9054 & n16818 ) ;
  assign n23227 = n8041 ^ n2781 ^ n1817 ;
  assign n23228 = n18825 ^ n5153 ^ n3488 ;
  assign n23229 = ( n1718 & n19354 ) | ( n1718 & n23228 ) | ( n19354 & n23228 ) ;
  assign n23230 = n23229 ^ n17344 ^ n3367 ;
  assign n23231 = ( ~n23226 & n23227 ) | ( ~n23226 & n23230 ) | ( n23227 & n23230 ) ;
  assign n23232 = ( ~n994 & n4049 ) | ( ~n994 & n8223 ) | ( n4049 & n8223 ) ;
  assign n23233 = ( n16038 & n18460 ) | ( n16038 & ~n22594 ) | ( n18460 & ~n22594 ) ;
  assign n23234 = n23233 ^ n17607 ^ n12486 ;
  assign n23235 = n14601 ^ n1710 ^ 1'b0 ;
  assign n23236 = ~n7192 & n23235 ;
  assign n23237 = n6327 ^ n5378 ^ 1'b0 ;
  assign n23238 = n17448 ^ n15866 ^ 1'b0 ;
  assign n23239 = n12586 ^ n9378 ^ n7405 ;
  assign n23240 = n12851 ^ n8730 ^ n950 ;
  assign n23241 = n17500 & n23240 ;
  assign n23242 = ( n12552 & ~n19735 ) | ( n12552 & n23241 ) | ( ~n19735 & n23241 ) ;
  assign n23243 = n12942 ^ n11445 ^ n3874 ;
  assign n23244 = ( n465 & n1191 ) | ( n465 & n10812 ) | ( n1191 & n10812 ) ;
  assign n23245 = n17421 ^ n9512 ^ n3444 ;
  assign n23246 = ( n4836 & n17191 ) | ( n4836 & ~n23245 ) | ( n17191 & ~n23245 ) ;
  assign n23248 = n10746 ^ n9769 ^ n1239 ;
  assign n23249 = ( n4570 & ~n16098 ) | ( n4570 & n23248 ) | ( ~n16098 & n23248 ) ;
  assign n23247 = ( ~n3740 & n22197 ) | ( ~n3740 & n22568 ) | ( n22197 & n22568 ) ;
  assign n23250 = n23249 ^ n23247 ^ n6173 ;
  assign n23251 = n5037 | n7691 ;
  assign n23252 = n23251 ^ n6587 ^ 1'b0 ;
  assign n23253 = n19508 ^ n6170 ^ 1'b0 ;
  assign n23254 = n17303 & n23253 ;
  assign n23257 = n18194 ^ n15799 ^ n5357 ;
  assign n23255 = n5600 | n11672 ;
  assign n23256 = ( ~n649 & n21727 ) | ( ~n649 & n23255 ) | ( n21727 & n23255 ) ;
  assign n23258 = n23257 ^ n23256 ^ n8370 ;
  assign n23264 = n19178 ^ n8585 ^ n7636 ;
  assign n23259 = n3133 ^ n2373 ^ n588 ;
  assign n23260 = n4246 | n23259 ;
  assign n23261 = n20213 ^ n14041 ^ n581 ;
  assign n23262 = ( ~n6054 & n16073 ) | ( ~n6054 & n23261 ) | ( n16073 & n23261 ) ;
  assign n23263 = ( n10449 & n23260 ) | ( n10449 & ~n23262 ) | ( n23260 & ~n23262 ) ;
  assign n23265 = n23264 ^ n23263 ^ n21284 ;
  assign n23266 = n17047 ^ n6310 ^ n3983 ;
  assign n23267 = n19096 ^ n17627 ^ 1'b0 ;
  assign n23270 = ( n582 & n17216 ) | ( n582 & ~n20365 ) | ( n17216 & ~n20365 ) ;
  assign n23268 = n16263 & ~n19753 ;
  assign n23269 = n23268 ^ n10243 ^ n6208 ;
  assign n23271 = n23270 ^ n23269 ^ n8350 ;
  assign n23272 = ( n1839 & n14457 ) | ( n1839 & n18577 ) | ( n14457 & n18577 ) ;
  assign n23273 = n17501 ^ n6733 ^ 1'b0 ;
  assign n23274 = ~n13493 & n23273 ;
  assign n23275 = ( n11961 & ~n13121 ) | ( n11961 & n23274 ) | ( ~n13121 & n23274 ) ;
  assign n23276 = ( n2875 & n7969 ) | ( n2875 & ~n23275 ) | ( n7969 & ~n23275 ) ;
  assign n23277 = n13665 ^ n10745 ^ n3704 ;
  assign n23278 = n22016 | n23277 ;
  assign n23279 = n23278 ^ n12048 ^ n10702 ;
  assign n23282 = n9465 ^ n6323 ^ n614 ;
  assign n23283 = n23282 ^ n14700 ^ n1545 ;
  assign n23280 = n7370 & ~n13042 ;
  assign n23281 = ~n1448 & n23280 ;
  assign n23284 = n23283 ^ n23281 ^ n1173 ;
  assign n23285 = ~n2736 & n2944 ;
  assign n23292 = n7015 & ~n22058 ;
  assign n23290 = n17684 ^ n13009 ^ n11737 ;
  assign n23291 = ( n20322 & n22816 ) | ( n20322 & n23290 ) | ( n22816 & n23290 ) ;
  assign n23293 = n23292 ^ n23291 ^ 1'b0 ;
  assign n23294 = n9465 | n23293 ;
  assign n23287 = n17461 ^ n5194 ^ 1'b0 ;
  assign n23288 = n23287 ^ n16842 ^ 1'b0 ;
  assign n23286 = ( ~n1365 & n9558 ) | ( ~n1365 & n9764 ) | ( n9558 & n9764 ) ;
  assign n23289 = n23288 ^ n23286 ^ n22527 ;
  assign n23295 = n23294 ^ n23289 ^ n13045 ;
  assign n23296 = n9435 ^ n6705 ^ 1'b0 ;
  assign n23297 = ( n4116 & n20235 ) | ( n4116 & n23296 ) | ( n20235 & n23296 ) ;
  assign n23300 = n22373 ^ n2718 ^ n959 ;
  assign n23301 = n12525 & n23300 ;
  assign n23302 = n23301 ^ n11062 ^ n8177 ;
  assign n23298 = ( n730 & ~n2709 ) | ( n730 & n9569 ) | ( ~n2709 & n9569 ) ;
  assign n23299 = ( n6941 & n10133 ) | ( n6941 & n23298 ) | ( n10133 & n23298 ) ;
  assign n23303 = n23302 ^ n23299 ^ n13792 ;
  assign n23304 = n6802 ^ n3613 ^ 1'b0 ;
  assign n23305 = n3287 & n23304 ;
  assign n23306 = n23305 ^ n9166 ^ 1'b0 ;
  assign n23307 = n23306 ^ n9904 ^ n4466 ;
  assign n23308 = n11156 ^ n10186 ^ n8623 ;
  assign n23309 = n23308 ^ n8648 ^ n3351 ;
  assign n23310 = n20244 ^ n6739 ^ n2682 ;
  assign n23311 = n23310 ^ n2273 ^ 1'b0 ;
  assign n23312 = ~n21613 & n23311 ;
  assign n23313 = n23312 ^ n18723 ^ 1'b0 ;
  assign n23314 = n10734 & ~n10795 ;
  assign n23315 = n22839 ^ n14860 ^ n9585 ;
  assign n23316 = n10307 ^ n9256 ^ 1'b0 ;
  assign n23317 = n23316 ^ n21396 ^ n20724 ;
  assign n23318 = n11514 ^ n3975 ^ n2757 ;
  assign n23319 = n23318 ^ n17022 ^ n1844 ;
  assign n23320 = n20603 ^ n5039 ^ n4622 ;
  assign n23321 = ( n2153 & n2820 ) | ( n2153 & ~n7947 ) | ( n2820 & ~n7947 ) ;
  assign n23322 = ( n743 & n7564 ) | ( n743 & ~n11916 ) | ( n7564 & ~n11916 ) ;
  assign n23323 = ( n4032 & ~n17480 ) | ( n4032 & n23322 ) | ( ~n17480 & n23322 ) ;
  assign n23324 = n20699 ^ n11096 ^ n3115 ;
  assign n23325 = n23324 ^ n12089 ^ n5083 ;
  assign n23327 = n3999 ^ n1139 ^ n328 ;
  assign n23326 = n18171 ^ n5454 ^ n4907 ;
  assign n23328 = n23327 ^ n23326 ^ n4488 ;
  assign n23329 = ( n7958 & ~n22343 ) | ( n7958 & n23328 ) | ( ~n22343 & n23328 ) ;
  assign n23330 = n14395 ^ n13511 ^ 1'b0 ;
  assign n23331 = n5800 ^ n5189 ^ 1'b0 ;
  assign n23332 = n23331 ^ n9682 ^ n8323 ;
  assign n23333 = ( n2305 & n23330 ) | ( n2305 & ~n23332 ) | ( n23330 & ~n23332 ) ;
  assign n23335 = n21830 ^ n9639 ^ n5946 ;
  assign n23334 = n15650 ^ n7642 ^ n791 ;
  assign n23336 = n23335 ^ n23334 ^ n7149 ;
  assign n23337 = n23336 ^ n20663 ^ n18828 ;
  assign n23338 = n7493 ^ n5691 ^ n910 ;
  assign n23339 = ( n5331 & n23059 ) | ( n5331 & ~n23338 ) | ( n23059 & ~n23338 ) ;
  assign n23341 = n3275 | n4762 ;
  assign n23342 = n624 | n23341 ;
  assign n23340 = n1712 ^ n333 ^ n301 ;
  assign n23343 = n23342 ^ n23340 ^ n10585 ;
  assign n23344 = ( ~n2475 & n10752 ) | ( ~n2475 & n23343 ) | ( n10752 & n23343 ) ;
  assign n23345 = ( n4692 & n23339 ) | ( n4692 & ~n23344 ) | ( n23339 & ~n23344 ) ;
  assign n23346 = n21424 ^ n14484 ^ n5129 ;
  assign n23347 = n23346 ^ n15215 ^ n12766 ;
  assign n23349 = ( n2382 & n14486 ) | ( n2382 & n22140 ) | ( n14486 & n22140 ) ;
  assign n23348 = n21630 ^ n3668 ^ n1205 ;
  assign n23350 = n23349 ^ n23348 ^ n18870 ;
  assign n23351 = n11430 & ~n22831 ;
  assign n23352 = n23351 ^ n18496 ^ 1'b0 ;
  assign n23353 = ( n8521 & n13207 ) | ( n8521 & ~n23352 ) | ( n13207 & ~n23352 ) ;
  assign n23354 = n23353 ^ n22538 ^ n2776 ;
  assign n23355 = ( ~n11950 & n14665 ) | ( ~n11950 & n21825 ) | ( n14665 & n21825 ) ;
  assign n23358 = n17041 & n19201 ;
  assign n23359 = n23358 ^ n8910 ^ n6096 ;
  assign n23356 = ( n532 & n2124 ) | ( n532 & ~n13135 ) | ( n2124 & ~n13135 ) ;
  assign n23357 = n23356 ^ n18005 ^ n13653 ;
  assign n23360 = n23359 ^ n23357 ^ n16974 ;
  assign n23362 = n6347 | n6708 ;
  assign n23361 = ~n9153 & n18804 ;
  assign n23363 = n23362 ^ n23361 ^ 1'b0 ;
  assign n23364 = n21570 ^ n12837 ^ 1'b0 ;
  assign n23365 = ~n21237 & n23364 ;
  assign n23366 = ( n513 & ~n3679 ) | ( n513 & n4399 ) | ( ~n3679 & n4399 ) ;
  assign n23367 = n23366 ^ n10712 ^ n1475 ;
  assign n23368 = ( n3594 & n6064 ) | ( n3594 & ~n6582 ) | ( n6064 & ~n6582 ) ;
  assign n23369 = ( n12001 & ~n23367 ) | ( n12001 & n23368 ) | ( ~n23367 & n23368 ) ;
  assign n23370 = n23369 ^ n6903 ^ 1'b0 ;
  assign n23371 = n5924 & ~n7300 ;
  assign n23372 = n8287 ^ n4706 ^ n3134 ;
  assign n23373 = n23372 ^ n15193 ^ n10544 ;
  assign n23374 = n23373 ^ n7904 ^ 1'b0 ;
  assign n23375 = n2651 | n5368 ;
  assign n23376 = n23375 ^ n3658 ^ 1'b0 ;
  assign n23377 = n23376 ^ n21092 ^ n8550 ;
  assign n23378 = n15689 ^ n10342 ^ n1299 ;
  assign n23379 = n23378 ^ n15714 ^ n12359 ;
  assign n23380 = n250 & n2976 ;
  assign n23381 = n23380 ^ n4525 ^ 1'b0 ;
  assign n23382 = ( n166 & n1373 ) | ( n166 & ~n3402 ) | ( n1373 & ~n3402 ) ;
  assign n23383 = n23382 ^ n19123 ^ n4230 ;
  assign n23384 = n8787 ^ n8371 ^ n2544 ;
  assign n23385 = ( ~n6621 & n8907 ) | ( ~n6621 & n23384 ) | ( n8907 & n23384 ) ;
  assign n23386 = ( ~n2233 & n2665 ) | ( ~n2233 & n16192 ) | ( n2665 & n16192 ) ;
  assign n23387 = n23386 ^ n6512 ^ n1036 ;
  assign n23388 = ( x25 & ~n8090 ) | ( x25 & n20157 ) | ( ~n8090 & n20157 ) ;
  assign n23389 = ~n5522 & n6672 ;
  assign n23390 = n23389 ^ n9074 ^ 1'b0 ;
  assign n23391 = n23390 ^ n16384 ^ n3055 ;
  assign n23392 = n15713 ^ n8620 ^ n8230 ;
  assign n23393 = n23392 ^ n9426 ^ n3158 ;
  assign n23394 = ( ~n3577 & n12751 ) | ( ~n3577 & n13207 ) | ( n12751 & n13207 ) ;
  assign n23395 = n23394 ^ n9848 ^ n9224 ;
  assign n23396 = n23395 ^ n18268 ^ n4878 ;
  assign n23397 = ( n5724 & n10845 ) | ( n5724 & ~n17062 ) | ( n10845 & ~n17062 ) ;
  assign n23398 = ( n14566 & n17268 ) | ( n14566 & n23397 ) | ( n17268 & n23397 ) ;
  assign n23399 = n10246 & ~n13757 ;
  assign n23400 = ~n7522 & n23399 ;
  assign n23402 = n22432 ^ n16683 ^ n2171 ;
  assign n23401 = n1805 | n3233 ;
  assign n23403 = n23402 ^ n23401 ^ n4912 ;
  assign n23404 = ( ~n234 & n9335 ) | ( ~n234 & n17555 ) | ( n9335 & n17555 ) ;
  assign n23405 = n23404 ^ n21225 ^ n1933 ;
  assign n23406 = n19624 ^ n5496 ^ n1074 ;
  assign n23407 = ( ~n5869 & n8944 ) | ( ~n5869 & n23406 ) | ( n8944 & n23406 ) ;
  assign n23408 = ( n10527 & n13316 ) | ( n10527 & n23407 ) | ( n13316 & n23407 ) ;
  assign n23409 = n23408 ^ n23048 ^ n17992 ;
  assign n23410 = n15932 ^ n2975 ^ x36 ;
  assign n23411 = n21188 ^ n13534 ^ n9397 ;
  assign n23412 = ( n3764 & n6111 ) | ( n3764 & n23411 ) | ( n6111 & n23411 ) ;
  assign n23413 = n22263 ^ n19784 ^ 1'b0 ;
  assign n23414 = n23413 ^ n11451 ^ n11161 ;
  assign n23415 = ( n1034 & ~n2824 ) | ( n1034 & n3870 ) | ( ~n2824 & n3870 ) ;
  assign n23416 = n19497 | n23415 ;
  assign n23417 = n23416 ^ n20838 ^ n6885 ;
  assign n23418 = n1723 & n3239 ;
  assign n23419 = n5686 & n15585 ;
  assign n23420 = n23419 ^ n11353 ^ n435 ;
  assign n23424 = ( n2470 & n8520 ) | ( n2470 & n10493 ) | ( n8520 & n10493 ) ;
  assign n23425 = n16083 ^ n15942 ^ n9707 ;
  assign n23426 = ( n21167 & n23424 ) | ( n21167 & ~n23425 ) | ( n23424 & ~n23425 ) ;
  assign n23421 = n14436 ^ n4423 ^ n2591 ;
  assign n23422 = ( n11688 & ~n13184 ) | ( n11688 & n20191 ) | ( ~n13184 & n20191 ) ;
  assign n23423 = ( n10616 & n23421 ) | ( n10616 & ~n23422 ) | ( n23421 & ~n23422 ) ;
  assign n23427 = n23426 ^ n23423 ^ n10103 ;
  assign n23428 = ( ~n1451 & n7544 ) | ( ~n1451 & n15487 ) | ( n7544 & n15487 ) ;
  assign n23429 = n23428 ^ n9851 ^ 1'b0 ;
  assign n23434 = n20923 ^ n12941 ^ n11709 ;
  assign n23430 = ( n2513 & ~n14812 ) | ( n2513 & n16621 ) | ( ~n14812 & n16621 ) ;
  assign n23431 = n23430 ^ n9396 ^ n1147 ;
  assign n23432 = n7040 ^ n2069 ^ 1'b0 ;
  assign n23433 = ( n5021 & n23431 ) | ( n5021 & n23432 ) | ( n23431 & n23432 ) ;
  assign n23435 = n23434 ^ n23433 ^ n16189 ;
  assign n23436 = n20635 ^ n15865 ^ n3379 ;
  assign n23437 = n23436 ^ n20295 ^ n10689 ;
  assign n23438 = n23437 ^ n10943 ^ n10729 ;
  assign n23439 = ~n436 & n19206 ;
  assign n23440 = ~n21368 & n23439 ;
  assign n23441 = n23440 ^ n8424 ^ n4959 ;
  assign n23442 = n7064 ^ n1857 ^ n1367 ;
  assign n23443 = n18219 ^ n15081 ^ n12426 ;
  assign n23444 = ( ~n4474 & n17326 ) | ( ~n4474 & n23443 ) | ( n17326 & n23443 ) ;
  assign n23445 = n23444 ^ n5242 ^ x51 ;
  assign n23446 = ( n1166 & n5559 ) | ( n1166 & ~n10401 ) | ( n5559 & ~n10401 ) ;
  assign n23447 = n23446 ^ n7315 ^ n6069 ;
  assign n23449 = ( n2306 & n2908 ) | ( n2306 & n5248 ) | ( n2908 & n5248 ) ;
  assign n23450 = n23449 ^ n4827 ^ n2058 ;
  assign n23451 = n10816 ^ n8061 ^ n7628 ;
  assign n23452 = ( ~n10683 & n23450 ) | ( ~n10683 & n23451 ) | ( n23450 & n23451 ) ;
  assign n23448 = n17991 ^ n13435 ^ n5791 ;
  assign n23453 = n23452 ^ n23448 ^ n13959 ;
  assign n23454 = ( n6568 & n15591 ) | ( n6568 & n18008 ) | ( n15591 & n18008 ) ;
  assign n23455 = n15930 ^ n2413 ^ n273 ;
  assign n23456 = n23455 ^ n11061 ^ 1'b0 ;
  assign n23457 = n23456 ^ n9084 ^ n8021 ;
  assign n23458 = ~n9891 & n23457 ;
  assign n23459 = n23458 ^ n10611 ^ 1'b0 ;
  assign n23460 = n11124 ^ n7469 ^ 1'b0 ;
  assign n23461 = n1284 & n23460 ;
  assign n23462 = x87 & n11421 ;
  assign n23463 = n23462 ^ n4384 ^ 1'b0 ;
  assign n23464 = ( ~n4765 & n6340 ) | ( ~n4765 & n7807 ) | ( n6340 & n7807 ) ;
  assign n23465 = ( n2063 & n9660 ) | ( n2063 & n23464 ) | ( n9660 & n23464 ) ;
  assign n23469 = ( n2728 & n5005 ) | ( n2728 & n17552 ) | ( n5005 & n17552 ) ;
  assign n23466 = ( n1511 & ~n6228 ) | ( n1511 & n10946 ) | ( ~n6228 & n10946 ) ;
  assign n23467 = n21312 & n23466 ;
  assign n23468 = n5887 & n23467 ;
  assign n23470 = n23469 ^ n23468 ^ n14711 ;
  assign n23473 = n12252 ^ n8070 ^ n1335 ;
  assign n23474 = n23473 ^ n8002 ^ n5252 ;
  assign n23475 = ( ~n1783 & n17973 ) | ( ~n1783 & n23474 ) | ( n17973 & n23474 ) ;
  assign n23476 = n23475 ^ n18100 ^ n10890 ;
  assign n23471 = n14628 ^ n11143 ^ 1'b0 ;
  assign n23472 = ( n1998 & n20288 ) | ( n1998 & ~n23471 ) | ( n20288 & ~n23471 ) ;
  assign n23477 = n23476 ^ n23472 ^ n1213 ;
  assign n23478 = n14337 ^ n13526 ^ n4333 ;
  assign n23479 = n11007 & ~n23478 ;
  assign n23480 = ( n7078 & n17276 ) | ( n7078 & ~n23479 ) | ( n17276 & ~n23479 ) ;
  assign n23481 = ( n1251 & n4171 ) | ( n1251 & n19588 ) | ( n4171 & n19588 ) ;
  assign n23482 = n23481 ^ n10849 ^ n183 ;
  assign n23483 = n23482 ^ n15395 ^ n10554 ;
  assign n23484 = n13125 ^ n11657 ^ n6694 ;
  assign n23485 = ( n17074 & n19632 ) | ( n17074 & ~n23484 ) | ( n19632 & ~n23484 ) ;
  assign n23486 = n19462 ^ n3591 ^ 1'b0 ;
  assign n23487 = n429 & ~n23486 ;
  assign n23488 = ( n2566 & n5314 ) | ( n2566 & ~n9602 ) | ( n5314 & ~n9602 ) ;
  assign n23489 = n9674 ^ n9360 ^ n442 ;
  assign n23490 = n9905 | n23489 ;
  assign n23491 = ( n4310 & ~n16272 ) | ( n4310 & n23490 ) | ( ~n16272 & n23490 ) ;
  assign n23492 = n23491 ^ n22369 ^ n15742 ;
  assign n23493 = n14752 ^ n4964 ^ n2823 ;
  assign n23494 = n21538 ^ n20466 ^ n4377 ;
  assign n23495 = n10609 ^ n9713 ^ n8927 ;
  assign n23496 = n19038 ^ n11771 ^ n8971 ;
  assign n23497 = n965 & n22179 ;
  assign n23498 = n23497 ^ n19723 ^ n7222 ;
  assign n23499 = n7608 ^ n5912 ^ n5078 ;
  assign n23500 = n8813 ^ n8203 ^ n1692 ;
  assign n23501 = n5781 & n11181 ;
  assign n23502 = n23500 & n23501 ;
  assign n23503 = ( n3709 & n23499 ) | ( n3709 & n23502 ) | ( n23499 & n23502 ) ;
  assign n23504 = ( n6088 & n20276 ) | ( n6088 & ~n21018 ) | ( n20276 & ~n21018 ) ;
  assign n23505 = n23504 ^ n18453 ^ n10787 ;
  assign n23506 = n5096 & ~n9942 ;
  assign n23507 = n16163 ^ n4790 ^ n2770 ;
  assign n23508 = ( n14854 & n23506 ) | ( n14854 & ~n23507 ) | ( n23506 & ~n23507 ) ;
  assign n23509 = n17968 ^ n13194 ^ n3178 ;
  assign n23510 = n12412 ^ n4306 ^ 1'b0 ;
  assign n23511 = ( n991 & n10883 ) | ( n991 & ~n17736 ) | ( n10883 & ~n17736 ) ;
  assign n23512 = ( ~n2025 & n5296 ) | ( ~n2025 & n8118 ) | ( n5296 & n8118 ) ;
  assign n23513 = n23512 ^ n2579 ^ 1'b0 ;
  assign n23514 = ~n3559 & n23513 ;
  assign n23515 = ( ~n9452 & n17940 ) | ( ~n9452 & n23514 ) | ( n17940 & n23514 ) ;
  assign n23516 = ( n10443 & n23511 ) | ( n10443 & n23515 ) | ( n23511 & n23515 ) ;
  assign n23517 = n22698 ^ n16090 ^ n6613 ;
  assign n23518 = n23517 ^ n3597 ^ n745 ;
  assign n23521 = n2591 ^ n955 ^ n839 ;
  assign n23520 = ( n194 & ~n5550 ) | ( n194 & n11648 ) | ( ~n5550 & n11648 ) ;
  assign n23522 = n23521 ^ n23520 ^ n13912 ;
  assign n23519 = n11243 ^ n7530 ^ n3046 ;
  assign n23523 = n23522 ^ n23519 ^ n21262 ;
  assign n23524 = ( n3986 & n11376 ) | ( n3986 & ~n20862 ) | ( n11376 & ~n20862 ) ;
  assign n23525 = n15552 ^ n15038 ^ n1918 ;
  assign n23526 = ( n10787 & ~n10887 ) | ( n10787 & n15153 ) | ( ~n10887 & n15153 ) ;
  assign n23527 = n16825 ^ n5533 ^ n1342 ;
  assign n23528 = n23527 ^ n18545 ^ n5259 ;
  assign n23529 = n15121 ^ n1511 ^ 1'b0 ;
  assign n23530 = ( ~n23526 & n23528 ) | ( ~n23526 & n23529 ) | ( n23528 & n23529 ) ;
  assign n23531 = n15170 ^ n748 ^ 1'b0 ;
  assign n23532 = ~n2353 & n23531 ;
  assign n23533 = ( ~n6342 & n13282 ) | ( ~n6342 & n17142 ) | ( n13282 & n17142 ) ;
  assign n23534 = n472 & ~n23533 ;
  assign n23535 = n23534 ^ n19611 ^ 1'b0 ;
  assign n23536 = ( ~n11426 & n23532 ) | ( ~n11426 & n23535 ) | ( n23532 & n23535 ) ;
  assign n23537 = ( n782 & ~n2667 ) | ( n782 & n15325 ) | ( ~n2667 & n15325 ) ;
  assign n23538 = n1486 | n11091 ;
  assign n23539 = n23538 ^ n216 ^ 1'b0 ;
  assign n23540 = ( n18488 & ~n23537 ) | ( n18488 & n23539 ) | ( ~n23537 & n23539 ) ;
  assign n23541 = n2250 | n18743 ;
  assign n23542 = n22688 & ~n23541 ;
  assign n23543 = n11363 ^ n2182 ^ 1'b0 ;
  assign n23544 = n23543 ^ n16432 ^ n6765 ;
  assign n23545 = n21759 ^ n14315 ^ 1'b0 ;
  assign n23546 = ( n15052 & ~n21536 ) | ( n15052 & n23545 ) | ( ~n21536 & n23545 ) ;
  assign n23547 = n4123 ^ n3414 ^ n2810 ;
  assign n23548 = ( n11093 & ~n16460 ) | ( n11093 & n23547 ) | ( ~n16460 & n23547 ) ;
  assign n23549 = n12331 ^ n7330 ^ n6170 ;
  assign n23550 = ( n9443 & n10431 ) | ( n9443 & n23549 ) | ( n10431 & n23549 ) ;
  assign n23551 = ( n6299 & n23269 ) | ( n6299 & n23550 ) | ( n23269 & n23550 ) ;
  assign n23552 = n15110 ^ n10613 ^ n8900 ;
  assign n23554 = n6276 & ~n7553 ;
  assign n23555 = n23554 ^ n696 ^ 1'b0 ;
  assign n23553 = n10060 ^ n7443 ^ 1'b0 ;
  assign n23556 = n23555 ^ n23553 ^ n12042 ;
  assign n23558 = n15307 ^ n4638 ^ n4099 ;
  assign n23557 = ( n7874 & ~n15696 ) | ( n7874 & n20723 ) | ( ~n15696 & n20723 ) ;
  assign n23559 = n23558 ^ n23557 ^ n2828 ;
  assign n23564 = n1965 | n7726 ;
  assign n23565 = n23564 ^ n1055 ^ 1'b0 ;
  assign n23562 = ~n5006 & n6369 ;
  assign n23563 = n23562 ^ n11645 ^ 1'b0 ;
  assign n23560 = n1584 & ~n7546 ;
  assign n23561 = n23560 ^ n21716 ^ n8578 ;
  assign n23566 = n23565 ^ n23563 ^ n23561 ;
  assign n23567 = n11439 ^ n10206 ^ n5808 ;
  assign n23568 = n13355 | n23567 ;
  assign n23569 = n23568 ^ n6283 ^ 1'b0 ;
  assign n23570 = ( n2066 & n8092 ) | ( n2066 & ~n9259 ) | ( n8092 & ~n9259 ) ;
  assign n23571 = n23570 ^ n9127 ^ n7416 ;
  assign n23572 = ( n13678 & ~n23569 ) | ( n13678 & n23571 ) | ( ~n23569 & n23571 ) ;
  assign n23573 = ( n3651 & n11081 ) | ( n3651 & ~n23572 ) | ( n11081 & ~n23572 ) ;
  assign n23574 = n23573 ^ n19217 ^ n528 ;
  assign n23575 = ( n11495 & n15370 ) | ( n11495 & n21470 ) | ( n15370 & n21470 ) ;
  assign n23576 = ( ~n482 & n11216 ) | ( ~n482 & n19687 ) | ( n11216 & n19687 ) ;
  assign n23577 = n13437 & n23576 ;
  assign n23578 = n12419 & n23577 ;
  assign n23579 = n11439 & ~n15653 ;
  assign n23580 = ~n2712 & n23579 ;
  assign n23581 = n18127 ^ n5161 ^ 1'b0 ;
  assign n23582 = ( n11553 & n23580 ) | ( n11553 & ~n23581 ) | ( n23580 & ~n23581 ) ;
  assign n23583 = ( ~n2342 & n13986 ) | ( ~n2342 & n18881 ) | ( n13986 & n18881 ) ;
  assign n23584 = n956 & ~n4499 ;
  assign n23585 = ( n3669 & n7763 ) | ( n3669 & n23584 ) | ( n7763 & n23584 ) ;
  assign n23586 = ( n12612 & ~n15746 ) | ( n12612 & n23585 ) | ( ~n15746 & n23585 ) ;
  assign n23587 = ( n2935 & ~n17363 ) | ( n2935 & n23586 ) | ( ~n17363 & n23586 ) ;
  assign n23588 = n23587 ^ n12109 ^ n11686 ;
  assign n23589 = ( n948 & ~n3272 ) | ( n948 & n8393 ) | ( ~n3272 & n8393 ) ;
  assign n23590 = ( n15942 & n18405 ) | ( n15942 & ~n23589 ) | ( n18405 & ~n23589 ) ;
  assign n23591 = n5610 ^ n3053 ^ n1104 ;
  assign n23594 = n17796 ^ n11076 ^ n10274 ;
  assign n23592 = n23452 ^ n22082 ^ n4374 ;
  assign n23593 = ~n1901 & n23592 ;
  assign n23595 = n23594 ^ n23593 ^ 1'b0 ;
  assign n23596 = n6309 ^ n1351 ^ 1'b0 ;
  assign n23597 = n5053 & ~n23596 ;
  assign n23598 = n23597 ^ n10275 ^ n5735 ;
  assign n23599 = ( ~n1282 & n8706 ) | ( ~n1282 & n12518 ) | ( n8706 & n12518 ) ;
  assign n23600 = ( n2932 & n21395 ) | ( n2932 & n23599 ) | ( n21395 & n23599 ) ;
  assign n23601 = ( n2536 & ~n23598 ) | ( n2536 & n23600 ) | ( ~n23598 & n23600 ) ;
  assign n23602 = n12433 | n16454 ;
  assign n23603 = n9570 ^ n1187 ^ 1'b0 ;
  assign n23604 = n23603 ^ n9224 ^ n1140 ;
  assign n23605 = n23604 ^ n23182 ^ n1074 ;
  assign n23606 = ( n3059 & n7671 ) | ( n3059 & n23605 ) | ( n7671 & n23605 ) ;
  assign n23607 = ( ~n692 & n10665 ) | ( ~n692 & n10877 ) | ( n10665 & n10877 ) ;
  assign n23608 = ( n10332 & n10590 ) | ( n10332 & ~n12597 ) | ( n10590 & ~n12597 ) ;
  assign n23609 = n23608 ^ n19004 ^ n1261 ;
  assign n23610 = n14764 ^ n9464 ^ n3698 ;
  assign n23611 = n15785 ^ n5694 ^ x70 ;
  assign n23612 = n23611 ^ n8907 ^ 1'b0 ;
  assign n23613 = ( n10394 & ~n23610 ) | ( n10394 & n23612 ) | ( ~n23610 & n23612 ) ;
  assign n23614 = ( ~n17869 & n23609 ) | ( ~n17869 & n23613 ) | ( n23609 & n23613 ) ;
  assign n23615 = n1104 & ~n14208 ;
  assign n23616 = n23615 ^ n15047 ^ 1'b0 ;
  assign n23617 = n2995 & ~n19378 ;
  assign n23618 = n23617 ^ n16874 ^ 1'b0 ;
  assign n23619 = n23618 ^ n20600 ^ n5826 ;
  assign n23622 = n1372 & ~n9519 ;
  assign n23620 = n12885 & ~n13820 ;
  assign n23621 = n23620 ^ n8869 ^ n4226 ;
  assign n23623 = n23622 ^ n23621 ^ n17060 ;
  assign n23627 = n14627 & ~n15099 ;
  assign n23628 = n23627 ^ n14227 ^ 1'b0 ;
  assign n23624 = n10488 | n13985 ;
  assign n23625 = ~n13487 & n23624 ;
  assign n23626 = n23625 ^ n9313 ^ 1'b0 ;
  assign n23629 = n23628 ^ n23626 ^ n13198 ;
  assign n23630 = n8533 ^ n5275 ^ 1'b0 ;
  assign n23631 = ( n6060 & n20438 ) | ( n6060 & n23630 ) | ( n20438 & n23630 ) ;
  assign n23632 = ( x9 & n4482 ) | ( x9 & ~n8610 ) | ( n4482 & ~n8610 ) ;
  assign n23633 = ( n783 & n913 ) | ( n783 & ~n2183 ) | ( n913 & ~n2183 ) ;
  assign n23634 = n23633 ^ n5150 ^ n258 ;
  assign n23635 = ( n1287 & ~n23632 ) | ( n1287 & n23634 ) | ( ~n23632 & n23634 ) ;
  assign n23636 = n1695 & ~n23635 ;
  assign n23637 = n14490 ^ n10992 ^ n6174 ;
  assign n23638 = ( n4933 & n8606 ) | ( n4933 & ~n13814 ) | ( n8606 & ~n13814 ) ;
  assign n23639 = n23638 ^ n15872 ^ n2055 ;
  assign n23640 = n4303 ^ n1103 ^ 1'b0 ;
  assign n23642 = n11279 ^ n10425 ^ n9909 ;
  assign n23643 = n23642 ^ n5910 ^ n1605 ;
  assign n23641 = n11522 ^ n10464 ^ n4774 ;
  assign n23644 = n23643 ^ n23641 ^ n20869 ;
  assign n23645 = ( n3373 & ~n9542 ) | ( n3373 & n10716 ) | ( ~n9542 & n10716 ) ;
  assign n23646 = ( n5294 & n11723 ) | ( n5294 & ~n23645 ) | ( n11723 & ~n23645 ) ;
  assign n23647 = n23646 ^ n15913 ^ n12671 ;
  assign n23648 = n17625 ^ n15174 ^ n10400 ;
  assign n23649 = n23648 ^ n18816 ^ n11902 ;
  assign n23650 = n8501 ^ n6918 ^ n3036 ;
  assign n23651 = n14861 ^ n14815 ^ x12 ;
  assign n23652 = n23651 ^ n22072 ^ n4270 ;
  assign n23654 = n21539 ^ n4134 ^ 1'b0 ;
  assign n23653 = ( n4610 & n14855 ) | ( n4610 & n21763 ) | ( n14855 & n21763 ) ;
  assign n23655 = n23654 ^ n23653 ^ n11193 ;
  assign n23656 = n2373 & n3307 ;
  assign n23657 = n5076 | n8502 ;
  assign n23658 = n7412 & ~n23657 ;
  assign n23659 = ( n4655 & n5026 ) | ( n4655 & n8783 ) | ( n5026 & n8783 ) ;
  assign n23660 = n23659 ^ n3145 ^ 1'b0 ;
  assign n23661 = ( n23656 & n23658 ) | ( n23656 & n23660 ) | ( n23658 & n23660 ) ;
  assign n23662 = n9528 ^ n7454 ^ n3554 ;
  assign n23663 = ~n16263 & n23662 ;
  assign n23664 = n23663 ^ n5554 ^ 1'b0 ;
  assign n23665 = n3648 | n23449 ;
  assign n23666 = ~n7813 & n23665 ;
  assign n23669 = n10990 ^ n7349 ^ n1339 ;
  assign n23667 = ~n16361 & n23382 ;
  assign n23668 = n23667 ^ n14077 ^ 1'b0 ;
  assign n23670 = n23669 ^ n23668 ^ n9523 ;
  assign n23671 = ( ~n8704 & n17824 ) | ( ~n8704 & n23670 ) | ( n17824 & n23670 ) ;
  assign n23672 = n6696 ^ n6640 ^ n4130 ;
  assign n23673 = n23672 ^ n5678 ^ n2731 ;
  assign n23674 = ( n14874 & n20276 ) | ( n14874 & ~n22215 ) | ( n20276 & ~n22215 ) ;
  assign n23675 = ( n3539 & n4315 ) | ( n3539 & n8604 ) | ( n4315 & n8604 ) ;
  assign n23676 = ( n9937 & n10867 ) | ( n9937 & n23675 ) | ( n10867 & n23675 ) ;
  assign n23677 = ( n7971 & n9749 ) | ( n7971 & n22258 ) | ( n9749 & n22258 ) ;
  assign n23678 = n23677 ^ n18475 ^ n5709 ;
  assign n23679 = ( n3446 & n7003 ) | ( n3446 & ~n12063 ) | ( n7003 & ~n12063 ) ;
  assign n23680 = n7879 & n10287 ;
  assign n23681 = ( ~n1531 & n8902 ) | ( ~n1531 & n14063 ) | ( n8902 & n14063 ) ;
  assign n23682 = n12549 | n23681 ;
  assign n23683 = n23682 ^ n6991 ^ 1'b0 ;
  assign n23684 = n1247 ^ n582 ^ 1'b0 ;
  assign n23685 = n23684 ^ n13821 ^ n4814 ;
  assign n23686 = ( n3403 & n5390 ) | ( n3403 & n11737 ) | ( n5390 & n11737 ) ;
  assign n23687 = n17729 & ~n18237 ;
  assign n23688 = ~n23686 & n23687 ;
  assign n23689 = ( n6623 & n10992 ) | ( n6623 & n12154 ) | ( n10992 & n12154 ) ;
  assign n23690 = n23689 ^ n5061 ^ x15 ;
  assign n23691 = ( ~n720 & n1341 ) | ( ~n720 & n1388 ) | ( n1341 & n1388 ) ;
  assign n23692 = ( n2031 & ~n12584 ) | ( n2031 & n23691 ) | ( ~n12584 & n23691 ) ;
  assign n23693 = ( ~n1248 & n2786 ) | ( ~n1248 & n4236 ) | ( n2786 & n4236 ) ;
  assign n23694 = ( ~n12502 & n13208 ) | ( ~n12502 & n23693 ) | ( n13208 & n23693 ) ;
  assign n23695 = ( n3589 & n14869 ) | ( n3589 & n15477 ) | ( n14869 & n15477 ) ;
  assign n23696 = n23506 ^ n17031 ^ n3533 ;
  assign n23697 = ( n2170 & n6807 ) | ( n2170 & ~n23696 ) | ( n6807 & ~n23696 ) ;
  assign n23698 = n7778 ^ n2272 ^ 1'b0 ;
  assign n23699 = ( n21607 & n23697 ) | ( n21607 & ~n23698 ) | ( n23697 & ~n23698 ) ;
  assign n23700 = ( n9794 & ~n17690 ) | ( n9794 & n21260 ) | ( ~n17690 & n21260 ) ;
  assign n23701 = n15583 ^ n9412 ^ n7344 ;
  assign n23702 = ( n14647 & ~n23489 ) | ( n14647 & n23701 ) | ( ~n23489 & n23701 ) ;
  assign n23704 = n279 & n5719 ;
  assign n23703 = ( n5069 & ~n9503 ) | ( n5069 & n19244 ) | ( ~n9503 & n19244 ) ;
  assign n23705 = n23704 ^ n23703 ^ n23446 ;
  assign n23706 = n2661 & ~n17873 ;
  assign n23707 = ~n22436 & n23706 ;
  assign n23715 = n8926 ^ n5368 ^ n3925 ;
  assign n23712 = ~n4089 & n8890 ;
  assign n23713 = n23712 ^ n10721 ^ 1'b0 ;
  assign n23714 = n23713 ^ n12475 ^ n3813 ;
  assign n23716 = n23715 ^ n23714 ^ n13891 ;
  assign n23717 = n21664 ^ n14124 ^ 1'b0 ;
  assign n23718 = ~n23716 & n23717 ;
  assign n23709 = n6437 ^ n2162 ^ n1620 ;
  assign n23708 = ( ~n10502 & n13702 ) | ( ~n10502 & n17965 ) | ( n13702 & n17965 ) ;
  assign n23710 = n23709 ^ n23708 ^ 1'b0 ;
  assign n23711 = ( ~n8758 & n16309 ) | ( ~n8758 & n23710 ) | ( n16309 & n23710 ) ;
  assign n23719 = n23718 ^ n23711 ^ n13779 ;
  assign n23720 = ( n6591 & n14369 ) | ( n6591 & n23408 ) | ( n14369 & n23408 ) ;
  assign n23721 = ( ~n6396 & n7407 ) | ( ~n6396 & n14945 ) | ( n7407 & n14945 ) ;
  assign n23722 = ~n21190 & n21255 ;
  assign n23723 = ( n4368 & n12448 ) | ( n4368 & ~n12942 ) | ( n12448 & ~n12942 ) ;
  assign n23724 = n12370 ^ n5143 ^ n2194 ;
  assign n23725 = n23724 ^ n4536 ^ n532 ;
  assign n23726 = n20475 ^ n14404 ^ n6660 ;
  assign n23732 = n14383 ^ n7015 ^ n4400 ;
  assign n23730 = n9136 ^ n7266 ^ n6050 ;
  assign n23727 = ( n1133 & n16231 ) | ( n1133 & ~n17384 ) | ( n16231 & ~n17384 ) ;
  assign n23728 = n4064 ^ n796 ^ 1'b0 ;
  assign n23729 = n23727 | n23728 ;
  assign n23731 = n23730 ^ n23729 ^ n19284 ;
  assign n23733 = n23732 ^ n23731 ^ n4807 ;
  assign n23734 = n19743 ^ n15794 ^ 1'b0 ;
  assign n23735 = ( n15526 & ~n23529 ) | ( n15526 & n23734 ) | ( ~n23529 & n23734 ) ;
  assign n23738 = n12050 ^ n566 ^ n204 ;
  assign n23736 = n20138 ^ n17090 ^ n14337 ;
  assign n23737 = ( n13798 & n19170 ) | ( n13798 & ~n23736 ) | ( n19170 & ~n23736 ) ;
  assign n23739 = n23738 ^ n23737 ^ n12784 ;
  assign n23740 = ( n2766 & ~n6387 ) | ( n2766 & n18406 ) | ( ~n6387 & n18406 ) ;
  assign n23741 = n23740 ^ n19585 ^ n6251 ;
  assign n23742 = n23741 ^ n23504 ^ n22146 ;
  assign n23743 = n15915 ^ n12565 ^ n7442 ;
  assign n23744 = n23743 ^ n8799 ^ n184 ;
  assign n23746 = ~n1141 & n1243 ;
  assign n23745 = n15374 ^ n7958 ^ n4212 ;
  assign n23747 = n23746 ^ n23745 ^ x79 ;
  assign n23748 = n23747 ^ n11251 ^ 1'b0 ;
  assign n23749 = ~n11529 & n23748 ;
  assign n23750 = ( n2340 & ~n5389 ) | ( n2340 & n10669 ) | ( ~n5389 & n10669 ) ;
  assign n23751 = n23750 ^ n21497 ^ n5568 ;
  assign n23752 = n5196 ^ n243 ^ 1'b0 ;
  assign n23753 = ( ~n8569 & n8971 ) | ( ~n8569 & n23752 ) | ( n8971 & n23752 ) ;
  assign n23754 = ( ~n4359 & n12766 ) | ( ~n4359 & n14366 ) | ( n12766 & n14366 ) ;
  assign n23755 = ( ~n8267 & n12255 ) | ( ~n8267 & n23754 ) | ( n12255 & n23754 ) ;
  assign n23756 = n17848 ^ n3392 ^ 1'b0 ;
  assign n23757 = ( n4313 & n23755 ) | ( n4313 & n23756 ) | ( n23755 & n23756 ) ;
  assign n23758 = ( n10069 & n17421 ) | ( n10069 & n19459 ) | ( n17421 & n19459 ) ;
  assign n23759 = n15353 ^ n7452 ^ n163 ;
  assign n23760 = n23759 ^ n22052 ^ n21371 ;
  assign n23761 = n16680 ^ n15904 ^ 1'b0 ;
  assign n23762 = ( n5398 & n17268 ) | ( n5398 & n20916 ) | ( n17268 & n20916 ) ;
  assign n23763 = ( n9570 & n16247 ) | ( n9570 & ~n17276 ) | ( n16247 & ~n17276 ) ;
  assign n23764 = n23763 ^ n14738 ^ 1'b0 ;
  assign n23765 = n23762 & n23764 ;
  assign n23766 = n571 & n4609 ;
  assign n23767 = n9985 ^ n6598 ^ n779 ;
  assign n23768 = ( ~n3381 & n23766 ) | ( ~n3381 & n23767 ) | ( n23766 & n23767 ) ;
  assign n23769 = n2201 | n6919 ;
  assign n23770 = ~n2309 & n23769 ;
  assign n23771 = n23770 ^ n21347 ^ n15424 ;
  assign n23772 = n8239 ^ n5494 ^ 1'b0 ;
  assign n23773 = ~n12106 & n23772 ;
  assign n23774 = n23773 ^ n16605 ^ n5149 ;
  assign n23775 = ( x99 & ~n2712 ) | ( x99 & n9212 ) | ( ~n2712 & n9212 ) ;
  assign n23776 = n7626 & n8621 ;
  assign n23777 = n2947 & n23776 ;
  assign n23778 = ( n2426 & n13720 ) | ( n2426 & n21109 ) | ( n13720 & n21109 ) ;
  assign n23779 = n13720 ^ n1580 ^ n189 ;
  assign n23781 = n10519 ^ n2753 ^ 1'b0 ;
  assign n23780 = ( n226 & n7442 ) | ( n226 & n11233 ) | ( n7442 & n11233 ) ;
  assign n23782 = n23781 ^ n23780 ^ n16280 ;
  assign n23783 = n18886 ^ n2388 ^ 1'b0 ;
  assign n23784 = ( ~n9391 & n14231 ) | ( ~n9391 & n19158 ) | ( n14231 & n19158 ) ;
  assign n23785 = n19270 ^ n5390 ^ 1'b0 ;
  assign n23786 = ( n1320 & n12086 ) | ( n1320 & ~n23785 ) | ( n12086 & ~n23785 ) ;
  assign n23787 = ( n2616 & n2766 ) | ( n2616 & ~n11912 ) | ( n2766 & ~n11912 ) ;
  assign n23788 = ( ~n15265 & n20059 ) | ( ~n15265 & n23787 ) | ( n20059 & n23787 ) ;
  assign n23789 = n4245 | n9694 ;
  assign n23790 = n21552 & ~n23789 ;
  assign n23791 = n21487 ^ n18101 ^ 1'b0 ;
  assign n23792 = n3940 | n23791 ;
  assign n23793 = n22344 ^ n16420 ^ n11140 ;
  assign n23794 = n7681 | n9424 ;
  assign n23795 = n14206 | n23794 ;
  assign n23796 = ( ~x59 & n3246 ) | ( ~x59 & n23795 ) | ( n3246 & n23795 ) ;
  assign n23797 = ( n1452 & n2726 ) | ( n1452 & ~n23796 ) | ( n2726 & ~n23796 ) ;
  assign n23798 = ( ~n4146 & n23793 ) | ( ~n4146 & n23797 ) | ( n23793 & n23797 ) ;
  assign n23799 = ( n2977 & n5290 ) | ( n2977 & ~n14241 ) | ( n5290 & ~n14241 ) ;
  assign n23800 = n15461 ^ n14656 ^ 1'b0 ;
  assign n23801 = ( n21411 & n22378 ) | ( n21411 & n23800 ) | ( n22378 & n23800 ) ;
  assign n23802 = n23799 & n23801 ;
  assign n23803 = n5109 & ~n7193 ;
  assign n23804 = n23803 ^ n6189 ^ 1'b0 ;
  assign n23805 = n23804 ^ n15954 ^ n504 ;
  assign n23806 = n15389 ^ n10321 ^ n1730 ;
  assign n23807 = ( n14792 & n23805 ) | ( n14792 & n23806 ) | ( n23805 & n23806 ) ;
  assign n23808 = ( n9968 & n17696 ) | ( n9968 & ~n20699 ) | ( n17696 & ~n20699 ) ;
  assign n23809 = ( n6405 & ~n9833 ) | ( n6405 & n16375 ) | ( ~n9833 & n16375 ) ;
  assign n23810 = n23809 ^ n9540 ^ n2538 ;
  assign n23811 = n23810 ^ n1280 ^ 1'b0 ;
  assign n23812 = ( ~n13619 & n23808 ) | ( ~n13619 & n23811 ) | ( n23808 & n23811 ) ;
  assign n23813 = ( n3127 & n7966 ) | ( n3127 & ~n11481 ) | ( n7966 & ~n11481 ) ;
  assign n23814 = ( n8854 & n10599 ) | ( n8854 & n23813 ) | ( n10599 & n23813 ) ;
  assign n23815 = n23814 ^ n11494 ^ n2040 ;
  assign n23816 = ( n1983 & n4433 ) | ( n1983 & n4864 ) | ( n4433 & n4864 ) ;
  assign n23817 = ( n4139 & n6889 ) | ( n4139 & n23816 ) | ( n6889 & n23816 ) ;
  assign n23818 = n23817 ^ n23105 ^ 1'b0 ;
  assign n23819 = n11511 ^ n6922 ^ n4987 ;
  assign n23820 = n20386 ^ n12037 ^ n6910 ;
  assign n23821 = n3835 ^ n2507 ^ n818 ;
  assign n23822 = n11982 ^ n567 ^ n282 ;
  assign n23823 = n23822 ^ n11853 ^ 1'b0 ;
  assign n23824 = ( n6838 & n14580 ) | ( n6838 & ~n23823 ) | ( n14580 & ~n23823 ) ;
  assign n23825 = n23824 ^ n18758 ^ n7837 ;
  assign n23826 = ( n5822 & n23821 ) | ( n5822 & n23825 ) | ( n23821 & n23825 ) ;
  assign n23827 = n13299 ^ n7794 ^ n1373 ;
  assign n23828 = ~n2933 & n13377 ;
  assign n23829 = n23828 ^ n17081 ^ n16054 ;
  assign n23830 = n14965 ^ n7416 ^ n3308 ;
  assign n23831 = n1502 & n23830 ;
  assign n23832 = ~n23475 & n23831 ;
  assign n23833 = n2634 & ~n23648 ;
  assign n23834 = n23833 ^ n6636 ^ 1'b0 ;
  assign n23835 = ( ~n4780 & n11215 ) | ( ~n4780 & n23834 ) | ( n11215 & n23834 ) ;
  assign n23836 = n22723 ^ n7117 ^ 1'b0 ;
  assign n23837 = ( n5490 & ~n11663 ) | ( n5490 & n19047 ) | ( ~n11663 & n19047 ) ;
  assign n23838 = n10153 ^ n1926 ^ 1'b0 ;
  assign n23839 = ( n697 & n5458 ) | ( n697 & n8383 ) | ( n5458 & n8383 ) ;
  assign n23840 = n23839 ^ n5351 ^ n2489 ;
  assign n23841 = n23840 ^ n8117 ^ n7717 ;
  assign n23842 = n3697 & ~n6278 ;
  assign n23843 = ~n3021 & n23842 ;
  assign n23844 = n11498 & n23843 ;
  assign n23845 = n13868 ^ n9334 ^ n199 ;
  assign n23850 = n2324 ^ n2147 ^ n1275 ;
  assign n23849 = ( ~n3454 & n13493 ) | ( ~n3454 & n16370 ) | ( n13493 & n16370 ) ;
  assign n23846 = n19793 ^ n16495 ^ n13036 ;
  assign n23847 = n15907 & n23846 ;
  assign n23848 = n22841 & n23847 ;
  assign n23851 = n23850 ^ n23849 ^ n23848 ;
  assign n23852 = n10741 ^ n6100 ^ 1'b0 ;
  assign n23853 = ~n17379 & n23852 ;
  assign n23854 = ( n1849 & n12904 ) | ( n1849 & ~n23853 ) | ( n12904 & ~n23853 ) ;
  assign n23855 = ( n10136 & n15339 ) | ( n10136 & ~n23854 ) | ( n15339 & ~n23854 ) ;
  assign n23856 = n15733 & n22955 ;
  assign n23857 = ( ~n7059 & n23718 ) | ( ~n7059 & n23856 ) | ( n23718 & n23856 ) ;
  assign n23858 = n17232 ^ n3304 ^ 1'b0 ;
  assign n23861 = n870 & ~n4218 ;
  assign n23862 = n23861 ^ n18148 ^ 1'b0 ;
  assign n23859 = n4780 ^ n4339 ^ n2574 ;
  assign n23860 = ( n9609 & n11015 ) | ( n9609 & ~n23859 ) | ( n11015 & ~n23859 ) ;
  assign n23863 = n23862 ^ n23860 ^ n15020 ;
  assign n23864 = ( n699 & n3594 ) | ( n699 & n19434 ) | ( n3594 & n19434 ) ;
  assign n23865 = n14358 ^ n4770 ^ 1'b0 ;
  assign n23866 = n16272 ^ n3817 ^ n3293 ;
  assign n23867 = ( n390 & n1608 ) | ( n390 & n7330 ) | ( n1608 & n7330 ) ;
  assign n23868 = ( ~n11723 & n22277 ) | ( ~n11723 & n23867 ) | ( n22277 & n23867 ) ;
  assign n23869 = n23868 ^ n17237 ^ n4862 ;
  assign n23870 = n23859 ^ n17638 ^ n13443 ;
  assign n23871 = ( n16154 & ~n23869 ) | ( n16154 & n23870 ) | ( ~n23869 & n23870 ) ;
  assign n23872 = ( n4236 & n10713 ) | ( n4236 & n11948 ) | ( n10713 & n11948 ) ;
  assign n23873 = n22421 ^ n19937 ^ n10449 ;
  assign n23874 = n8966 ^ n2260 ^ n1179 ;
  assign n23875 = ( n4094 & n9757 ) | ( n4094 & n23874 ) | ( n9757 & n23874 ) ;
  assign n23876 = n8988 ^ n5960 ^ n5180 ;
  assign n23877 = ( n1055 & ~n14384 ) | ( n1055 & n23876 ) | ( ~n14384 & n23876 ) ;
  assign n23878 = n19155 ^ n15808 ^ n1630 ;
  assign n23879 = n23878 ^ n20289 ^ 1'b0 ;
  assign n23880 = n19952 ^ n6416 ^ n249 ;
  assign n23881 = ( n6066 & n6598 ) | ( n6066 & ~n13756 ) | ( n6598 & ~n13756 ) ;
  assign n23882 = ( n1693 & n4817 ) | ( n1693 & n11652 ) | ( n4817 & n11652 ) ;
  assign n23883 = n19737 ^ n10923 ^ n3255 ;
  assign n23884 = ( n2823 & n14369 ) | ( n2823 & ~n23883 ) | ( n14369 & ~n23883 ) ;
  assign n23885 = ( n6534 & n11959 ) | ( n6534 & ~n23884 ) | ( n11959 & ~n23884 ) ;
  assign n23886 = ( n22358 & n23882 ) | ( n22358 & n23885 ) | ( n23882 & n23885 ) ;
  assign n23887 = n6223 ^ n1008 ^ 1'b0 ;
  assign n23888 = ( n423 & ~n6068 ) | ( n423 & n23887 ) | ( ~n6068 & n23887 ) ;
  assign n23889 = n129 & ~n14908 ;
  assign n23890 = n13937 & n23889 ;
  assign n23891 = ( n201 & ~n12379 ) | ( n201 & n23890 ) | ( ~n12379 & n23890 ) ;
  assign n23892 = n10207 ^ n7565 ^ n3925 ;
  assign n23893 = ( n7568 & ~n21188 ) | ( n7568 & n22664 ) | ( ~n21188 & n22664 ) ;
  assign n23894 = n23893 ^ n23658 ^ n7522 ;
  assign n23895 = ( ~n1628 & n7434 ) | ( ~n1628 & n16118 ) | ( n7434 & n16118 ) ;
  assign n23896 = ~n15448 & n23895 ;
  assign n23902 = ~n721 & n1595 ;
  assign n23903 = n23902 ^ n406 ^ 1'b0 ;
  assign n23899 = n985 | n5161 ;
  assign n23900 = n23899 ^ n18273 ^ 1'b0 ;
  assign n23898 = n3482 | n14117 ;
  assign n23901 = n23900 ^ n23898 ^ 1'b0 ;
  assign n23897 = ~n6278 & n7196 ;
  assign n23904 = n23903 ^ n23901 ^ n23897 ;
  assign n23905 = ( n268 & ~n14956 ) | ( n268 & n23904 ) | ( ~n14956 & n23904 ) ;
  assign n23906 = ( n7528 & n16156 ) | ( n7528 & ~n20927 ) | ( n16156 & ~n20927 ) ;
  assign n23912 = n8764 | n13281 ;
  assign n23907 = n18171 ^ n11722 ^ n2018 ;
  assign n23908 = ( ~n10093 & n10584 ) | ( ~n10093 & n23907 ) | ( n10584 & n23907 ) ;
  assign n23909 = ( n10809 & ~n14457 ) | ( n10809 & n23908 ) | ( ~n14457 & n23908 ) ;
  assign n23910 = ( n5853 & n13610 ) | ( n5853 & n23909 ) | ( n13610 & n23909 ) ;
  assign n23911 = n23910 ^ n16526 ^ n15334 ;
  assign n23913 = n23912 ^ n23911 ^ n3338 ;
  assign n23914 = ( n5351 & n8211 ) | ( n5351 & n12466 ) | ( n8211 & n12466 ) ;
  assign n23915 = ( n12491 & n19223 ) | ( n12491 & ~n23914 ) | ( n19223 & ~n23914 ) ;
  assign n23916 = n23915 ^ n3263 ^ n466 ;
  assign n23917 = n23916 ^ n18585 ^ n14664 ;
  assign n23918 = ( n304 & ~n1815 ) | ( n304 & n6400 ) | ( ~n1815 & n6400 ) ;
  assign n23919 = ( n513 & n22538 ) | ( n513 & n23918 ) | ( n22538 & n23918 ) ;
  assign n23920 = ( n3781 & n6608 ) | ( n3781 & n13901 ) | ( n6608 & n13901 ) ;
  assign n23921 = n19636 ^ n16231 ^ n14584 ;
  assign n23922 = ( n220 & ~n14302 ) | ( n220 & n14455 ) | ( ~n14302 & n14455 ) ;
  assign n23923 = n1838 | n22957 ;
  assign n23924 = ( n977 & ~n18933 ) | ( n977 & n23923 ) | ( ~n18933 & n23923 ) ;
  assign n23925 = n23075 ^ n15933 ^ n6267 ;
  assign n23926 = ( ~n23922 & n23924 ) | ( ~n23922 & n23925 ) | ( n23924 & n23925 ) ;
  assign n23927 = ( n879 & n6027 ) | ( n879 & ~n21508 ) | ( n6027 & ~n21508 ) ;
  assign n23928 = n9853 & ~n23927 ;
  assign n23929 = n254 & n5922 ;
  assign n23930 = n23929 ^ n4631 ^ 1'b0 ;
  assign n23933 = n10121 ^ n3239 ^ n1291 ;
  assign n23931 = n12700 ^ n10993 ^ n466 ;
  assign n23932 = ( ~n3698 & n18165 ) | ( ~n3698 & n23931 ) | ( n18165 & n23931 ) ;
  assign n23934 = n23933 ^ n23932 ^ n7171 ;
  assign n23935 = n23934 ^ n8125 ^ n5240 ;
  assign n23936 = ( n14011 & ~n23930 ) | ( n14011 & n23935 ) | ( ~n23930 & n23935 ) ;
  assign n23937 = ( ~n1083 & n23805 ) | ( ~n1083 & n23936 ) | ( n23805 & n23936 ) ;
  assign n23938 = n23937 ^ n11499 ^ 1'b0 ;
  assign n23939 = n3905 & ~n23938 ;
  assign n23940 = n23939 ^ n14208 ^ n9611 ;
  assign n23941 = n23914 ^ n17055 ^ n15203 ;
  assign n23942 = n19473 ^ n7196 ^ n534 ;
  assign n23943 = n23942 ^ n4024 ^ n1758 ;
  assign n23949 = ( n1270 & n1494 ) | ( n1270 & n12149 ) | ( n1494 & n12149 ) ;
  assign n23948 = ( n6168 & ~n9242 ) | ( n6168 & n10397 ) | ( ~n9242 & n10397 ) ;
  assign n23946 = n7317 ^ n1750 ^ 1'b0 ;
  assign n23944 = n15928 ^ n13607 ^ 1'b0 ;
  assign n23945 = ( n8798 & n12326 ) | ( n8798 & n23944 ) | ( n12326 & n23944 ) ;
  assign n23947 = n23946 ^ n23945 ^ n13151 ;
  assign n23950 = n23949 ^ n23948 ^ n23947 ;
  assign n23953 = n16804 ^ n15848 ^ n2402 ;
  assign n23954 = n8286 & ~n23953 ;
  assign n23955 = ( n2013 & ~n21574 ) | ( n2013 & n23954 ) | ( ~n21574 & n23954 ) ;
  assign n23951 = n11272 ^ n3025 ^ n596 ;
  assign n23952 = n23951 ^ n8164 ^ n2976 ;
  assign n23956 = n23955 ^ n23952 ^ n1643 ;
  assign n23957 = ( n2892 & n9863 ) | ( n2892 & n16824 ) | ( n9863 & n16824 ) ;
  assign n23958 = n14224 ^ n6688 ^ n4244 ;
  assign n23959 = n20747 & n23958 ;
  assign n23960 = ~n3832 & n23959 ;
  assign n23961 = ( n3601 & n6807 ) | ( n3601 & ~n12304 ) | ( n6807 & ~n12304 ) ;
  assign n23962 = n781 | n21634 ;
  assign n23963 = n1013 & ~n23962 ;
  assign n23964 = n23963 ^ n19289 ^ n14664 ;
  assign n23965 = n1261 & ~n9512 ;
  assign n23966 = ~n3052 & n23965 ;
  assign n23967 = ( ~n13902 & n22259 ) | ( ~n13902 & n23966 ) | ( n22259 & n23966 ) ;
  assign n23968 = ( ~n23961 & n23964 ) | ( ~n23961 & n23967 ) | ( n23964 & n23967 ) ;
  assign n23969 = n7715 & ~n22625 ;
  assign n23970 = n23969 ^ n5822 ^ n2902 ;
  assign n23973 = n8407 ^ n1026 ^ 1'b0 ;
  assign n23972 = ( n7417 & ~n7802 ) | ( n7417 & n10130 ) | ( ~n7802 & n10130 ) ;
  assign n23971 = ( n1114 & n9553 ) | ( n1114 & ~n20330 ) | ( n9553 & ~n20330 ) ;
  assign n23974 = n23973 ^ n23972 ^ n23971 ;
  assign n23975 = n12521 ^ n8033 ^ n4772 ;
  assign n23976 = ( n2899 & n20732 ) | ( n2899 & n23975 ) | ( n20732 & n23975 ) ;
  assign n23977 = n10500 ^ n8124 ^ n2035 ;
  assign n23978 = n23977 ^ n23245 ^ n19690 ;
  assign n23979 = n18447 ^ n5065 ^ n4096 ;
  assign n23980 = n23979 ^ n21364 ^ 1'b0 ;
  assign n23981 = n23980 ^ n19731 ^ n12044 ;
  assign n23982 = n23981 ^ n19710 ^ n15468 ;
  assign n23983 = ~n1809 & n7371 ;
  assign n23984 = ( ~n1592 & n6134 ) | ( ~n1592 & n23983 ) | ( n6134 & n23983 ) ;
  assign n23985 = ~n14878 & n23984 ;
  assign n23986 = n23985 ^ n5009 ^ 1'b0 ;
  assign n23987 = ( n7358 & n8528 ) | ( n7358 & n8624 ) | ( n8528 & n8624 ) ;
  assign n23988 = n23987 ^ n16582 ^ n3907 ;
  assign n23989 = ( n881 & n7763 ) | ( n881 & ~n14419 ) | ( n7763 & ~n14419 ) ;
  assign n23993 = ( ~n1209 & n2378 ) | ( ~n1209 & n6304 ) | ( n2378 & n6304 ) ;
  assign n23990 = n16515 ^ n15587 ^ x0 ;
  assign n23991 = n23990 ^ n5684 ^ 1'b0 ;
  assign n23992 = n5780 & ~n23991 ;
  assign n23994 = n23993 ^ n23992 ^ n16429 ;
  assign n23995 = ( ~n6956 & n23989 ) | ( ~n6956 & n23994 ) | ( n23989 & n23994 ) ;
  assign n24000 = ( n5106 & ~n5120 ) | ( n5106 & n15726 ) | ( ~n5120 & n15726 ) ;
  assign n24001 = n751 & ~n24000 ;
  assign n24002 = n24001 ^ n3999 ^ 1'b0 ;
  assign n23996 = n23973 ^ n20804 ^ n7640 ;
  assign n23997 = n20313 & ~n23996 ;
  assign n23998 = n3232 & n23997 ;
  assign n23999 = ( n2328 & n13684 ) | ( n2328 & ~n23998 ) | ( n13684 & ~n23998 ) ;
  assign n24003 = n24002 ^ n23999 ^ n22907 ;
  assign n24004 = ( ~n7910 & n16091 ) | ( ~n7910 & n23539 ) | ( n16091 & n23539 ) ;
  assign n24005 = n1687 ^ x3 ^ 1'b0 ;
  assign n24006 = ( ~n3922 & n20795 ) | ( ~n3922 & n24005 ) | ( n20795 & n24005 ) ;
  assign n24008 = n12171 ^ n5833 ^ 1'b0 ;
  assign n24007 = n8052 ^ n6437 ^ n879 ;
  assign n24009 = n24008 ^ n24007 ^ n2850 ;
  assign n24010 = n22859 ^ n2874 ^ 1'b0 ;
  assign n24011 = ( n2222 & ~n3757 ) | ( n2222 & n16681 ) | ( ~n3757 & n16681 ) ;
  assign n24012 = n24011 ^ n23228 ^ n19322 ;
  assign n24013 = n19956 ^ n18483 ^ n13616 ;
  assign n24014 = n24013 ^ n13499 ^ n11814 ;
  assign n24015 = n18299 | n24014 ;
  assign n24016 = n9888 ^ n2735 ^ n1203 ;
  assign n24017 = ( ~n933 & n1480 ) | ( ~n933 & n4866 ) | ( n1480 & n4866 ) ;
  assign n24018 = ( n7168 & n8530 ) | ( n7168 & ~n24017 ) | ( n8530 & ~n24017 ) ;
  assign n24019 = n13733 ^ n12658 ^ n2245 ;
  assign n24020 = ( n391 & ~n9317 ) | ( n391 & n24019 ) | ( ~n9317 & n24019 ) ;
  assign n24021 = n3565 & ~n16275 ;
  assign n24022 = n24021 ^ n3715 ^ 1'b0 ;
  assign n24023 = n12530 | n24022 ;
  assign n24024 = n10047 ^ n3992 ^ n3243 ;
  assign n24025 = n17706 ^ n4951 ^ 1'b0 ;
  assign n24026 = n18011 & n24025 ;
  assign n24027 = n24026 ^ n17379 ^ 1'b0 ;
  assign n24028 = ( n6872 & n18511 ) | ( n6872 & n22575 ) | ( n18511 & n22575 ) ;
  assign n24029 = n15618 ^ n3580 ^ 1'b0 ;
  assign n24030 = n14793 & ~n24029 ;
  assign n24031 = n24030 ^ n23572 ^ n8230 ;
  assign n24032 = ( n5522 & n14301 ) | ( n5522 & ~n24031 ) | ( n14301 & ~n24031 ) ;
  assign n24033 = n20276 ^ n20084 ^ n11566 ;
  assign n24034 = ( ~n2977 & n5765 ) | ( ~n2977 & n14713 ) | ( n5765 & n14713 ) ;
  assign n24035 = n24034 ^ n23475 ^ n988 ;
  assign n24036 = n24035 ^ n9164 ^ n6602 ;
  assign n24041 = n11267 ^ n5898 ^ n2257 ;
  assign n24037 = ( n11570 & n13760 ) | ( n11570 & n14075 ) | ( n13760 & n14075 ) ;
  assign n24038 = n24037 ^ n11071 ^ n5042 ;
  assign n24039 = ( ~n2665 & n7652 ) | ( ~n2665 & n24038 ) | ( n7652 & n24038 ) ;
  assign n24040 = n24039 ^ n11523 ^ n10050 ;
  assign n24042 = n24041 ^ n24040 ^ 1'b0 ;
  assign n24043 = n10375 | n24042 ;
  assign n24044 = ( ~n8361 & n24036 ) | ( ~n8361 & n24043 ) | ( n24036 & n24043 ) ;
  assign n24045 = n14185 ^ n5054 ^ 1'b0 ;
  assign n24046 = ( n4222 & n14689 ) | ( n4222 & ~n24045 ) | ( n14689 & ~n24045 ) ;
  assign n24047 = ( n10130 & n14505 ) | ( n10130 & ~n15892 ) | ( n14505 & ~n15892 ) ;
  assign n24048 = ( n2869 & n3136 ) | ( n2869 & ~n8251 ) | ( n3136 & ~n8251 ) ;
  assign n24049 = n6061 ^ n1634 ^ 1'b0 ;
  assign n24050 = n1960 & n24049 ;
  assign n24051 = n24050 ^ n22756 ^ n12950 ;
  assign n24052 = ( ~n4836 & n7140 ) | ( ~n4836 & n19502 ) | ( n7140 & n19502 ) ;
  assign n24053 = ( ~n2466 & n9830 ) | ( ~n2466 & n24052 ) | ( n9830 & n24052 ) ;
  assign n24056 = n464 & ~n8478 ;
  assign n24054 = ( n2188 & n3242 ) | ( n2188 & ~n3673 ) | ( n3242 & ~n3673 ) ;
  assign n24055 = ( n7402 & n13606 ) | ( n7402 & ~n24054 ) | ( n13606 & ~n24054 ) ;
  assign n24057 = n24056 ^ n24055 ^ 1'b0 ;
  assign n24060 = n23259 ^ n19565 ^ 1'b0 ;
  assign n24058 = n23914 ^ n8446 ^ n1098 ;
  assign n24059 = ( ~n9621 & n20881 ) | ( ~n9621 & n24058 ) | ( n20881 & n24058 ) ;
  assign n24061 = n24060 ^ n24059 ^ n3888 ;
  assign n24062 = ( n10091 & ~n18401 ) | ( n10091 & n23434 ) | ( ~n18401 & n23434 ) ;
  assign n24063 = n24062 ^ n18512 ^ n18274 ;
  assign n24064 = ( ~n18092 & n24061 ) | ( ~n18092 & n24063 ) | ( n24061 & n24063 ) ;
  assign n24065 = n23016 ^ n2541 ^ 1'b0 ;
  assign n24066 = n17824 & n24065 ;
  assign n24067 = ( ~n8588 & n15820 ) | ( ~n8588 & n19237 ) | ( n15820 & n19237 ) ;
  assign n24070 = n7979 ^ n2483 ^ n1291 ;
  assign n24071 = ( x75 & ~n7228 ) | ( x75 & n24070 ) | ( ~n7228 & n24070 ) ;
  assign n24068 = ( n6328 & n10143 ) | ( n6328 & ~n17587 ) | ( n10143 & ~n17587 ) ;
  assign n24069 = ( n2224 & n17847 ) | ( n2224 & ~n24068 ) | ( n17847 & ~n24068 ) ;
  assign n24072 = n24071 ^ n24069 ^ 1'b0 ;
  assign n24073 = ~n2686 & n24072 ;
  assign n24074 = n9829 ^ n6991 ^ 1'b0 ;
  assign n24075 = n22750 ^ n1787 ^ n1772 ;
  assign n24076 = ( n7391 & n14488 ) | ( n7391 & n23887 ) | ( n14488 & n23887 ) ;
  assign n24077 = n23339 ^ n13887 ^ 1'b0 ;
  assign n24078 = ( n3715 & n9938 ) | ( n3715 & n14201 ) | ( n9938 & n14201 ) ;
  assign n24079 = n9372 ^ n5722 ^ n329 ;
  assign n24080 = ( ~n2598 & n20920 ) | ( ~n2598 & n23887 ) | ( n20920 & n23887 ) ;
  assign n24081 = n24080 ^ n22555 ^ n3559 ;
  assign n24082 = n10992 & n19344 ;
  assign n24083 = ( n8559 & ~n12290 ) | ( n8559 & n18193 ) | ( ~n12290 & n18193 ) ;
  assign n24084 = ( n6411 & n10873 ) | ( n6411 & ~n19117 ) | ( n10873 & ~n19117 ) ;
  assign n24085 = ( n8613 & n9379 ) | ( n8613 & n24084 ) | ( n9379 & n24084 ) ;
  assign n24086 = n24085 ^ n22664 ^ n12437 ;
  assign n24087 = ( n368 & ~n6708 ) | ( n368 & n24086 ) | ( ~n6708 & n24086 ) ;
  assign n24088 = ( n5875 & n10360 ) | ( n5875 & n11447 ) | ( n10360 & n11447 ) ;
  assign n24089 = ( ~n1020 & n8875 ) | ( ~n1020 & n24088 ) | ( n8875 & n24088 ) ;
  assign n24090 = n6093 ^ n3230 ^ n1056 ;
  assign n24091 = ( x115 & n1213 ) | ( x115 & ~n1345 ) | ( n1213 & ~n1345 ) ;
  assign n24092 = n24091 ^ n13996 ^ n3290 ;
  assign n24093 = ( n11608 & ~n24090 ) | ( n11608 & n24092 ) | ( ~n24090 & n24092 ) ;
  assign n24094 = n11132 ^ n8721 ^ n7273 ;
  assign n24095 = n19177 ^ n15834 ^ n9482 ;
  assign n24096 = n13667 & n24095 ;
  assign n24097 = n24096 ^ n19139 ^ 1'b0 ;
  assign n24098 = ( n4440 & n13904 ) | ( n4440 & ~n20744 ) | ( n13904 & ~n20744 ) ;
  assign n24100 = ( x82 & n13028 ) | ( x82 & ~n15042 ) | ( n13028 & ~n15042 ) ;
  assign n24101 = ( n13086 & n14588 ) | ( n13086 & n24100 ) | ( n14588 & n24100 ) ;
  assign n24099 = n17380 ^ n14309 ^ 1'b0 ;
  assign n24102 = n24101 ^ n24099 ^ n4325 ;
  assign n24103 = ( n5172 & n7087 ) | ( n5172 & n8653 ) | ( n7087 & n8653 ) ;
  assign n24104 = n21914 | n24103 ;
  assign n24105 = n23012 ^ n7152 ^ n429 ;
  assign n24106 = n7626 ^ n7047 ^ n4311 ;
  assign n24107 = n24106 ^ n5161 ^ n1063 ;
  assign n24108 = n17178 ^ n16817 ^ n15746 ;
  assign n24109 = ( ~n9634 & n18379 ) | ( ~n9634 & n24108 ) | ( n18379 & n24108 ) ;
  assign n24110 = ~n18448 & n24109 ;
  assign n24111 = n6517 | n24110 ;
  assign n24112 = ~n2928 & n18091 ;
  assign n24114 = n8138 ^ n2339 ^ n807 ;
  assign n24113 = ( n320 & ~n432 ) | ( n320 & n18204 ) | ( ~n432 & n18204 ) ;
  assign n24115 = n24114 ^ n24113 ^ n9430 ;
  assign n24117 = n5800 & ~n9853 ;
  assign n24118 = ~n761 & n24117 ;
  assign n24119 = ( n6096 & n12658 ) | ( n6096 & ~n24118 ) | ( n12658 & ~n24118 ) ;
  assign n24116 = ( n745 & n11029 ) | ( n745 & ~n16237 ) | ( n11029 & ~n16237 ) ;
  assign n24120 = n24119 ^ n24116 ^ n2399 ;
  assign n24121 = n21440 ^ n18706 ^ n17208 ;
  assign n24122 = n9089 & n17867 ;
  assign n24123 = n24122 ^ n3230 ^ n1577 ;
  assign n24124 = n24123 ^ n14642 ^ n4285 ;
  assign n24125 = n16455 ^ n10183 ^ n2885 ;
  assign n24126 = ( ~n12534 & n19794 ) | ( ~n12534 & n24125 ) | ( n19794 & n24125 ) ;
  assign n24127 = ( n380 & ~n2779 ) | ( n380 & n16931 ) | ( ~n2779 & n16931 ) ;
  assign n24128 = ( n16081 & n20233 ) | ( n16081 & n24127 ) | ( n20233 & n24127 ) ;
  assign n24131 = ( n352 & n3571 ) | ( n352 & n9556 ) | ( n3571 & n9556 ) ;
  assign n24130 = ( n7924 & n8274 ) | ( n7924 & ~n11466 ) | ( n8274 & ~n11466 ) ;
  assign n24132 = n24131 ^ n24130 ^ n21420 ;
  assign n24129 = n2642 & ~n20095 ;
  assign n24133 = n24132 ^ n24129 ^ n10162 ;
  assign n24134 = ~n24128 & n24133 ;
  assign n24135 = n24134 ^ n12058 ^ 1'b0 ;
  assign n24136 = n17844 ^ n2109 ^ 1'b0 ;
  assign n24137 = n22815 & ~n24136 ;
  assign n24138 = ( n2121 & ~n7240 ) | ( n2121 & n16318 ) | ( ~n7240 & n16318 ) ;
  assign n24139 = ( n2730 & ~n14976 ) | ( n2730 & n21908 ) | ( ~n14976 & n21908 ) ;
  assign n24140 = n24139 ^ n18221 ^ n17234 ;
  assign n24141 = ( n482 & ~n8172 ) | ( n482 & n22239 ) | ( ~n8172 & n22239 ) ;
  assign n24142 = ( ~n9073 & n12443 ) | ( ~n9073 & n24141 ) | ( n12443 & n24141 ) ;
  assign n24143 = n9671 ^ n3541 ^ n3073 ;
  assign n24146 = ( ~n691 & n2276 ) | ( ~n691 & n15812 ) | ( n2276 & n15812 ) ;
  assign n24144 = ( n960 & ~n3371 ) | ( n960 & n6093 ) | ( ~n3371 & n6093 ) ;
  assign n24145 = n11809 | n24144 ;
  assign n24147 = n24146 ^ n24145 ^ 1'b0 ;
  assign n24148 = ( n3042 & ~n6274 ) | ( n3042 & n7390 ) | ( ~n6274 & n7390 ) ;
  assign n24149 = n24148 ^ n19445 ^ n13193 ;
  assign n24150 = ~n2504 & n22932 ;
  assign n24151 = ~n15951 & n24150 ;
  assign n24152 = ( ~n1874 & n3773 ) | ( ~n1874 & n5157 ) | ( n3773 & n5157 ) ;
  assign n24153 = ( n15024 & n18500 ) | ( n15024 & ~n24152 ) | ( n18500 & ~n24152 ) ;
  assign n24154 = ( x19 & ~n809 ) | ( x19 & n8731 ) | ( ~n809 & n8731 ) ;
  assign n24155 = ( n186 & n24153 ) | ( n186 & ~n24154 ) | ( n24153 & ~n24154 ) ;
  assign n24156 = n7552 & ~n24155 ;
  assign n24157 = n24156 ^ n16990 ^ 1'b0 ;
  assign n24158 = ( n2477 & n7214 ) | ( n2477 & ~n11998 ) | ( n7214 & ~n11998 ) ;
  assign n24159 = ( x122 & n1057 ) | ( x122 & n24158 ) | ( n1057 & n24158 ) ;
  assign n24160 = ( n203 & n4096 ) | ( n203 & ~n24159 ) | ( n4096 & ~n24159 ) ;
  assign n24161 = ( ~n11494 & n16235 ) | ( ~n11494 & n19111 ) | ( n16235 & n19111 ) ;
  assign n24162 = n24161 ^ n15300 ^ n3742 ;
  assign n24163 = n6313 ^ n4414 ^ n3107 ;
  assign n24164 = ( n2476 & n6956 ) | ( n2476 & n24163 ) | ( n6956 & n24163 ) ;
  assign n24165 = n24164 ^ n7615 ^ n249 ;
  assign n24166 = n20217 ^ n17242 ^ n6299 ;
  assign n24167 = n24166 ^ n12235 ^ n8595 ;
  assign n24168 = ( n1610 & n5781 ) | ( n1610 & n23610 ) | ( n5781 & n23610 ) ;
  assign n24169 = n24168 ^ n13598 ^ 1'b0 ;
  assign n24170 = n24169 ^ n13668 ^ n9391 ;
  assign n24171 = ( n19712 & n20573 ) | ( n19712 & ~n24170 ) | ( n20573 & ~n24170 ) ;
  assign n24172 = ( x18 & ~n7072 ) | ( x18 & n24171 ) | ( ~n7072 & n24171 ) ;
  assign n24173 = n6752 ^ n6280 ^ n2073 ;
  assign n24174 = n24173 ^ n5930 ^ n1951 ;
  assign n24175 = ( n1322 & n5125 ) | ( n1322 & ~n8378 ) | ( n5125 & ~n8378 ) ;
  assign n24176 = ( n4461 & n16426 ) | ( n4461 & n18268 ) | ( n16426 & n18268 ) ;
  assign n24178 = ( n5395 & n5599 ) | ( n5395 & n9688 ) | ( n5599 & n9688 ) ;
  assign n24179 = n24178 ^ n23415 ^ n6029 ;
  assign n24177 = ~n5621 & n9152 ;
  assign n24180 = n24179 ^ n24177 ^ 1'b0 ;
  assign n24181 = n2403 & ~n21864 ;
  assign n24182 = n24181 ^ n3956 ^ 1'b0 ;
  assign n24186 = n8294 ^ n1898 ^ n648 ;
  assign n24187 = n24186 ^ n8932 ^ n8546 ;
  assign n24183 = ( ~n5831 & n7180 ) | ( ~n5831 & n13164 ) | ( n7180 & n13164 ) ;
  assign n24184 = ( ~n6223 & n15930 ) | ( ~n6223 & n24183 ) | ( n15930 & n24183 ) ;
  assign n24185 = ~n5351 & n24184 ;
  assign n24188 = n24187 ^ n24185 ^ n17416 ;
  assign n24189 = ( n8029 & ~n24182 ) | ( n8029 & n24188 ) | ( ~n24182 & n24188 ) ;
  assign n24190 = n22704 ^ n16094 ^ 1'b0 ;
  assign n24191 = n8990 & n24190 ;
  assign n24192 = n24191 ^ n7927 ^ n4122 ;
  assign n24199 = n13222 ^ n2077 ^ n676 ;
  assign n24197 = n23555 ^ n11522 ^ n4348 ;
  assign n24198 = ( n7976 & n23846 ) | ( n7976 & ~n24197 ) | ( n23846 & ~n24197 ) ;
  assign n24193 = n8445 ^ n5682 ^ n3380 ;
  assign n24194 = n24193 ^ n14632 ^ n384 ;
  assign n24195 = ( ~n1093 & n2335 ) | ( ~n1093 & n24194 ) | ( n2335 & n24194 ) ;
  assign n24196 = ~n1204 & n24195 ;
  assign n24200 = n24199 ^ n24198 ^ n24196 ;
  assign n24201 = n19271 ^ n14749 ^ n5931 ;
  assign n24202 = ( n6614 & ~n21351 ) | ( n6614 & n24201 ) | ( ~n21351 & n24201 ) ;
  assign n24203 = n18565 ^ n7987 ^ n6481 ;
  assign n24204 = n24203 ^ n18151 ^ n14204 ;
  assign n24205 = ~n6016 & n18180 ;
  assign n24206 = n1958 & n4005 ;
  assign n24207 = n21988 ^ n9381 ^ 1'b0 ;
  assign n24208 = ( n16092 & n24206 ) | ( n16092 & ~n24207 ) | ( n24206 & ~n24207 ) ;
  assign n24212 = ( n14739 & n20825 ) | ( n14739 & n22982 ) | ( n20825 & n22982 ) ;
  assign n24209 = n2724 | n6099 ;
  assign n24210 = n6330 & n24209 ;
  assign n24211 = ( ~n18689 & n19212 ) | ( ~n18689 & n24210 ) | ( n19212 & n24210 ) ;
  assign n24213 = n24212 ^ n24211 ^ n7556 ;
  assign n24215 = ( n885 & n4769 ) | ( n885 & n12814 ) | ( n4769 & n12814 ) ;
  assign n24214 = n13198 & ~n22064 ;
  assign n24216 = n24215 ^ n24214 ^ 1'b0 ;
  assign n24217 = n16610 ^ n8315 ^ n3371 ;
  assign n24218 = ( n1629 & ~n24216 ) | ( n1629 & n24217 ) | ( ~n24216 & n24217 ) ;
  assign n24219 = n24218 ^ n14629 ^ n2541 ;
  assign n24220 = ( n2399 & n14467 ) | ( n2399 & ~n24219 ) | ( n14467 & ~n24219 ) ;
  assign n24221 = n15919 ^ n4170 ^ n1311 ;
  assign n24222 = n24221 ^ n9837 ^ n7346 ;
  assign n24223 = ( n4514 & n22547 ) | ( n4514 & n24222 ) | ( n22547 & n24222 ) ;
  assign n24224 = n21950 ^ n9507 ^ 1'b0 ;
  assign n24225 = n4203 | n24224 ;
  assign n24226 = n24225 ^ n15799 ^ 1'b0 ;
  assign n24227 = n17658 ^ n9360 ^ 1'b0 ;
  assign n24228 = ( n2820 & ~n9036 ) | ( n2820 & n24227 ) | ( ~n9036 & n24227 ) ;
  assign n24229 = n24228 ^ n2449 ^ n1661 ;
  assign n24230 = n9600 & n11548 ;
  assign n24231 = n24230 ^ n11764 ^ 1'b0 ;
  assign n24232 = n24231 ^ n13256 ^ n12460 ;
  assign n24233 = ( n2934 & ~n10386 ) | ( n2934 & n13139 ) | ( ~n10386 & n13139 ) ;
  assign n24234 = n14088 ^ n6219 ^ n4867 ;
  assign n24235 = ( n233 & ~n7839 ) | ( n233 & n24234 ) | ( ~n7839 & n24234 ) ;
  assign n24236 = n24233 | n24235 ;
  assign n24237 = n1668 | n24236 ;
  assign n24238 = n17869 ^ n6457 ^ n5865 ;
  assign n24239 = ( ~n13840 & n22394 ) | ( ~n13840 & n24238 ) | ( n22394 & n24238 ) ;
  assign n24240 = n8072 | n9533 ;
  assign n24241 = n24240 ^ n6775 ^ 1'b0 ;
  assign n24242 = ( n5144 & n24239 ) | ( n5144 & n24241 ) | ( n24239 & n24241 ) ;
  assign n24243 = n23437 ^ n8567 ^ n3103 ;
  assign n24244 = ( n3467 & n6029 ) | ( n3467 & n9479 ) | ( n6029 & n9479 ) ;
  assign n24247 = n11655 ^ n9722 ^ n8033 ;
  assign n24245 = n16620 ^ n14809 ^ n4060 ;
  assign n24246 = ( ~n775 & n2247 ) | ( ~n775 & n24245 ) | ( n2247 & n24245 ) ;
  assign n24248 = n24247 ^ n24246 ^ n22277 ;
  assign n24249 = n9682 ^ n3521 ^ n148 ;
  assign n24250 = n9613 ^ n9479 ^ n3153 ;
  assign n24251 = ~n7796 & n24250 ;
  assign n24252 = n24251 ^ n19158 ^ 1'b0 ;
  assign n24253 = ( ~n22799 & n24249 ) | ( ~n22799 & n24252 ) | ( n24249 & n24252 ) ;
  assign n24255 = n10230 ^ n7935 ^ n796 ;
  assign n24254 = n2438 | n8690 ;
  assign n24256 = n24255 ^ n24254 ^ n9431 ;
  assign n24257 = n18686 ^ n14006 ^ n3999 ;
  assign n24258 = ( n10065 & ~n18566 ) | ( n10065 & n24257 ) | ( ~n18566 & n24257 ) ;
  assign n24259 = n12319 ^ n6567 ^ 1'b0 ;
  assign n24260 = ( n8369 & n9827 ) | ( n8369 & ~n10904 ) | ( n9827 & ~n10904 ) ;
  assign n24262 = n13598 ^ n647 ^ 1'b0 ;
  assign n24261 = n9270 ^ n6206 ^ 1'b0 ;
  assign n24263 = n24262 ^ n24261 ^ n7765 ;
  assign n24264 = n3830 ^ n1227 ^ 1'b0 ;
  assign n24265 = ( n6748 & n8757 ) | ( n6748 & ~n20313 ) | ( n8757 & ~n20313 ) ;
  assign n24266 = n24265 ^ n11466 ^ n2288 ;
  assign n24267 = ( n1554 & n8530 ) | ( n1554 & ~n10265 ) | ( n8530 & ~n10265 ) ;
  assign n24268 = ( n4540 & n4967 ) | ( n4540 & ~n24267 ) | ( n4967 & ~n24267 ) ;
  assign n24269 = n19728 ^ n16745 ^ n15584 ;
  assign n24270 = n19228 ^ n13096 ^ n8706 ;
  assign n24271 = ( n9947 & n17336 ) | ( n9947 & ~n24270 ) | ( n17336 & ~n24270 ) ;
  assign n24272 = ( n7763 & n14290 ) | ( n7763 & n14379 ) | ( n14290 & n14379 ) ;
  assign n24273 = ( n9767 & n19632 ) | ( n9767 & n24272 ) | ( n19632 & n24272 ) ;
  assign n24274 = n24273 ^ n11718 ^ 1'b0 ;
  assign n24275 = n21585 & ~n24274 ;
  assign n24278 = n17583 ^ n10688 ^ n9712 ;
  assign n24276 = n17175 ^ n5291 ^ n3351 ;
  assign n24277 = ( n2869 & n7543 ) | ( n2869 & ~n24276 ) | ( n7543 & ~n24276 ) ;
  assign n24279 = n24278 ^ n24277 ^ n21482 ;
  assign n24280 = n22270 ^ n22096 ^ n16658 ;
  assign n24281 = n20475 ^ n19217 ^ n18149 ;
  assign n24283 = ( n5423 & n5441 ) | ( n5423 & n11166 ) | ( n5441 & n11166 ) ;
  assign n24282 = ( n3497 & n5014 ) | ( n3497 & ~n12772 ) | ( n5014 & ~n12772 ) ;
  assign n24284 = n24283 ^ n24282 ^ n13480 ;
  assign n24285 = ( n3441 & ~n5900 ) | ( n3441 & n6328 ) | ( ~n5900 & n6328 ) ;
  assign n24286 = n24285 ^ n9745 ^ n6214 ;
  assign n24287 = n17377 ^ n3737 ^ 1'b0 ;
  assign n24288 = n19321 | n24287 ;
  assign n24289 = ( n3874 & n6121 ) | ( n3874 & ~n6748 ) | ( n6121 & ~n6748 ) ;
  assign n24290 = n24289 ^ n6493 ^ n367 ;
  assign n24291 = ( n7311 & n14757 ) | ( n7311 & n24290 ) | ( n14757 & n24290 ) ;
  assign n24292 = n24291 ^ n9201 ^ 1'b0 ;
  assign n24293 = ( n510 & n592 ) | ( n510 & n718 ) | ( n592 & n718 ) ;
  assign n24294 = ( n7761 & n21231 ) | ( n7761 & n24293 ) | ( n21231 & n24293 ) ;
  assign n24295 = n13566 ^ n3354 ^ 1'b0 ;
  assign n24296 = n21011 ^ n13760 ^ n4959 ;
  assign n24297 = n18056 ^ n10076 ^ n2861 ;
  assign n24298 = ( ~n3953 & n8814 ) | ( ~n3953 & n11424 ) | ( n8814 & n11424 ) ;
  assign n24299 = n10452 & ~n24298 ;
  assign n24300 = n10295 ^ n2932 ^ n666 ;
  assign n24301 = n24300 ^ n14908 ^ n3225 ;
  assign n24302 = n3317 & n24301 ;
  assign n24303 = ( n2581 & n12515 ) | ( n2581 & n24302 ) | ( n12515 & n24302 ) ;
  assign n24304 = ( n24297 & n24299 ) | ( n24297 & ~n24303 ) | ( n24299 & ~n24303 ) ;
  assign n24305 = ( n10132 & n24296 ) | ( n10132 & ~n24304 ) | ( n24296 & ~n24304 ) ;
  assign n24306 = ( ~n10780 & n10820 ) | ( ~n10780 & n15670 ) | ( n10820 & n15670 ) ;
  assign n24307 = ( n4883 & ~n6787 ) | ( n4883 & n24306 ) | ( ~n6787 & n24306 ) ;
  assign n24308 = n15297 ^ n3727 ^ n2088 ;
  assign n24309 = ~n2701 & n24308 ;
  assign n24310 = n24309 ^ n7871 ^ 1'b0 ;
  assign n24311 = ~n5423 & n17676 ;
  assign n24313 = n8496 | n10779 ;
  assign n24314 = ~n481 & n24313 ;
  assign n24315 = ~n7502 & n24314 ;
  assign n24312 = ~n6792 & n23466 ;
  assign n24316 = n24315 ^ n24312 ^ n21760 ;
  assign n24317 = ( n696 & n6075 ) | ( n696 & n16577 ) | ( n6075 & n16577 ) ;
  assign n24318 = n24317 ^ n3549 ^ n1417 ;
  assign n24319 = n23108 ^ n14609 ^ n12548 ;
  assign n24320 = n13794 ^ n9004 ^ n595 ;
  assign n24321 = n23533 ^ n19762 ^ n6079 ;
  assign n24322 = ( n1612 & n17698 ) | ( n1612 & ~n21479 ) | ( n17698 & ~n21479 ) ;
  assign n24330 = ~n516 & n6563 ;
  assign n24324 = ( n2031 & n3057 ) | ( n2031 & n7625 ) | ( n3057 & n7625 ) ;
  assign n24323 = n11124 & n19721 ;
  assign n24325 = n24324 ^ n24323 ^ 1'b0 ;
  assign n24326 = ~n11553 & n24325 ;
  assign n24327 = n24326 ^ n18017 ^ 1'b0 ;
  assign n24328 = n24327 ^ n17796 ^ n7164 ;
  assign n24329 = n24328 ^ n16587 ^ n13447 ;
  assign n24331 = n24330 ^ n24329 ^ n17606 ;
  assign n24332 = n15160 ^ n6095 ^ n3036 ;
  assign n24333 = ( n13697 & n23185 ) | ( n13697 & n23944 ) | ( n23185 & n23944 ) ;
  assign n24334 = ~n24332 & n24333 ;
  assign n24335 = n24334 ^ n24037 ^ 1'b0 ;
  assign n24337 = n10855 ^ n5417 ^ n3289 ;
  assign n24336 = ( n2617 & ~n3630 ) | ( n2617 & n9418 ) | ( ~n3630 & n9418 ) ;
  assign n24338 = n24337 ^ n24336 ^ n14863 ;
  assign n24339 = n23331 ^ n8530 ^ n4684 ;
  assign n24340 = ( n1659 & n14309 ) | ( n1659 & n24339 ) | ( n14309 & n24339 ) ;
  assign n24341 = ( ~n5281 & n19727 ) | ( ~n5281 & n22658 ) | ( n19727 & n22658 ) ;
  assign n24342 = n24341 ^ n19876 ^ n19211 ;
  assign n24343 = n24342 ^ n2550 ^ n714 ;
  assign n24344 = ( n7206 & n7307 ) | ( n7206 & n10124 ) | ( n7307 & n10124 ) ;
  assign n24345 = n24344 ^ n23989 ^ n5121 ;
  assign n24346 = ( n18225 & ~n19896 ) | ( n18225 & n24345 ) | ( ~n19896 & n24345 ) ;
  assign n24349 = ( n1027 & n5630 ) | ( n1027 & n9938 ) | ( n5630 & n9938 ) ;
  assign n24348 = n6733 ^ n2303 ^ 1'b0 ;
  assign n24347 = n23452 ^ n19390 ^ 1'b0 ;
  assign n24350 = n24349 ^ n24348 ^ n24347 ;
  assign n24351 = n18431 ^ n12121 ^ n8046 ;
  assign n24352 = n23787 ^ n11592 ^ n2052 ;
  assign n24353 = ( n5693 & n16656 ) | ( n5693 & ~n24352 ) | ( n16656 & ~n24352 ) ;
  assign n24354 = ~n15156 & n24353 ;
  assign n24355 = n4413 & n24354 ;
  assign n24356 = n20960 ^ n15483 ^ 1'b0 ;
  assign n24357 = n11671 & ~n24356 ;
  assign n24359 = n16283 ^ n14530 ^ n9885 ;
  assign n24358 = ( ~n2507 & n10674 ) | ( ~n2507 & n23047 ) | ( n10674 & n23047 ) ;
  assign n24360 = n24359 ^ n24358 ^ n506 ;
  assign n24361 = n24360 ^ n13267 ^ n4142 ;
  assign n24362 = n18368 ^ n6172 ^ 1'b0 ;
  assign n24363 = n24362 ^ n15002 ^ n13345 ;
  assign n24364 = n12531 ^ n6040 ^ 1'b0 ;
  assign n24365 = n20045 ^ n7696 ^ n3808 ;
  assign n24366 = ( n14480 & ~n16296 ) | ( n14480 & n16755 ) | ( ~n16296 & n16755 ) ;
  assign n24367 = n24366 ^ n12053 ^ n4929 ;
  assign n24368 = n24367 ^ n7189 ^ 1'b0 ;
  assign n24369 = ( ~n22258 & n24365 ) | ( ~n22258 & n24368 ) | ( n24365 & n24368 ) ;
  assign n24370 = n24369 ^ n10249 ^ n7951 ;
  assign n24371 = n12426 ^ n11679 ^ n10298 ;
  assign n24372 = ( n6497 & n19980 ) | ( n6497 & n21157 ) | ( n19980 & n21157 ) ;
  assign n24373 = ( n18247 & ~n24371 ) | ( n18247 & n24372 ) | ( ~n24371 & n24372 ) ;
  assign n24374 = n6764 ^ n1195 ^ 1'b0 ;
  assign n24375 = n7179 & n24374 ;
  assign n24376 = n24375 ^ n5020 ^ 1'b0 ;
  assign n24377 = ~n4222 & n5090 ;
  assign n24378 = n21864 & n24377 ;
  assign n24379 = n8155 ^ n8033 ^ n3241 ;
  assign n24380 = n10525 | n24379 ;
  assign n24381 = n24378 & ~n24380 ;
  assign n24382 = ( n7670 & ~n9475 ) | ( n7670 & n13958 ) | ( ~n9475 & n13958 ) ;
  assign n24383 = n5304 ^ n2451 ^ n1452 ;
  assign n24384 = ( n5277 & ~n24382 ) | ( n5277 & n24383 ) | ( ~n24382 & n24383 ) ;
  assign n24385 = n2485 | n20515 ;
  assign n24386 = n23331 ^ n2029 ^ n868 ;
  assign n24387 = ( n153 & n2343 ) | ( n153 & ~n24386 ) | ( n2343 & ~n24386 ) ;
  assign n24388 = ~n8883 & n24387 ;
  assign n24389 = ( n4356 & n12614 ) | ( n4356 & n13265 ) | ( n12614 & n13265 ) ;
  assign n24390 = n10598 | n23152 ;
  assign n24391 = ( n2757 & n3666 ) | ( n2757 & ~n24390 ) | ( n3666 & ~n24390 ) ;
  assign n24392 = ( n13643 & n20208 ) | ( n13643 & n24391 ) | ( n20208 & n24391 ) ;
  assign n24393 = n3609 | n16823 ;
  assign n24394 = n24392 & ~n24393 ;
  assign n24395 = ( ~n287 & n6571 ) | ( ~n287 & n17005 ) | ( n6571 & n17005 ) ;
  assign n24396 = n4166 & ~n13221 ;
  assign n24397 = n24395 & n24396 ;
  assign n24398 = n17154 ^ n11032 ^ n9951 ;
  assign n24399 = n5536 ^ n2291 ^ n978 ;
  assign n24400 = n24399 ^ n10099 ^ n2659 ;
  assign n24401 = ( n6955 & n20194 ) | ( n6955 & n24400 ) | ( n20194 & n24400 ) ;
  assign n24402 = n22014 ^ n17956 ^ n16851 ;
  assign n24403 = ( n14219 & n16864 ) | ( n14219 & ~n22143 ) | ( n16864 & ~n22143 ) ;
  assign n24404 = n21984 ^ n4287 ^ 1'b0 ;
  assign n24405 = n24404 ^ n19425 ^ n6812 ;
  assign n24406 = n22625 ^ n20755 ^ n16681 ;
  assign n24407 = ( n4175 & ~n10979 ) | ( n4175 & n15104 ) | ( ~n10979 & n15104 ) ;
  assign n24408 = ( ~n11585 & n16236 ) | ( ~n11585 & n21470 ) | ( n16236 & n21470 ) ;
  assign n24409 = ( n7508 & ~n18963 ) | ( n7508 & n24408 ) | ( ~n18963 & n24408 ) ;
  assign n24411 = n4582 ^ n1311 ^ 1'b0 ;
  assign n24412 = n4426 & n24411 ;
  assign n24410 = ( n7481 & n9424 ) | ( n7481 & n18589 ) | ( n9424 & n18589 ) ;
  assign n24413 = n24412 ^ n24410 ^ n18504 ;
  assign n24414 = n2459 ^ n2172 ^ 1'b0 ;
  assign n24415 = n24413 & ~n24414 ;
  assign n24416 = n20443 & ~n20455 ;
  assign n24417 = n24416 ^ n7411 ^ 1'b0 ;
  assign n24418 = n22366 ^ n12319 ^ n7605 ;
  assign n24419 = ( n540 & ~n5516 ) | ( n540 & n6125 ) | ( ~n5516 & n6125 ) ;
  assign n24420 = ( ~n1624 & n14739 ) | ( ~n1624 & n24419 ) | ( n14739 & n24419 ) ;
  assign n24421 = ~n1431 & n24420 ;
  assign n24422 = n17801 ^ n7297 ^ n2268 ;
  assign n24423 = ( n917 & n7777 ) | ( n917 & n18739 ) | ( n7777 & n18739 ) ;
  assign n24425 = ( n6672 & ~n10753 ) | ( n6672 & n18674 ) | ( ~n10753 & n18674 ) ;
  assign n24424 = n7562 & n24252 ;
  assign n24426 = n24425 ^ n24424 ^ 1'b0 ;
  assign n24427 = ( n15038 & ~n24423 ) | ( n15038 & n24426 ) | ( ~n24423 & n24426 ) ;
  assign n24428 = n12910 ^ n11605 ^ n2941 ;
  assign n24429 = n20930 ^ n20079 ^ n19498 ;
  assign n24430 = ( n9688 & ~n19800 ) | ( n9688 & n21218 ) | ( ~n19800 & n21218 ) ;
  assign n24431 = ( n1580 & ~n13329 ) | ( n1580 & n24430 ) | ( ~n13329 & n24430 ) ;
  assign n24432 = n24431 ^ n23291 ^ n2589 ;
  assign n24433 = ( n4370 & n6073 ) | ( n4370 & ~n8712 ) | ( n6073 & ~n8712 ) ;
  assign n24434 = n24433 ^ n17496 ^ n11149 ;
  assign n24435 = n4362 & n6563 ;
  assign n24436 = n1157 & n24435 ;
  assign n24437 = ~n7263 & n24436 ;
  assign n24438 = n17695 ^ n7090 ^ n3182 ;
  assign n24440 = ( n643 & n3196 ) | ( n643 & n10855 ) | ( n3196 & n10855 ) ;
  assign n24439 = n7874 ^ n235 ^ x75 ;
  assign n24441 = n24440 ^ n24439 ^ n6358 ;
  assign n24442 = n24441 ^ n18016 ^ 1'b0 ;
  assign n24443 = n3777 & n17527 ;
  assign n24444 = ( ~n5419 & n6020 ) | ( ~n5419 & n21218 ) | ( n6020 & n21218 ) ;
  assign n24445 = ( n3484 & n7375 ) | ( n3484 & n24444 ) | ( n7375 & n24444 ) ;
  assign n24446 = n24445 ^ n16212 ^ n484 ;
  assign n24447 = ~n2690 & n6427 ;
  assign n24448 = ~n15242 & n24447 ;
  assign n24449 = n20362 ^ n2928 ^ n2359 ;
  assign n24450 = ( ~n3033 & n10561 ) | ( ~n3033 & n17570 ) | ( n10561 & n17570 ) ;
  assign n24451 = ( ~n21284 & n24449 ) | ( ~n21284 & n24450 ) | ( n24449 & n24450 ) ;
  assign n24452 = n14473 ^ n13876 ^ n13697 ;
  assign n24459 = n2167 & n3758 ;
  assign n24460 = n22040 & n24459 ;
  assign n24458 = ( n1349 & n17706 ) | ( n1349 & ~n19410 ) | ( n17706 & ~n19410 ) ;
  assign n24457 = ( n1573 & n2757 ) | ( n1573 & n7255 ) | ( n2757 & n7255 ) ;
  assign n24461 = n24460 ^ n24458 ^ n24457 ;
  assign n24454 = ( n7113 & n7587 ) | ( n7113 & ~n9349 ) | ( n7587 & ~n9349 ) ;
  assign n24455 = n24454 ^ n6991 ^ n5343 ;
  assign n24453 = n9012 ^ n4197 ^ 1'b0 ;
  assign n24456 = n24455 ^ n24453 ^ n14042 ;
  assign n24462 = n24461 ^ n24456 ^ n24358 ;
  assign n24463 = n4152 & n8163 ;
  assign n24465 = n13130 ^ n5096 ^ n3591 ;
  assign n24464 = n3306 & n21918 ;
  assign n24466 = n24465 ^ n24464 ^ 1'b0 ;
  assign n24467 = ( n11381 & n16462 ) | ( n11381 & n24466 ) | ( n16462 & n24466 ) ;
  assign n24468 = ( ~n3598 & n12525 ) | ( ~n3598 & n19473 ) | ( n12525 & n19473 ) ;
  assign n24469 = n15636 ^ n9712 ^ n3303 ;
  assign n24470 = n22624 ^ n21716 ^ n1703 ;
  assign n24471 = ( n16174 & n24469 ) | ( n16174 & ~n24470 ) | ( n24469 & ~n24470 ) ;
  assign n24472 = n6289 & ~n9335 ;
  assign n24473 = n24472 ^ n19753 ^ 1'b0 ;
  assign n24474 = n24473 ^ n14861 ^ n7206 ;
  assign n24475 = ( ~n10636 & n12376 ) | ( ~n10636 & n16899 ) | ( n12376 & n16899 ) ;
  assign n24476 = ( n20231 & ~n24474 ) | ( n20231 & n24475 ) | ( ~n24474 & n24475 ) ;
  assign n24477 = ( n7603 & n14290 ) | ( n7603 & ~n20517 ) | ( n14290 & ~n20517 ) ;
  assign n24478 = ( n4498 & ~n4850 ) | ( n4498 & n12802 ) | ( ~n4850 & n12802 ) ;
  assign n24479 = n24478 ^ n15119 ^ n10680 ;
  assign n24480 = n14786 ^ n12515 ^ n302 ;
  assign n24481 = n24480 ^ n16061 ^ n14641 ;
  assign n24482 = ( n7794 & n22293 ) | ( n7794 & n24481 ) | ( n22293 & n24481 ) ;
  assign n24483 = n4430 ^ n4162 ^ n3316 ;
  assign n24484 = ( n4435 & n24482 ) | ( n4435 & ~n24483 ) | ( n24482 & ~n24483 ) ;
  assign n24485 = n24484 ^ n10411 ^ n5578 ;
  assign n24487 = ( n905 & n18180 ) | ( n905 & n22434 ) | ( n18180 & n22434 ) ;
  assign n24488 = ( n16543 & ~n22545 ) | ( n16543 & n24487 ) | ( ~n22545 & n24487 ) ;
  assign n24486 = n17434 ^ n10013 ^ n4071 ;
  assign n24489 = n24488 ^ n24486 ^ n16430 ;
  assign n24490 = ( ~n5233 & n8151 ) | ( ~n5233 & n14356 ) | ( n8151 & n14356 ) ;
  assign n24491 = ( n195 & n21361 ) | ( n195 & ~n23506 ) | ( n21361 & ~n23506 ) ;
  assign n24492 = ( n7519 & n24490 ) | ( n7519 & ~n24491 ) | ( n24490 & ~n24491 ) ;
  assign n24493 = n322 | n3271 ;
  assign n24494 = n24493 ^ n4925 ^ n1016 ;
  assign n24495 = ( n5644 & n17893 ) | ( n5644 & ~n23175 ) | ( n17893 & ~n23175 ) ;
  assign n24496 = ( n9134 & ~n24494 ) | ( n9134 & n24495 ) | ( ~n24494 & n24495 ) ;
  assign n24497 = ( ~n8588 & n9364 ) | ( ~n8588 & n15862 ) | ( n9364 & n15862 ) ;
  assign n24498 = n24497 ^ n14633 ^ 1'b0 ;
  assign n24499 = ( n2922 & n13827 ) | ( n2922 & n24498 ) | ( n13827 & n24498 ) ;
  assign n24500 = n5251 & n9895 ;
  assign n24501 = ( n202 & n8485 ) | ( n202 & n12660 ) | ( n8485 & n12660 ) ;
  assign n24502 = ( n351 & n4631 ) | ( n351 & n24501 ) | ( n4631 & n24501 ) ;
  assign n24503 = n11356 ^ n6473 ^ n5143 ;
  assign n24504 = n15923 ^ n1499 ^ 1'b0 ;
  assign n24505 = n1589 & n24504 ;
  assign n24506 = n24505 ^ n18383 ^ n5692 ;
  assign n24507 = n24506 ^ n15389 ^ n4625 ;
  assign n24508 = n23059 ^ n2553 ^ n1497 ;
  assign n24509 = n24508 ^ n1157 ^ n280 ;
  assign n24510 = n14781 ^ n12630 ^ n4223 ;
  assign n24511 = n24510 ^ n21289 ^ n823 ;
  assign n24512 = n16491 ^ n8603 ^ n3982 ;
  assign n24513 = ( n6966 & n9066 ) | ( n6966 & n20969 ) | ( n9066 & n20969 ) ;
  assign n24514 = n24513 ^ n10745 ^ x118 ;
  assign n24515 = ( n19268 & n20388 ) | ( n19268 & ~n24514 ) | ( n20388 & ~n24514 ) ;
  assign n24516 = n1711 | n20402 ;
  assign n24517 = n24516 ^ n14449 ^ 1'b0 ;
  assign n24518 = ( n2703 & n6318 ) | ( n2703 & n6372 ) | ( n6318 & n6372 ) ;
  assign n24519 = n21799 & ~n24518 ;
  assign n24520 = n418 & n24519 ;
  assign n24521 = ( n11371 & n12348 ) | ( n11371 & n24488 ) | ( n12348 & n24488 ) ;
  assign n24525 = n7730 ^ n5026 ^ n656 ;
  assign n24522 = ( n2874 & n4576 ) | ( n2874 & ~n7807 ) | ( n4576 & ~n7807 ) ;
  assign n24523 = ( n10668 & ~n21629 ) | ( n10668 & n24522 ) | ( ~n21629 & n24522 ) ;
  assign n24524 = n24523 ^ n8354 ^ n7490 ;
  assign n24526 = n24525 ^ n24524 ^ n22872 ;
  assign n24527 = n24526 ^ n12087 ^ n10836 ;
  assign n24528 = ( ~n3196 & n5470 ) | ( ~n3196 & n23555 ) | ( n5470 & n23555 ) ;
  assign n24529 = ( n1331 & ~n7382 ) | ( n1331 & n24528 ) | ( ~n7382 & n24528 ) ;
  assign n24530 = n18496 & n24529 ;
  assign n24531 = n24530 ^ n15344 ^ 1'b0 ;
  assign n24532 = n24531 ^ n13566 ^ n11280 ;
  assign n24533 = n6559 ^ n4611 ^ n555 ;
  assign n24538 = ( ~n1503 & n9529 ) | ( ~n1503 & n9540 ) | ( n9529 & n9540 ) ;
  assign n24536 = ~n2629 & n10264 ;
  assign n24534 = ( n11111 & ~n12115 ) | ( n11111 & n18918 ) | ( ~n12115 & n18918 ) ;
  assign n24535 = n24534 ^ n24298 ^ n5914 ;
  assign n24537 = n24536 ^ n24535 ^ n599 ;
  assign n24539 = n24538 ^ n24537 ^ n23885 ;
  assign n24540 = n22528 ^ n12397 ^ n384 ;
  assign n24541 = ( n5153 & n12945 ) | ( n5153 & ~n24171 ) | ( n12945 & ~n24171 ) ;
  assign n24542 = n22356 ^ n14826 ^ 1'b0 ;
  assign n24543 = n23158 ^ n12569 ^ 1'b0 ;
  assign n24544 = n5000 & ~n24543 ;
  assign n24545 = ~n18531 & n24544 ;
  assign n24546 = n24545 ^ n6513 ^ 1'b0 ;
  assign n24547 = n6726 ^ n4663 ^ 1'b0 ;
  assign n24548 = ( n1584 & n18492 ) | ( n1584 & ~n24547 ) | ( n18492 & ~n24547 ) ;
  assign n24549 = n23745 ^ n3332 ^ n1477 ;
  assign n24550 = ( n6536 & ~n17706 ) | ( n6536 & n24549 ) | ( ~n17706 & n24549 ) ;
  assign n24551 = n17403 ^ n7133 ^ 1'b0 ;
  assign n24552 = ( n1712 & ~n22539 ) | ( n1712 & n22822 ) | ( ~n22539 & n22822 ) ;
  assign n24553 = n4690 ^ n2987 ^ n2247 ;
  assign n24554 = ( n2022 & n8156 ) | ( n2022 & n11082 ) | ( n8156 & n11082 ) ;
  assign n24555 = n8659 ^ n7168 ^ n5378 ;
  assign n24556 = n24555 ^ n21613 ^ n840 ;
  assign n24557 = ~n3876 & n23316 ;
  assign n24558 = n24557 ^ n12086 ^ 1'b0 ;
  assign n24559 = n14789 | n24558 ;
  assign n24561 = n13880 ^ n11760 ^ n2476 ;
  assign n24562 = n24561 ^ n13281 ^ n3035 ;
  assign n24563 = n24562 ^ n20136 ^ n16147 ;
  assign n24560 = ~n7137 & n20241 ;
  assign n24564 = n24563 ^ n24560 ^ 1'b0 ;
  assign n24565 = ( n6403 & ~n14490 ) | ( n6403 & n14583 ) | ( ~n14490 & n14583 ) ;
  assign n24566 = n24565 ^ n3375 ^ n334 ;
  assign n24567 = n17462 ^ n13415 ^ n11552 ;
  assign n24568 = n8529 ^ n1764 ^ n258 ;
  assign n24569 = ( n490 & n1478 ) | ( n490 & ~n4553 ) | ( n1478 & ~n4553 ) ;
  assign n24570 = ( n10811 & ~n24568 ) | ( n10811 & n24569 ) | ( ~n24568 & n24569 ) ;
  assign n24571 = n15923 ^ n13649 ^ n564 ;
  assign n24572 = n15193 | n24571 ;
  assign n24573 = ( ~n285 & n859 ) | ( ~n285 & n17574 ) | ( n859 & n17574 ) ;
  assign n24574 = n15827 ^ n6171 ^ 1'b0 ;
  assign n24575 = n22383 & ~n24574 ;
  assign n24576 = ( ~n11521 & n20422 ) | ( ~n11521 & n24575 ) | ( n20422 & n24575 ) ;
  assign n24577 = n24576 ^ n12331 ^ 1'b0 ;
  assign n24578 = ( n4018 & n7334 ) | ( n4018 & ~n10583 ) | ( n7334 & ~n10583 ) ;
  assign n24579 = n4993 | n24399 ;
  assign n24580 = n24579 ^ n24108 ^ 1'b0 ;
  assign n24581 = ( ~n10157 & n24578 ) | ( ~n10157 & n24580 ) | ( n24578 & n24580 ) ;
  assign n24582 = n1393 & n5092 ;
  assign n24583 = n24582 ^ n20277 ^ 1'b0 ;
  assign n24586 = ( n3817 & n3935 ) | ( n3817 & ~n5015 ) | ( n3935 & ~n5015 ) ;
  assign n24587 = n12614 ^ n5685 ^ n3726 ;
  assign n24588 = n24587 ^ n18391 ^ 1'b0 ;
  assign n24589 = ~n24586 & n24588 ;
  assign n24584 = ( n2490 & ~n15207 ) | ( n2490 & n20258 ) | ( ~n15207 & n20258 ) ;
  assign n24585 = n24584 ^ n22881 ^ 1'b0 ;
  assign n24590 = n24589 ^ n24585 ^ n3954 ;
  assign n24591 = n22035 ^ n15466 ^ n5946 ;
  assign n24592 = n17610 ^ n15848 ^ n10060 ;
  assign n24593 = ( n1858 & n5549 ) | ( n1858 & n6270 ) | ( n5549 & n6270 ) ;
  assign n24594 = n24593 ^ n18520 ^ n8648 ;
  assign n24595 = ~n24592 & n24594 ;
  assign n24596 = ( ~n4398 & n12643 ) | ( ~n4398 & n12784 ) | ( n12643 & n12784 ) ;
  assign n24597 = ( n11257 & n13876 ) | ( n11257 & n24596 ) | ( n13876 & n24596 ) ;
  assign n24598 = ( ~n3788 & n11942 ) | ( ~n3788 & n17379 ) | ( n11942 & n17379 ) ;
  assign n24599 = ( n1817 & n12574 ) | ( n1817 & ~n24598 ) | ( n12574 & ~n24598 ) ;
  assign n24600 = n24599 ^ n14448 ^ n4977 ;
  assign n24602 = n1707 ^ n1462 ^ n907 ;
  assign n24601 = n8446 ^ n5795 ^ n4567 ;
  assign n24603 = n24602 ^ n24601 ^ n375 ;
  assign n24604 = n24603 ^ n419 ^ 1'b0 ;
  assign n24605 = n17717 & ~n24604 ;
  assign n24606 = ~n3411 & n8380 ;
  assign n24607 = n24606 ^ n677 ^ 1'b0 ;
  assign n24608 = n24607 ^ n15220 ^ 1'b0 ;
  assign n24609 = n9423 & ~n24608 ;
  assign n24610 = n7907 & n10994 ;
  assign n24611 = ( ~n1881 & n2209 ) | ( ~n1881 & n7314 ) | ( n2209 & n7314 ) ;
  assign n24612 = n24611 ^ n23558 ^ n4808 ;
  assign n24613 = ( n11209 & n20578 ) | ( n11209 & ~n24612 ) | ( n20578 & ~n24612 ) ;
  assign n24617 = ( n6366 & n11768 ) | ( n6366 & n14776 ) | ( n11768 & n14776 ) ;
  assign n24618 = ( n8686 & ~n9588 ) | ( n8686 & n24617 ) | ( ~n9588 & n24617 ) ;
  assign n24614 = n23277 ^ n14273 ^ n6199 ;
  assign n24615 = n24614 ^ n14733 ^ n2273 ;
  assign n24616 = ( n11814 & n15724 ) | ( n11814 & n24615 ) | ( n15724 & n24615 ) ;
  assign n24619 = n24618 ^ n24616 ^ n24461 ;
  assign n24620 = n12460 ^ n8599 ^ n5905 ;
  assign n24621 = n23090 ^ n18119 ^ n15281 ;
  assign n24622 = ( n20009 & n24620 ) | ( n20009 & n24621 ) | ( n24620 & n24621 ) ;
  assign n24623 = ( n3729 & ~n14938 ) | ( n3729 & n20541 ) | ( ~n14938 & n20541 ) ;
  assign n24624 = ( n5241 & ~n18934 ) | ( n5241 & n24623 ) | ( ~n18934 & n24623 ) ;
  assign n24626 = n3358 | n16910 ;
  assign n24625 = ~n8834 & n10601 ;
  assign n24627 = n24626 ^ n24625 ^ n3593 ;
  assign n24628 = n24627 ^ n16969 ^ n14208 ;
  assign n24629 = ( ~n12264 & n18768 ) | ( ~n12264 & n24628 ) | ( n18768 & n24628 ) ;
  assign n24630 = n16653 ^ n4485 ^ n3175 ;
  assign n24631 = n17121 ^ n3172 ^ n1700 ;
  assign n24632 = n24631 ^ n15936 ^ n630 ;
  assign n24633 = ( n7891 & n8310 ) | ( n7891 & ~n17105 ) | ( n8310 & ~n17105 ) ;
  assign n24634 = ( ~n3441 & n5309 ) | ( ~n3441 & n7737 ) | ( n5309 & n7737 ) ;
  assign n24635 = ( n3022 & ~n15592 ) | ( n3022 & n24634 ) | ( ~n15592 & n24634 ) ;
  assign n24636 = ( n4015 & n24633 ) | ( n4015 & n24635 ) | ( n24633 & n24635 ) ;
  assign n24637 = ( n660 & n2427 ) | ( n660 & ~n16253 ) | ( n2427 & ~n16253 ) ;
  assign n24638 = n24637 ^ n9171 ^ n2906 ;
  assign n24639 = n11077 ^ n10704 ^ n6482 ;
  assign n24640 = n5599 & n24639 ;
  assign n24641 = n13999 ^ n9202 ^ n7076 ;
  assign n24642 = ( x10 & n15683 ) | ( x10 & ~n24641 ) | ( n15683 & ~n24641 ) ;
  assign n24643 = ( ~n1644 & n22489 ) | ( ~n1644 & n24642 ) | ( n22489 & n24642 ) ;
  assign n24644 = n23287 ^ n19519 ^ n9343 ;
  assign n24645 = n4062 ^ n4007 ^ n3765 ;
  assign n24646 = ( n2600 & n2837 ) | ( n2600 & ~n12387 ) | ( n2837 & ~n12387 ) ;
  assign n24647 = n516 & n24646 ;
  assign n24648 = ( n7243 & ~n9833 ) | ( n7243 & n24647 ) | ( ~n9833 & n24647 ) ;
  assign n24649 = ( n24644 & n24645 ) | ( n24644 & ~n24648 ) | ( n24645 & ~n24648 ) ;
  assign n24650 = ~n6812 & n17463 ;
  assign n24651 = ( n983 & n1876 ) | ( n983 & n6928 ) | ( n1876 & n6928 ) ;
  assign n24652 = n24651 ^ n3070 ^ n2489 ;
  assign n24653 = n21371 ^ n4765 ^ 1'b0 ;
  assign n24654 = ~n24652 & n24653 ;
  assign n24655 = ( ~n15799 & n24650 ) | ( ~n15799 & n24654 ) | ( n24650 & n24654 ) ;
  assign n24656 = ( n422 & ~n8616 ) | ( n422 & n11879 ) | ( ~n8616 & n11879 ) ;
  assign n24657 = n9149 | n18871 ;
  assign n24658 = n24657 ^ n1021 ^ 1'b0 ;
  assign n24659 = ( n905 & ~n17075 ) | ( n905 & n24658 ) | ( ~n17075 & n24658 ) ;
  assign n24660 = n18912 ^ n8510 ^ 1'b0 ;
  assign n24661 = ( n720 & n17291 ) | ( n720 & n22669 ) | ( n17291 & n22669 ) ;
  assign n24662 = ( n1482 & ~n11258 ) | ( n1482 & n24661 ) | ( ~n11258 & n24661 ) ;
  assign n24663 = n20814 ^ n11814 ^ n11099 ;
  assign n24664 = n24663 ^ n21784 ^ n2410 ;
  assign n24665 = ( n939 & n11955 ) | ( n939 & ~n23416 ) | ( n11955 & ~n23416 ) ;
  assign n24666 = n10280 ^ n5469 ^ n5400 ;
  assign n24667 = ~n11346 & n24666 ;
  assign n24668 = ( n1438 & n10809 ) | ( n1438 & n11382 ) | ( n10809 & n11382 ) ;
  assign n24669 = ( n2267 & n8094 ) | ( n2267 & ~n24668 ) | ( n8094 & ~n24668 ) ;
  assign n24670 = n24669 ^ n21682 ^ n5831 ;
  assign n24671 = n7428 ^ n1172 ^ 1'b0 ;
  assign n24672 = n18857 & ~n24671 ;
  assign n24673 = n908 & ~n12792 ;
  assign n24674 = n24673 ^ n4019 ^ 1'b0 ;
  assign n24675 = n24672 & n24674 ;
  assign n24676 = ~n4151 & n9609 ;
  assign n24677 = n24676 ^ n8581 ^ n6088 ;
  assign n24678 = ( n5578 & ~n15985 ) | ( n5578 & n24677 ) | ( ~n15985 & n24677 ) ;
  assign n24679 = ( ~n1084 & n7212 ) | ( ~n1084 & n24678 ) | ( n7212 & n24678 ) ;
  assign n24680 = n18885 | n21883 ;
  assign n24681 = n24679 | n24680 ;
  assign n24682 = n21143 ^ n12140 ^ n1490 ;
  assign n24683 = n24682 ^ n22249 ^ n15814 ;
  assign n24684 = n24330 ^ n21454 ^ n19832 ;
  assign n24685 = ( n2156 & n6114 ) | ( n2156 & ~n24684 ) | ( n6114 & ~n24684 ) ;
  assign n24686 = n3325 ^ x101 ^ 1'b0 ;
  assign n24687 = ( ~n3883 & n7654 ) | ( ~n3883 & n24686 ) | ( n7654 & n24686 ) ;
  assign n24688 = ( ~n9412 & n11129 ) | ( ~n9412 & n24687 ) | ( n11129 & n24687 ) ;
  assign n24689 = ( n1361 & n18373 ) | ( n1361 & n20986 ) | ( n18373 & n20986 ) ;
  assign n24690 = ( n7201 & n24688 ) | ( n7201 & n24689 ) | ( n24688 & n24689 ) ;
  assign n24691 = ( n4972 & n12630 ) | ( n4972 & ~n17824 ) | ( n12630 & ~n17824 ) ;
  assign n24692 = ( n14215 & n20355 ) | ( n14215 & n24691 ) | ( n20355 & n24691 ) ;
  assign n24693 = n12768 ^ n6913 ^ 1'b0 ;
  assign n24694 = n24692 & n24693 ;
  assign n24695 = ( n2085 & n4858 ) | ( n2085 & n24694 ) | ( n4858 & n24694 ) ;
  assign n24696 = n20089 ^ n13966 ^ n5802 ;
  assign n24697 = n6636 ^ n2808 ^ n2269 ;
  assign n24698 = n6007 | n10623 ;
  assign n24699 = n24698 ^ n21201 ^ 1'b0 ;
  assign n24700 = n20797 | n24699 ;
  assign n24701 = n24700 ^ n22931 ^ n14703 ;
  assign n24702 = ( n11558 & ~n24697 ) | ( n11558 & n24701 ) | ( ~n24697 & n24701 ) ;
  assign n24703 = ( ~n7592 & n9929 ) | ( ~n7592 & n11393 ) | ( n9929 & n11393 ) ;
  assign n24704 = n24703 ^ n14614 ^ n926 ;
  assign n24705 = ( n8344 & ~n17640 ) | ( n8344 & n24704 ) | ( ~n17640 & n24704 ) ;
  assign n24708 = ( n2414 & n13552 ) | ( n2414 & ~n18778 ) | ( n13552 & ~n18778 ) ;
  assign n24706 = ( n6404 & n10775 ) | ( n6404 & n13090 ) | ( n10775 & n13090 ) ;
  assign n24707 = ( n15101 & n19457 ) | ( n15101 & n24706 ) | ( n19457 & n24706 ) ;
  assign n24709 = n24708 ^ n24707 ^ n430 ;
  assign n24710 = n21227 | n22637 ;
  assign n24711 = n23378 | n24710 ;
  assign n24712 = n14404 & n16977 ;
  assign n24713 = n16574 & n24712 ;
  assign n24714 = ( n2607 & n4075 ) | ( n2607 & n15911 ) | ( n4075 & n15911 ) ;
  assign n24715 = ( n7344 & ~n19485 ) | ( n7344 & n23567 ) | ( ~n19485 & n23567 ) ;
  assign n24716 = ( n14211 & ~n24714 ) | ( n14211 & n24715 ) | ( ~n24714 & n24715 ) ;
  assign n24717 = ( n2481 & n16804 ) | ( n2481 & n24478 ) | ( n16804 & n24478 ) ;
  assign n24718 = n24717 ^ n2315 ^ 1'b0 ;
  assign n24719 = ( n2798 & ~n2816 ) | ( n2798 & n12032 ) | ( ~n2816 & n12032 ) ;
  assign n24720 = n7099 | n24719 ;
  assign n24721 = n24720 ^ n16245 ^ 1'b0 ;
  assign n24722 = n24721 ^ n8403 ^ n7175 ;
  assign n24723 = n24718 & n24722 ;
  assign n24724 = n24723 ^ n19037 ^ n14669 ;
  assign n24725 = ( ~n10169 & n13159 ) | ( ~n10169 & n15005 ) | ( n13159 & n15005 ) ;
  assign n24726 = ( n785 & ~n1331 ) | ( n785 & n2152 ) | ( ~n1331 & n2152 ) ;
  assign n24727 = n24725 & n24726 ;
  assign n24728 = ( ~n17815 & n21002 ) | ( ~n17815 & n24727 ) | ( n21002 & n24727 ) ;
  assign n24729 = ( n444 & n5327 ) | ( n444 & ~n22912 ) | ( n5327 & ~n22912 ) ;
  assign n24730 = n24729 ^ n20542 ^ 1'b0 ;
  assign n24731 = ( n6094 & n8300 ) | ( n6094 & ~n8794 ) | ( n8300 & ~n8794 ) ;
  assign n24732 = n24731 ^ n7104 ^ n995 ;
  assign n24733 = n16199 ^ n9686 ^ 1'b0 ;
  assign n24734 = ~n15714 & n24733 ;
  assign n24735 = n24734 ^ n20302 ^ n16587 ;
  assign n24736 = n19489 | n22606 ;
  assign n24737 = n19271 & ~n24736 ;
  assign n24739 = ( x13 & n7765 ) | ( x13 & n18500 ) | ( n7765 & n18500 ) ;
  assign n24738 = n14306 ^ n14275 ^ n14270 ;
  assign n24740 = n24739 ^ n24738 ^ n5632 ;
  assign n24741 = x21 & n24740 ;
  assign n24744 = n2664 ^ n435 ^ 1'b0 ;
  assign n24745 = ( n11749 & n21052 ) | ( n11749 & n24744 ) | ( n21052 & n24744 ) ;
  assign n24746 = ( ~n2657 & n14337 ) | ( ~n2657 & n24745 ) | ( n14337 & n24745 ) ;
  assign n24742 = n19926 ^ n3088 ^ n1525 ;
  assign n24743 = ( n5126 & n8645 ) | ( n5126 & n24742 ) | ( n8645 & n24742 ) ;
  assign n24747 = n24746 ^ n24743 ^ n6764 ;
  assign n24748 = ( n7156 & ~n16714 ) | ( n7156 & n19492 ) | ( ~n16714 & n19492 ) ;
  assign n24749 = n24748 ^ n19214 ^ n852 ;
  assign n24750 = n19037 ^ n10861 ^ n8506 ;
  assign n24751 = ( n4401 & ~n8445 ) | ( n4401 & n24041 ) | ( ~n8445 & n24041 ) ;
  assign n24752 = ( ~x46 & n18380 ) | ( ~x46 & n24751 ) | ( n18380 & n24751 ) ;
  assign n24753 = ( n3772 & n8370 ) | ( n3772 & ~n24752 ) | ( n8370 & ~n24752 ) ;
  assign n24754 = n14662 ^ n6399 ^ n3630 ;
  assign n24756 = n18889 ^ n4223 ^ n4083 ;
  assign n24757 = ( n8054 & ~n20851 ) | ( n8054 & n24756 ) | ( ~n20851 & n24756 ) ;
  assign n24755 = ( n3916 & n4075 ) | ( n3916 & ~n11267 ) | ( n4075 & ~n11267 ) ;
  assign n24758 = n24757 ^ n24755 ^ n17574 ;
  assign n24759 = n16245 ^ n10944 ^ n2162 ;
  assign n24760 = ( n5149 & n10800 ) | ( n5149 & ~n12448 ) | ( n10800 & ~n12448 ) ;
  assign n24761 = n24760 ^ n6352 ^ 1'b0 ;
  assign n24762 = ( ~n9028 & n24759 ) | ( ~n9028 & n24761 ) | ( n24759 & n24761 ) ;
  assign n24763 = ( n491 & n8462 ) | ( n491 & n24247 ) | ( n8462 & n24247 ) ;
  assign n24764 = ( n21987 & ~n23472 ) | ( n21987 & n24763 ) | ( ~n23472 & n24763 ) ;
  assign n24765 = ( x34 & n690 ) | ( x34 & n4624 ) | ( n690 & n4624 ) ;
  assign n24766 = ( n15658 & ~n16542 ) | ( n15658 & n24765 ) | ( ~n16542 & n24765 ) ;
  assign n24767 = n21430 ^ n14185 ^ n9851 ;
  assign n24768 = ( ~n1130 & n4544 ) | ( ~n1130 & n14997 ) | ( n4544 & n14997 ) ;
  assign n24769 = ( n3186 & n11071 ) | ( n3186 & n16962 ) | ( n11071 & n16962 ) ;
  assign n24770 = ( ~n1456 & n3013 ) | ( ~n1456 & n10010 ) | ( n3013 & n10010 ) ;
  assign n24771 = n24770 ^ n22082 ^ n1190 ;
  assign n24772 = ( ~n9987 & n19381 ) | ( ~n9987 & n24771 ) | ( n19381 & n24771 ) ;
  assign n24774 = n2751 & ~n19459 ;
  assign n24775 = n6606 & n24774 ;
  assign n24773 = ( n1792 & ~n3957 ) | ( n1792 & n19449 ) | ( ~n3957 & n19449 ) ;
  assign n24776 = n24775 ^ n24773 ^ n16515 ;
  assign n24777 = n24776 ^ n11053 ^ n10994 ;
  assign n24778 = ( ~n2442 & n15464 ) | ( ~n2442 & n23200 ) | ( n15464 & n23200 ) ;
  assign n24779 = n11700 ^ n8483 ^ 1'b0 ;
  assign n24780 = ( ~n9038 & n24231 ) | ( ~n9038 & n24779 ) | ( n24231 & n24779 ) ;
  assign n24781 = n5871 & ~n8184 ;
  assign n24782 = n24781 ^ n11884 ^ 1'b0 ;
  assign n24784 = ( ~n443 & n5245 ) | ( ~n443 & n20028 ) | ( n5245 & n20028 ) ;
  assign n24783 = n11974 & ~n17781 ;
  assign n24785 = n24784 ^ n24783 ^ 1'b0 ;
  assign n24786 = ( ~n3318 & n12385 ) | ( ~n3318 & n21045 ) | ( n12385 & n21045 ) ;
  assign n24790 = n11468 ^ n1420 ^ 1'b0 ;
  assign n24787 = n12232 ^ n4869 ^ n2977 ;
  assign n24788 = n24787 ^ n10677 ^ n8702 ;
  assign n24789 = n24788 ^ n10268 ^ n8115 ;
  assign n24791 = n24790 ^ n24789 ^ n5312 ;
  assign n24792 = n17873 ^ n8243 ^ n542 ;
  assign n24793 = n5223 ^ n793 ^ 1'b0 ;
  assign n24794 = n5166 & ~n24793 ;
  assign n24795 = n24794 ^ n2806 ^ 1'b0 ;
  assign n24796 = n15596 ^ n3196 ^ 1'b0 ;
  assign n24797 = n16134 & n24796 ;
  assign n24798 = n24797 ^ n795 ^ 1'b0 ;
  assign n24799 = n19277 | n24798 ;
  assign n24800 = ( n5174 & ~n24795 ) | ( n5174 & n24799 ) | ( ~n24795 & n24799 ) ;
  assign n24803 = ( n2853 & n5831 ) | ( n2853 & ~n9229 ) | ( n5831 & ~n9229 ) ;
  assign n24801 = ( ~n4439 & n9533 ) | ( ~n4439 & n14952 ) | ( n9533 & n14952 ) ;
  assign n24802 = ( n405 & n21221 ) | ( n405 & ~n24801 ) | ( n21221 & ~n24801 ) ;
  assign n24804 = n24803 ^ n24802 ^ n2937 ;
  assign n24805 = ( n2438 & n8241 ) | ( n2438 & ~n18119 ) | ( n8241 & ~n18119 ) ;
  assign n24806 = n24805 ^ n5285 ^ n264 ;
  assign n24807 = n13936 ^ n7945 ^ n4847 ;
  assign n24808 = ( n12329 & n24806 ) | ( n12329 & ~n24807 ) | ( n24806 & ~n24807 ) ;
  assign n24809 = n9722 ^ n6407 ^ n1696 ;
  assign n24810 = n24809 ^ n17698 ^ n3179 ;
  assign n24811 = ( ~n2882 & n17548 ) | ( ~n2882 & n24810 ) | ( n17548 & n24810 ) ;
  assign n24813 = n21423 ^ n10502 ^ n8180 ;
  assign n24812 = n7271 ^ n4587 ^ 1'b0 ;
  assign n24814 = n24813 ^ n24812 ^ n7897 ;
  assign n24815 = n22625 ^ n9920 ^ n4325 ;
  assign n24816 = ( n7196 & ~n7338 ) | ( n7196 & n24815 ) | ( ~n7338 & n24815 ) ;
  assign n24817 = n9115 ^ n5799 ^ n1727 ;
  assign n24818 = ( n676 & n19303 ) | ( n676 & n20398 ) | ( n19303 & n20398 ) ;
  assign n24820 = ( n681 & n6208 ) | ( n681 & n19492 ) | ( n6208 & n19492 ) ;
  assign n24819 = n11739 ^ n8279 ^ 1'b0 ;
  assign n24821 = n24820 ^ n24819 ^ n24469 ;
  assign n24822 = n10240 & ~n10380 ;
  assign n24823 = n19077 ^ n3323 ^ 1'b0 ;
  assign n24824 = n18256 ^ n7369 ^ n1654 ;
  assign n24825 = ( n722 & n13496 ) | ( n722 & ~n24824 ) | ( n13496 & ~n24824 ) ;
  assign n24826 = n24825 ^ n7910 ^ 1'b0 ;
  assign n24827 = ~n24823 & n24826 ;
  assign n24828 = ( n1693 & ~n13307 ) | ( n1693 & n22780 ) | ( ~n13307 & n22780 ) ;
  assign n24829 = ( n4002 & n15773 ) | ( n4002 & n22527 ) | ( n15773 & n22527 ) ;
  assign n24830 = ( ~n5754 & n24828 ) | ( ~n5754 & n24829 ) | ( n24828 & n24829 ) ;
  assign n24831 = n16081 ^ n8926 ^ n605 ;
  assign n24832 = n5648 | n24831 ;
  assign n24833 = n14439 ^ n9720 ^ n3476 ;
  assign n24834 = n24833 ^ n19139 ^ n13531 ;
  assign n24835 = ( n6277 & n24832 ) | ( n6277 & n24834 ) | ( n24832 & n24834 ) ;
  assign n24838 = n18404 ^ n13304 ^ n7068 ;
  assign n24836 = n5398 ^ n4018 ^ 1'b0 ;
  assign n24837 = n24836 ^ n8251 ^ 1'b0 ;
  assign n24839 = n24838 ^ n24837 ^ n2769 ;
  assign n24840 = n19492 ^ n17425 ^ n313 ;
  assign n24841 = n6282 ^ n4374 ^ n3295 ;
  assign n24842 = n23446 ^ n15020 ^ n11014 ;
  assign n24843 = ( x45 & ~n1226 ) | ( x45 & n24842 ) | ( ~n1226 & n24842 ) ;
  assign n24844 = n24843 ^ n11226 ^ 1'b0 ;
  assign n24845 = n24844 ^ n8691 ^ n360 ;
  assign n24846 = n14447 ^ n8775 ^ 1'b0 ;
  assign n24847 = ~n24845 & n24846 ;
  assign n24848 = n8262 ^ n4135 ^ 1'b0 ;
  assign n24849 = ( ~n2178 & n9000 ) | ( ~n2178 & n13636 ) | ( n9000 & n13636 ) ;
  assign n24850 = n24849 ^ n10262 ^ n361 ;
  assign n24851 = ( n13025 & n15057 ) | ( n13025 & ~n19561 ) | ( n15057 & ~n19561 ) ;
  assign n24852 = ( ~n1461 & n2539 ) | ( ~n1461 & n12730 ) | ( n2539 & n12730 ) ;
  assign n24853 = ( x98 & n1022 ) | ( x98 & ~n1695 ) | ( n1022 & ~n1695 ) ;
  assign n24854 = ( n4206 & n14162 ) | ( n4206 & n24853 ) | ( n14162 & n24853 ) ;
  assign n24855 = n24854 ^ n16262 ^ n11138 ;
  assign n24856 = ( n3870 & n11220 ) | ( n3870 & n24855 ) | ( n11220 & n24855 ) ;
  assign n24857 = ( ~n10098 & n21784 ) | ( ~n10098 & n24856 ) | ( n21784 & n24856 ) ;
  assign n24858 = n12377 | n12436 ;
  assign n24859 = n24858 ^ n18207 ^ n13274 ;
  assign n24860 = n5125 & ~n12480 ;
  assign n24861 = n24860 ^ n11622 ^ 1'b0 ;
  assign n24862 = n24861 ^ n14522 ^ n7931 ;
  assign n24863 = ~n2966 & n5860 ;
  assign n24864 = n24863 ^ n2113 ^ 1'b0 ;
  assign n24865 = n8827 ^ n4508 ^ 1'b0 ;
  assign n24866 = n2542 & n24865 ;
  assign n24867 = n12803 ^ n6520 ^ 1'b0 ;
  assign n24868 = ( ~n24864 & n24866 ) | ( ~n24864 & n24867 ) | ( n24866 & n24867 ) ;
  assign n24869 = ( n411 & ~n9708 ) | ( n411 & n14164 ) | ( ~n9708 & n14164 ) ;
  assign n24870 = n7384 & n8990 ;
  assign n24871 = n24870 ^ n14073 ^ 1'b0 ;
  assign n24872 = ( n1460 & n2975 ) | ( n1460 & ~n6439 ) | ( n2975 & ~n6439 ) ;
  assign n24873 = n24872 ^ n23670 ^ n11807 ;
  assign n24876 = n7596 ^ n3138 ^ n962 ;
  assign n24875 = ( n1842 & n3931 ) | ( n1842 & ~n19183 ) | ( n3931 & ~n19183 ) ;
  assign n24874 = ( n3576 & n7151 ) | ( n3576 & ~n11576 ) | ( n7151 & ~n11576 ) ;
  assign n24877 = n24876 ^ n24875 ^ n24874 ;
  assign n24878 = ( n1158 & ~n3884 ) | ( n1158 & n15967 ) | ( ~n3884 & n15967 ) ;
  assign n24879 = ( n4906 & n9942 ) | ( n4906 & n18736 ) | ( n9942 & n18736 ) ;
  assign n24880 = n24879 ^ n19300 ^ n18096 ;
  assign n24881 = ( ~n17755 & n19909 ) | ( ~n17755 & n24880 ) | ( n19909 & n24880 ) ;
  assign n24882 = n22276 ^ n20432 ^ n12479 ;
  assign n24883 = n5476 & n7191 ;
  assign n24884 = n24883 ^ n18087 ^ 1'b0 ;
  assign n24885 = n24884 ^ n15093 ^ 1'b0 ;
  assign n24886 = n18061 ^ n9631 ^ n8875 ;
  assign n24888 = n11696 ^ n3281 ^ 1'b0 ;
  assign n24889 = ~n7335 & n24888 ;
  assign n24890 = ( n1112 & ~n14562 ) | ( n1112 & n24889 ) | ( ~n14562 & n24889 ) ;
  assign n24887 = ( ~n2717 & n11418 ) | ( ~n2717 & n21849 ) | ( n11418 & n21849 ) ;
  assign n24891 = n24890 ^ n24887 ^ n10587 ;
  assign n24892 = ( n8954 & n24886 ) | ( n8954 & n24891 ) | ( n24886 & n24891 ) ;
  assign n24897 = ( ~n7118 & n8793 ) | ( ~n7118 & n8952 ) | ( n8793 & n8952 ) ;
  assign n24893 = ( n142 & n3201 ) | ( n142 & n11130 ) | ( n3201 & n11130 ) ;
  assign n24894 = ( ~n2899 & n11047 ) | ( ~n2899 & n24893 ) | ( n11047 & n24893 ) ;
  assign n24895 = ( n3145 & ~n18645 ) | ( n3145 & n20728 ) | ( ~n18645 & n20728 ) ;
  assign n24896 = ( n16335 & n24894 ) | ( n16335 & ~n24895 ) | ( n24894 & ~n24895 ) ;
  assign n24898 = n24897 ^ n24896 ^ n8016 ;
  assign n24899 = n10393 ^ n8886 ^ n8643 ;
  assign n24900 = ~n3966 & n12048 ;
  assign n24901 = n24900 ^ n18282 ^ 1'b0 ;
  assign n24902 = n24901 ^ n9132 ^ 1'b0 ;
  assign n24903 = n24899 | n24902 ;
  assign n24904 = ( ~x66 & n8268 ) | ( ~x66 & n19086 ) | ( n8268 & n19086 ) ;
  assign n24905 = n14820 ^ n7148 ^ n4508 ;
  assign n24906 = ( n19289 & n24904 ) | ( n19289 & ~n24905 ) | ( n24904 & ~n24905 ) ;
  assign n24907 = ( n2314 & n13574 ) | ( n2314 & n24906 ) | ( n13574 & n24906 ) ;
  assign n24908 = ( n2820 & ~n10052 ) | ( n2820 & n13199 ) | ( ~n10052 & n13199 ) ;
  assign n24909 = n8303 ^ n3314 ^ 1'b0 ;
  assign n24910 = n24908 & ~n24909 ;
  assign n24911 = n24910 ^ n10700 ^ n4346 ;
  assign n24912 = n24911 ^ n24706 ^ n7153 ;
  assign n24913 = ( n7153 & n9728 ) | ( n7153 & n17427 ) | ( n9728 & n17427 ) ;
  assign n24914 = n24913 ^ n10391 ^ 1'b0 ;
  assign n24915 = ( ~x52 & n5802 ) | ( ~x52 & n24914 ) | ( n5802 & n24914 ) ;
  assign n24917 = ( n3462 & n6528 ) | ( n3462 & ~n8575 ) | ( n6528 & ~n8575 ) ;
  assign n24916 = ( n4544 & n7211 ) | ( n4544 & n22496 ) | ( n7211 & n22496 ) ;
  assign n24918 = n24917 ^ n24916 ^ n23187 ;
  assign n24919 = n24918 ^ n20447 ^ n14885 ;
  assign n24920 = n17198 ^ n13655 ^ n13162 ;
  assign n24921 = ( n8505 & ~n14392 ) | ( n8505 & n21205 ) | ( ~n14392 & n21205 ) ;
  assign n24922 = ~n3457 & n14891 ;
  assign n24923 = ~n4620 & n24922 ;
  assign n24924 = ( ~n2097 & n24921 ) | ( ~n2097 & n24923 ) | ( n24921 & n24923 ) ;
  assign n24925 = n18925 ^ n15513 ^ n7266 ;
  assign n24926 = n9470 & n24925 ;
  assign n24927 = n13584 & n24926 ;
  assign n24928 = n22880 ^ n11639 ^ n9208 ;
  assign n24929 = ( n12881 & n15270 ) | ( n12881 & n24928 ) | ( n15270 & n24928 ) ;
  assign n24930 = ( n19095 & n21422 ) | ( n19095 & ~n24813 ) | ( n21422 & ~n24813 ) ;
  assign n24931 = ( n731 & n19765 ) | ( n731 & n21991 ) | ( n19765 & n21991 ) ;
  assign n24933 = ( n2767 & ~n9024 ) | ( n2767 & n16270 ) | ( ~n9024 & n16270 ) ;
  assign n24934 = n24933 ^ n3142 ^ n1308 ;
  assign n24932 = ( n3952 & ~n5338 ) | ( n3952 & n17112 ) | ( ~n5338 & n17112 ) ;
  assign n24935 = n24934 ^ n24932 ^ n6396 ;
  assign n24936 = n15282 ^ n12071 ^ n8389 ;
  assign n24937 = n16133 ^ n7461 ^ n2858 ;
  assign n24938 = ( n6546 & n9776 ) | ( n6546 & ~n24937 ) | ( n9776 & ~n24937 ) ;
  assign n24939 = n3610 & ~n6829 ;
  assign n24940 = n24939 ^ n21884 ^ 1'b0 ;
  assign n24941 = n24522 ^ n9902 ^ n1636 ;
  assign n24942 = n24941 ^ n17096 ^ n10446 ;
  assign n24943 = ( n1737 & n5149 ) | ( n1737 & n16073 ) | ( n5149 & n16073 ) ;
  assign n24944 = ( ~n13598 & n14918 ) | ( ~n13598 & n24943 ) | ( n14918 & n24943 ) ;
  assign n24945 = n4387 & ~n10534 ;
  assign n24946 = n15536 ^ n5466 ^ n3469 ;
  assign n24947 = n24946 ^ n20078 ^ n12158 ;
  assign n24948 = ( n492 & ~n3154 ) | ( n492 & n14028 ) | ( ~n3154 & n14028 ) ;
  assign n24950 = n10874 ^ x52 ^ 1'b0 ;
  assign n24949 = n21354 ^ n15225 ^ n3029 ;
  assign n24951 = n24950 ^ n24949 ^ n17985 ;
  assign n24952 = n24951 ^ n17261 ^ n2756 ;
  assign n24953 = n22824 ^ n7780 ^ 1'b0 ;
  assign n24954 = n18689 ^ n3822 ^ 1'b0 ;
  assign n24955 = ( n15343 & ~n24953 ) | ( n15343 & n24954 ) | ( ~n24953 & n24954 ) ;
  assign n24963 = n20987 ^ n14732 ^ n3802 ;
  assign n24964 = n24963 ^ n2314 ^ n1552 ;
  assign n24961 = ( ~n1983 & n16931 ) | ( ~n1983 & n17123 ) | ( n16931 & n17123 ) ;
  assign n24962 = n24961 ^ n10153 ^ n213 ;
  assign n24959 = ~n7379 & n9143 ;
  assign n24958 = n23037 ^ n8802 ^ n919 ;
  assign n24960 = n24959 ^ n24958 ^ n7667 ;
  assign n24965 = n24964 ^ n24962 ^ n24960 ;
  assign n24956 = n15669 ^ n11879 ^ n4049 ;
  assign n24957 = n24956 ^ n11038 ^ n10954 ;
  assign n24966 = n24965 ^ n24957 ^ n23621 ;
  assign n24967 = n9994 & ~n11981 ;
  assign n24968 = n4483 & n24967 ;
  assign n24969 = n8581 ^ n4130 ^ 1'b0 ;
  assign n24970 = ( n5508 & ~n16357 ) | ( n5508 & n24969 ) | ( ~n16357 & n24969 ) ;
  assign n24971 = n21952 ^ n8942 ^ n8754 ;
  assign n24972 = n12531 ^ n11537 ^ n11315 ;
  assign n24973 = n24972 ^ n22418 ^ n3051 ;
  assign n24974 = ( n7022 & n10676 ) | ( n7022 & ~n14604 ) | ( n10676 & ~n14604 ) ;
  assign n24977 = ( ~n247 & n1367 ) | ( ~n247 & n16635 ) | ( n1367 & n16635 ) ;
  assign n24975 = ( ~n1881 & n4043 ) | ( ~n1881 & n4660 ) | ( n4043 & n4660 ) ;
  assign n24976 = ( n13466 & n19747 ) | ( n13466 & n24975 ) | ( n19747 & n24975 ) ;
  assign n24978 = n24977 ^ n24976 ^ 1'b0 ;
  assign n24979 = ( n4171 & n9764 ) | ( n4171 & n23816 ) | ( n9764 & n23816 ) ;
  assign n24980 = n20225 ^ n7917 ^ n1893 ;
  assign n24981 = ( n10925 & ~n11684 ) | ( n10925 & n14233 ) | ( ~n11684 & n14233 ) ;
  assign n24982 = n24981 ^ n16299 ^ n13745 ;
  assign n24983 = n24982 ^ n10051 ^ 1'b0 ;
  assign n24984 = ( n1252 & ~n1449 ) | ( n1252 & n3888 ) | ( ~n1449 & n3888 ) ;
  assign n24985 = n24984 ^ n15598 ^ 1'b0 ;
  assign n24986 = ( ~n871 & n3089 ) | ( ~n871 & n6941 ) | ( n3089 & n6941 ) ;
  assign n24987 = n24986 ^ n2724 ^ 1'b0 ;
  assign n24988 = n24987 ^ n3029 ^ n491 ;
  assign n24989 = n8635 | n9552 ;
  assign n24990 = n19731 ^ n8754 ^ n1410 ;
  assign n24991 = ( n708 & ~n8447 ) | ( n708 & n15218 ) | ( ~n8447 & n15218 ) ;
  assign n24992 = ( n8548 & n9200 ) | ( n8548 & ~n23977 ) | ( n9200 & ~n23977 ) ;
  assign n24993 = ~n4886 & n24992 ;
  assign n24994 = n10427 & n24993 ;
  assign n24995 = ( ~n8844 & n13435 ) | ( ~n8844 & n15524 ) | ( n13435 & n15524 ) ;
  assign n24996 = ( n24991 & ~n24994 ) | ( n24991 & n24995 ) | ( ~n24994 & n24995 ) ;
  assign n24997 = n18696 ^ n11071 ^ n452 ;
  assign n24998 = n7118 ^ n2179 ^ 1'b0 ;
  assign n24999 = n22800 ^ n22645 ^ 1'b0 ;
  assign n25000 = n10302 | n24999 ;
  assign n25001 = n12314 ^ n1538 ^ n905 ;
  assign n25002 = n3727 & n25001 ;
  assign n25003 = ( n1171 & ~n9663 ) | ( n1171 & n24194 ) | ( ~n9663 & n24194 ) ;
  assign n25004 = n25003 ^ n10163 ^ n8250 ;
  assign n25005 = ( n1739 & ~n2431 ) | ( n1739 & n8408 ) | ( ~n2431 & n8408 ) ;
  assign n25006 = ( ~n15394 & n19350 ) | ( ~n15394 & n25005 ) | ( n19350 & n25005 ) ;
  assign n25007 = n24091 ^ n5646 ^ n1364 ;
  assign n25008 = n21296 ^ n8635 ^ n3987 ;
  assign n25009 = ( n12109 & n25007 ) | ( n12109 & ~n25008 ) | ( n25007 & ~n25008 ) ;
  assign n25010 = ( n11288 & n11440 ) | ( n11288 & ~n24199 ) | ( n11440 & ~n24199 ) ;
  assign n25011 = ( n2963 & n5838 ) | ( n2963 & n11144 ) | ( n5838 & n11144 ) ;
  assign n25012 = n25011 ^ n6107 ^ n4072 ;
  assign n25013 = ( n17637 & n24513 ) | ( n17637 & n25012 ) | ( n24513 & n25012 ) ;
  assign n25014 = ( n20048 & ~n21286 ) | ( n20048 & n25013 ) | ( ~n21286 & n25013 ) ;
  assign n25015 = n16908 ^ n5579 ^ n1492 ;
  assign n25016 = n2942 | n18483 ;
  assign n25017 = n25016 ^ n6849 ^ 1'b0 ;
  assign n25018 = n1983 | n10717 ;
  assign n25019 = ( n15776 & n25017 ) | ( n15776 & ~n25018 ) | ( n25017 & ~n25018 ) ;
  assign n25020 = n25019 ^ n594 ^ n284 ;
  assign n25021 = n3328 & n17133 ;
  assign n25022 = n25021 ^ n20947 ^ 1'b0 ;
  assign n25023 = n19671 ^ n16483 ^ n15352 ;
  assign n25024 = ( ~n5522 & n11809 ) | ( ~n5522 & n23094 ) | ( n11809 & n23094 ) ;
  assign n25025 = n4966 & ~n13860 ;
  assign n25026 = n25025 ^ n4096 ^ 1'b0 ;
  assign n25027 = n25026 ^ n4992 ^ n709 ;
  assign n25028 = ( n3531 & n3547 ) | ( n3531 & n3939 ) | ( n3547 & n3939 ) ;
  assign n25029 = n4210 | n25028 ;
  assign n25030 = n25029 ^ n5625 ^ n258 ;
  assign n25031 = n23130 & n25030 ;
  assign n25032 = n25031 ^ n1154 ^ 1'b0 ;
  assign n25033 = ( n15108 & ~n25027 ) | ( n15108 & n25032 ) | ( ~n25027 & n25032 ) ;
  assign n25034 = n4857 & n18912 ;
  assign n25035 = n25034 ^ n8991 ^ 1'b0 ;
  assign n25036 = ( n3752 & n17262 ) | ( n3752 & ~n25035 ) | ( n17262 & ~n25035 ) ;
  assign n25037 = ~n1594 & n17784 ;
  assign n25038 = n25037 ^ n21736 ^ n2355 ;
  assign n25039 = n12314 & ~n15929 ;
  assign n25040 = ~n13729 & n25039 ;
  assign n25041 = n25040 ^ n914 ^ 1'b0 ;
  assign n25042 = ( n3381 & n12454 ) | ( n3381 & n25041 ) | ( n12454 & n25041 ) ;
  assign n25043 = n13882 ^ n9582 ^ n1854 ;
  assign n25044 = n25043 ^ n10659 ^ n2824 ;
  assign n25045 = ~n442 & n5517 ;
  assign n25046 = n607 & n13242 ;
  assign n25047 = n25045 & n25046 ;
  assign n25048 = ( ~n3983 & n16674 ) | ( ~n3983 & n23416 ) | ( n16674 & n23416 ) ;
  assign n25049 = n18776 ^ n17830 ^ n13164 ;
  assign n25050 = ( n4438 & n25048 ) | ( n4438 & n25049 ) | ( n25048 & n25049 ) ;
  assign n25051 = ( ~n361 & n10149 ) | ( ~n361 & n25050 ) | ( n10149 & n25050 ) ;
  assign n25052 = ( n4152 & ~n15783 ) | ( n4152 & n22690 ) | ( ~n15783 & n22690 ) ;
  assign n25053 = n4605 ^ n4269 ^ n3106 ;
  assign n25054 = n14051 ^ n4321 ^ 1'b0 ;
  assign n25055 = ( n15395 & n25053 ) | ( n15395 & n25054 ) | ( n25053 & n25054 ) ;
  assign n25056 = ( n261 & n14717 ) | ( n261 & ~n25055 ) | ( n14717 & ~n25055 ) ;
  assign n25057 = ( ~n3031 & n13037 ) | ( ~n3031 & n24387 ) | ( n13037 & n24387 ) ;
  assign n25058 = ( n1494 & ~n9654 ) | ( n1494 & n20614 ) | ( ~n9654 & n20614 ) ;
  assign n25059 = ( n9684 & n19062 ) | ( n9684 & n25058 ) | ( n19062 & n25058 ) ;
  assign n25060 = n17609 ^ n6409 ^ n6111 ;
  assign n25061 = n25060 ^ n14842 ^ n13483 ;
  assign n25062 = ( n17154 & n25059 ) | ( n17154 & n25061 ) | ( n25059 & n25061 ) ;
  assign n25063 = n19059 ^ n3197 ^ n3020 ;
  assign n25064 = n17543 | n18347 ;
  assign n25065 = ( n6146 & n8621 ) | ( n6146 & ~n25064 ) | ( n8621 & ~n25064 ) ;
  assign n25066 = ( n3447 & n3885 ) | ( n3447 & n25065 ) | ( n3885 & n25065 ) ;
  assign n25067 = ( n3442 & ~n8070 ) | ( n3442 & n21534 ) | ( ~n8070 & n21534 ) ;
  assign n25068 = ( n2868 & n3529 ) | ( n2868 & n5049 ) | ( n3529 & n5049 ) ;
  assign n25069 = ( n4910 & n16094 ) | ( n4910 & n25068 ) | ( n16094 & n25068 ) ;
  assign n25070 = ( ~n3055 & n25067 ) | ( ~n3055 & n25069 ) | ( n25067 & n25069 ) ;
  assign n25071 = n12816 & n15055 ;
  assign n25072 = ~n13163 & n25071 ;
  assign n25073 = n19216 ^ n982 ^ 1'b0 ;
  assign n25074 = ( n3503 & n9491 ) | ( n3503 & n21391 ) | ( n9491 & n21391 ) ;
  assign n25075 = ( ~n180 & n2781 ) | ( ~n180 & n6407 ) | ( n2781 & n6407 ) ;
  assign n25076 = n22610 ^ n10496 ^ n9491 ;
  assign n25077 = n25076 ^ n9314 ^ n850 ;
  assign n25078 = ( n3720 & ~n25075 ) | ( n3720 & n25077 ) | ( ~n25075 & n25077 ) ;
  assign n25079 = n15294 ^ n4570 ^ n1726 ;
  assign n25080 = n25079 ^ n3379 ^ n3358 ;
  assign n25081 = n23384 ^ n19418 ^ n7325 ;
  assign n25082 = n16591 ^ n16223 ^ n5286 ;
  assign n25083 = ( n9451 & n15973 ) | ( n9451 & ~n25082 ) | ( n15973 & ~n25082 ) ;
  assign n25084 = ~n3247 & n7776 ;
  assign n25085 = n25084 ^ n14666 ^ 1'b0 ;
  assign n25086 = n15935 ^ n15647 ^ n3762 ;
  assign n25087 = n25086 ^ n16558 ^ n5619 ;
  assign n25088 = ( n11455 & n20699 ) | ( n11455 & n25087 ) | ( n20699 & n25087 ) ;
  assign n25089 = n16364 ^ n4922 ^ n2002 ;
  assign n25090 = ~n5497 & n18356 ;
  assign n25091 = n5998 & n25090 ;
  assign n25092 = ( n15358 & n25089 ) | ( n15358 & ~n25091 ) | ( n25089 & ~n25091 ) ;
  assign n25096 = n6310 ^ n5383 ^ n2481 ;
  assign n25095 = ( n13799 & n16594 ) | ( n13799 & n19931 ) | ( n16594 & n19931 ) ;
  assign n25093 = n16103 ^ n9204 ^ 1'b0 ;
  assign n25094 = n25093 ^ n8015 ^ 1'b0 ;
  assign n25097 = n25096 ^ n25095 ^ n25094 ;
  assign n25098 = n22756 ^ n3778 ^ x82 ;
  assign n25099 = ( ~n10887 & n11073 ) | ( ~n10887 & n18376 ) | ( n11073 & n18376 ) ;
  assign n25100 = n25099 ^ n18032 ^ n3565 ;
  assign n25102 = ( ~x13 & n6532 ) | ( ~x13 & n15579 ) | ( n6532 & n15579 ) ;
  assign n25101 = ( n17775 & n19168 ) | ( n17775 & ~n23415 ) | ( n19168 & ~n23415 ) ;
  assign n25103 = n25102 ^ n25101 ^ n4696 ;
  assign n25104 = n9682 ^ n2703 ^ 1'b0 ;
  assign n25105 = n25104 ^ n19318 ^ n8528 ;
  assign n25106 = ( n1841 & ~n13652 ) | ( n1841 & n18228 ) | ( ~n13652 & n18228 ) ;
  assign n25107 = ~n9059 & n25106 ;
  assign n25108 = n25107 ^ n5584 ^ 1'b0 ;
  assign n25109 = ~n1354 & n1586 ;
  assign n25110 = ~n3867 & n25109 ;
  assign n25111 = ~n13487 & n25110 ;
  assign n25112 = n14440 ^ x58 ^ 1'b0 ;
  assign n25113 = n25112 ^ n18221 ^ n14711 ;
  assign n25114 = ( n855 & ~n3033 ) | ( n855 & n25005 ) | ( ~n3033 & n25005 ) ;
  assign n25115 = ( n10649 & n10658 ) | ( n10649 & ~n20531 ) | ( n10658 & ~n20531 ) ;
  assign n25116 = ( ~n2686 & n12781 ) | ( ~n2686 & n25115 ) | ( n12781 & n25115 ) ;
  assign n25117 = ( n8478 & ~n8968 ) | ( n8478 & n25104 ) | ( ~n8968 & n25104 ) ;
  assign n25118 = n23458 ^ n19176 ^ n4082 ;
  assign n25119 = ( ~n7854 & n13305 ) | ( ~n7854 & n24290 ) | ( n13305 & n24290 ) ;
  assign n25120 = ( n13685 & n15282 ) | ( n13685 & ~n25119 ) | ( n15282 & ~n25119 ) ;
  assign n25121 = n7407 & n19863 ;
  assign n25122 = ~n13471 & n25121 ;
  assign n25123 = ( n9322 & ~n18045 ) | ( n9322 & n25122 ) | ( ~n18045 & n25122 ) ;
  assign n25124 = n18119 ^ n17210 ^ n15589 ;
  assign n25125 = n25124 ^ n8006 ^ 1'b0 ;
  assign n25126 = ~n1632 & n25125 ;
  assign n25127 = n18273 ^ n8220 ^ n3949 ;
  assign n25128 = n13754 ^ n6571 ^ 1'b0 ;
  assign n25129 = ( n547 & n2515 ) | ( n547 & n11470 ) | ( n2515 & n11470 ) ;
  assign n25130 = ( n3068 & ~n18227 ) | ( n3068 & n21292 ) | ( ~n18227 & n21292 ) ;
  assign n25131 = n4997 & n5788 ;
  assign n25132 = ~n386 & n25131 ;
  assign n25139 = ( n362 & n2935 ) | ( n362 & ~n7280 ) | ( n2935 & ~n7280 ) ;
  assign n25136 = n14918 ^ n3505 ^ 1'b0 ;
  assign n25137 = n6251 & n25136 ;
  assign n25133 = n5180 ^ n5172 ^ n5079 ;
  assign n25134 = n1255 & ~n25133 ;
  assign n25135 = n25134 ^ n16933 ^ n10131 ;
  assign n25138 = n25137 ^ n25135 ^ n3563 ;
  assign n25140 = n25139 ^ n25138 ^ n7494 ;
  assign n25141 = n19752 ^ n5894 ^ n1057 ;
  assign n25142 = ( n2569 & n23199 ) | ( n2569 & ~n25141 ) | ( n23199 & ~n25141 ) ;
  assign n25143 = ( ~n3301 & n14714 ) | ( ~n3301 & n18215 ) | ( n14714 & n18215 ) ;
  assign n25144 = ( n6593 & n13564 ) | ( n6593 & n24273 ) | ( n13564 & n24273 ) ;
  assign n25145 = n8877 ^ n3831 ^ n266 ;
  assign n25146 = n25145 ^ n9877 ^ n4437 ;
  assign n25147 = ( n5066 & n19223 ) | ( n5066 & n22713 ) | ( n19223 & n22713 ) ;
  assign n25149 = ( n4599 & n9706 ) | ( n4599 & ~n9836 ) | ( n9706 & ~n9836 ) ;
  assign n25148 = ~n2201 & n18399 ;
  assign n25150 = n25149 ^ n25148 ^ 1'b0 ;
  assign n25153 = ( n7133 & ~n10126 ) | ( n7133 & n20603 ) | ( ~n10126 & n20603 ) ;
  assign n25154 = n8798 ^ n7046 ^ n5059 ;
  assign n25155 = n25154 ^ n21565 ^ n9545 ;
  assign n25156 = ( n3233 & n25153 ) | ( n3233 & n25155 ) | ( n25153 & n25155 ) ;
  assign n25157 = n25156 ^ n5910 ^ n2432 ;
  assign n25151 = ( ~n1804 & n5213 ) | ( ~n1804 & n16673 ) | ( n5213 & n16673 ) ;
  assign n25152 = ( ~n1874 & n13395 ) | ( ~n1874 & n25151 ) | ( n13395 & n25151 ) ;
  assign n25158 = n25157 ^ n25152 ^ n12072 ;
  assign n25159 = n25158 ^ n15324 ^ n10890 ;
  assign n25160 = n25159 ^ n13681 ^ 1'b0 ;
  assign n25162 = n2791 | n12294 ;
  assign n25163 = n25162 ^ n14396 ^ 1'b0 ;
  assign n25161 = n9342 ^ n8744 ^ n3907 ;
  assign n25164 = n25163 ^ n25161 ^ n5783 ;
  assign n25165 = n22703 ^ n21170 ^ n13362 ;
  assign n25166 = ( n16880 & n25164 ) | ( n16880 & ~n25165 ) | ( n25164 & ~n25165 ) ;
  assign n25167 = n14993 ^ n5840 ^ n5349 ;
  assign n25168 = ( n4317 & ~n16299 ) | ( n4317 & n21473 ) | ( ~n16299 & n21473 ) ;
  assign n25169 = ( n9956 & ~n10196 ) | ( n9956 & n16563 ) | ( ~n10196 & n16563 ) ;
  assign n25170 = n8572 | n25169 ;
  assign n25171 = n8720 & ~n25170 ;
  assign n25172 = n25171 ^ n19376 ^ n6798 ;
  assign n25173 = n13601 ^ n5524 ^ n3623 ;
  assign n25174 = ( n4172 & ~n16019 ) | ( n4172 & n25173 ) | ( ~n16019 & n25173 ) ;
  assign n25175 = n23620 ^ n19445 ^ 1'b0 ;
  assign n25176 = n5556 ^ n4342 ^ 1'b0 ;
  assign n25177 = n11447 ^ n3975 ^ n575 ;
  assign n25178 = n25177 ^ n3553 ^ n1198 ;
  assign n25179 = ( n14175 & n15240 ) | ( n14175 & n23346 ) | ( n15240 & n23346 ) ;
  assign n25180 = n18078 ^ n11175 ^ n7028 ;
  assign n25181 = n2592 ^ n1662 ^ 1'b0 ;
  assign n25182 = ~n2113 & n25181 ;
  assign n25183 = n25182 ^ n17985 ^ n8470 ;
  assign n25184 = ( n20834 & ~n22334 ) | ( n20834 & n25183 ) | ( ~n22334 & n25183 ) ;
  assign n25185 = n23907 ^ n7883 ^ n588 ;
  assign n25186 = ~n6850 & n17791 ;
  assign n25187 = ~n14841 & n25186 ;
  assign n25188 = ( n2437 & n25185 ) | ( n2437 & ~n25187 ) | ( n25185 & ~n25187 ) ;
  assign n25189 = ( n659 & ~n7817 ) | ( n659 & n12224 ) | ( ~n7817 & n12224 ) ;
  assign n25190 = n19037 ^ n3624 ^ n3031 ;
  assign n25191 = n25190 ^ n20491 ^ n12909 ;
  assign n25192 = n25191 ^ n9269 ^ 1'b0 ;
  assign n25193 = n25189 & ~n25192 ;
  assign n25194 = ( n5936 & n11644 ) | ( n5936 & n20523 ) | ( n11644 & n20523 ) ;
  assign n25195 = n10787 ^ n10042 ^ 1'b0 ;
  assign n25196 = n10703 ^ n8060 ^ n1673 ;
  assign n25200 = n22104 ^ n2708 ^ 1'b0 ;
  assign n25197 = n12631 ^ n2173 ^ n571 ;
  assign n25198 = n25197 ^ n23175 ^ n21759 ;
  assign n25199 = ( n3068 & n15343 ) | ( n3068 & n25198 ) | ( n15343 & n25198 ) ;
  assign n25201 = n25200 ^ n25199 ^ n6705 ;
  assign n25202 = ( n4043 & n18383 ) | ( n4043 & n18565 ) | ( n18383 & n18565 ) ;
  assign n25203 = n25202 ^ n18405 ^ n12053 ;
  assign n25204 = n25203 ^ n5137 ^ n3134 ;
  assign n25205 = n3213 ^ n3052 ^ 1'b0 ;
  assign n25206 = n2967 | n25205 ;
  assign n25207 = ( ~n3644 & n5428 ) | ( ~n3644 & n8271 ) | ( n5428 & n8271 ) ;
  assign n25208 = n14904 ^ n11683 ^ n8813 ;
  assign n25209 = n16260 & n25208 ;
  assign n25213 = ( n11268 & n17578 ) | ( n11268 & n19876 ) | ( n17578 & n19876 ) ;
  assign n25210 = ( ~n7686 & n11733 ) | ( ~n7686 & n22459 ) | ( n11733 & n22459 ) ;
  assign n25211 = n25210 ^ n6536 ^ n2986 ;
  assign n25212 = n25211 ^ n12700 ^ n7282 ;
  assign n25214 = n25213 ^ n25212 ^ n9265 ;
  assign n25215 = n22620 ^ n692 ^ 1'b0 ;
  assign n25216 = ( n1724 & ~n3672 ) | ( n1724 & n10216 ) | ( ~n3672 & n10216 ) ;
  assign n25217 = n25216 ^ n5916 ^ n1835 ;
  assign n25218 = ( ~n7278 & n25215 ) | ( ~n7278 & n25217 ) | ( n25215 & n25217 ) ;
  assign n25219 = ( n3556 & ~n17552 ) | ( n3556 & n18541 ) | ( ~n17552 & n18541 ) ;
  assign n25220 = n21819 ^ n3104 ^ x25 ;
  assign n25221 = n23545 ^ n7954 ^ n7842 ;
  assign n25222 = ( n13444 & ~n14734 ) | ( n13444 & n25221 ) | ( ~n14734 & n25221 ) ;
  assign n25223 = n25222 ^ n13544 ^ 1'b0 ;
  assign n25224 = ( n1118 & n6256 ) | ( n1118 & ~n20552 ) | ( n6256 & ~n20552 ) ;
  assign n25225 = ~n6349 & n9283 ;
  assign n25226 = n25224 & n25225 ;
  assign n25227 = ( n4472 & n5253 ) | ( n4472 & n10506 ) | ( n5253 & n10506 ) ;
  assign n25228 = n25227 ^ n3992 ^ 1'b0 ;
  assign n25229 = ( n11565 & n22760 ) | ( n11565 & ~n25228 ) | ( n22760 & ~n25228 ) ;
  assign n25230 = ( n25223 & n25226 ) | ( n25223 & ~n25229 ) | ( n25226 & ~n25229 ) ;
  assign n25231 = n25230 ^ n15663 ^ n15133 ;
  assign n25233 = n8671 ^ n7606 ^ n5535 ;
  assign n25232 = n8825 | n11249 ;
  assign n25234 = n25233 ^ n25232 ^ 1'b0 ;
  assign n25235 = n25234 ^ n7400 ^ n6460 ;
  assign n25236 = n11609 & n18912 ;
  assign n25237 = n25236 ^ n18793 ^ n12178 ;
  assign n25238 = n8302 ^ n8297 ^ n1968 ;
  assign n25239 = x82 & n16404 ;
  assign n25240 = n8255 & n25239 ;
  assign n25241 = n20700 ^ n11908 ^ n2378 ;
  assign n25242 = ( n5427 & n25240 ) | ( n5427 & ~n25241 ) | ( n25240 & ~n25241 ) ;
  assign n25244 = n11761 ^ n7262 ^ n2941 ;
  assign n25245 = ( n13252 & n18172 ) | ( n13252 & ~n25244 ) | ( n18172 & ~n25244 ) ;
  assign n25243 = ( n9717 & n14075 ) | ( n9717 & n17029 ) | ( n14075 & n17029 ) ;
  assign n25246 = n25245 ^ n25243 ^ n15841 ;
  assign n25247 = n25246 ^ n7688 ^ n5701 ;
  assign n25249 = ( ~n1789 & n1820 ) | ( ~n1789 & n9488 ) | ( n1820 & n9488 ) ;
  assign n25248 = ( n7341 & n7477 ) | ( n7341 & ~n16385 ) | ( n7477 & ~n16385 ) ;
  assign n25250 = n25249 ^ n25248 ^ n12634 ;
  assign n25252 = n25152 ^ n22493 ^ x17 ;
  assign n25251 = n3536 & n4802 ;
  assign n25253 = n25252 ^ n25251 ^ 1'b0 ;
  assign n25254 = n23431 ^ n11590 ^ 1'b0 ;
  assign n25255 = ~n8272 & n25254 ;
  assign n25256 = n7597 & n25255 ;
  assign n25257 = n25256 ^ n2669 ^ 1'b0 ;
  assign n25258 = ( ~n16499 & n19174 ) | ( ~n16499 & n25257 ) | ( n19174 & n25257 ) ;
  assign n25259 = n24975 ^ n9178 ^ 1'b0 ;
  assign n25260 = ( n1570 & ~n17914 ) | ( n1570 & n25259 ) | ( ~n17914 & n25259 ) ;
  assign n25261 = n19455 ^ n16725 ^ n15877 ;
  assign n25262 = n25261 ^ n17938 ^ n16101 ;
  assign n25263 = ( ~n1633 & n6704 ) | ( ~n1633 & n12097 ) | ( n6704 & n12097 ) ;
  assign n25264 = n25263 ^ n20425 ^ n5851 ;
  assign n25266 = n5296 ^ n4250 ^ n1549 ;
  assign n25265 = n4882 ^ n1780 ^ n945 ;
  assign n25267 = n25266 ^ n25265 ^ n572 ;
  assign n25268 = ( x86 & n2045 ) | ( x86 & ~n6404 ) | ( n2045 & ~n6404 ) ;
  assign n25269 = n25268 ^ n23185 ^ n5384 ;
  assign n25270 = ( ~n19271 & n20692 ) | ( ~n19271 & n25104 ) | ( n20692 & n25104 ) ;
  assign n25271 = n10432 ^ n8223 ^ 1'b0 ;
  assign n25272 = n11343 & n25271 ;
  assign n25274 = ( ~n7365 & n10360 ) | ( ~n7365 & n11503 ) | ( n10360 & n11503 ) ;
  assign n25275 = n25274 ^ n22557 ^ n11230 ;
  assign n25273 = n22676 ^ n21258 ^ n7194 ;
  assign n25276 = n25275 ^ n25273 ^ n14931 ;
  assign n25277 = n8727 ^ n4161 ^ n1598 ;
  assign n25278 = n4857 & ~n25277 ;
  assign n25279 = n25276 & n25278 ;
  assign n25280 = n9720 ^ n7206 ^ n3752 ;
  assign n25281 = n22005 ^ n7224 ^ n2873 ;
  assign n25282 = n21584 ^ n10344 ^ 1'b0 ;
  assign n25284 = n22812 ^ n17542 ^ n994 ;
  assign n25283 = ( n6041 & ~n6125 ) | ( n6041 & n20034 ) | ( ~n6125 & n20034 ) ;
  assign n25285 = n25284 ^ n25283 ^ n25215 ;
  assign n25286 = n7488 ^ n4346 ^ n1068 ;
  assign n25287 = n25286 ^ n19174 ^ n7362 ;
  assign n25288 = n6809 ^ n1639 ^ 1'b0 ;
  assign n25289 = n8294 | n25288 ;
  assign n25290 = n11578 ^ n8168 ^ n687 ;
  assign n25291 = n25290 ^ n7136 ^ n5242 ;
  assign n25292 = n25291 ^ n20499 ^ n16436 ;
  assign n25293 = ( n25287 & n25289 ) | ( n25287 & ~n25292 ) | ( n25289 & ~n25292 ) ;
  assign n25295 = n20760 ^ n11573 ^ n1201 ;
  assign n25294 = n22493 ^ n20218 ^ n13958 ;
  assign n25296 = n25295 ^ n25294 ^ n12143 ;
  assign n25297 = ( ~n10990 & n16070 ) | ( ~n10990 & n25296 ) | ( n16070 & n25296 ) ;
  assign n25298 = n25297 ^ n10673 ^ n7377 ;
  assign n25299 = ( n1629 & ~n7403 ) | ( n1629 & n7671 ) | ( ~n7403 & n7671 ) ;
  assign n25300 = ( n2203 & n5579 ) | ( n2203 & ~n8119 ) | ( n5579 & ~n8119 ) ;
  assign n25301 = n25300 ^ n11462 ^ 1'b0 ;
  assign n25302 = ( n10982 & n20289 ) | ( n10982 & n22343 ) | ( n20289 & n22343 ) ;
  assign n25303 = n25302 ^ n3011 ^ 1'b0 ;
  assign n25307 = n21574 ^ n15092 ^ n10561 ;
  assign n25304 = n19460 ^ n6899 ^ n577 ;
  assign n25305 = ( ~n7513 & n15843 ) | ( ~n7513 & n25304 ) | ( n15843 & n25304 ) ;
  assign n25306 = n550 | n25305 ;
  assign n25308 = n25307 ^ n25306 ^ 1'b0 ;
  assign n25309 = n20005 ^ n19820 ^ n1988 ;
  assign n25310 = n8099 & ~n21950 ;
  assign n25311 = n19969 ^ n14997 ^ n1080 ;
  assign n25312 = n9714 ^ n6794 ^ n4602 ;
  assign n25313 = ( n4137 & n6660 ) | ( n4137 & n9892 ) | ( n6660 & n9892 ) ;
  assign n25314 = n25313 ^ n4273 ^ x125 ;
  assign n25321 = ( n973 & ~n4486 ) | ( n973 & n8178 ) | ( ~n4486 & n8178 ) ;
  assign n25320 = ( ~n1981 & n2658 ) | ( ~n1981 & n12190 ) | ( n2658 & n12190 ) ;
  assign n25322 = n25321 ^ n25320 ^ n22437 ;
  assign n25319 = n25134 ^ n13674 ^ n13080 ;
  assign n25315 = n2198 & n7850 ;
  assign n25316 = n7477 & n25315 ;
  assign n25317 = ~n7248 & n8802 ;
  assign n25318 = n25316 & n25317 ;
  assign n25323 = n25322 ^ n25319 ^ n25318 ;
  assign n25324 = n24212 ^ n9333 ^ 1'b0 ;
  assign n25325 = n15295 ^ n14011 ^ 1'b0 ;
  assign n25326 = ( n2732 & ~n10328 ) | ( n2732 & n24461 ) | ( ~n10328 & n24461 ) ;
  assign n25327 = ( ~n6219 & n10686 ) | ( ~n6219 & n24041 ) | ( n10686 & n24041 ) ;
  assign n25328 = n18725 ^ n13520 ^ n1130 ;
  assign n25329 = ( n14654 & n25327 ) | ( n14654 & ~n25328 ) | ( n25327 & ~n25328 ) ;
  assign n25330 = n1571 | n5123 ;
  assign n25331 = n14248 & ~n25330 ;
  assign n25332 = n25331 ^ n22375 ^ 1'b0 ;
  assign n25333 = n4714 & ~n25332 ;
  assign n25334 = ( n8768 & ~n24580 ) | ( n8768 & n25333 ) | ( ~n24580 & n25333 ) ;
  assign n25335 = ( n1745 & ~n12932 ) | ( n1745 & n25334 ) | ( ~n12932 & n25334 ) ;
  assign n25336 = ( n6121 & n10126 ) | ( n6121 & n17222 ) | ( n10126 & n17222 ) ;
  assign n25337 = ( n8509 & ~n11805 ) | ( n8509 & n25336 ) | ( ~n11805 & n25336 ) ;
  assign n25338 = ~n11229 & n11560 ;
  assign n25339 = n5113 & ~n8297 ;
  assign n25340 = n25339 ^ n22400 ^ n172 ;
  assign n25341 = ( n2654 & ~n6547 ) | ( n2654 & n9168 ) | ( ~n6547 & n9168 ) ;
  assign n25342 = ( ~n1733 & n10080 ) | ( ~n1733 & n25341 ) | ( n10080 & n25341 ) ;
  assign n25343 = ( n10576 & ~n13622 ) | ( n10576 & n25342 ) | ( ~n13622 & n25342 ) ;
  assign n25344 = ( n4905 & n14773 ) | ( n4905 & ~n21017 ) | ( n14773 & ~n21017 ) ;
  assign n25345 = n25344 ^ n2170 ^ n915 ;
  assign n25346 = n12648 ^ n4183 ^ n3822 ;
  assign n25347 = n25346 ^ n18791 ^ n13037 ;
  assign n25348 = n23149 ^ n20467 ^ n8664 ;
  assign n25349 = ( n1434 & n9554 ) | ( n1434 & n17797 ) | ( n9554 & n17797 ) ;
  assign n25350 = ( n12051 & ~n12238 ) | ( n12051 & n15552 ) | ( ~n12238 & n15552 ) ;
  assign n25351 = ( n9715 & n25349 ) | ( n9715 & n25350 ) | ( n25349 & n25350 ) ;
  assign n25352 = n2945 & n9487 ;
  assign n25353 = n25352 ^ n6959 ^ 1'b0 ;
  assign n25354 = n25353 ^ n13528 ^ 1'b0 ;
  assign n25355 = ( ~n11835 & n25173 ) | ( ~n11835 & n25354 ) | ( n25173 & n25354 ) ;
  assign n25356 = ( n11356 & n20120 ) | ( n11356 & ~n25355 ) | ( n20120 & ~n25355 ) ;
  assign n25357 = ( n11559 & ~n13603 ) | ( n11559 & n25356 ) | ( ~n13603 & n25356 ) ;
  assign n25358 = ( n2253 & ~n6551 ) | ( n2253 & n11583 ) | ( ~n6551 & n11583 ) ;
  assign n25359 = n21639 ^ n3335 ^ 1'b0 ;
  assign n25360 = n25358 & ~n25359 ;
  assign n25361 = ( ~n6053 & n20877 ) | ( ~n6053 & n25344 ) | ( n20877 & n25344 ) ;
  assign n25362 = n4948 ^ n4141 ^ 1'b0 ;
  assign n25363 = ( n3817 & n11682 ) | ( n3817 & n17206 ) | ( n11682 & n17206 ) ;
  assign n25364 = ( n3973 & n12730 ) | ( n3973 & ~n25363 ) | ( n12730 & ~n25363 ) ;
  assign n25365 = n24278 ^ n463 ^ 1'b0 ;
  assign n25366 = n23804 | n25365 ;
  assign n25367 = ( n25362 & n25364 ) | ( n25362 & ~n25366 ) | ( n25364 & ~n25366 ) ;
  assign n25368 = ( n15876 & n21221 ) | ( n15876 & n25367 ) | ( n21221 & n25367 ) ;
  assign n25369 = ( n498 & n11060 ) | ( n498 & n22658 ) | ( n11060 & n22658 ) ;
  assign n25370 = n15894 ^ n10114 ^ n1341 ;
  assign n25371 = n19641 ^ n11187 ^ n3099 ;
  assign n25372 = ( ~n1293 & n25370 ) | ( ~n1293 & n25371 ) | ( n25370 & n25371 ) ;
  assign n25373 = ( ~n10672 & n25369 ) | ( ~n10672 & n25372 ) | ( n25369 & n25372 ) ;
  assign n25374 = n23740 ^ n13751 ^ n7685 ;
  assign n25375 = ( n3081 & ~n3536 ) | ( n3081 & n22082 ) | ( ~n3536 & n22082 ) ;
  assign n25376 = ( n12747 & ~n16804 ) | ( n12747 & n25375 ) | ( ~n16804 & n25375 ) ;
  assign n25377 = n25376 ^ n16625 ^ 1'b0 ;
  assign n25378 = ~n9643 & n18114 ;
  assign n25379 = n10026 & ~n16095 ;
  assign n25380 = ~n11570 & n25379 ;
  assign n25381 = n17587 ^ n10465 ^ n7485 ;
  assign n25382 = ( ~n5728 & n10991 ) | ( ~n5728 & n23603 ) | ( n10991 & n23603 ) ;
  assign n25383 = ( n6098 & ~n20419 ) | ( n6098 & n25382 ) | ( ~n20419 & n25382 ) ;
  assign n25384 = ( ~n16634 & n17169 ) | ( ~n16634 & n25383 ) | ( n17169 & n25383 ) ;
  assign n25385 = n25384 ^ n19793 ^ n18859 ;
  assign n25386 = ( ~n10393 & n25381 ) | ( ~n10393 & n25385 ) | ( n25381 & n25385 ) ;
  assign n25387 = n7392 ^ n2825 ^ n1330 ;
  assign n25388 = n25387 ^ n17668 ^ n15354 ;
  assign n25389 = n25388 ^ n9375 ^ n225 ;
  assign n25390 = ( ~n3184 & n11581 ) | ( ~n3184 & n18714 ) | ( n11581 & n18714 ) ;
  assign n25391 = n25390 ^ n12155 ^ 1'b0 ;
  assign n25392 = ( n778 & n1384 ) | ( n778 & n25391 ) | ( n1384 & n25391 ) ;
  assign n25393 = n2767 & ~n6968 ;
  assign n25394 = n17685 & n25393 ;
  assign n25395 = ( n7753 & n20102 ) | ( n7753 & n25394 ) | ( n20102 & n25394 ) ;
  assign n25399 = n13600 ^ n4488 ^ n819 ;
  assign n25400 = n25399 ^ n9608 ^ 1'b0 ;
  assign n25401 = ~n2929 & n25400 ;
  assign n25397 = ( n917 & ~n2287 ) | ( n917 & n2674 ) | ( ~n2287 & n2674 ) ;
  assign n25398 = n22859 & ~n25397 ;
  assign n25396 = n19488 ^ n17135 ^ n7081 ;
  assign n25402 = n25401 ^ n25398 ^ n25396 ;
  assign n25403 = n25402 ^ n10761 ^ n3373 ;
  assign n25404 = ( n8865 & n17275 ) | ( n8865 & n25403 ) | ( n17275 & n25403 ) ;
  assign n25405 = n14165 ^ n8110 ^ x107 ;
  assign n25406 = n25405 ^ n1417 ^ 1'b0 ;
  assign n25410 = n16586 ^ n14334 ^ n13314 ;
  assign n25407 = ( n380 & n1771 ) | ( n380 & ~n3835 ) | ( n1771 & ~n3835 ) ;
  assign n25408 = ( ~n1334 & n6806 ) | ( ~n1334 & n25407 ) | ( n6806 & n25407 ) ;
  assign n25409 = ( n1399 & ~n9652 ) | ( n1399 & n25408 ) | ( ~n9652 & n25408 ) ;
  assign n25411 = n25410 ^ n25409 ^ n14558 ;
  assign n25412 = n19339 ^ n14414 ^ n4230 ;
  assign n25413 = n25412 ^ n24040 ^ n7336 ;
  assign n25414 = ( ~n4415 & n6281 ) | ( ~n4415 & n24921 ) | ( n6281 & n24921 ) ;
  assign n25415 = n9654 & n13799 ;
  assign n25416 = n25414 & n25415 ;
  assign n25417 = n21326 ^ n7686 ^ n6136 ;
  assign n25418 = n25417 ^ n9348 ^ 1'b0 ;
  assign n25419 = n991 & ~n25418 ;
  assign n25420 = ( x117 & n11555 ) | ( x117 & n17940 ) | ( n11555 & n17940 ) ;
  assign n25421 = ( n19417 & ~n24837 ) | ( n19417 & n25420 ) | ( ~n24837 & n25420 ) ;
  assign n25422 = n25421 ^ n24238 ^ 1'b0 ;
  assign n25429 = x38 | n4423 ;
  assign n25423 = n6872 ^ n2928 ^ n1121 ;
  assign n25424 = n2309 | n4983 ;
  assign n25425 = n6812 & ~n25424 ;
  assign n25426 = n25425 ^ n8230 ^ 1'b0 ;
  assign n25427 = ( n6300 & n25423 ) | ( n6300 & ~n25426 ) | ( n25423 & ~n25426 ) ;
  assign n25428 = n25427 ^ n20939 ^ 1'b0 ;
  assign n25430 = n25429 ^ n25428 ^ n25268 ;
  assign n25431 = ( n1569 & ~n12128 ) | ( n1569 & n14304 ) | ( ~n12128 & n14304 ) ;
  assign n25432 = ( n4158 & n4514 ) | ( n4158 & n12779 ) | ( n4514 & n12779 ) ;
  assign n25433 = ( n14347 & ~n15524 ) | ( n14347 & n22347 ) | ( ~n15524 & n22347 ) ;
  assign n25434 = ( n409 & n2983 ) | ( n409 & n14022 ) | ( n2983 & n14022 ) ;
  assign n25435 = ( ~n1750 & n11869 ) | ( ~n1750 & n14450 ) | ( n11869 & n14450 ) ;
  assign n25436 = ( n22176 & n25434 ) | ( n22176 & ~n25435 ) | ( n25434 & ~n25435 ) ;
  assign n25437 = ( ~n10310 & n11309 ) | ( ~n10310 & n11349 ) | ( n11309 & n11349 ) ;
  assign n25438 = ( n2902 & ~n14832 ) | ( n2902 & n25437 ) | ( ~n14832 & n25437 ) ;
  assign n25439 = n1023 & ~n25438 ;
  assign n25440 = ~n22460 & n25439 ;
  assign n25441 = n6964 & n14321 ;
  assign n25442 = n10222 ^ n7755 ^ 1'b0 ;
  assign n25443 = n991 & n25442 ;
  assign n25444 = n25443 ^ n4571 ^ 1'b0 ;
  assign n25445 = n5228 & n25444 ;
  assign n25446 = ( n4038 & ~n8716 ) | ( n4038 & n25445 ) | ( ~n8716 & n25445 ) ;
  assign n25447 = n25210 ^ n23421 ^ n15719 ;
  assign n25448 = n3020 & n6034 ;
  assign n25449 = ~n1933 & n22201 ;
  assign n25450 = ( ~n4916 & n25448 ) | ( ~n4916 & n25449 ) | ( n25448 & n25449 ) ;
  assign n25451 = n20517 ^ n20033 ^ 1'b0 ;
  assign n25452 = n11288 & ~n17723 ;
  assign n25453 = n25451 & n25452 ;
  assign n25454 = n19226 ^ n18269 ^ n12388 ;
  assign n25455 = n10811 ^ n5703 ^ n2509 ;
  assign n25456 = ( n2947 & n13531 ) | ( n2947 & ~n25455 ) | ( n13531 & ~n25455 ) ;
  assign n25457 = ( ~n8626 & n20162 ) | ( ~n8626 & n25456 ) | ( n20162 & n25456 ) ;
  assign n25458 = n5224 ^ n1075 ^ 1'b0 ;
  assign n25459 = ( n10538 & ~n11749 ) | ( n10538 & n22043 ) | ( ~n11749 & n22043 ) ;
  assign n25460 = n16515 ^ n11970 ^ n9745 ;
  assign n25461 = ( ~n13600 & n14828 ) | ( ~n13600 & n25460 ) | ( n14828 & n25460 ) ;
  assign n25462 = n9471 ^ n6959 ^ n426 ;
  assign n25463 = n4926 & n5228 ;
  assign n25464 = n25462 & n25463 ;
  assign n25465 = ( n19198 & ~n21797 ) | ( n19198 & n25464 ) | ( ~n21797 & n25464 ) ;
  assign n25466 = ~n1065 & n2197 ;
  assign n25467 = n25466 ^ n20081 ^ 1'b0 ;
  assign n25472 = n20955 ^ n15757 ^ n13546 ;
  assign n25468 = n21190 ^ n14041 ^ n6427 ;
  assign n25469 = n25468 ^ n19947 ^ n10474 ;
  assign n25470 = n25469 ^ n11674 ^ n2417 ;
  assign n25471 = n16388 | n25470 ;
  assign n25473 = n25472 ^ n25471 ^ 1'b0 ;
  assign n25474 = n23128 ^ n9804 ^ n1869 ;
  assign n25475 = n25474 ^ n11293 ^ n4697 ;
  assign n25476 = n7763 & n17540 ;
  assign n25477 = ~n24505 & n25476 ;
  assign n25478 = n25477 ^ n7019 ^ 1'b0 ;
  assign n25479 = ~n25475 & n25478 ;
  assign n25480 = ~n7609 & n11723 ;
  assign n25481 = n25480 ^ n22528 ^ 1'b0 ;
  assign n25482 = ( n12387 & n13324 ) | ( n12387 & ~n25481 ) | ( n13324 & ~n25481 ) ;
  assign n25483 = ( n1730 & ~n18793 ) | ( n1730 & n24493 ) | ( ~n18793 & n24493 ) ;
  assign n25484 = ( n923 & n9173 ) | ( n923 & ~n21039 ) | ( n9173 & ~n21039 ) ;
  assign n25485 = ( n17493 & n21585 ) | ( n17493 & ~n23012 ) | ( n21585 & ~n23012 ) ;
  assign n25486 = n14530 ^ n10223 ^ n2243 ;
  assign n25487 = ( n9005 & n9337 ) | ( n9005 & n25486 ) | ( n9337 & n25486 ) ;
  assign n25488 = n23114 ^ n18894 ^ n896 ;
  assign n25489 = n5281 ^ n4613 ^ n3280 ;
  assign n25490 = ( n13825 & n24308 ) | ( n13825 & ~n25489 ) | ( n24308 & ~n25489 ) ;
  assign n25491 = ( n2456 & n11688 ) | ( n2456 & n21621 ) | ( n11688 & n21621 ) ;
  assign n25492 = ( n5807 & ~n25490 ) | ( n5807 & n25491 ) | ( ~n25490 & n25491 ) ;
  assign n25493 = ( ~n2849 & n12302 ) | ( ~n2849 & n25492 ) | ( n12302 & n25492 ) ;
  assign n25494 = n25493 ^ n16805 ^ n6083 ;
  assign n25495 = ( n21663 & n25096 ) | ( n21663 & ~n25494 ) | ( n25096 & ~n25494 ) ;
  assign n25498 = n3946 ^ n2388 ^ 1'b0 ;
  assign n25499 = ~n1477 & n25498 ;
  assign n25496 = ( n5059 & n12546 ) | ( n5059 & n18481 ) | ( n12546 & n18481 ) ;
  assign n25497 = n25496 ^ n18499 ^ n15875 ;
  assign n25500 = n25499 ^ n25497 ^ n2012 ;
  assign n25501 = n19354 ^ n14183 ^ n11958 ;
  assign n25502 = ( n4949 & n15008 ) | ( n4949 & ~n18026 ) | ( n15008 & ~n18026 ) ;
  assign n25503 = ( n19695 & n21545 ) | ( n19695 & n25502 ) | ( n21545 & n25502 ) ;
  assign n25509 = ( ~n845 & n12371 ) | ( ~n845 & n16368 ) | ( n12371 & n16368 ) ;
  assign n25508 = n5229 & ~n14435 ;
  assign n25510 = n25509 ^ n25508 ^ 1'b0 ;
  assign n25504 = ( ~n1954 & n3739 ) | ( ~n1954 & n9533 ) | ( n3739 & n9533 ) ;
  assign n25505 = n12091 | n25504 ;
  assign n25506 = n1199 & ~n25505 ;
  assign n25507 = ( n6501 & n22421 ) | ( n6501 & ~n25506 ) | ( n22421 & ~n25506 ) ;
  assign n25511 = n25510 ^ n25507 ^ n16002 ;
  assign n25512 = n25511 ^ n19645 ^ n2458 ;
  assign n25513 = n21574 ^ n8555 ^ n4887 ;
  assign n25514 = n25513 ^ n22164 ^ n12501 ;
  assign n25515 = n25514 ^ n14333 ^ n13307 ;
  assign n25516 = ( n7183 & n19519 ) | ( n7183 & n22827 ) | ( n19519 & n22827 ) ;
  assign n25517 = n25516 ^ n2045 ^ 1'b0 ;
  assign n25518 = ( n3192 & ~n9956 ) | ( n3192 & n13023 ) | ( ~n9956 & n13023 ) ;
  assign n25519 = ( n4775 & n16301 ) | ( n4775 & n25518 ) | ( n16301 & n25518 ) ;
  assign n25520 = n22376 & n25519 ;
  assign n25521 = n25520 ^ n24014 ^ n9658 ;
  assign n25522 = n12252 ^ n4628 ^ n2638 ;
  assign n25523 = n25522 ^ n24455 ^ n2142 ;
  assign n25525 = n22061 ^ n6208 ^ n4181 ;
  assign n25524 = n20444 ^ n9230 ^ n985 ;
  assign n25526 = n25525 ^ n25524 ^ n8096 ;
  assign n25527 = n12414 ^ n8345 ^ n7325 ;
  assign n25528 = n12189 ^ n10590 ^ n465 ;
  assign n25529 = n25528 ^ n5201 ^ n5012 ;
  assign n25530 = ( n21075 & n25527 ) | ( n21075 & ~n25529 ) | ( n25527 & ~n25529 ) ;
  assign n25531 = ( ~n339 & n20793 ) | ( ~n339 & n24410 ) | ( n20793 & n24410 ) ;
  assign n25532 = n9716 ^ n3339 ^ n3257 ;
  assign n25533 = n25532 ^ n22632 ^ 1'b0 ;
  assign n25534 = n1485 & n25533 ;
  assign n25535 = ( n5049 & ~n6470 ) | ( n5049 & n9381 ) | ( ~n6470 & n9381 ) ;
  assign n25536 = ( n3548 & n4622 ) | ( n3548 & ~n25535 ) | ( n4622 & ~n25535 ) ;
  assign n25537 = n25536 ^ n15705 ^ 1'b0 ;
  assign n25538 = ( n7355 & n12137 ) | ( n7355 & ~n22577 ) | ( n12137 & ~n22577 ) ;
  assign n25539 = n6582 ^ n2285 ^ n1625 ;
  assign n25540 = n25539 ^ n23809 ^ n7539 ;
  assign n25541 = ( n10747 & ~n25538 ) | ( n10747 & n25540 ) | ( ~n25538 & n25540 ) ;
  assign n25542 = ( n2188 & n4944 ) | ( n2188 & n15838 ) | ( n4944 & n15838 ) ;
  assign n25543 = n8981 ^ n5288 ^ n4068 ;
  assign n25544 = n25543 ^ n19180 ^ n10492 ;
  assign n25545 = ( n4015 & ~n25542 ) | ( n4015 & n25544 ) | ( ~n25542 & n25544 ) ;
  assign n25546 = ( n3800 & n13947 ) | ( n3800 & ~n20552 ) | ( n13947 & ~n20552 ) ;
  assign n25547 = n25546 ^ n6774 ^ n6237 ;
  assign n25548 = ( n2437 & ~n18017 ) | ( n2437 & n25547 ) | ( ~n18017 & n25547 ) ;
  assign n25549 = ( n11969 & n22220 ) | ( n11969 & ~n23084 ) | ( n22220 & ~n23084 ) ;
  assign n25550 = ( n2101 & ~n12192 ) | ( n2101 & n24374 ) | ( ~n12192 & n24374 ) ;
  assign n25551 = n18280 ^ n13541 ^ n7308 ;
  assign n25554 = n13089 ^ n1068 ^ n161 ;
  assign n25552 = n7347 | n10403 ;
  assign n25553 = n4794 & ~n25552 ;
  assign n25555 = n25554 ^ n25553 ^ n13410 ;
  assign n25556 = n1454 & ~n16621 ;
  assign n25557 = n2387 & n25556 ;
  assign n25558 = n25557 ^ n5234 ^ 1'b0 ;
  assign n25559 = n2195 & ~n25558 ;
  assign n25560 = ( n2100 & ~n15853 ) | ( n2100 & n19731 ) | ( ~n15853 & n19731 ) ;
  assign n25561 = n24050 ^ n9813 ^ n1905 ;
  assign n25562 = n15514 ^ n13082 ^ 1'b0 ;
  assign n25568 = n5658 ^ n882 ^ 1'b0 ;
  assign n25569 = n25568 ^ n22640 ^ n21828 ;
  assign n25566 = ( n2453 & n12402 ) | ( n2453 & ~n16198 ) | ( n12402 & ~n16198 ) ;
  assign n25563 = n4076 ^ n2437 ^ n955 ;
  assign n25564 = n6394 & ~n25563 ;
  assign n25565 = ( n5990 & n17661 ) | ( n5990 & ~n25564 ) | ( n17661 & ~n25564 ) ;
  assign n25567 = n25566 ^ n25565 ^ n5372 ;
  assign n25570 = n25569 ^ n25567 ^ n4004 ;
  assign n25573 = n23406 ^ n17745 ^ n2991 ;
  assign n25571 = n5740 ^ n1722 ^ n1525 ;
  assign n25572 = n4108 & ~n25571 ;
  assign n25574 = n25573 ^ n25572 ^ n14714 ;
  assign n25575 = n21156 ^ n16486 ^ n3272 ;
  assign n25576 = n1747 | n11841 ;
  assign n25577 = n25575 | n25576 ;
  assign n25578 = ( ~n399 & n12739 ) | ( ~n399 & n12954 ) | ( n12739 & n12954 ) ;
  assign n25579 = ( ~n2274 & n8333 ) | ( ~n2274 & n14216 ) | ( n8333 & n14216 ) ;
  assign n25580 = ( n2265 & n5024 ) | ( n2265 & n8033 ) | ( n5024 & n8033 ) ;
  assign n25581 = ( n7332 & ~n13428 ) | ( n7332 & n25580 ) | ( ~n13428 & n25580 ) ;
  assign n25582 = ( ~n717 & n14306 ) | ( ~n717 & n25581 ) | ( n14306 & n25581 ) ;
  assign n25583 = ( n10103 & n25579 ) | ( n10103 & n25582 ) | ( n25579 & n25582 ) ;
  assign n25584 = n25583 ^ n6974 ^ n6413 ;
  assign n25585 = ( n2906 & n5299 ) | ( n2906 & ~n11862 ) | ( n5299 & ~n11862 ) ;
  assign n25586 = n25585 ^ n6224 ^ 1'b0 ;
  assign n25587 = ( n556 & n14656 ) | ( n556 & n25586 ) | ( n14656 & n25586 ) ;
  assign n25588 = n24336 ^ n14478 ^ n13062 ;
  assign n25589 = n5743 | n14204 ;
  assign n25590 = ( n4961 & n13542 ) | ( n4961 & ~n25589 ) | ( n13542 & ~n25589 ) ;
  assign n25591 = n25590 ^ n9017 ^ n6318 ;
  assign n25592 = n2095 & ~n11916 ;
  assign n25593 = ~n16198 & n25592 ;
  assign n25594 = ( n5583 & ~n25591 ) | ( n5583 & n25593 ) | ( ~n25591 & n25593 ) ;
  assign n25595 = ( n3039 & ~n3774 ) | ( n3039 & n7407 ) | ( ~n3774 & n7407 ) ;
  assign n25596 = ( n14607 & ~n14684 ) | ( n14607 & n25595 ) | ( ~n14684 & n25595 ) ;
  assign n25597 = n25596 ^ n1925 ^ 1'b0 ;
  assign n25598 = n6753 | n20359 ;
  assign n25599 = n25598 ^ n11891 ^ 1'b0 ;
  assign n25600 = ( n1445 & n9001 ) | ( n1445 & ~n21268 ) | ( n9001 & ~n21268 ) ;
  assign n25601 = ( n2095 & n7638 ) | ( n2095 & ~n24347 ) | ( n7638 & ~n24347 ) ;
  assign n25602 = ( n5039 & n25600 ) | ( n5039 & ~n25601 ) | ( n25600 & ~n25601 ) ;
  assign n25603 = ~n12773 & n22649 ;
  assign n25604 = n4134 & n8907 ;
  assign n25605 = n25604 ^ n23176 ^ 1'b0 ;
  assign n25606 = ( ~n8630 & n25603 ) | ( ~n8630 & n25605 ) | ( n25603 & n25605 ) ;
  assign n25607 = ~n10918 & n16462 ;
  assign n25608 = n25607 ^ n20225 ^ n11643 ;
  assign n25609 = ( n5743 & ~n13426 ) | ( n5743 & n22464 ) | ( ~n13426 & n22464 ) ;
  assign n25610 = ( ~n2450 & n2730 ) | ( ~n2450 & n6668 ) | ( n2730 & n6668 ) ;
  assign n25611 = n152 & ~n15295 ;
  assign n25612 = ~n647 & n25611 ;
  assign n25613 = ( n806 & n2894 ) | ( n806 & n5224 ) | ( n2894 & n5224 ) ;
  assign n25614 = ( n11385 & n12648 ) | ( n11385 & n19532 ) | ( n12648 & n19532 ) ;
  assign n25615 = n25614 ^ n15240 ^ n947 ;
  assign n25616 = ( n1037 & n25613 ) | ( n1037 & ~n25615 ) | ( n25613 & ~n25615 ) ;
  assign n25617 = ( n25610 & n25612 ) | ( n25610 & n25616 ) | ( n25612 & n25616 ) ;
  assign n25618 = n2816 & ~n3580 ;
  assign n25619 = n10854 ^ n9268 ^ n8715 ;
  assign n25621 = ( n256 & n2425 ) | ( n256 & n10492 ) | ( n2425 & n10492 ) ;
  assign n25620 = n4656 & n20793 ;
  assign n25622 = n25621 ^ n25620 ^ 1'b0 ;
  assign n25623 = n8491 ^ n8304 ^ 1'b0 ;
  assign n25624 = n9330 & n25623 ;
  assign n25625 = ( n1718 & ~n11257 ) | ( n1718 & n15366 ) | ( ~n11257 & n15366 ) ;
  assign n25626 = n25625 ^ n24563 ^ n6047 ;
  assign n25628 = n25472 ^ n10001 ^ n8189 ;
  assign n25627 = ( n9333 & ~n22585 ) | ( n9333 & n24838 ) | ( ~n22585 & n24838 ) ;
  assign n25629 = n25628 ^ n25627 ^ n7106 ;
  assign n25630 = ( ~n1817 & n4913 ) | ( ~n1817 & n7935 ) | ( n4913 & n7935 ) ;
  assign n25631 = n25630 ^ n15386 ^ n11435 ;
  assign n25632 = n2895 & ~n23563 ;
  assign n25633 = ( ~n1964 & n3180 ) | ( ~n1964 & n6443 ) | ( n3180 & n6443 ) ;
  assign n25634 = n7729 ^ n4985 ^ n2890 ;
  assign n25635 = ( n22696 & ~n25633 ) | ( n22696 & n25634 ) | ( ~n25633 & n25634 ) ;
  assign n25636 = ( n3709 & n7192 ) | ( n3709 & ~n9171 ) | ( n7192 & ~n9171 ) ;
  assign n25637 = ( n259 & n1308 ) | ( n259 & n2137 ) | ( n1308 & n2137 ) ;
  assign n25638 = ~n17269 & n20658 ;
  assign n25639 = n25638 ^ n16634 ^ 1'b0 ;
  assign n25640 = n5429 & n20673 ;
  assign n25641 = n25640 ^ n2046 ^ 1'b0 ;
  assign n25642 = n22861 ^ n13415 ^ n11024 ;
  assign n25643 = n25642 ^ n15927 ^ n4879 ;
  assign n25644 = ( n1970 & n15077 ) | ( n1970 & ~n23622 ) | ( n15077 & ~n23622 ) ;
  assign n25645 = ( ~n7489 & n22211 ) | ( ~n7489 & n25644 ) | ( n22211 & n25644 ) ;
  assign n25646 = n22803 ^ n20565 ^ n11710 ;
  assign n25647 = n25646 ^ n13915 ^ n1397 ;
  assign n25648 = n8681 & n9808 ;
  assign n25649 = n11610 ^ n7532 ^ n5497 ;
  assign n25650 = ~n13737 & n25649 ;
  assign n25651 = n25648 & n25650 ;
  assign n25652 = n25651 ^ n6064 ^ n2260 ;
  assign n25653 = n23153 ^ n720 ^ 1'b0 ;
  assign n25655 = ( n522 & n4160 ) | ( n522 & ~n13904 ) | ( n4160 & ~n13904 ) ;
  assign n25654 = n17113 ^ n9719 ^ n1506 ;
  assign n25656 = n25655 ^ n25654 ^ n224 ;
  assign n25657 = n6045 | n22214 ;
  assign n25658 = ( ~n19465 & n25656 ) | ( ~n19465 & n25657 ) | ( n25656 & n25657 ) ;
  assign n25659 = n20036 ^ n18336 ^ n3139 ;
  assign n25661 = n5372 | n9304 ;
  assign n25662 = n25661 ^ n2450 ^ 1'b0 ;
  assign n25660 = n7855 & ~n15882 ;
  assign n25663 = n25662 ^ n25660 ^ 1'b0 ;
  assign n25664 = n20715 ^ n17183 ^ n16189 ;
  assign n25665 = n25664 ^ n4270 ^ 1'b0 ;
  assign n25666 = n11442 & n25665 ;
  assign n25668 = ( n3988 & ~n8929 ) | ( n3988 & n16277 ) | ( ~n8929 & n16277 ) ;
  assign n25667 = ( ~n2208 & n2568 ) | ( ~n2208 & n12695 ) | ( n2568 & n12695 ) ;
  assign n25669 = n25668 ^ n25667 ^ n10318 ;
  assign n25670 = ( n536 & n10931 ) | ( n536 & n25669 ) | ( n10931 & n25669 ) ;
  assign n25671 = ( ~n8640 & n11559 ) | ( ~n8640 & n14553 ) | ( n11559 & n14553 ) ;
  assign n25672 = n233 | n25671 ;
  assign n25673 = n25672 ^ n1115 ^ 1'b0 ;
  assign n25674 = n12887 ^ n2349 ^ 1'b0 ;
  assign n25675 = ~n14782 & n25674 ;
  assign n25676 = n22009 ^ n4212 ^ n3533 ;
  assign n25677 = ( n14092 & n25675 ) | ( n14092 & ~n25676 ) | ( n25675 & ~n25676 ) ;
  assign n25678 = n15174 ^ n6259 ^ n5761 ;
  assign n25679 = n17316 ^ n13224 ^ n331 ;
  assign n25680 = n20428 ^ n8382 ^ n2656 ;
  assign n25681 = n25680 ^ n2898 ^ 1'b0 ;
  assign n25682 = ( n10720 & ~n14861 ) | ( n10720 & n19793 ) | ( ~n14861 & n19793 ) ;
  assign n25683 = ( n4608 & n18747 ) | ( n4608 & ~n25682 ) | ( n18747 & ~n25682 ) ;
  assign n25684 = ( ~n6858 & n22268 ) | ( ~n6858 & n25683 ) | ( n22268 & n25683 ) ;
  assign n25685 = n25684 ^ n16462 ^ n14358 ;
  assign n25686 = ( ~n3970 & n5794 ) | ( ~n3970 & n8399 ) | ( n5794 & n8399 ) ;
  assign n25687 = n4360 | n25686 ;
  assign n25688 = n5682 ^ n1735 ^ n315 ;
  assign n25689 = ( n16236 & n19271 ) | ( n16236 & ~n25688 ) | ( n19271 & ~n25688 ) ;
  assign n25690 = n18483 ^ n2610 ^ n832 ;
  assign n25691 = ~n6582 & n25690 ;
  assign n25692 = n25691 ^ n6342 ^ 1'b0 ;
  assign n25693 = ( n8156 & ~n22567 ) | ( n8156 & n23549 ) | ( ~n22567 & n23549 ) ;
  assign n25694 = ( n3091 & ~n24127 ) | ( n3091 & n24861 ) | ( ~n24127 & n24861 ) ;
  assign n25695 = n5000 ^ n4482 ^ n3622 ;
  assign n25696 = n25695 ^ n21701 ^ n8940 ;
  assign n25697 = n8564 ^ n8233 ^ n4726 ;
  assign n25698 = ( ~n3654 & n17349 ) | ( ~n3654 & n25697 ) | ( n17349 & n25697 ) ;
  assign n25699 = n19594 ^ n11677 ^ n7228 ;
  assign n25700 = n25699 ^ n17888 ^ n8865 ;
  assign n25701 = n5021 ^ n4165 ^ n1183 ;
  assign n25702 = n25701 ^ n1729 ^ n1354 ;
  assign n25703 = n24919 ^ n17688 ^ 1'b0 ;
  assign n25704 = n6157 | n25703 ;
  assign n25705 = n12095 ^ n4163 ^ 1'b0 ;
  assign n25706 = n19005 | n25705 ;
  assign n25707 = n17375 ^ n6041 ^ n3982 ;
  assign n25708 = n503 & ~n7860 ;
  assign n25709 = ( n13745 & ~n17786 ) | ( n13745 & n18182 ) | ( ~n17786 & n18182 ) ;
  assign n25710 = n25709 ^ n14432 ^ n148 ;
  assign n25711 = ( n16022 & n19409 ) | ( n16022 & n25710 ) | ( n19409 & n25710 ) ;
  assign n25712 = ( n10808 & n20542 ) | ( n10808 & ~n25711 ) | ( n20542 & ~n25711 ) ;
  assign n25713 = ( n3548 & n6511 ) | ( n3548 & n9834 ) | ( n6511 & n9834 ) ;
  assign n25714 = ( n2884 & n4438 ) | ( n2884 & ~n25713 ) | ( n4438 & ~n25713 ) ;
  assign n25715 = n25714 ^ n17900 ^ n5906 ;
  assign n25716 = ( n25708 & n25712 ) | ( n25708 & ~n25715 ) | ( n25712 & ~n25715 ) ;
  assign n25717 = n24041 ^ n11146 ^ n2239 ;
  assign n25718 = n16982 ^ n13015 ^ n1665 ;
  assign n25719 = n7761 & n25718 ;
  assign n25720 = n25719 ^ n11424 ^ 1'b0 ;
  assign n25721 = n15675 ^ n7688 ^ n3483 ;
  assign n25722 = ( ~n1027 & n25720 ) | ( ~n1027 & n25721 ) | ( n25720 & n25721 ) ;
  assign n25724 = n18914 ^ n16714 ^ n5675 ;
  assign n25723 = n24038 ^ n18364 ^ n7972 ;
  assign n25725 = n25724 ^ n25723 ^ n14870 ;
  assign n25726 = ( n10484 & n13554 ) | ( n10484 & ~n24207 ) | ( n13554 & ~n24207 ) ;
  assign n25727 = n9936 ^ n440 ^ 1'b0 ;
  assign n25728 = n25727 ^ n12597 ^ n10770 ;
  assign n25729 = n22811 ^ n10235 ^ n5222 ;
  assign n25730 = ( n2439 & n9651 ) | ( n2439 & ~n18379 ) | ( n9651 & ~n18379 ) ;
  assign n25731 = n4655 & ~n25730 ;
  assign n25732 = n25731 ^ n15504 ^ n3290 ;
  assign n25733 = ( n2196 & n10349 ) | ( n2196 & ~n14855 ) | ( n10349 & ~n14855 ) ;
  assign n25734 = n14332 ^ n4899 ^ 1'b0 ;
  assign n25735 = ~n1252 & n25734 ;
  assign n25736 = n25735 ^ n16634 ^ n6559 ;
  assign n25737 = ( ~n7280 & n25733 ) | ( ~n7280 & n25736 ) | ( n25733 & n25736 ) ;
  assign n25738 = n25266 ^ x83 ^ 1'b0 ;
  assign n25739 = n13387 | n25738 ;
  assign n25740 = n25739 ^ n25713 ^ n4302 ;
  assign n25741 = ( n4438 & ~n11051 ) | ( n4438 & n14751 ) | ( ~n11051 & n14751 ) ;
  assign n25742 = ( n2382 & ~n6743 ) | ( n2382 & n25741 ) | ( ~n6743 & n25741 ) ;
  assign n25743 = ( n4259 & n9882 ) | ( n4259 & n11146 ) | ( n9882 & n11146 ) ;
  assign n25744 = n25743 ^ n6413 ^ 1'b0 ;
  assign n25745 = n25744 ^ n16794 ^ n11828 ;
  assign n25746 = n2607 ^ n1336 ^ n1231 ;
  assign n25747 = ( n10868 & ~n16475 ) | ( n10868 & n25746 ) | ( ~n16475 & n25746 ) ;
  assign n25748 = ( n10053 & ~n16360 ) | ( n10053 & n25747 ) | ( ~n16360 & n25747 ) ;
  assign n25749 = n9628 ^ n8804 ^ n3629 ;
  assign n25750 = ( ~n691 & n20367 ) | ( ~n691 & n21473 ) | ( n20367 & n21473 ) ;
  assign n25751 = ( n283 & ~n3723 ) | ( n283 & n25750 ) | ( ~n3723 & n25750 ) ;
  assign n25752 = ( n1587 & n4518 ) | ( n1587 & n5738 ) | ( n4518 & n5738 ) ;
  assign n25753 = n16739 ^ n4251 ^ n3189 ;
  assign n25754 = n25753 ^ n20284 ^ n555 ;
  assign n25755 = ( n632 & ~n25752 ) | ( n632 & n25754 ) | ( ~n25752 & n25754 ) ;
  assign n25756 = n22233 ^ n7790 ^ n5122 ;
  assign n25757 = n15348 ^ n3008 ^ 1'b0 ;
  assign n25758 = n2054 & n4997 ;
  assign n25759 = ~n25757 & n25758 ;
  assign n25760 = ( x66 & n15156 ) | ( x66 & ~n15794 ) | ( n15156 & ~n15794 ) ;
  assign n25761 = ( n5721 & n14863 ) | ( n5721 & ~n25760 ) | ( n14863 & ~n25760 ) ;
  assign n25762 = n13527 ^ n1772 ^ n1164 ;
  assign n25763 = n25762 ^ n17249 ^ n14990 ;
  assign n25766 = ( n14847 & n16000 ) | ( n14847 & ~n16134 ) | ( n16000 & ~n16134 ) ;
  assign n25764 = ( n1143 & n1976 ) | ( n1143 & n20272 ) | ( n1976 & n20272 ) ;
  assign n25765 = ( n5906 & n18301 ) | ( n5906 & ~n25764 ) | ( n18301 & ~n25764 ) ;
  assign n25767 = n25766 ^ n25765 ^ 1'b0 ;
  assign n25768 = n25767 ^ n19123 ^ n12007 ;
  assign n25769 = n8350 ^ n3719 ^ 1'b0 ;
  assign n25770 = ~n9478 & n25769 ;
  assign n25771 = n25770 ^ n12220 ^ x14 ;
  assign n25775 = n4392 | n12367 ;
  assign n25776 = ~n5904 & n25775 ;
  assign n25777 = n12095 & n25776 ;
  assign n25772 = n16585 ^ n6276 ^ n3698 ;
  assign n25773 = n25772 ^ n18139 ^ 1'b0 ;
  assign n25774 = n5885 & n25773 ;
  assign n25778 = n25777 ^ n25774 ^ n7206 ;
  assign n25779 = n1794 & ~n12887 ;
  assign n25780 = n25779 ^ n3447 ^ 1'b0 ;
  assign n25781 = n25780 ^ n19282 ^ n11746 ;
  assign n25782 = n25781 ^ n18256 ^ n9683 ;
  assign n25783 = ( n3555 & n9861 ) | ( n3555 & ~n25782 ) | ( n9861 & ~n25782 ) ;
  assign n25784 = n21372 ^ n11739 ^ n4211 ;
  assign n25785 = n1311 | n25784 ;
  assign n25786 = n25785 ^ n8538 ^ 1'b0 ;
  assign n25787 = n9701 & ~n21286 ;
  assign n25788 = n25787 ^ n10223 ^ 1'b0 ;
  assign n25789 = ( n3266 & ~n10273 ) | ( n3266 & n14788 ) | ( ~n10273 & n14788 ) ;
  assign n25790 = n21810 & ~n25789 ;
  assign n25791 = n21425 ^ n20477 ^ n7564 ;
  assign n25793 = n23257 ^ n19934 ^ n1689 ;
  assign n25792 = ~n13228 & n17295 ;
  assign n25794 = n25793 ^ n25792 ^ n18799 ;
  assign n25795 = ~n1679 & n7851 ;
  assign n25796 = n6102 & n25795 ;
  assign n25797 = ~n1797 & n25796 ;
  assign n25798 = n25797 ^ n17292 ^ n1904 ;
  assign n25799 = ( n1021 & n11424 ) | ( n1021 & n23933 ) | ( n11424 & n23933 ) ;
  assign n25800 = n18642 ^ n10061 ^ 1'b0 ;
  assign n25801 = n25800 ^ n16312 ^ n14845 ;
  assign n25802 = n19454 ^ n11240 ^ n7764 ;
  assign n25803 = ( ~n25799 & n25801 ) | ( ~n25799 & n25802 ) | ( n25801 & n25802 ) ;
  assign n25805 = ( n4617 & n5950 ) | ( n4617 & n9557 ) | ( n5950 & n9557 ) ;
  assign n25806 = n25805 ^ n14106 ^ n9268 ;
  assign n25807 = ( n10219 & ~n23620 ) | ( n10219 & n25806 ) | ( ~n23620 & n25806 ) ;
  assign n25804 = ( n710 & n11306 ) | ( n710 & ~n18205 ) | ( n11306 & ~n18205 ) ;
  assign n25808 = n25807 ^ n25804 ^ n13074 ;
  assign n25809 = ( n3419 & n17804 ) | ( n3419 & n22539 ) | ( n17804 & n22539 ) ;
  assign n25813 = n11671 ^ n8101 ^ 1'b0 ;
  assign n25810 = n12529 ^ n8889 ^ n8506 ;
  assign n25811 = ( n7875 & n13164 ) | ( n7875 & ~n25810 ) | ( n13164 & ~n25810 ) ;
  assign n25812 = n25811 ^ n17290 ^ n7262 ;
  assign n25814 = n25813 ^ n25812 ^ n23598 ;
  assign n25815 = n25814 ^ n23589 ^ 1'b0 ;
  assign n25816 = n25815 ^ n2846 ^ 1'b0 ;
  assign n25817 = ~n2923 & n3507 ;
  assign n25818 = n25817 ^ n12966 ^ 1'b0 ;
  assign n25819 = ( ~n3229 & n18230 ) | ( ~n3229 & n20343 ) | ( n18230 & n20343 ) ;
  assign n25820 = n25819 ^ n13778 ^ 1'b0 ;
  assign n25821 = n4995 & n25820 ;
  assign n25822 = ( n4309 & n4872 ) | ( n4309 & ~n8694 ) | ( n4872 & ~n8694 ) ;
  assign n25823 = n2114 | n17624 ;
  assign n25824 = n3520 | n3591 ;
  assign n25825 = n25824 ^ n22364 ^ 1'b0 ;
  assign n25826 = ( ~n8881 & n8946 ) | ( ~n8881 & n11466 ) | ( n8946 & n11466 ) ;
  assign n25827 = ( n7115 & ~n25825 ) | ( n7115 & n25826 ) | ( ~n25825 & n25826 ) ;
  assign n25828 = n7157 ^ n887 ^ n332 ;
  assign n25829 = ( ~n7938 & n12096 ) | ( ~n7938 & n25828 ) | ( n12096 & n25828 ) ;
  assign n25830 = ( n19722 & n23059 ) | ( n19722 & ~n24529 ) | ( n23059 & ~n24529 ) ;
  assign n25831 = n14837 ^ n11583 ^ n1684 ;
  assign n25834 = n3022 & ~n5625 ;
  assign n25835 = n9044 & n25834 ;
  assign n25832 = n10088 ^ n8140 ^ n845 ;
  assign n25833 = n6184 | n25832 ;
  assign n25836 = n25835 ^ n25833 ^ 1'b0 ;
  assign n25837 = n25509 ^ n13686 ^ n5305 ;
  assign n25839 = ( n8026 & n17709 ) | ( n8026 & n21338 ) | ( n17709 & n21338 ) ;
  assign n25840 = ( n11408 & ~n23430 ) | ( n11408 & n25839 ) | ( ~n23430 & n25839 ) ;
  assign n25838 = n9416 ^ n1608 ^ 1'b0 ;
  assign n25841 = n25840 ^ n25838 ^ n15530 ;
  assign n25842 = n2892 & n15684 ;
  assign n25843 = ( ~n3601 & n11325 ) | ( ~n3601 & n14964 ) | ( n11325 & n14964 ) ;
  assign n25844 = n18768 ^ n11686 ^ n11439 ;
  assign n25845 = ( n3467 & n10925 ) | ( n3467 & ~n15949 ) | ( n10925 & ~n15949 ) ;
  assign n25846 = n10366 & ~n25845 ;
  assign n25847 = n5109 & n25846 ;
  assign n25848 = ~n2652 & n25847 ;
  assign n25849 = ( n7057 & n8985 ) | ( n7057 & ~n25848 ) | ( n8985 & ~n25848 ) ;
  assign n25850 = ( n734 & ~n25844 ) | ( n734 & n25849 ) | ( ~n25844 & n25849 ) ;
  assign n25851 = n22798 ^ n21081 ^ n8064 ;
  assign n25852 = n12130 ^ n6622 ^ 1'b0 ;
  assign n25853 = n7062 | n25852 ;
  assign n25854 = ( n8441 & ~n19159 ) | ( n8441 & n19381 ) | ( ~n19159 & n19381 ) ;
  assign n25858 = n15713 ^ n10452 ^ n3699 ;
  assign n25855 = n18146 ^ n6152 ^ n2880 ;
  assign n25856 = n1340 & ~n7879 ;
  assign n25857 = ~n25855 & n25856 ;
  assign n25859 = n25858 ^ n25857 ^ n21728 ;
  assign n25861 = n10394 ^ n6961 ^ n2698 ;
  assign n25860 = n10447 ^ n10369 ^ n1515 ;
  assign n25862 = n25861 ^ n25860 ^ n24531 ;
  assign n25863 = n20401 ^ n12812 ^ n2487 ;
  assign n25864 = ( ~n1291 & n7039 ) | ( ~n1291 & n12811 ) | ( n7039 & n12811 ) ;
  assign n25865 = ( n19863 & n19889 ) | ( n19863 & n25864 ) | ( n19889 & n25864 ) ;
  assign n25866 = ( n22455 & ~n25863 ) | ( n22455 & n25865 ) | ( ~n25863 & n25865 ) ;
  assign n25867 = ( ~n418 & n1662 ) | ( ~n418 & n3718 ) | ( n1662 & n3718 ) ;
  assign n25868 = n17621 ^ n15347 ^ n10750 ;
  assign n25869 = n25868 ^ n18483 ^ n14096 ;
  assign n25870 = ( n14505 & n25867 ) | ( n14505 & n25869 ) | ( n25867 & n25869 ) ;
  assign n25871 = n19968 ^ n19790 ^ n6818 ;
  assign n25872 = ~n20254 & n25871 ;
  assign n25873 = n3936 & n25872 ;
  assign n25874 = n9412 & ~n13175 ;
  assign n25875 = ~n3935 & n25874 ;
  assign n25876 = n25875 ^ n13010 ^ n7129 ;
  assign n25877 = ( n13303 & ~n21535 ) | ( n13303 & n25876 ) | ( ~n21535 & n25876 ) ;
  assign n25878 = ( n2470 & ~n25873 ) | ( n2470 & n25877 ) | ( ~n25873 & n25877 ) ;
  assign n25879 = n9717 ^ n4121 ^ n3938 ;
  assign n25880 = n25879 ^ n14312 ^ n6197 ;
  assign n25881 = n2227 | n15211 ;
  assign n25882 = n9175 | n25881 ;
  assign n25883 = n17957 ^ n12915 ^ n7530 ;
  assign n25884 = n25883 ^ n8974 ^ n1026 ;
  assign n25885 = n23817 ^ n16588 ^ n6716 ;
  assign n25886 = n25885 ^ n18922 ^ n4274 ;
  assign n25888 = n7840 ^ n3149 ^ 1'b0 ;
  assign n25889 = ~n3465 & n25888 ;
  assign n25887 = ( n11055 & n12133 ) | ( n11055 & n22126 ) | ( n12133 & n22126 ) ;
  assign n25890 = n25889 ^ n25887 ^ n1309 ;
  assign n25891 = n2402 & ~n15986 ;
  assign n25892 = n25891 ^ x99 ^ 1'b0 ;
  assign n25893 = ( n20983 & n24789 ) | ( n20983 & n25892 ) | ( n24789 & n25892 ) ;
  assign n25894 = n13036 ^ n8239 ^ n2114 ;
  assign n25895 = n12150 ^ n11584 ^ n5249 ;
  assign n25896 = n22087 ^ n21601 ^ n430 ;
  assign n25897 = ( n5103 & n8707 ) | ( n5103 & ~n25896 ) | ( n8707 & ~n25896 ) ;
  assign n25898 = n25897 ^ n3123 ^ 1'b0 ;
  assign n25899 = n24809 & ~n25898 ;
  assign n25900 = n6982 | n13986 ;
  assign n25901 = n9379 & ~n25900 ;
  assign n25902 = ( n1479 & ~n5476 ) | ( n1479 & n22863 ) | ( ~n5476 & n22863 ) ;
  assign n25903 = n22663 ^ n17245 ^ n10957 ;
  assign n25904 = n24478 ^ n18204 ^ n5115 ;
  assign n25905 = ( n9027 & n14233 ) | ( n9027 & ~n17207 ) | ( n14233 & ~n17207 ) ;
  assign n25906 = ( n992 & n10619 ) | ( n992 & ~n25905 ) | ( n10619 & ~n25905 ) ;
  assign n25907 = n25906 ^ n16910 ^ n1063 ;
  assign n25908 = n3323 ^ n1751 ^ n1369 ;
  assign n25909 = n919 & n3476 ;
  assign n25910 = ( x96 & n2378 ) | ( x96 & ~n8363 ) | ( n2378 & ~n8363 ) ;
  assign n25911 = ( ~n8622 & n21554 ) | ( ~n8622 & n25910 ) | ( n21554 & n25910 ) ;
  assign n25912 = ( n25908 & ~n25909 ) | ( n25908 & n25911 ) | ( ~n25909 & n25911 ) ;
  assign n25913 = ( n2402 & n5838 ) | ( n2402 & ~n13431 ) | ( n5838 & ~n13431 ) ;
  assign n25914 = n7702 ^ n1663 ^ 1'b0 ;
  assign n25915 = n6024 & n25914 ;
  assign n25916 = n25913 & n25915 ;
  assign n25917 = n8002 | n8035 ;
  assign n25918 = n25917 ^ n9985 ^ n6762 ;
  assign n25919 = ( n18325 & ~n23227 ) | ( n18325 & n25918 ) | ( ~n23227 & n25918 ) ;
  assign n25922 = n10101 ^ n7352 ^ n3628 ;
  assign n25920 = ~n4352 & n5462 ;
  assign n25921 = n25920 ^ n2509 ^ n1538 ;
  assign n25923 = n25922 ^ n25921 ^ n7198 ;
  assign n25924 = n13115 ^ n8305 ^ n2795 ;
  assign n25925 = ( n16905 & ~n25923 ) | ( n16905 & n25924 ) | ( ~n25923 & n25924 ) ;
  assign n25928 = n11921 ^ n7548 ^ 1'b0 ;
  assign n25929 = ~n12131 & n25928 ;
  assign n25927 = ( n14320 & n14710 ) | ( n14320 & n22732 ) | ( n14710 & n22732 ) ;
  assign n25926 = ( n7361 & n10887 ) | ( n7361 & n18624 ) | ( n10887 & n18624 ) ;
  assign n25930 = n25929 ^ n25927 ^ n25926 ;
  assign n25931 = ( n13048 & n18720 ) | ( n13048 & n19424 ) | ( n18720 & n19424 ) ;
  assign n25932 = ( n6309 & n11762 ) | ( n6309 & ~n24368 ) | ( n11762 & ~n24368 ) ;
  assign n25933 = n18406 ^ n13624 ^ n9399 ;
  assign n25934 = ( ~n3122 & n7511 ) | ( ~n3122 & n10358 ) | ( n7511 & n10358 ) ;
  assign n25935 = ( ~n12497 & n25933 ) | ( ~n12497 & n25934 ) | ( n25933 & n25934 ) ;
  assign n25936 = n25363 ^ n22251 ^ n757 ;
  assign n25937 = n12211 ^ n7338 ^ n3982 ;
  assign n25938 = n14757 ^ n3259 ^ 1'b0 ;
  assign n25939 = ( n4050 & n15581 ) | ( n4050 & ~n25938 ) | ( n15581 & ~n25938 ) ;
  assign n25940 = ( ~n6978 & n25937 ) | ( ~n6978 & n25939 ) | ( n25937 & n25939 ) ;
  assign n25941 = n9415 ^ n1943 ^ 1'b0 ;
  assign n25942 = n17485 & n25746 ;
  assign n25943 = n23752 ^ n6877 ^ n5639 ;
  assign n25944 = ( ~n898 & n20276 ) | ( ~n898 & n25943 ) | ( n20276 & n25943 ) ;
  assign n25945 = n10238 ^ n3734 ^ 1'b0 ;
  assign n25946 = ( n1400 & n21269 ) | ( n1400 & n25945 ) | ( n21269 & n25945 ) ;
  assign n25949 = ( n6004 & ~n13143 ) | ( n6004 & n16091 ) | ( ~n13143 & n16091 ) ;
  assign n25948 = ( ~n7778 & n7988 ) | ( ~n7778 & n8845 ) | ( n7988 & n8845 ) ;
  assign n25947 = n15658 ^ n13571 ^ n907 ;
  assign n25950 = n25949 ^ n25948 ^ n25947 ;
  assign n25951 = n25950 ^ n22448 ^ n9934 ;
  assign n25952 = n25259 ^ n10191 ^ n6338 ;
  assign n25953 = n23944 ^ n10591 ^ n7209 ;
  assign n25954 = ~n1434 & n12213 ;
  assign n25955 = n5195 & n25954 ;
  assign n25956 = n25955 ^ n15993 ^ n10619 ;
  assign n25957 = n25956 ^ n14905 ^ n2780 ;
  assign n25960 = n24751 ^ n12983 ^ n7478 ;
  assign n25961 = ( n1738 & n4539 ) | ( n1738 & ~n25960 ) | ( n4539 & ~n25960 ) ;
  assign n25958 = n19922 ^ n19162 ^ n4294 ;
  assign n25959 = n25958 ^ n15656 ^ n13736 ;
  assign n25962 = n25961 ^ n25959 ^ n1172 ;
  assign n25963 = n24070 ^ n14864 ^ n12368 ;
  assign n25964 = ( n4118 & n10439 ) | ( n4118 & n15115 ) | ( n10439 & n15115 ) ;
  assign n25965 = ( n2326 & n12242 ) | ( n2326 & ~n25964 ) | ( n12242 & ~n25964 ) ;
  assign n25966 = n25965 ^ n5146 ^ 1'b0 ;
  assign n25967 = n25963 | n25966 ;
  assign n25968 = ( n4317 & ~n4711 ) | ( n4317 & n18245 ) | ( ~n4711 & n18245 ) ;
  assign n25969 = ~n9789 & n19849 ;
  assign n25970 = n25968 & n25969 ;
  assign n25971 = ( n220 & n6163 ) | ( n220 & n7766 ) | ( n6163 & n7766 ) ;
  assign n25972 = n17138 ^ n10319 ^ n7379 ;
  assign n25973 = n20023 ^ n10942 ^ 1'b0 ;
  assign n25974 = ( n25971 & n25972 ) | ( n25971 & ~n25973 ) | ( n25972 & ~n25973 ) ;
  assign n25975 = n24589 ^ n13834 ^ 1'b0 ;
  assign n25976 = ( n356 & n6922 ) | ( n356 & ~n10611 ) | ( n6922 & ~n10611 ) ;
  assign n25977 = n25695 ^ n16028 ^ 1'b0 ;
  assign n25978 = ( n4470 & n15432 ) | ( n4470 & n17086 ) | ( n15432 & n17086 ) ;
  assign n25979 = n3184 & n16824 ;
  assign n25980 = ~n25978 & n25979 ;
  assign n25981 = n18646 ^ n7877 ^ n4065 ;
  assign n25982 = n25981 ^ n19635 ^ 1'b0 ;
  assign n25983 = n11652 | n25982 ;
  assign n25984 = n5715 & n20157 ;
  assign n25985 = n8623 & n25984 ;
  assign n25986 = n25985 ^ n15012 ^ n3658 ;
  assign n25987 = n16248 ^ n8628 ^ 1'b0 ;
  assign n25988 = n13404 & n25987 ;
  assign n25990 = n11148 ^ n6559 ^ n4540 ;
  assign n25991 = ( n5897 & ~n8823 ) | ( n5897 & n25990 ) | ( ~n8823 & n25990 ) ;
  assign n25989 = n24618 ^ n4422 ^ n3657 ;
  assign n25992 = n25991 ^ n25989 ^ 1'b0 ;
  assign n25993 = ( n11493 & n13716 ) | ( n11493 & ~n22426 ) | ( n13716 & ~n22426 ) ;
  assign n25994 = n25993 ^ n23095 ^ n7314 ;
  assign n25995 = n25994 ^ n16061 ^ n405 ;
  assign n25996 = n12095 ^ n7890 ^ n7337 ;
  assign n25997 = n24474 & ~n25996 ;
  assign n25998 = n25997 ^ n13856 ^ 1'b0 ;
  assign n25999 = ( n2923 & ~n10059 ) | ( n2923 & n25998 ) | ( ~n10059 & n25998 ) ;
  assign n26000 = ( ~n1047 & n10386 ) | ( ~n1047 & n21211 ) | ( n10386 & n21211 ) ;
  assign n26001 = ( n4285 & n10809 ) | ( n4285 & n25331 ) | ( n10809 & n25331 ) ;
  assign n26002 = ( n4814 & ~n17425 ) | ( n4814 & n26001 ) | ( ~n17425 & n26001 ) ;
  assign n26003 = n7115 | n9058 ;
  assign n26004 = n26003 ^ n1243 ^ 1'b0 ;
  assign n26005 = n3352 & n26004 ;
  assign n26006 = n25948 ^ n11014 ^ 1'b0 ;
  assign n26008 = n2152 | n18368 ;
  assign n26007 = n13741 ^ n7983 ^ n3677 ;
  assign n26009 = n26008 ^ n26007 ^ n7131 ;
  assign n26010 = n24960 ^ n11269 ^ n2448 ;
  assign n26011 = n11250 ^ n4667 ^ n748 ;
  assign n26012 = n26011 ^ n21810 ^ n13437 ;
  assign n26013 = ( n1232 & n3410 ) | ( n1232 & ~n14435 ) | ( n3410 & ~n14435 ) ;
  assign n26014 = n26013 ^ n24058 ^ n3028 ;
  assign n26015 = ( ~n1044 & n9949 ) | ( ~n1044 & n12769 ) | ( n9949 & n12769 ) ;
  assign n26016 = ( n5308 & n12133 ) | ( n5308 & ~n26015 ) | ( n12133 & ~n26015 ) ;
  assign n26017 = n21973 ^ n21048 ^ n11622 ;
  assign n26018 = ( n15551 & n26016 ) | ( n15551 & ~n26017 ) | ( n26016 & ~n26017 ) ;
  assign n26019 = ( x95 & ~n1006 ) | ( x95 & n17940 ) | ( ~n1006 & n17940 ) ;
  assign n26020 = n11396 & n26019 ;
  assign n26021 = n26018 & n26020 ;
  assign n26022 = ( n17532 & n26014 ) | ( n17532 & n26021 ) | ( n26014 & n26021 ) ;
  assign n26024 = n18927 ^ n4578 ^ 1'b0 ;
  assign n26025 = n1752 & n26024 ;
  assign n26026 = ( n1786 & n5720 ) | ( n1786 & n26025 ) | ( n5720 & n26025 ) ;
  assign n26027 = ( n923 & n25383 ) | ( n923 & ~n26026 ) | ( n25383 & ~n26026 ) ;
  assign n26023 = ( n2457 & n5870 ) | ( n2457 & ~n15174 ) | ( n5870 & ~n15174 ) ;
  assign n26028 = n26027 ^ n26023 ^ 1'b0 ;
  assign n26029 = ~n26022 & n26028 ;
  assign n26030 = ( n748 & n2660 ) | ( n748 & n3703 ) | ( n2660 & n3703 ) ;
  assign n26031 = ( n6047 & n22227 ) | ( n6047 & ~n26030 ) | ( n22227 & ~n26030 ) ;
  assign n26032 = n26031 ^ n8092 ^ n4110 ;
  assign n26033 = n17245 ^ n6807 ^ n2893 ;
  assign n26034 = n10984 ^ n8820 ^ n7995 ;
  assign n26035 = ( n17527 & ~n18931 ) | ( n17527 & n26034 ) | ( ~n18931 & n26034 ) ;
  assign n26036 = ( n19462 & ~n26033 ) | ( n19462 & n26035 ) | ( ~n26033 & n26035 ) ;
  assign n26037 = n12089 ^ n5485 ^ 1'b0 ;
  assign n26038 = n12835 & n26037 ;
  assign n26039 = ( n4383 & n15405 ) | ( n4383 & ~n26038 ) | ( n15405 & ~n26038 ) ;
  assign n26040 = n26039 ^ n21387 ^ n5135 ;
  assign n26041 = ( n5520 & ~n8101 ) | ( n5520 & n12076 ) | ( ~n8101 & n12076 ) ;
  assign n26042 = ( ~n7767 & n8089 ) | ( ~n7767 & n14122 ) | ( n8089 & n14122 ) ;
  assign n26043 = n4104 | n6666 ;
  assign n26044 = n2151 & ~n26043 ;
  assign n26045 = ( ~n12576 & n21074 ) | ( ~n12576 & n26044 ) | ( n21074 & n26044 ) ;
  assign n26049 = ( n15634 & ~n16226 ) | ( n15634 & n22888 ) | ( ~n16226 & n22888 ) ;
  assign n26046 = n11614 ^ n4709 ^ n1140 ;
  assign n26047 = ( n1594 & n5395 ) | ( n1594 & n26046 ) | ( n5395 & n26046 ) ;
  assign n26048 = n26047 ^ n22829 ^ n3736 ;
  assign n26050 = n26049 ^ n26048 ^ n18086 ;
  assign n26051 = n18396 ^ n2530 ^ n1100 ;
  assign n26052 = ( n5151 & ~n7836 ) | ( n5151 & n14905 ) | ( ~n7836 & n14905 ) ;
  assign n26053 = n26052 ^ n12770 ^ x50 ;
  assign n26054 = ( n4471 & n17677 ) | ( n4471 & ~n24972 ) | ( n17677 & ~n24972 ) ;
  assign n26055 = n10196 ^ n8310 ^ x36 ;
  assign n26056 = ( n10409 & n15266 ) | ( n10409 & ~n26055 ) | ( n15266 & ~n26055 ) ;
  assign n26057 = ( ~n5025 & n9896 ) | ( ~n5025 & n21341 ) | ( n9896 & n21341 ) ;
  assign n26058 = n26057 ^ n20333 ^ n12172 ;
  assign n26059 = ( n5375 & ~n16969 ) | ( n5375 & n26058 ) | ( ~n16969 & n26058 ) ;
  assign n26060 = n26059 ^ n10746 ^ n7843 ;
  assign n26061 = ( n7044 & n12253 ) | ( n7044 & n21756 ) | ( n12253 & n21756 ) ;
  assign n26062 = ( n6290 & ~n7626 ) | ( n6290 & n14476 ) | ( ~n7626 & n14476 ) ;
  assign n26063 = ( ~n10033 & n11309 ) | ( ~n10033 & n26062 ) | ( n11309 & n26062 ) ;
  assign n26065 = n1778 & n12504 ;
  assign n26064 = n6862 & n19389 ;
  assign n26066 = n26065 ^ n26064 ^ 1'b0 ;
  assign n26067 = n25933 ^ n5643 ^ n2918 ;
  assign n26068 = n24617 ^ n21164 ^ n16296 ;
  assign n26071 = n12199 ^ n9290 ^ n6176 ;
  assign n26069 = ( n3502 & ~n5719 ) | ( n3502 & n16028 ) | ( ~n5719 & n16028 ) ;
  assign n26070 = n26069 ^ n14544 ^ 1'b0 ;
  assign n26072 = n26071 ^ n26070 ^ n7262 ;
  assign n26073 = ( n6523 & ~n10166 ) | ( n6523 & n13081 ) | ( ~n10166 & n13081 ) ;
  assign n26074 = ( n461 & n12478 ) | ( n461 & n18677 ) | ( n12478 & n18677 ) ;
  assign n26075 = n26074 ^ n17523 ^ n6251 ;
  assign n26076 = ~n678 & n11041 ;
  assign n26077 = ~n4819 & n19096 ;
  assign n26078 = ~n26076 & n26077 ;
  assign n26079 = ( n10647 & n22256 ) | ( n10647 & ~n26078 ) | ( n22256 & ~n26078 ) ;
  assign n26080 = ( n588 & n848 ) | ( n588 & n3419 ) | ( n848 & n3419 ) ;
  assign n26081 = ( n6384 & ~n6992 ) | ( n6384 & n22907 ) | ( ~n6992 & n22907 ) ;
  assign n26082 = n26081 ^ n21984 ^ n21973 ;
  assign n26083 = ( n2566 & n26080 ) | ( n2566 & ~n26082 ) | ( n26080 & ~n26082 ) ;
  assign n26084 = n24660 ^ n21601 ^ 1'b0 ;
  assign n26085 = n1821 & n26084 ;
  assign n26086 = ( n1799 & n3901 ) | ( n1799 & ~n7934 ) | ( n3901 & ~n7934 ) ;
  assign n26087 = n26086 ^ n11725 ^ n5373 ;
  assign n26093 = ( n1041 & n4827 ) | ( n1041 & n4869 ) | ( n4827 & n4869 ) ;
  assign n26094 = ( n1821 & n23378 ) | ( n1821 & ~n26093 ) | ( n23378 & ~n26093 ) ;
  assign n26088 = ( n2110 & n6002 ) | ( n2110 & n7626 ) | ( n6002 & n7626 ) ;
  assign n26089 = ~n11419 & n26088 ;
  assign n26090 = n26089 ^ n8400 ^ 1'b0 ;
  assign n26091 = ( x2 & n11191 ) | ( x2 & n26090 ) | ( n11191 & n26090 ) ;
  assign n26092 = ( n2753 & n12036 ) | ( n2753 & n26091 ) | ( n12036 & n26091 ) ;
  assign n26095 = n26094 ^ n26092 ^ n3979 ;
  assign n26096 = ( ~n2648 & n4384 ) | ( ~n2648 & n22892 ) | ( n4384 & n22892 ) ;
  assign n26097 = ( n5739 & n15701 ) | ( n5739 & ~n26096 ) | ( n15701 & ~n26096 ) ;
  assign n26098 = n17962 ^ n4454 ^ n4229 ;
  assign n26099 = n26098 ^ n19783 ^ x46 ;
  assign n26100 = n3733 | n26099 ;
  assign n26101 = ( n6486 & n11937 ) | ( n6486 & ~n14867 ) | ( n11937 & ~n14867 ) ;
  assign n26102 = ( ~x107 & n847 ) | ( ~x107 & n3416 ) | ( n847 & n3416 ) ;
  assign n26103 = n2469 & ~n9040 ;
  assign n26104 = n26103 ^ n1033 ^ 1'b0 ;
  assign n26105 = ~n26102 & n26104 ;
  assign n26106 = n26105 ^ n15705 ^ 1'b0 ;
  assign n26107 = n26106 ^ n14566 ^ n11835 ;
  assign n26108 = n26107 ^ n20284 ^ 1'b0 ;
  assign n26109 = ( n3964 & n19699 ) | ( n3964 & n20085 ) | ( n19699 & n20085 ) ;
  assign n26113 = ( n2091 & n6689 ) | ( n2091 & ~n8096 ) | ( n6689 & ~n8096 ) ;
  assign n26110 = n22599 ^ n1760 ^ x101 ;
  assign n26111 = n26110 ^ n23846 ^ n15216 ;
  assign n26112 = n8051 & ~n26111 ;
  assign n26114 = n26113 ^ n26112 ^ 1'b0 ;
  assign n26115 = n2334 | n16508 ;
  assign n26116 = n1541 | n26115 ;
  assign n26117 = n16038 ^ n15266 ^ 1'b0 ;
  assign n26118 = n26116 & n26117 ;
  assign n26119 = n17847 ^ n12280 ^ n363 ;
  assign n26120 = n9781 ^ n8648 ^ n2609 ;
  assign n26121 = n24131 ^ n139 ^ 1'b0 ;
  assign n26122 = ( n1036 & n7244 ) | ( n1036 & ~n12700 ) | ( n7244 & ~n12700 ) ;
  assign n26123 = n22379 ^ n15408 ^ n3298 ;
  assign n26124 = ( n9929 & ~n10423 ) | ( n9929 & n26123 ) | ( ~n10423 & n26123 ) ;
  assign n26125 = n22216 ^ n5557 ^ 1'b0 ;
  assign n26126 = ( ~n7746 & n16390 ) | ( ~n7746 & n23143 ) | ( n16390 & n23143 ) ;
  assign n26127 = ( n8396 & n16283 ) | ( n8396 & ~n26126 ) | ( n16283 & ~n26126 ) ;
  assign n26128 = ( n5505 & n10105 ) | ( n5505 & ~n26127 ) | ( n10105 & ~n26127 ) ;
  assign n26129 = ( n624 & n8777 ) | ( n624 & n26128 ) | ( n8777 & n26128 ) ;
  assign n26130 = n26129 ^ n15271 ^ 1'b0 ;
  assign n26131 = ~n13239 & n26130 ;
  assign n26132 = n9543 & n10615 ;
  assign n26133 = n2574 | n19865 ;
  assign n26134 = n6800 & ~n7456 ;
  assign n26135 = ( n3067 & n9562 ) | ( n3067 & ~n20152 ) | ( n9562 & ~n20152 ) ;
  assign n26136 = ( n13301 & n13916 ) | ( n13301 & n26135 ) | ( n13916 & n26135 ) ;
  assign n26137 = n26136 ^ n25753 ^ n19554 ;
  assign n26138 = n11270 ^ n2371 ^ 1'b0 ;
  assign n26139 = n22345 ^ n18743 ^ 1'b0 ;
  assign n26140 = n26138 & n26139 ;
  assign n26141 = n16590 ^ n15463 ^ n7467 ;
  assign n26142 = n12373 ^ n6119 ^ n3877 ;
  assign n26143 = ( n2175 & n15416 ) | ( n2175 & n26142 ) | ( n15416 & n26142 ) ;
  assign n26144 = n1408 & n21611 ;
  assign n26145 = n26144 ^ n15185 ^ 1'b0 ;
  assign n26146 = ( n4979 & n6956 ) | ( n4979 & n7576 ) | ( n6956 & n7576 ) ;
  assign n26147 = ~n19150 & n19287 ;
  assign n26148 = ( ~n18149 & n26146 ) | ( ~n18149 & n26147 ) | ( n26146 & n26147 ) ;
  assign n26149 = ( n8545 & n11639 ) | ( n8545 & n12881 ) | ( n11639 & n12881 ) ;
  assign n26150 = n2151 & n6974 ;
  assign n26151 = n26150 ^ n18020 ^ n15055 ;
  assign n26152 = ( n3389 & n4838 ) | ( n3389 & n24148 ) | ( n4838 & n24148 ) ;
  assign n26154 = n8785 ^ n7959 ^ n5277 ;
  assign n26153 = n25013 ^ n12974 ^ n6162 ;
  assign n26155 = n26154 ^ n26153 ^ n4558 ;
  assign n26156 = n21720 ^ n17552 ^ n7449 ;
  assign n26157 = n26156 ^ n25155 ^ n19287 ;
  assign n26158 = n18316 ^ n15513 ^ 1'b0 ;
  assign n26159 = n908 | n26158 ;
  assign n26160 = ( ~n244 & n3044 ) | ( ~n244 & n23373 ) | ( n3044 & n23373 ) ;
  assign n26161 = n21572 ^ n14383 ^ 1'b0 ;
  assign n26164 = n23878 ^ n5108 ^ n3367 ;
  assign n26162 = n1002 & ~n1340 ;
  assign n26163 = ~n20410 & n26162 ;
  assign n26165 = n26164 ^ n26163 ^ n14178 ;
  assign n26166 = ( n2250 & ~n9044 ) | ( n2250 & n14841 ) | ( ~n9044 & n14841 ) ;
  assign n26167 = n19271 & n26166 ;
  assign n26168 = ( n8622 & ~n18677 ) | ( n8622 & n26167 ) | ( ~n18677 & n26167 ) ;
  assign n26169 = ( ~n10218 & n14818 ) | ( ~n10218 & n23085 ) | ( n14818 & n23085 ) ;
  assign n26170 = n6883 & ~n25037 ;
  assign n26171 = ( ~n180 & n6610 ) | ( ~n180 & n26170 ) | ( n6610 & n26170 ) ;
  assign n26172 = n26171 ^ n15839 ^ 1'b0 ;
  assign n26175 = ( n258 & n9721 ) | ( n258 & n24144 ) | ( n9721 & n24144 ) ;
  assign n26176 = n26175 ^ n5369 ^ n2457 ;
  assign n26177 = n26176 ^ n7244 ^ n373 ;
  assign n26173 = n4620 & n17289 ;
  assign n26174 = n26173 ^ n12800 ^ n6504 ;
  assign n26178 = n26177 ^ n26174 ^ n16060 ;
  assign n26179 = n22013 ^ n11715 ^ n3055 ;
  assign n26180 = n13784 ^ n13170 ^ n6313 ;
  assign n26181 = n26180 ^ n188 ^ 1'b0 ;
  assign n26182 = ( ~n1844 & n4334 ) | ( ~n1844 & n12140 ) | ( n4334 & n12140 ) ;
  assign n26183 = n26182 ^ n8164 ^ n4024 ;
  assign n26184 = ( n11626 & ~n18161 ) | ( n11626 & n26183 ) | ( ~n18161 & n26183 ) ;
  assign n26185 = n1945 & n16569 ;
  assign n26186 = n26185 ^ n10187 ^ 1'b0 ;
  assign n26187 = n25806 ^ n25486 ^ n4036 ;
  assign n26188 = ( n7387 & ~n13097 ) | ( n7387 & n13318 ) | ( ~n13097 & n13318 ) ;
  assign n26189 = ( n7017 & ~n20447 ) | ( n7017 & n26188 ) | ( ~n20447 & n26188 ) ;
  assign n26190 = n13056 ^ n9553 ^ 1'b0 ;
  assign n26191 = n26190 ^ n24721 ^ n5637 ;
  assign n26192 = ( n11077 & ~n17677 ) | ( n11077 & n26191 ) | ( ~n17677 & n26191 ) ;
  assign n26194 = n17208 ^ n9340 ^ n744 ;
  assign n26195 = n26194 ^ n19350 ^ n8674 ;
  assign n26193 = ( n4892 & n6733 ) | ( n4892 & n6840 ) | ( n6733 & n6840 ) ;
  assign n26196 = n26195 ^ n26193 ^ n10868 ;
  assign n26197 = n20534 ^ n20277 ^ n9058 ;
  assign n26198 = ~n3031 & n3884 ;
  assign n26199 = n1473 & n26198 ;
  assign n26200 = ( n8156 & n9025 ) | ( n8156 & n26199 ) | ( n9025 & n26199 ) ;
  assign n26201 = n9955 & n26200 ;
  assign n26202 = n15399 ^ n10408 ^ n7650 ;
  assign n26203 = n22143 | n22884 ;
  assign n26204 = ( n3441 & n26202 ) | ( n3441 & ~n26203 ) | ( n26202 & ~n26203 ) ;
  assign n26205 = n25017 ^ n3159 ^ n2731 ;
  assign n26206 = ( n9143 & n12157 ) | ( n9143 & n26205 ) | ( n12157 & n26205 ) ;
  assign n26207 = n23839 ^ n20064 ^ n17442 ;
  assign n26208 = ( n26204 & ~n26206 ) | ( n26204 & n26207 ) | ( ~n26206 & n26207 ) ;
  assign n26209 = ( ~n11639 & n14278 ) | ( ~n11639 & n26104 ) | ( n14278 & n26104 ) ;
  assign n26210 = ( n817 & ~n17268 ) | ( n817 & n26209 ) | ( ~n17268 & n26209 ) ;
  assign n26211 = n8652 & n24374 ;
  assign n26212 = n22670 & n26211 ;
  assign n26213 = n22944 ^ n2695 ^ n1819 ;
  assign n26214 = n26213 ^ n16536 ^ n9001 ;
  assign n26215 = n26214 ^ n14908 ^ n5004 ;
  assign n26216 = ~n13888 & n26215 ;
  assign n26217 = ~n5326 & n26216 ;
  assign n26218 = n26217 ^ n19993 ^ 1'b0 ;
  assign n26219 = n10698 | n14903 ;
  assign n26220 = n23327 ^ n9360 ^ n3750 ;
  assign n26221 = ( ~n5110 & n5657 ) | ( ~n5110 & n26220 ) | ( n5657 & n26220 ) ;
  assign n26223 = n15541 ^ n4596 ^ n1879 ;
  assign n26222 = ( ~n2538 & n10065 ) | ( ~n2538 & n23746 ) | ( n10065 & n23746 ) ;
  assign n26224 = n26223 ^ n26222 ^ n6427 ;
  assign n26225 = ( n12790 & n22139 ) | ( n12790 & n24128 ) | ( n22139 & n24128 ) ;
  assign n26226 = n24853 ^ n18698 ^ n4670 ;
  assign n26227 = ~n7388 & n12558 ;
  assign n26228 = ~n26226 & n26227 ;
  assign n26229 = ( n12106 & n13494 ) | ( n12106 & ~n26228 ) | ( n13494 & ~n26228 ) ;
  assign n26230 = ( n1052 & ~n22150 ) | ( n1052 & n26229 ) | ( ~n22150 & n26229 ) ;
  assign n26231 = n26230 ^ n9149 ^ n5385 ;
  assign n26232 = n11337 ^ n7129 ^ 1'b0 ;
  assign n26233 = ( n16101 & ~n22999 ) | ( n16101 & n26232 ) | ( ~n22999 & n26232 ) ;
  assign n26234 = ( ~n2983 & n10117 ) | ( ~n2983 & n10630 ) | ( n10117 & n10630 ) ;
  assign n26235 = ( ~n8662 & n24382 ) | ( ~n8662 & n26234 ) | ( n24382 & n26234 ) ;
  assign n26236 = n3519 ^ x19 ^ 1'b0 ;
  assign n26237 = n26235 & n26236 ;
  assign n26239 = n21074 ^ n14045 ^ n9523 ;
  assign n26238 = n2343 | n16147 ;
  assign n26240 = n26239 ^ n26238 ^ 1'b0 ;
  assign n26241 = ~n3745 & n26240 ;
  assign n26242 = n8098 & n26241 ;
  assign n26243 = n7724 ^ n6947 ^ n4176 ;
  assign n26244 = n26243 ^ n13935 ^ n6916 ;
  assign n26245 = ( n11700 & ~n24374 ) | ( n11700 & n26244 ) | ( ~n24374 & n26244 ) ;
  assign n26246 = n24598 ^ n23050 ^ 1'b0 ;
  assign n26247 = n1694 & n26246 ;
  assign n26248 = ( ~n18885 & n19372 ) | ( ~n18885 & n26247 ) | ( n19372 & n26247 ) ;
  assign n26249 = n24894 ^ n8247 ^ n3104 ;
  assign n26250 = n18691 ^ n12236 ^ n7717 ;
  assign n26251 = n26250 ^ n22078 ^ n18108 ;
  assign n26252 = n18933 ^ n10704 ^ n7498 ;
  assign n26253 = ( ~n6686 & n18640 ) | ( ~n6686 & n26252 ) | ( n18640 & n26252 ) ;
  assign n26254 = n9466 ^ x76 ^ 1'b0 ;
  assign n26255 = n3364 | n26254 ;
  assign n26256 = n17894 | n26255 ;
  assign n26257 = n13165 & n25802 ;
  assign n26258 = n26257 ^ n26055 ^ 1'b0 ;
  assign n26259 = n21948 ^ n9322 ^ n1467 ;
  assign n26260 = n26259 ^ n22512 ^ n4717 ;
  assign n26262 = n11933 ^ n7769 ^ n3528 ;
  assign n26261 = ( n9883 & ~n12605 ) | ( n9883 & n21423 ) | ( ~n12605 & n21423 ) ;
  assign n26263 = n26262 ^ n26261 ^ n12070 ;
  assign n26264 = n18760 ^ n9249 ^ n6109 ;
  assign n26265 = ~n20956 & n26113 ;
  assign n26266 = ~n7759 & n26265 ;
  assign n26267 = ( n17025 & ~n26264 ) | ( n17025 & n26266 ) | ( ~n26264 & n26266 ) ;
  assign n26268 = ( n5235 & ~n16817 ) | ( n5235 & n17060 ) | ( ~n16817 & n17060 ) ;
  assign n26269 = ( n7283 & n12521 ) | ( n7283 & n25382 ) | ( n12521 & n25382 ) ;
  assign n26270 = n26269 ^ n9232 ^ n2342 ;
  assign n26271 = n26270 ^ n5578 ^ 1'b0 ;
  assign n26272 = ( ~n1162 & n1677 ) | ( ~n1162 & n15201 ) | ( n1677 & n15201 ) ;
  assign n26273 = n26272 ^ n15468 ^ n1429 ;
  assign n26274 = n26273 ^ n15587 ^ n13056 ;
  assign n26275 = n16628 ^ n12648 ^ n11800 ;
  assign n26276 = ~n22995 & n26275 ;
  assign n26277 = n26276 ^ n15258 ^ 1'b0 ;
  assign n26278 = n26277 ^ n17901 ^ n7522 ;
  assign n26279 = n10510 ^ n9833 ^ 1'b0 ;
  assign n26280 = n26279 ^ n12708 ^ n10469 ;
  assign n26281 = n26280 ^ n16188 ^ n13381 ;
  assign n26282 = ( n3427 & n24285 ) | ( n3427 & n25510 ) | ( n24285 & n25510 ) ;
  assign n26283 = n449 & n14867 ;
  assign n26284 = n26283 ^ n16140 ^ 1'b0 ;
  assign n26285 = n22392 & ~n26284 ;
  assign n26286 = n26285 ^ n11346 ^ 1'b0 ;
  assign n26289 = n14734 ^ n10560 ^ n1408 ;
  assign n26287 = ( n3044 & n9891 ) | ( n3044 & n13018 ) | ( n9891 & n13018 ) ;
  assign n26288 = n12738 | n26287 ;
  assign n26290 = n26289 ^ n26288 ^ 1'b0 ;
  assign n26291 = n26290 ^ n19847 ^ n145 ;
  assign n26292 = n839 & n4973 ;
  assign n26293 = n18787 & n26292 ;
  assign n26294 = ( n1940 & n26291 ) | ( n1940 & n26293 ) | ( n26291 & n26293 ) ;
  assign n26295 = ( ~n4087 & n6981 ) | ( ~n4087 & n26294 ) | ( n6981 & n26294 ) ;
  assign n26297 = n4474 | n19519 ;
  assign n26298 = n16288 & ~n26297 ;
  assign n26296 = n16753 ^ n9642 ^ n9043 ;
  assign n26299 = n26298 ^ n26296 ^ n4232 ;
  assign n26300 = ( n2492 & ~n3500 ) | ( n2492 & n6137 ) | ( ~n3500 & n6137 ) ;
  assign n26301 = n26300 ^ n11584 ^ n1059 ;
  assign n26302 = ( n9061 & n10055 ) | ( n9061 & n17481 ) | ( n10055 & n17481 ) ;
  assign n26303 = ( n7514 & ~n23411 ) | ( n7514 & n26302 ) | ( ~n23411 & n26302 ) ;
  assign n26304 = n1201 ^ n1137 ^ 1'b0 ;
  assign n26305 = ( n4694 & n6690 ) | ( n4694 & n26304 ) | ( n6690 & n26304 ) ;
  assign n26306 = n26305 ^ n19047 ^ n7755 ;
  assign n26308 = ( n2500 & n20615 ) | ( n2500 & n22479 ) | ( n20615 & n22479 ) ;
  assign n26307 = ( n7876 & ~n9889 ) | ( n7876 & n9981 ) | ( ~n9889 & n9981 ) ;
  assign n26309 = n26308 ^ n26307 ^ n15808 ;
  assign n26310 = ( n14714 & n21912 ) | ( n14714 & ~n26309 ) | ( n21912 & ~n26309 ) ;
  assign n26311 = n17108 ^ n12260 ^ n9449 ;
  assign n26312 = n19341 & ~n26311 ;
  assign n26313 = n17242 & n26312 ;
  assign n26314 = n22707 ^ n9896 ^ 1'b0 ;
  assign n26315 = n6853 | n26314 ;
  assign n26316 = ( ~n204 & n2124 ) | ( ~n204 & n5261 ) | ( n2124 & n5261 ) ;
  assign n26317 = n3031 | n18397 ;
  assign n26318 = ( n1623 & n8983 ) | ( n1623 & n26317 ) | ( n8983 & n26317 ) ;
  assign n26319 = n8754 ^ n5088 ^ n3815 ;
  assign n26320 = n2880 ^ n2747 ^ n1847 ;
  assign n26321 = n11934 & ~n20700 ;
  assign n26322 = ~n9484 & n26321 ;
  assign n26323 = ( n26319 & n26320 ) | ( n26319 & ~n26322 ) | ( n26320 & ~n26322 ) ;
  assign n26324 = n15439 ^ n3719 ^ n944 ;
  assign n26325 = ( n8702 & ~n12231 ) | ( n8702 & n26324 ) | ( ~n12231 & n26324 ) ;
  assign n26326 = n10234 ^ n2037 ^ n1150 ;
  assign n26327 = ( n23101 & ~n26325 ) | ( n23101 & n26326 ) | ( ~n26325 & n26326 ) ;
  assign n26328 = n10619 ^ n2858 ^ 1'b0 ;
  assign n26329 = ( ~n3648 & n8682 ) | ( ~n3648 & n23698 ) | ( n8682 & n23698 ) ;
  assign n26330 = ( n2580 & ~n26328 ) | ( n2580 & n26329 ) | ( ~n26328 & n26329 ) ;
  assign n26331 = n26330 ^ n24439 ^ 1'b0 ;
  assign n26332 = ( ~n2265 & n4751 ) | ( ~n2265 & n6265 ) | ( n4751 & n6265 ) ;
  assign n26333 = ( n4717 & n4801 ) | ( n4717 & n11039 ) | ( n4801 & n11039 ) ;
  assign n26334 = n26333 ^ n7622 ^ n3602 ;
  assign n26335 = n4426 & ~n7470 ;
  assign n26336 = n7991 ^ n5887 ^ 1'b0 ;
  assign n26337 = ( n8906 & n26335 ) | ( n8906 & n26336 ) | ( n26335 & n26336 ) ;
  assign n26338 = ( n11502 & ~n14403 ) | ( n11502 & n26337 ) | ( ~n14403 & n26337 ) ;
  assign n26342 = n8603 ^ n4642 ^ n4045 ;
  assign n26343 = n26342 ^ n9602 ^ n2004 ;
  assign n26339 = ( n508 & n13363 ) | ( n508 & n19802 ) | ( n13363 & n19802 ) ;
  assign n26340 = ( ~n12655 & n25760 ) | ( ~n12655 & n26339 ) | ( n25760 & n26339 ) ;
  assign n26341 = ( n3259 & ~n12567 ) | ( n3259 & n26340 ) | ( ~n12567 & n26340 ) ;
  assign n26344 = n26343 ^ n26341 ^ n8104 ;
  assign n26345 = n8059 ^ n7761 ^ 1'b0 ;
  assign n26346 = ( n5124 & ~n14542 ) | ( n5124 & n26345 ) | ( ~n14542 & n26345 ) ;
  assign n26347 = n698 & n16866 ;
  assign n26349 = n1562 & n9549 ;
  assign n26348 = n18876 ^ n14442 ^ n212 ;
  assign n26350 = n26349 ^ n26348 ^ n4755 ;
  assign n26354 = n17880 ^ n9863 ^ n5893 ;
  assign n26352 = n347 & ~n19544 ;
  assign n26353 = ( n7010 & n19047 ) | ( n7010 & n26352 ) | ( n19047 & n26352 ) ;
  assign n26351 = ( n6143 & ~n16734 ) | ( n6143 & n20707 ) | ( ~n16734 & n20707 ) ;
  assign n26355 = n26354 ^ n26353 ^ n26351 ;
  assign n26356 = ( n9138 & ~n18729 ) | ( n9138 & n26355 ) | ( ~n18729 & n26355 ) ;
  assign n26357 = ~n17598 & n22493 ;
  assign n26358 = n10924 | n22585 ;
  assign n26359 = ( n25686 & n26357 ) | ( n25686 & n26358 ) | ( n26357 & n26358 ) ;
  assign n26360 = n20001 ^ n6547 ^ 1'b0 ;
  assign n26361 = n16973 ^ n789 ^ 1'b0 ;
  assign n26362 = n26360 & n26361 ;
  assign n26363 = n12611 | n15127 ;
  assign n26364 = n15424 & ~n26363 ;
  assign n26365 = ( ~n4499 & n12006 ) | ( ~n4499 & n19794 ) | ( n12006 & n19794 ) ;
  assign n26366 = n10723 & n15972 ;
  assign n26367 = n26366 ^ n11035 ^ 1'b0 ;
  assign n26368 = n26367 ^ n11491 ^ n288 ;
  assign n26370 = n12433 | n17008 ;
  assign n26371 = n26370 ^ n24647 ^ 1'b0 ;
  assign n26369 = ( n2860 & ~n7547 ) | ( n2860 & n23158 ) | ( ~n7547 & n23158 ) ;
  assign n26372 = n26371 ^ n26369 ^ n14446 ;
  assign n26373 = n22414 ^ n16408 ^ n1913 ;
  assign n26374 = n6736 ^ n3467 ^ n2487 ;
  assign n26375 = ( n5353 & n10395 ) | ( n5353 & ~n26374 ) | ( n10395 & ~n26374 ) ;
  assign n26376 = n18535 ^ n14472 ^ 1'b0 ;
  assign n26377 = ~n18613 & n26376 ;
  assign n26378 = n26377 ^ n26358 ^ n7078 ;
  assign n26379 = n13708 ^ n1427 ^ 1'b0 ;
  assign n26380 = n15665 & n26379 ;
  assign n26381 = n26380 ^ n12791 ^ 1'b0 ;
  assign n26382 = n9538 | n26381 ;
  assign n26383 = ( ~n3379 & n8340 ) | ( ~n3379 & n14413 ) | ( n8340 & n14413 ) ;
  assign n26384 = n26383 ^ n12500 ^ 1'b0 ;
  assign n26385 = ~n13311 & n26384 ;
  assign n26386 = n22106 ^ n2414 ^ n1260 ;
  assign n26387 = n15628 ^ n3489 ^ n3429 ;
  assign n26388 = ( n16163 & ~n26386 ) | ( n16163 & n26387 ) | ( ~n26386 & n26387 ) ;
  assign n26389 = ( ~n8980 & n9647 ) | ( ~n8980 & n22550 ) | ( n9647 & n22550 ) ;
  assign n26390 = ( n3461 & n4860 ) | ( n3461 & n14817 ) | ( n4860 & n14817 ) ;
  assign n26391 = ( n26377 & ~n26389 ) | ( n26377 & n26390 ) | ( ~n26389 & n26390 ) ;
  assign n26392 = ( n16835 & ~n19178 ) | ( n16835 & n26391 ) | ( ~n19178 & n26391 ) ;
  assign n26393 = ( n1814 & n3180 ) | ( n1814 & ~n15670 ) | ( n3180 & ~n15670 ) ;
  assign n26394 = ( n5761 & ~n10271 ) | ( n5761 & n10656 ) | ( ~n10271 & n10656 ) ;
  assign n26395 = n26394 ^ n4135 ^ n3111 ;
  assign n26396 = n26395 ^ n21367 ^ n10539 ;
  assign n26397 = ( ~n3719 & n3907 ) | ( ~n3719 & n24349 ) | ( n3907 & n24349 ) ;
  assign n26398 = n26397 ^ n25766 ^ 1'b0 ;
  assign n26399 = ~n15493 & n26398 ;
  assign n26400 = ( n10179 & n26396 ) | ( n10179 & ~n26399 ) | ( n26396 & ~n26399 ) ;
  assign n26401 = ( n6592 & n26393 ) | ( n6592 & ~n26400 ) | ( n26393 & ~n26400 ) ;
  assign n26402 = n23893 ^ n19366 ^ n18031 ;
  assign n26403 = n14603 ^ n10921 ^ n5151 ;
  assign n26404 = n2629 | n11733 ;
  assign n26405 = n1940 & n11392 ;
  assign n26406 = ( n4748 & ~n18046 ) | ( n4748 & n26405 ) | ( ~n18046 & n26405 ) ;
  assign n26407 = ( n12032 & n26404 ) | ( n12032 & n26406 ) | ( n26404 & n26406 ) ;
  assign n26408 = ( n10971 & n18432 ) | ( n10971 & ~n26407 ) | ( n18432 & ~n26407 ) ;
  assign n26409 = n2404 & n9400 ;
  assign n26410 = n26409 ^ n12015 ^ 1'b0 ;
  assign n26411 = n9991 ^ n609 ^ 1'b0 ;
  assign n26412 = n26410 & ~n26411 ;
  assign n26413 = ( n3623 & ~n7755 ) | ( n3623 & n23108 ) | ( ~n7755 & n23108 ) ;
  assign n26414 = ( n2283 & n25813 ) | ( n2283 & n26413 ) | ( n25813 & n26413 ) ;
  assign n26415 = n25793 ^ n16396 ^ n2336 ;
  assign n26416 = ( ~n1401 & n4670 ) | ( ~n1401 & n9947 ) | ( n4670 & n9947 ) ;
  assign n26417 = n2823 & ~n9297 ;
  assign n26418 = n11147 ^ n8327 ^ n7161 ;
  assign n26419 = ( n4842 & n26417 ) | ( n4842 & ~n26418 ) | ( n26417 & ~n26418 ) ;
  assign n26420 = ( ~n1687 & n17235 ) | ( ~n1687 & n21509 ) | ( n17235 & n21509 ) ;
  assign n26421 = n26420 ^ n6252 ^ n1786 ;
  assign n26422 = ( n5084 & ~n8519 ) | ( n5084 & n17578 ) | ( ~n8519 & n17578 ) ;
  assign n26423 = ~n5691 & n26422 ;
  assign n26424 = n26423 ^ n313 ^ 1'b0 ;
  assign n26425 = ( n1684 & ~n26421 ) | ( n1684 & n26424 ) | ( ~n26421 & n26424 ) ;
  assign n26426 = n13746 & n17379 ;
  assign n26428 = n9603 ^ n2417 ^ 1'b0 ;
  assign n26427 = n9197 ^ n4304 ^ n1306 ;
  assign n26429 = n26428 ^ n26427 ^ n23481 ;
  assign n26430 = ~n5035 & n7120 ;
  assign n26431 = n26430 ^ n15309 ^ 1'b0 ;
  assign n26432 = ( n1006 & n7671 ) | ( n1006 & n19473 ) | ( n7671 & n19473 ) ;
  assign n26433 = ( n2670 & n5654 ) | ( n2670 & ~n25772 ) | ( n5654 & ~n25772 ) ;
  assign n26434 = n21765 ^ n486 ^ 1'b0 ;
  assign n26435 = n8618 & ~n18505 ;
  assign n26436 = n16471 & n26435 ;
  assign n26437 = ( n21231 & n26434 ) | ( n21231 & n26436 ) | ( n26434 & n26436 ) ;
  assign n26438 = ( n2396 & n19452 ) | ( n2396 & ~n19510 ) | ( n19452 & ~n19510 ) ;
  assign n26439 = n8304 ^ n989 ^ x40 ;
  assign n26440 = n26439 ^ n14914 ^ n12369 ;
  assign n26441 = n26440 ^ n6521 ^ n769 ;
  assign n26442 = ( n20124 & n26438 ) | ( n20124 & n26441 ) | ( n26438 & n26441 ) ;
  assign n26443 = ( n10668 & n16013 ) | ( n10668 & ~n21082 ) | ( n16013 & ~n21082 ) ;
  assign n26444 = ( ~n4801 & n8807 ) | ( ~n4801 & n26443 ) | ( n8807 & n26443 ) ;
  assign n26445 = n8996 ^ n4850 ^ n2552 ;
  assign n26446 = n20712 ^ n6556 ^ n3293 ;
  assign n26447 = ( ~n7449 & n11726 ) | ( ~n7449 & n15676 ) | ( n11726 & n15676 ) ;
  assign n26448 = ( n26445 & n26446 ) | ( n26445 & n26447 ) | ( n26446 & n26447 ) ;
  assign n26449 = ~n4650 & n12642 ;
  assign n26450 = n26449 ^ n22649 ^ n17940 ;
  assign n26451 = n19540 ^ n3018 ^ 1'b0 ;
  assign n26452 = n4130 & ~n26451 ;
  assign n26453 = n19991 ^ n12517 ^ n11069 ;
  assign n26454 = ( ~n14432 & n26452 ) | ( ~n14432 & n26453 ) | ( n26452 & n26453 ) ;
  assign n26455 = ( n465 & ~n1417 ) | ( n465 & n25873 ) | ( ~n1417 & n25873 ) ;
  assign n26456 = n556 & ~n6281 ;
  assign n26457 = ~n26455 & n26456 ;
  assign n26458 = n16563 ^ n14356 ^ n2842 ;
  assign n26459 = n10773 ^ n10760 ^ n2276 ;
  assign n26460 = n26459 ^ n8884 ^ 1'b0 ;
  assign n26461 = ( n2119 & n15800 ) | ( n2119 & n25649 ) | ( n15800 & n25649 ) ;
  assign n26462 = ( ~n671 & n6122 ) | ( ~n671 & n26461 ) | ( n6122 & n26461 ) ;
  assign n26463 = n25766 ^ n6406 ^ n4064 ;
  assign n26464 = n26463 ^ n15902 ^ n7081 ;
  assign n26465 = ( n914 & n6575 ) | ( n914 & ~n15276 ) | ( n6575 & ~n15276 ) ;
  assign n26466 = n3416 ^ n2467 ^ 1'b0 ;
  assign n26467 = ~n439 & n19438 ;
  assign n26468 = n26467 ^ n15535 ^ 1'b0 ;
  assign n26469 = n16044 ^ n8821 ^ n6598 ;
  assign n26470 = ( ~n1984 & n19014 ) | ( ~n1984 & n24579 ) | ( n19014 & n24579 ) ;
  assign n26471 = ( n1409 & n1476 ) | ( n1409 & ~n16427 ) | ( n1476 & ~n16427 ) ;
  assign n26477 = n2183 & ~n11889 ;
  assign n26472 = n6134 ^ n2091 ^ 1'b0 ;
  assign n26473 = n26472 ^ n7576 ^ n6148 ;
  assign n26474 = n26473 ^ n4764 ^ 1'b0 ;
  assign n26475 = n26474 ^ n8911 ^ 1'b0 ;
  assign n26476 = n26475 ^ n21046 ^ n9853 ;
  assign n26478 = n26477 ^ n26476 ^ n22385 ;
  assign n26479 = n20456 ^ n19806 ^ n19430 ;
  assign n26480 = n21597 ^ n14333 ^ n10581 ;
  assign n26482 = n10204 ^ n2034 ^ n1838 ;
  assign n26481 = n19825 & n20816 ;
  assign n26483 = n26482 ^ n26481 ^ 1'b0 ;
  assign n26484 = n22322 ^ n1608 ^ 1'b0 ;
  assign n26485 = n19476 & n26484 ;
  assign n26486 = n26485 ^ n19149 ^ n2026 ;
  assign n26487 = n21719 ^ n13248 ^ n1340 ;
  assign n26488 = ~n8707 & n10653 ;
  assign n26489 = ~n10621 & n11437 ;
  assign n26490 = n5472 & n26489 ;
  assign n26491 = n26488 & ~n26490 ;
  assign n26492 = n2988 & n26491 ;
  assign n26493 = n23799 & ~n26492 ;
  assign n26494 = ( ~n201 & n532 ) | ( ~n201 & n15558 ) | ( n532 & n15558 ) ;
  assign n26495 = n19997 ^ n16997 ^ n13987 ;
  assign n26496 = ( n1047 & n7771 ) | ( n1047 & n26495 ) | ( n7771 & n26495 ) ;
  assign n26497 = n13282 ^ n9922 ^ n4162 ;
  assign n26498 = n11305 ^ n4014 ^ n1052 ;
  assign n26499 = n3806 | n18862 ;
  assign n26500 = n24826 | n26499 ;
  assign n26501 = n4124 ^ n2636 ^ 1'b0 ;
  assign n26502 = n15442 | n26501 ;
  assign n26503 = ( ~n7907 & n9435 ) | ( ~n7907 & n24824 ) | ( n9435 & n24824 ) ;
  assign n26504 = n3426 & ~n18793 ;
  assign n26505 = n26504 ^ n23878 ^ 1'b0 ;
  assign n26506 = n17075 ^ n12389 ^ n10708 ;
  assign n26507 = ( ~n26503 & n26505 ) | ( ~n26503 & n26506 ) | ( n26505 & n26506 ) ;
  assign n26508 = n13121 ^ n7667 ^ n3771 ;
  assign n26509 = n26508 ^ n19368 ^ 1'b0 ;
  assign n26510 = ( n3994 & n19856 ) | ( n3994 & n26509 ) | ( n19856 & n26509 ) ;
  assign n26511 = n6821 | n26510 ;
  assign n26517 = n8809 ^ n6896 ^ n2228 ;
  assign n26513 = n7658 ^ n4871 ^ n3469 ;
  assign n26512 = n15466 & ~n25354 ;
  assign n26514 = n26513 ^ n26512 ^ 1'b0 ;
  assign n26515 = n2404 & n26514 ;
  assign n26516 = n26515 ^ n2265 ^ 1'b0 ;
  assign n26518 = n26517 ^ n26516 ^ n24677 ;
  assign n26519 = ( n422 & n11286 ) | ( n422 & ~n12077 ) | ( n11286 & ~n12077 ) ;
  assign n26520 = ( n2667 & n10073 ) | ( n2667 & n26519 ) | ( n10073 & n26519 ) ;
  assign n26521 = n16612 & n17578 ;
  assign n26522 = ( n5331 & n11581 ) | ( n5331 & n15254 ) | ( n11581 & n15254 ) ;
  assign n26523 = ( n11168 & n26521 ) | ( n11168 & ~n26522 ) | ( n26521 & ~n26522 ) ;
  assign n26524 = ( n1741 & n7176 ) | ( n1741 & ~n9713 ) | ( n7176 & ~n9713 ) ;
  assign n26525 = n26524 ^ n25631 ^ n4623 ;
  assign n26526 = ( n4452 & n7665 ) | ( n4452 & ~n16533 ) | ( n7665 & ~n16533 ) ;
  assign n26527 = n26526 ^ n19624 ^ n10139 ;
  assign n26534 = ~n2132 & n14187 ;
  assign n26531 = n14062 ^ n6348 ^ n805 ;
  assign n26532 = ( n5429 & n7753 ) | ( n5429 & ~n26531 ) | ( n7753 & ~n26531 ) ;
  assign n26533 = n26532 ^ n1806 ^ n465 ;
  assign n26528 = n23175 ^ n18857 ^ 1'b0 ;
  assign n26529 = ~n10971 & n26528 ;
  assign n26530 = ( ~n6436 & n22444 ) | ( ~n6436 & n26529 ) | ( n22444 & n26529 ) ;
  assign n26535 = n26534 ^ n26533 ^ n26530 ;
  assign n26536 = n11474 ^ n6398 ^ n4519 ;
  assign n26537 = n7467 ^ n2444 ^ n582 ;
  assign n26538 = ( n1928 & n26536 ) | ( n1928 & ~n26537 ) | ( n26536 & ~n26537 ) ;
  assign n26539 = ( n4948 & n18957 ) | ( n4948 & ~n23190 ) | ( n18957 & ~n23190 ) ;
  assign n26540 = n17778 ^ n10531 ^ n7122 ;
  assign n26541 = ( n793 & ~n14263 ) | ( n793 & n18661 ) | ( ~n14263 & n18661 ) ;
  assign n26542 = ( n8311 & n21260 ) | ( n8311 & ~n26541 ) | ( n21260 & ~n26541 ) ;
  assign n26543 = ( n14803 & n26540 ) | ( n14803 & n26542 ) | ( n26540 & n26542 ) ;
  assign n26544 = ( n2524 & n3652 ) | ( n2524 & n23632 ) | ( n3652 & n23632 ) ;
  assign n26545 = n21433 ^ n9717 ^ 1'b0 ;
  assign n26546 = n22535 | n26545 ;
  assign n26547 = n10572 ^ n7170 ^ n6665 ;
  assign n26548 = n23765 ^ n7489 ^ 1'b0 ;
  assign n26549 = ~n26547 & n26548 ;
  assign n26550 = n13481 ^ n10020 ^ n8280 ;
  assign n26551 = n17594 ^ n6065 ^ n255 ;
  assign n26552 = ( n512 & ~n7174 ) | ( n512 & n18113 ) | ( ~n7174 & n18113 ) ;
  assign n26553 = n22854 ^ n11672 ^ n7709 ;
  assign n26554 = ( ~n1380 & n3627 ) | ( ~n1380 & n8100 ) | ( n3627 & n8100 ) ;
  assign n26555 = n26554 ^ n15089 ^ n11624 ;
  assign n26556 = n26555 ^ n24235 ^ n20275 ;
  assign n26557 = n20431 ^ n14554 ^ n6444 ;
  assign n26561 = ( n6073 & n8490 ) | ( n6073 & ~n13902 ) | ( n8490 & ~n13902 ) ;
  assign n26558 = n19544 ^ n5528 ^ 1'b0 ;
  assign n26559 = n18857 & ~n26558 ;
  assign n26560 = ~n4440 & n26559 ;
  assign n26562 = n26561 ^ n26560 ^ n21621 ;
  assign n26563 = n20616 ^ n14725 ^ n3541 ;
  assign n26564 = ( n26557 & n26562 ) | ( n26557 & n26563 ) | ( n26562 & n26563 ) ;
  assign n26565 = n9949 ^ n8510 ^ n3179 ;
  assign n26566 = n4372 ^ n1754 ^ n750 ;
  assign n26567 = ( n2595 & n9747 ) | ( n2595 & ~n26566 ) | ( n9747 & ~n26566 ) ;
  assign n26568 = n26567 ^ n8850 ^ 1'b0 ;
  assign n26569 = n26568 ^ n3583 ^ n1179 ;
  assign n26570 = n21803 ^ n19838 ^ n5206 ;
  assign n26571 = n26570 ^ n12716 ^ 1'b0 ;
  assign n26572 = n8242 ^ n5246 ^ 1'b0 ;
  assign n26573 = ( n9328 & n17637 ) | ( n9328 & ~n26572 ) | ( n17637 & ~n26572 ) ;
  assign n26574 = ( n7314 & n12462 ) | ( n7314 & n13526 ) | ( n12462 & n13526 ) ;
  assign n26575 = ( n8986 & n11728 ) | ( n8986 & ~n14174 ) | ( n11728 & ~n14174 ) ;
  assign n26576 = n26575 ^ n26490 ^ n20064 ;
  assign n26577 = ( n882 & n7094 ) | ( n882 & n20587 ) | ( n7094 & n20587 ) ;
  assign n26578 = n26577 ^ n15084 ^ n251 ;
  assign n26579 = n26578 ^ n12786 ^ n3577 ;
  assign n26585 = ~n4782 & n26561 ;
  assign n26580 = ( n7691 & ~n10936 ) | ( n7691 & n21969 ) | ( ~n10936 & n21969 ) ;
  assign n26581 = n26580 ^ n22555 ^ n1074 ;
  assign n26582 = n17721 | n26581 ;
  assign n26583 = n6566 & ~n26582 ;
  assign n26584 = n26583 ^ n17809 ^ n14167 ;
  assign n26586 = n26585 ^ n26584 ^ n14554 ;
  assign n26587 = ( n9453 & n17287 ) | ( n9453 & ~n19544 ) | ( n17287 & ~n19544 ) ;
  assign n26588 = ( ~n1813 & n12837 ) | ( ~n1813 & n26587 ) | ( n12837 & n26587 ) ;
  assign n26589 = ( n3480 & n20816 ) | ( n3480 & ~n26588 ) | ( n20816 & ~n26588 ) ;
  assign n26590 = ( ~n9090 & n11548 ) | ( ~n9090 & n11971 ) | ( n11548 & n11971 ) ;
  assign n26591 = n12273 & n18703 ;
  assign n26592 = n26590 & n26591 ;
  assign n26593 = ( n17673 & ~n25353 ) | ( n17673 & n26592 ) | ( ~n25353 & n26592 ) ;
  assign n26594 = ( n3097 & ~n3482 ) | ( n3097 & n7787 ) | ( ~n3482 & n7787 ) ;
  assign n26595 = n26594 ^ n982 ^ n414 ;
  assign n26596 = n26595 ^ n16075 ^ n671 ;
  assign n26597 = ( n2964 & n15395 ) | ( n2964 & n25491 ) | ( n15395 & n25491 ) ;
  assign n26598 = n23611 ^ n13993 ^ n4596 ;
  assign n26599 = ( ~n1506 & n21244 ) | ( ~n1506 & n26598 ) | ( n21244 & n26598 ) ;
  assign n26600 = ( n699 & ~n1331 ) | ( n699 & n18097 ) | ( ~n1331 & n18097 ) ;
  assign n26601 = n16073 ^ n9590 ^ n6420 ;
  assign n26611 = ( ~n9738 & n10015 ) | ( ~n9738 & n21480 ) | ( n10015 & n21480 ) ;
  assign n26603 = ( ~n1825 & n14687 ) | ( ~n1825 & n16702 ) | ( n14687 & n16702 ) ;
  assign n26602 = n3837 & ~n6336 ;
  assign n26604 = n26603 ^ n26602 ^ 1'b0 ;
  assign n26608 = n23144 ^ n14160 ^ n1727 ;
  assign n26605 = ( ~n5847 & n7607 ) | ( ~n5847 & n12696 ) | ( n7607 & n12696 ) ;
  assign n26606 = ( n11604 & n18299 ) | ( n11604 & ~n26605 ) | ( n18299 & ~n26605 ) ;
  assign n26607 = n26606 ^ n19089 ^ n15439 ;
  assign n26609 = n26608 ^ n26607 ^ n5902 ;
  assign n26610 = ( n4834 & n26604 ) | ( n4834 & ~n26609 ) | ( n26604 & ~n26609 ) ;
  assign n26612 = n26611 ^ n26610 ^ n4527 ;
  assign n26617 = ( ~n3000 & n17008 ) | ( ~n3000 & n17448 ) | ( n17008 & n17448 ) ;
  assign n26613 = ~n2819 & n14389 ;
  assign n26614 = n12595 ^ n5989 ^ 1'b0 ;
  assign n26615 = ( n11657 & n26613 ) | ( n11657 & n26614 ) | ( n26613 & n26614 ) ;
  assign n26616 = ~n21907 & n26615 ;
  assign n26618 = n26617 ^ n26616 ^ 1'b0 ;
  assign n26621 = n9229 & ~n9392 ;
  assign n26622 = n26621 ^ n6373 ^ 1'b0 ;
  assign n26623 = n5622 & n9729 ;
  assign n26624 = ~n26622 & n26623 ;
  assign n26625 = n26624 ^ n11000 ^ n7349 ;
  assign n26619 = n14639 ^ n388 ^ 1'b0 ;
  assign n26620 = n5816 & ~n26619 ;
  assign n26626 = n26625 ^ n26620 ^ n8172 ;
  assign n26627 = n19701 ^ n16983 ^ n12804 ;
  assign n26628 = n13682 ^ n10076 ^ n3507 ;
  assign n26629 = ( ~n7382 & n20435 ) | ( ~n7382 & n26628 ) | ( n20435 & n26628 ) ;
  assign n26631 = n25076 ^ n13127 ^ 1'b0 ;
  assign n26632 = ~n1884 & n26631 ;
  assign n26630 = n24019 ^ n16380 ^ n1932 ;
  assign n26633 = n26632 ^ n26630 ^ n26540 ;
  assign n26634 = n19917 ^ n10394 ^ n3583 ;
  assign n26635 = n4544 & n26634 ;
  assign n26636 = ( n12379 & n26633 ) | ( n12379 & ~n26635 ) | ( n26633 & ~n26635 ) ;
  assign n26637 = ~n14157 & n16402 ;
  assign n26638 = ( n4246 & ~n15445 ) | ( n4246 & n26637 ) | ( ~n15445 & n26637 ) ;
  assign n26641 = ( n4500 & ~n6192 ) | ( n4500 & n17763 ) | ( ~n6192 & n17763 ) ;
  assign n26640 = ( n5857 & n18411 ) | ( n5857 & n18619 ) | ( n18411 & n18619 ) ;
  assign n26639 = ~n6395 & n18971 ;
  assign n26642 = n26641 ^ n26640 ^ n26639 ;
  assign n26643 = n19551 ^ n18468 ^ n10654 ;
  assign n26644 = n23533 ^ n3696 ^ 1'b0 ;
  assign n26645 = ~n9339 & n26644 ;
  assign n26646 = ( x91 & n7556 ) | ( x91 & n11936 ) | ( n7556 & n11936 ) ;
  assign n26647 = n9122 & n13248 ;
  assign n26648 = n26646 & n26647 ;
  assign n26649 = ( n788 & ~n4748 ) | ( n788 & n13882 ) | ( ~n4748 & n13882 ) ;
  assign n26650 = n26649 ^ n16136 ^ n8278 ;
  assign n26651 = n20988 ^ n2074 ^ n1722 ;
  assign n26652 = ~n1076 & n7968 ;
  assign n26653 = ~n967 & n26652 ;
  assign n26654 = n23490 ^ n10822 ^ n490 ;
  assign n26655 = ~n26374 & n26654 ;
  assign n26656 = n26653 & n26655 ;
  assign n26657 = ( n8367 & ~n11956 ) | ( n8367 & n26656 ) | ( ~n11956 & n26656 ) ;
  assign n26658 = n21436 ^ n14700 ^ n4497 ;
  assign n26659 = ( n4110 & n8022 ) | ( n4110 & n23809 ) | ( n8022 & n23809 ) ;
  assign n26660 = ( n6966 & n13353 ) | ( n6966 & ~n26659 ) | ( n13353 & ~n26659 ) ;
  assign n26661 = ( ~n962 & n1776 ) | ( ~n962 & n8320 ) | ( n1776 & n8320 ) ;
  assign n26662 = ( n2518 & n15076 ) | ( n2518 & ~n22859 ) | ( n15076 & ~n22859 ) ;
  assign n26663 = n26662 ^ n1626 ^ 1'b0 ;
  assign n26664 = n12580 & ~n26663 ;
  assign n26665 = n26664 ^ n7759 ^ n6587 ;
  assign n26666 = n17394 ^ n15087 ^ 1'b0 ;
  assign n26667 = ( n2038 & n18152 ) | ( n2038 & ~n25224 ) | ( n18152 & ~n25224 ) ;
  assign n26673 = n10590 ^ n8716 ^ n1896 ;
  assign n26672 = n7077 & n15407 ;
  assign n26674 = n26673 ^ n26672 ^ 1'b0 ;
  assign n26668 = ( n7074 & n18117 ) | ( n7074 & ~n20157 ) | ( n18117 & ~n20157 ) ;
  assign n26669 = n13290 & ~n26668 ;
  assign n26670 = ~n2920 & n26669 ;
  assign n26671 = n26670 ^ n24825 ^ n6107 ;
  assign n26675 = n26674 ^ n26671 ^ n23935 ;
  assign n26676 = n15753 ^ n2354 ^ 1'b0 ;
  assign n26677 = n4914 | n26676 ;
  assign n26678 = ( n2311 & n2938 ) | ( n2311 & n26677 ) | ( n2938 & n26677 ) ;
  assign n26679 = ~n2898 & n12170 ;
  assign n26680 = n26679 ^ n22724 ^ 1'b0 ;
  assign n26681 = n26680 ^ n7647 ^ n5416 ;
  assign n26682 = n14288 ^ n9390 ^ 1'b0 ;
  assign n26683 = ~n10643 & n26682 ;
  assign n26684 = n20837 ^ n13702 ^ n5917 ;
  assign n26685 = ( n7054 & n10913 ) | ( n7054 & ~n16271 ) | ( n10913 & ~n16271 ) ;
  assign n26686 = ( n734 & n1558 ) | ( n734 & n14609 ) | ( n1558 & n14609 ) ;
  assign n26687 = n14310 ^ n5773 ^ n3353 ;
  assign n26688 = n24686 ^ n9181 ^ n5576 ;
  assign n26689 = ~n16334 & n17897 ;
  assign n26690 = ~n26688 & n26689 ;
  assign n26691 = n26690 ^ n10945 ^ n5725 ;
  assign n26692 = n23701 ^ n16904 ^ n2658 ;
  assign n26693 = n26692 ^ n9533 ^ 1'b0 ;
  assign n26694 = n10726 ^ n9373 ^ n2737 ;
  assign n26695 = n26694 ^ n3134 ^ 1'b0 ;
  assign n26696 = n26693 & n26695 ;
  assign n26697 = ( n4802 & n7585 ) | ( n4802 & n14881 ) | ( n7585 & n14881 ) ;
  assign n26698 = ( n14484 & n15638 ) | ( n14484 & ~n20343 ) | ( n15638 & ~n20343 ) ;
  assign n26699 = n26698 ^ n16950 ^ n8302 ;
  assign n26700 = ( n10588 & ~n13629 ) | ( n10588 & n19895 ) | ( ~n13629 & n19895 ) ;
  assign n26701 = n26561 ^ n25249 ^ n4939 ;
  assign n26702 = n26701 ^ n20043 ^ n16719 ;
  assign n26703 = n2140 ^ n1052 ^ 1'b0 ;
  assign n26704 = ( n9486 & ~n22023 ) | ( n9486 & n26703 ) | ( ~n22023 & n26703 ) ;
  assign n26705 = ( n10190 & n14460 ) | ( n10190 & ~n24721 ) | ( n14460 & ~n24721 ) ;
  assign n26706 = n22617 ^ n19228 ^ n9416 ;
  assign n26707 = n15800 ^ n3988 ^ 1'b0 ;
  assign n26708 = n7246 & n26707 ;
  assign n26709 = n13868 & ~n19665 ;
  assign n26710 = n26709 ^ n19470 ^ 1'b0 ;
  assign n26711 = n16711 ^ n15372 ^ n4344 ;
  assign n26712 = n26711 ^ n17328 ^ n15339 ;
  assign n26713 = n17751 ^ n9319 ^ n5570 ;
  assign n26714 = n7341 ^ n4380 ^ n2498 ;
  assign n26715 = n26714 ^ n16070 ^ n5458 ;
  assign n26716 = ( ~n22895 & n26713 ) | ( ~n22895 & n26715 ) | ( n26713 & n26715 ) ;
  assign n26717 = ( ~n1308 & n7118 ) | ( ~n1308 & n16056 ) | ( n7118 & n16056 ) ;
  assign n26718 = n26717 ^ n7187 ^ 1'b0 ;
  assign n26720 = ( n1103 & n7193 ) | ( n1103 & ~n14516 ) | ( n7193 & ~n14516 ) ;
  assign n26719 = ( n3360 & n5680 ) | ( n3360 & ~n23633 ) | ( n5680 & ~n23633 ) ;
  assign n26721 = n26720 ^ n26719 ^ 1'b0 ;
  assign n26722 = n6686 & ~n26173 ;
  assign n26723 = n3020 & n7106 ;
  assign n26724 = n20795 & n26723 ;
  assign n26725 = n13561 ^ n12343 ^ 1'b0 ;
  assign n26726 = ( n2722 & n4836 ) | ( n2722 & ~n25305 ) | ( n4836 & ~n25305 ) ;
  assign n26727 = n26726 ^ n20795 ^ 1'b0 ;
  assign n26728 = n16199 ^ n7280 ^ n406 ;
  assign n26729 = n26728 ^ n13277 ^ n2219 ;
  assign n26730 = n18016 ^ n854 ^ 1'b0 ;
  assign n26731 = ( n591 & n3591 ) | ( n591 & ~n11205 ) | ( n3591 & ~n11205 ) ;
  assign n26732 = ( n10775 & ~n14896 ) | ( n10775 & n26731 ) | ( ~n14896 & n26731 ) ;
  assign n26733 = n10942 ^ n7305 ^ n4896 ;
  assign n26734 = ( n12435 & ~n15767 ) | ( n12435 & n26733 ) | ( ~n15767 & n26733 ) ;
  assign n26735 = ( n20868 & n26732 ) | ( n20868 & ~n26734 ) | ( n26732 & ~n26734 ) ;
  assign n26736 = ( n5011 & n10268 ) | ( n5011 & ~n24118 ) | ( n10268 & ~n24118 ) ;
  assign n26737 = ( n1176 & n5860 ) | ( n1176 & n15374 ) | ( n5860 & n15374 ) ;
  assign n26738 = ( n20467 & n26736 ) | ( n20467 & n26737 ) | ( n26736 & n26737 ) ;
  assign n26739 = ( n16597 & ~n23642 ) | ( n16597 & n26738 ) | ( ~n23642 & n26738 ) ;
  assign n26740 = n147 & n15547 ;
  assign n26741 = n26740 ^ n5296 ^ 1'b0 ;
  assign n26742 = n26741 ^ n10252 ^ n8842 ;
  assign n26743 = n18117 ^ n10108 ^ 1'b0 ;
  assign n26744 = n16691 & ~n26743 ;
  assign n26745 = ( n4077 & n10402 ) | ( n4077 & n23083 ) | ( n10402 & n23083 ) ;
  assign n26746 = n8629 & n26745 ;
  assign n26747 = n2185 & ~n8177 ;
  assign n26748 = n26746 & n26747 ;
  assign n26749 = n12292 ^ n9212 ^ n5918 ;
  assign n26750 = n26749 ^ n18432 ^ n16082 ;
  assign n26751 = ( ~n4598 & n10442 ) | ( ~n4598 & n11206 ) | ( n10442 & n11206 ) ;
  assign n26752 = ( ~n7088 & n23532 ) | ( ~n7088 & n26751 ) | ( n23532 & n26751 ) ;
  assign n26753 = n17181 ^ n6491 ^ n6454 ;
  assign n26754 = ( n3383 & ~n24812 ) | ( n3383 & n26753 ) | ( ~n24812 & n26753 ) ;
  assign n26755 = ( n2001 & n7749 ) | ( n2001 & n22005 ) | ( n7749 & n22005 ) ;
  assign n26756 = n26755 ^ n6890 ^ n1516 ;
  assign n26757 = n16744 | n26756 ;
  assign n26758 = ( ~n9941 & n13856 ) | ( ~n9941 & n16057 ) | ( n13856 & n16057 ) ;
  assign n26759 = ( ~n7723 & n10183 ) | ( ~n7723 & n13439 ) | ( n10183 & n13439 ) ;
  assign n26760 = ( ~n1026 & n5142 ) | ( ~n1026 & n26759 ) | ( n5142 & n26759 ) ;
  assign n26761 = ~n19809 & n26760 ;
  assign n26763 = ( n12800 & ~n17657 ) | ( n12800 & n18149 ) | ( ~n17657 & n18149 ) ;
  assign n26762 = n24169 ^ n19086 ^ n6976 ;
  assign n26764 = n26763 ^ n26762 ^ n3604 ;
  assign n26766 = ( n1941 & n8162 ) | ( n1941 & n8960 ) | ( n8162 & n8960 ) ;
  assign n26767 = n26766 ^ n2510 ^ 1'b0 ;
  assign n26768 = n22617 | n26767 ;
  assign n26765 = ( ~n8954 & n9962 ) | ( ~n8954 & n11555 ) | ( n9962 & n11555 ) ;
  assign n26769 = n26768 ^ n26765 ^ n742 ;
  assign n26771 = ( n3636 & n4224 ) | ( n3636 & ~n10230 ) | ( n4224 & ~n10230 ) ;
  assign n26772 = n26771 ^ n11087 ^ n3709 ;
  assign n26773 = n26772 ^ n14942 ^ n7310 ;
  assign n26774 = n26773 ^ n20482 ^ n17010 ;
  assign n26770 = ( n4390 & ~n13759 ) | ( n4390 & n18048 ) | ( ~n13759 & n18048 ) ;
  assign n26775 = n26774 ^ n26770 ^ n11318 ;
  assign n26776 = ( n1592 & n7148 ) | ( n1592 & ~n13242 ) | ( n7148 & ~n13242 ) ;
  assign n26777 = n18545 ^ n2689 ^ 1'b0 ;
  assign n26778 = n26776 | n26777 ;
  assign n26779 = n17658 ^ n14313 ^ n10077 ;
  assign n26781 = n16931 ^ n13243 ^ n7917 ;
  assign n26780 = n10940 ^ n5900 ^ n4717 ;
  assign n26782 = n26781 ^ n26780 ^ n15736 ;
  assign n26785 = n14119 ^ n12570 ^ n5783 ;
  assign n26783 = n4129 | n16352 ;
  assign n26784 = n26783 ^ n11413 ^ n2596 ;
  assign n26786 = n26785 ^ n26784 ^ n10408 ;
  assign n26787 = ( n18514 & n23656 ) | ( n18514 & n26510 ) | ( n23656 & n26510 ) ;
  assign n26788 = ( n9741 & n12433 ) | ( n9741 & n15423 ) | ( n12433 & n15423 ) ;
  assign n26789 = ( ~n3081 & n11088 ) | ( ~n3081 & n26788 ) | ( n11088 & n26788 ) ;
  assign n26790 = n1647 & ~n2206 ;
  assign n26791 = n26790 ^ n575 ^ 1'b0 ;
  assign n26792 = ( n555 & n9284 ) | ( n555 & ~n26791 ) | ( n9284 & ~n26791 ) ;
  assign n26793 = n26792 ^ n20296 ^ n15973 ;
  assign n26794 = n26793 ^ n7660 ^ n323 ;
  assign n26795 = n8966 ^ n6871 ^ n5775 ;
  assign n26796 = ( n3876 & n5078 ) | ( n3876 & ~n10672 ) | ( n5078 & ~n10672 ) ;
  assign n26797 = n19232 ^ n17494 ^ n3409 ;
  assign n26798 = ( ~n26795 & n26796 ) | ( ~n26795 & n26797 ) | ( n26796 & n26797 ) ;
  assign n26799 = n23509 ^ n1775 ^ 1'b0 ;
  assign n26800 = n22677 & n26799 ;
  assign n26801 = n24339 ^ n9639 ^ 1'b0 ;
  assign n26802 = n16423 | n26801 ;
  assign n26803 = ( n6843 & n8095 ) | ( n6843 & n20929 ) | ( n8095 & n20929 ) ;
  assign n26804 = n19524 ^ n17816 ^ 1'b0 ;
  assign n26805 = ( ~n4590 & n12051 ) | ( ~n4590 & n26804 ) | ( n12051 & n26804 ) ;
  assign n26806 = n7697 & n13851 ;
  assign n26807 = ( n8520 & ~n25255 ) | ( n8520 & n26806 ) | ( ~n25255 & n26806 ) ;
  assign n26808 = ( n3505 & n9949 ) | ( n3505 & n26807 ) | ( n9949 & n26807 ) ;
  assign n26814 = n15188 ^ n14862 ^ n152 ;
  assign n26811 = n16057 ^ n9462 ^ n1939 ;
  assign n26812 = ( ~n1376 & n2920 ) | ( ~n1376 & n26811 ) | ( n2920 & n26811 ) ;
  assign n26809 = n17934 ^ n7571 ^ 1'b0 ;
  assign n26810 = n26809 ^ n7171 ^ x32 ;
  assign n26813 = n26812 ^ n26810 ^ n13411 ;
  assign n26815 = n26814 ^ n26813 ^ n4162 ;
  assign n26816 = ( ~n7605 & n14315 ) | ( ~n7605 & n22600 ) | ( n14315 & n22600 ) ;
  assign n26817 = ( ~n826 & n13036 ) | ( ~n826 & n16452 ) | ( n13036 & n16452 ) ;
  assign n26818 = ( n12419 & ~n15442 ) | ( n12419 & n26817 ) | ( ~n15442 & n26817 ) ;
  assign n26819 = ( n6027 & ~n15334 ) | ( n6027 & n17268 ) | ( ~n15334 & n17268 ) ;
  assign n26820 = n11868 ^ n11391 ^ n7229 ;
  assign n26821 = n25855 ^ n14357 ^ n3536 ;
  assign n26822 = ( n11531 & n16340 ) | ( n11531 & n26821 ) | ( n16340 & n26821 ) ;
  assign n26823 = ( ~n4838 & n17755 ) | ( ~n4838 & n26822 ) | ( n17755 & n26822 ) ;
  assign n26824 = ( ~n9183 & n26820 ) | ( ~n9183 & n26823 ) | ( n26820 & n26823 ) ;
  assign n26825 = n26824 ^ n17655 ^ n15896 ;
  assign n26826 = n6862 ^ n4862 ^ n1739 ;
  assign n26827 = n26826 ^ n22813 ^ n17813 ;
  assign n26828 = n26827 ^ n14803 ^ n7572 ;
  assign n26829 = ( ~n3549 & n11965 ) | ( ~n3549 & n25716 ) | ( n11965 & n25716 ) ;
  assign n26830 = ( n3324 & ~n8050 ) | ( n3324 & n11139 ) | ( ~n8050 & n11139 ) ;
  assign n26831 = ( ~n15628 & n17188 ) | ( ~n15628 & n26830 ) | ( n17188 & n26830 ) ;
  assign n26832 = n18553 ^ n14326 ^ n5662 ;
  assign n26833 = ( n3851 & ~n5962 ) | ( n3851 & n12932 ) | ( ~n5962 & n12932 ) ;
  assign n26834 = ( ~n6318 & n26832 ) | ( ~n6318 & n26833 ) | ( n26832 & n26833 ) ;
  assign n26835 = ( n2580 & n19491 ) | ( n2580 & n21668 ) | ( n19491 & n21668 ) ;
  assign n26836 = n19119 ^ n12036 ^ n2478 ;
  assign n26838 = n4087 ^ n3570 ^ n2984 ;
  assign n26837 = n4174 & n18807 ;
  assign n26839 = n26838 ^ n26837 ^ 1'b0 ;
  assign n26840 = n7745 | n12108 ;
  assign n26841 = n26840 ^ n13597 ^ 1'b0 ;
  assign n26842 = ~n6605 & n26129 ;
  assign n26845 = ( n464 & n3025 ) | ( n464 & ~n7244 ) | ( n3025 & ~n7244 ) ;
  assign n26843 = n2372 | n5935 ;
  assign n26844 = n7669 & ~n26843 ;
  assign n26846 = n26845 ^ n26844 ^ n4282 ;
  assign n26847 = ( ~n1634 & n2222 ) | ( ~n1634 & n21727 ) | ( n2222 & n21727 ) ;
  assign n26848 = ( n8062 & ~n8465 ) | ( n8062 & n14334 ) | ( ~n8465 & n14334 ) ;
  assign n26849 = ( n24215 & n26847 ) | ( n24215 & ~n26848 ) | ( n26847 & ~n26848 ) ;
  assign n26850 = ( n326 & n12014 ) | ( n326 & ~n26849 ) | ( n12014 & ~n26849 ) ;
  assign n26851 = n26850 ^ n9829 ^ n1357 ;
  assign n26852 = ( ~n7370 & n18323 ) | ( ~n7370 & n26851 ) | ( n18323 & n26851 ) ;
  assign n26853 = n25959 ^ n9170 ^ n1318 ;
  assign n26854 = ( n1034 & n14278 ) | ( n1034 & ~n26853 ) | ( n14278 & ~n26853 ) ;
  assign n26855 = n23569 ^ n22265 ^ n2695 ;
  assign n26856 = ( n5078 & n9198 ) | ( n5078 & ~n16979 ) | ( n9198 & ~n16979 ) ;
  assign n26857 = n26856 ^ n14371 ^ n10068 ;
  assign n26858 = ( n20410 & n26855 ) | ( n20410 & ~n26857 ) | ( n26855 & ~n26857 ) ;
  assign n26859 = ( n5154 & ~n14973 ) | ( n5154 & n21951 ) | ( ~n14973 & n21951 ) ;
  assign n26860 = ( n3748 & n19986 ) | ( n3748 & n26859 ) | ( n19986 & n26859 ) ;
  assign n26861 = ~n4232 & n11678 ;
  assign n26862 = n26861 ^ n8033 ^ 1'b0 ;
  assign n26863 = n21568 & ~n26862 ;
  assign n26864 = n26863 ^ n17455 ^ 1'b0 ;
  assign n26865 = n2714 & n13077 ;
  assign n26866 = n26865 ^ n19851 ^ 1'b0 ;
  assign n26867 = n11193 ^ n1258 ^ 1'b0 ;
  assign n26868 = n17845 & n26867 ;
  assign n26869 = ( n18421 & ~n20782 ) | ( n18421 & n26868 ) | ( ~n20782 & n26868 ) ;
  assign n26870 = ( n14915 & n23697 ) | ( n14915 & n25292 ) | ( n23697 & n25292 ) ;
  assign n26871 = n12529 ^ n4758 ^ n1981 ;
  assign n26872 = n11913 & n26871 ;
  assign n26873 = ~n19071 & n26872 ;
  assign n26874 = ( ~n3709 & n8381 ) | ( ~n3709 & n26873 ) | ( n8381 & n26873 ) ;
  assign n26875 = n25223 ^ n8838 ^ n7731 ;
  assign n26876 = ( n1148 & ~n21224 ) | ( n1148 & n23458 ) | ( ~n21224 & n23458 ) ;
  assign n26877 = ( n13978 & ~n15454 ) | ( n13978 & n21361 ) | ( ~n15454 & n21361 ) ;
  assign n26878 = n26877 ^ n20844 ^ n3254 ;
  assign n26879 = n8516 ^ n8057 ^ 1'b0 ;
  assign n26880 = n7919 & ~n26879 ;
  assign n26881 = ( n2727 & ~n9193 ) | ( n2727 & n26880 ) | ( ~n9193 & n26880 ) ;
  assign n26882 = n16176 ^ n14539 ^ n13046 ;
  assign n26883 = ( n7792 & n11015 ) | ( n7792 & n26882 ) | ( n11015 & n26882 ) ;
  assign n26884 = ( n8455 & n24474 ) | ( n8455 & ~n26883 ) | ( n24474 & ~n26883 ) ;
  assign n26885 = n13277 ^ n9303 ^ n7799 ;
  assign n26886 = ( ~n3369 & n15975 ) | ( ~n3369 & n26885 ) | ( n15975 & n26885 ) ;
  assign n26887 = n6944 & ~n18717 ;
  assign n26888 = n22839 & n26887 ;
  assign n26889 = ( n602 & n4810 ) | ( n602 & ~n8396 ) | ( n4810 & ~n8396 ) ;
  assign n26890 = n13562 ^ n7617 ^ x1 ;
  assign n26891 = ( n12766 & n13546 ) | ( n12766 & ~n18315 ) | ( n13546 & ~n18315 ) ;
  assign n26892 = n26891 ^ n18737 ^ n14292 ;
  assign n26893 = n25124 ^ n10904 ^ n3263 ;
  assign n26894 = ( ~n2075 & n3124 ) | ( ~n2075 & n16139 ) | ( n3124 & n16139 ) ;
  assign n26895 = n25958 ^ n5113 ^ n1369 ;
  assign n26896 = n7660 ^ n4669 ^ n3161 ;
  assign n26897 = ~n3154 & n3827 ;
  assign n26898 = ~n13958 & n26897 ;
  assign n26899 = n8256 | n26898 ;
  assign n26900 = n10359 & ~n26899 ;
  assign n26901 = ( n1544 & n3357 ) | ( n1544 & n4140 ) | ( n3357 & n4140 ) ;
  assign n26902 = ( n26896 & n26900 ) | ( n26896 & n26901 ) | ( n26900 & n26901 ) ;
  assign n26903 = ( n12467 & n17408 ) | ( n12467 & n26406 ) | ( n17408 & n26406 ) ;
  assign n26904 = n3223 & ~n26903 ;
  assign n26905 = n3657 ^ n419 ^ 1'b0 ;
  assign n26906 = n21241 & n26905 ;
  assign n26907 = ~n2422 & n10416 ;
  assign n26908 = ~n26906 & n26907 ;
  assign n26909 = n24721 ^ n14435 ^ n5469 ;
  assign n26910 = ( n1707 & n6602 ) | ( n1707 & n26909 ) | ( n6602 & n26909 ) ;
  assign n26911 = ( n1784 & n4287 ) | ( n1784 & n4783 ) | ( n4287 & n4783 ) ;
  assign n26912 = ( n6432 & n15265 ) | ( n6432 & n19929 ) | ( n15265 & n19929 ) ;
  assign n26913 = n26912 ^ n15221 ^ n9265 ;
  assign n26914 = ( n475 & n1926 ) | ( n475 & n11077 ) | ( n1926 & n11077 ) ;
  assign n26915 = n26914 ^ n25744 ^ 1'b0 ;
  assign n26916 = ( ~n5487 & n25683 ) | ( ~n5487 & n25686 ) | ( n25683 & n25686 ) ;
  assign n26917 = n26916 ^ n24789 ^ n12909 ;
  assign n26918 = n19013 ^ n8595 ^ n5391 ;
  assign n26919 = ( ~n9482 & n9737 ) | ( ~n9482 & n26918 ) | ( n9737 & n26918 ) ;
  assign n26920 = n3877 | n11916 ;
  assign n26921 = n4887 & n8280 ;
  assign n26922 = n26921 ^ n12995 ^ 1'b0 ;
  assign n26923 = n26922 ^ n24770 ^ n18161 ;
  assign n26924 = n26923 ^ n1027 ^ 1'b0 ;
  assign n26925 = ( n868 & n12617 ) | ( n868 & ~n13420 ) | ( n12617 & ~n13420 ) ;
  assign n26926 = n26925 ^ n8462 ^ n801 ;
  assign n26927 = n1637 | n9323 ;
  assign n26929 = ( n3300 & n8663 ) | ( n3300 & n10643 ) | ( n8663 & n10643 ) ;
  assign n26928 = n13794 & ~n18455 ;
  assign n26930 = n26929 ^ n26928 ^ n13160 ;
  assign n26931 = n22297 ^ n1926 ^ x97 ;
  assign n26932 = n9431 & ~n20957 ;
  assign n26933 = ( n20770 & ~n26931 ) | ( n20770 & n26932 ) | ( ~n26931 & n26932 ) ;
  assign n26934 = n20514 ^ n1157 ^ n809 ;
  assign n26935 = ( n14564 & n15394 ) | ( n14564 & n21199 ) | ( n15394 & n21199 ) ;
  assign n26936 = ( ~n1475 & n3018 ) | ( ~n1475 & n13261 ) | ( n3018 & n13261 ) ;
  assign n26937 = ~n4600 & n13667 ;
  assign n26938 = n11850 & n26937 ;
  assign n26939 = ( n3199 & n7629 ) | ( n3199 & ~n26938 ) | ( n7629 & ~n26938 ) ;
  assign n26940 = n757 & n10787 ;
  assign n26941 = n26940 ^ n1626 ^ 1'b0 ;
  assign n26942 = n1670 & ~n26941 ;
  assign n26943 = ( ~n14719 & n15845 ) | ( ~n14719 & n26942 ) | ( n15845 & n26942 ) ;
  assign n26944 = n194 & ~n21201 ;
  assign n26945 = n26943 & n26944 ;
  assign n26946 = ( n14830 & ~n21810 ) | ( n14830 & n26945 ) | ( ~n21810 & n26945 ) ;
  assign n26947 = n26946 ^ n19585 ^ n6343 ;
  assign n26948 = ( ~n3411 & n3752 ) | ( ~n3411 & n11617 ) | ( n3752 & n11617 ) ;
  assign n26949 = n11213 ^ n7358 ^ n1715 ;
  assign n26950 = ~n13750 & n26949 ;
  assign n26951 = n26950 ^ n23654 ^ 1'b0 ;
  assign n26952 = ( n19364 & n26948 ) | ( n19364 & n26951 ) | ( n26948 & n26951 ) ;
  assign n26953 = ~n322 & n5136 ;
  assign n26954 = n417 & n26953 ;
  assign n26956 = ( n1840 & n5416 ) | ( n1840 & n6926 ) | ( n5416 & n6926 ) ;
  assign n26955 = n18051 & ~n21207 ;
  assign n26957 = n26956 ^ n26955 ^ 1'b0 ;
  assign n26958 = n6149 ^ n3993 ^ n894 ;
  assign n26959 = ( ~n11771 & n14648 ) | ( ~n11771 & n26958 ) | ( n14648 & n26958 ) ;
  assign n26960 = ( ~n15919 & n21442 ) | ( ~n15919 & n26959 ) | ( n21442 & n26959 ) ;
  assign n26961 = ( ~n3126 & n12751 ) | ( ~n3126 & n20804 ) | ( n12751 & n20804 ) ;
  assign n26962 = ( n11491 & n26439 ) | ( n11491 & n26961 ) | ( n26439 & n26961 ) ;
  assign n26963 = ( ~n555 & n2947 ) | ( ~n555 & n19843 ) | ( n2947 & n19843 ) ;
  assign n26964 = n26963 ^ n21653 ^ n15396 ;
  assign n26965 = ( n6947 & ~n7450 ) | ( n6947 & n8373 ) | ( ~n7450 & n8373 ) ;
  assign n26966 = n8250 ^ n7190 ^ 1'b0 ;
  assign n26967 = ~n26965 & n26966 ;
  assign n26968 = ( n15856 & n23573 ) | ( n15856 & ~n26967 ) | ( n23573 & ~n26967 ) ;
  assign n26969 = ( n1782 & n1918 ) | ( n1782 & ~n15375 ) | ( n1918 & ~n15375 ) ;
  assign n26970 = n26969 ^ n3601 ^ 1'b0 ;
  assign n26972 = ~n4654 & n8233 ;
  assign n26973 = n26972 ^ n2250 ^ 1'b0 ;
  assign n26974 = ( n2556 & n8378 ) | ( n2556 & ~n26973 ) | ( n8378 & ~n26973 ) ;
  assign n26971 = n26088 ^ n9577 ^ n3779 ;
  assign n26975 = n26974 ^ n26971 ^ n7508 ;
  assign n26976 = n11804 ^ n2309 ^ n775 ;
  assign n26977 = n26976 ^ n3280 ^ 1'b0 ;
  assign n26978 = ( n11868 & n18119 ) | ( n11868 & ~n20275 ) | ( n18119 & ~n20275 ) ;
  assign n26979 = n22962 ^ n6491 ^ 1'b0 ;
  assign n26980 = n6307 | n26979 ;
  assign n26981 = ( ~n26977 & n26978 ) | ( ~n26977 & n26980 ) | ( n26978 & n26980 ) ;
  assign n26982 = n17266 ^ n13239 ^ n6458 ;
  assign n26983 = ( ~n10029 & n12387 ) | ( ~n10029 & n26982 ) | ( n12387 & n26982 ) ;
  assign n26984 = ( n4673 & n7858 ) | ( n4673 & n26983 ) | ( n7858 & n26983 ) ;
  assign n26985 = n18364 ^ n17837 ^ 1'b0 ;
  assign n26986 = ~n24144 & n26985 ;
  assign n26987 = ( ~n4980 & n5793 ) | ( ~n4980 & n12353 ) | ( n5793 & n12353 ) ;
  assign n26988 = n4791 | n10174 ;
  assign n26989 = n26987 | n26988 ;
  assign n26991 = n14990 ^ n13056 ^ n189 ;
  assign n26990 = n3043 | n3552 ;
  assign n26992 = n26991 ^ n26990 ^ 1'b0 ;
  assign n26993 = n26992 ^ n25027 ^ n2940 ;
  assign n26994 = n7313 | n11019 ;
  assign n26995 = n26994 ^ n19336 ^ 1'b0 ;
  assign n26996 = n10216 ^ n7614 ^ n2026 ;
  assign n26997 = n11703 | n26996 ;
  assign n26998 = n3612 & ~n26997 ;
  assign n26999 = n26998 ^ n20207 ^ 1'b0 ;
  assign n27000 = ( n23373 & n26995 ) | ( n23373 & n26999 ) | ( n26995 & n26999 ) ;
  assign n27001 = ( n617 & ~n10218 ) | ( n617 & n11258 ) | ( ~n10218 & n11258 ) ;
  assign n27002 = n27001 ^ n4394 ^ n497 ;
  assign n27003 = n27002 ^ n18540 ^ n9315 ;
  assign n27004 = n27003 ^ n6823 ^ n1475 ;
  assign n27005 = ( n2081 & ~n5257 ) | ( n2081 & n7041 ) | ( ~n5257 & n7041 ) ;
  assign n27006 = n5830 & n8252 ;
  assign n27007 = ~n27005 & n27006 ;
  assign n27008 = n27007 ^ n26641 ^ n4809 ;
  assign n27010 = n5446 & ~n7079 ;
  assign n27011 = ~n9870 & n27010 ;
  assign n27009 = ( n3558 & n10650 ) | ( n3558 & n20640 ) | ( n10650 & n20640 ) ;
  assign n27012 = n27011 ^ n27009 ^ n15277 ;
  assign n27013 = n19814 ^ n6024 ^ n4801 ;
  assign n27014 = n27013 ^ n8954 ^ n1112 ;
  assign n27015 = n2553 & n20552 ;
  assign n27016 = ~n1516 & n27015 ;
  assign n27017 = ( n444 & ~n13925 ) | ( n444 & n27016 ) | ( ~n13925 & n27016 ) ;
  assign n27018 = ( n14534 & n18605 ) | ( n14534 & n27017 ) | ( n18605 & n27017 ) ;
  assign n27020 = ~n6062 & n20045 ;
  assign n27021 = n27020 ^ n3369 ^ 1'b0 ;
  assign n27019 = n1286 & ~n4091 ;
  assign n27022 = n27021 ^ n27019 ^ 1'b0 ;
  assign n27023 = ( n4960 & n9091 ) | ( n4960 & ~n15669 ) | ( n9091 & ~n15669 ) ;
  assign n27024 = n27023 ^ n25511 ^ n9529 ;
  assign n27027 = ( ~n195 & n1277 ) | ( ~n195 & n7260 ) | ( n1277 & n7260 ) ;
  assign n27028 = n27027 ^ n12241 ^ 1'b0 ;
  assign n27025 = n12506 ^ n9997 ^ n499 ;
  assign n27026 = n13538 & n27025 ;
  assign n27029 = n27028 ^ n27026 ^ n2246 ;
  assign n27030 = ( x114 & ~n14903 ) | ( x114 & n22010 ) | ( ~n14903 & n22010 ) ;
  assign n27031 = ( n1755 & ~n20924 ) | ( n1755 & n27030 ) | ( ~n20924 & n27030 ) ;
  assign n27032 = n732 & ~n7629 ;
  assign n27033 = ~n19299 & n27032 ;
  assign n27034 = ( ~n11300 & n18418 ) | ( ~n11300 & n27033 ) | ( n18418 & n27033 ) ;
  assign n27035 = n8092 & ~n22053 ;
  assign n27036 = ( n10216 & n13581 ) | ( n10216 & ~n16823 ) | ( n13581 & ~n16823 ) ;
  assign n27037 = n27036 ^ n26740 ^ n22981 ;
  assign n27038 = n4663 & n9042 ;
  assign n27039 = n7322 ^ n611 ^ 1'b0 ;
  assign n27040 = n27039 ^ n7660 ^ 1'b0 ;
  assign n27041 = n4494 & ~n18349 ;
  assign n27042 = n27041 ^ n21611 ^ n8917 ;
  assign n27043 = ( n21198 & ~n27040 ) | ( n21198 & n27042 ) | ( ~n27040 & n27042 ) ;
  assign n27044 = n20688 | n27043 ;
  assign n27045 = n27044 ^ n13089 ^ 1'b0 ;
  assign n27046 = n4570 & ~n27045 ;
  assign n27047 = n15029 ^ n4165 ^ 1'b0 ;
  assign n27048 = n6489 & ~n27047 ;
  assign n27049 = ( n9175 & n9517 ) | ( n9175 & ~n17848 ) | ( n9517 & ~n17848 ) ;
  assign n27050 = ~n639 & n6374 ;
  assign n27051 = ( n5456 & n11610 ) | ( n5456 & ~n27050 ) | ( n11610 & ~n27050 ) ;
  assign n27056 = n20095 ^ n16124 ^ n11925 ;
  assign n27057 = n12273 & ~n27056 ;
  assign n27058 = ~n9259 & n27057 ;
  assign n27055 = ( n2645 & n8788 ) | ( n2645 & n11910 ) | ( n8788 & n11910 ) ;
  assign n27052 = n21316 & ~n22040 ;
  assign n27053 = ( n477 & ~n7419 ) | ( n477 & n27052 ) | ( ~n7419 & n27052 ) ;
  assign n27054 = n27053 ^ n22280 ^ 1'b0 ;
  assign n27059 = n27058 ^ n27055 ^ n27054 ;
  assign n27060 = ( ~n8935 & n14001 ) | ( ~n8935 & n14898 ) | ( n14001 & n14898 ) ;
  assign n27061 = n16734 & ~n20082 ;
  assign n27062 = ( ~n709 & n903 ) | ( ~n709 & n7918 ) | ( n903 & n7918 ) ;
  assign n27063 = ( ~n7863 & n25139 ) | ( ~n7863 & n27062 ) | ( n25139 & n27062 ) ;
  assign n27064 = n6163 | n9306 ;
  assign n27065 = n17574 ^ n17139 ^ 1'b0 ;
  assign n27066 = n2607 & ~n27065 ;
  assign n27067 = n15210 ^ n11919 ^ n3625 ;
  assign n27068 = n23114 ^ n18205 ^ n7266 ;
  assign n27069 = ( n2069 & n27067 ) | ( n2069 & ~n27068 ) | ( n27067 & ~n27068 ) ;
  assign n27070 = n25630 ^ n18297 ^ n10359 ;
  assign n27071 = n7529 ^ n3352 ^ n2030 ;
  assign n27072 = ( n1052 & n11681 ) | ( n1052 & ~n27071 ) | ( n11681 & ~n27071 ) ;
  assign n27073 = n27072 ^ n25805 ^ n2293 ;
  assign n27074 = ( n4559 & n16927 ) | ( n4559 & n19519 ) | ( n16927 & n19519 ) ;
  assign n27075 = ( ~n5508 & n7642 ) | ( ~n5508 & n15902 ) | ( n7642 & n15902 ) ;
  assign n27076 = ( n9343 & ~n14432 ) | ( n9343 & n16587 ) | ( ~n14432 & n16587 ) ;
  assign n27077 = n27076 ^ n8557 ^ n4206 ;
  assign n27078 = ( ~n12517 & n27075 ) | ( ~n12517 & n27077 ) | ( n27075 & n27077 ) ;
  assign n27079 = ( n13737 & ~n16070 ) | ( n13737 & n19089 ) | ( ~n16070 & n19089 ) ;
  assign n27080 = ( n15967 & n20250 ) | ( n15967 & ~n23747 ) | ( n20250 & ~n23747 ) ;
  assign n27081 = n16196 | n27080 ;
  assign n27082 = ( n6256 & n10583 ) | ( n6256 & ~n22283 ) | ( n10583 & ~n22283 ) ;
  assign n27083 = n24654 ^ n22782 ^ n6765 ;
  assign n27084 = n27083 ^ n4376 ^ 1'b0 ;
  assign n27086 = ( x103 & ~n9257 ) | ( x103 & n11252 ) | ( ~n9257 & n11252 ) ;
  assign n27087 = ( n11891 & ~n19241 ) | ( n11891 & n27086 ) | ( ~n19241 & n27086 ) ;
  assign n27085 = n16845 ^ n12507 ^ n8765 ;
  assign n27088 = n27087 ^ n27085 ^ n1126 ;
  assign n27089 = n26898 ^ n5745 ^ n671 ;
  assign n27090 = ( ~n7885 & n16078 ) | ( ~n7885 & n27089 ) | ( n16078 & n27089 ) ;
  assign n27091 = n25491 ^ n22550 ^ n3876 ;
  assign n27092 = ( n3424 & n19923 ) | ( n3424 & n23214 ) | ( n19923 & n23214 ) ;
  assign n27093 = n17744 ^ n17504 ^ n11857 ;
  assign n27094 = n27093 ^ n2116 ^ 1'b0 ;
  assign n27095 = n25628 ^ n12523 ^ n285 ;
  assign n27096 = n27095 ^ n7693 ^ n4739 ;
  assign n27097 = n12052 & ~n20456 ;
  assign n27098 = ( n3449 & ~n6183 ) | ( n3449 & n18478 ) | ( ~n6183 & n18478 ) ;
  assign n27099 = n27098 ^ n13599 ^ 1'b0 ;
  assign n27100 = n4396 & n27099 ;
  assign n27101 = ( n7356 & n12032 ) | ( n7356 & n17604 ) | ( n12032 & n17604 ) ;
  assign n27102 = n27101 ^ n26353 ^ n20743 ;
  assign n27103 = n18002 & ~n25631 ;
  assign n27104 = ~n27102 & n27103 ;
  assign n27105 = n3424 & n13106 ;
  assign n27106 = ( x92 & n426 ) | ( x92 & n554 ) | ( n426 & n554 ) ;
  assign n27107 = n27106 ^ n19204 ^ n12926 ;
  assign n27108 = n20190 ^ n13925 ^ 1'b0 ;
  assign n27109 = n17382 ^ n13177 ^ n2099 ;
  assign n27110 = n16035 ^ n14976 ^ n1322 ;
  assign n27111 = ( n1582 & n2756 ) | ( n1582 & ~n17020 ) | ( n2756 & ~n17020 ) ;
  assign n27112 = n11259 ^ n8556 ^ n3387 ;
  assign n27113 = ( n9766 & n10908 ) | ( n9766 & n27112 ) | ( n10908 & n27112 ) ;
  assign n27114 = n27113 ^ n19269 ^ n3314 ;
  assign n27115 = n3767 ^ n2062 ^ 1'b0 ;
  assign n27116 = n17316 & n27115 ;
  assign n27117 = n17125 ^ n4192 ^ 1'b0 ;
  assign n27118 = n22053 & n27117 ;
  assign n27119 = n23290 ^ n23064 ^ n8376 ;
  assign n27120 = ~n21437 & n26293 ;
  assign n27121 = ~n1426 & n14111 ;
  assign n27122 = n27121 ^ n7079 ^ 1'b0 ;
  assign n27123 = ( ~n5768 & n25538 ) | ( ~n5768 & n27122 ) | ( n25538 & n27122 ) ;
  assign n27124 = n10989 ^ n7224 ^ n3251 ;
  assign n27125 = n27124 ^ n4983 ^ 1'b0 ;
  assign n27126 = n22345 ^ n16028 ^ n1765 ;
  assign n27127 = n27126 ^ n17028 ^ n2219 ;
  assign n27130 = n13004 ^ n3134 ^ n2124 ;
  assign n27128 = ( n3749 & n19925 ) | ( n3749 & n23557 ) | ( n19925 & n23557 ) ;
  assign n27129 = ( n2154 & n25875 ) | ( n2154 & n27128 ) | ( n25875 & n27128 ) ;
  assign n27131 = n27130 ^ n27129 ^ n3677 ;
  assign n27132 = ( n1731 & n4767 ) | ( n1731 & ~n27131 ) | ( n4767 & ~n27131 ) ;
  assign n27133 = n22735 ^ n20238 ^ n15795 ;
  assign n27134 = n12232 ^ n1195 ^ n1059 ;
  assign n27135 = n13538 | n21127 ;
  assign n27136 = n27134 | n27135 ;
  assign n27137 = n11884 ^ n368 ^ 1'b0 ;
  assign n27138 = n17252 ^ n10672 ^ n7349 ;
  assign n27139 = n9269 & ~n12442 ;
  assign n27140 = ( n7201 & n11204 ) | ( n7201 & n27139 ) | ( n11204 & n27139 ) ;
  assign n27141 = n24088 ^ n23185 ^ n14535 ;
  assign n27142 = n21085 ^ n20209 ^ n4850 ;
  assign n27143 = ( ~n7731 & n7769 ) | ( ~n7731 & n11620 ) | ( n7769 & n11620 ) ;
  assign n27150 = n23973 ^ n13953 ^ n13411 ;
  assign n27148 = n12696 ^ n10425 ^ n5490 ;
  assign n27149 = n27148 ^ n25777 ^ n12992 ;
  assign n27146 = x62 & n612 ;
  assign n27144 = n1298 & ~n10655 ;
  assign n27145 = n27144 ^ n15175 ^ 1'b0 ;
  assign n27147 = n27146 ^ n27145 ^ n16933 ;
  assign n27151 = n27150 ^ n27149 ^ n27147 ;
  assign n27154 = ( n9548 & n9685 ) | ( n9548 & ~n10078 ) | ( n9685 & ~n10078 ) ;
  assign n27152 = n12396 ^ n7737 ^ 1'b0 ;
  assign n27153 = ( n3247 & n5896 ) | ( n3247 & ~n27152 ) | ( n5896 & ~n27152 ) ;
  assign n27155 = n27154 ^ n27153 ^ n9789 ;
  assign n27156 = ( n578 & ~n3642 ) | ( n578 & n26524 ) | ( ~n3642 & n26524 ) ;
  assign n27157 = ( ~n14654 & n15229 ) | ( ~n14654 & n27156 ) | ( n15229 & n27156 ) ;
  assign n27158 = n13985 ^ n12423 ^ n6813 ;
  assign n27159 = n10480 ^ n6420 ^ n5007 ;
  assign n27160 = ( n14793 & ~n27158 ) | ( n14793 & n27159 ) | ( ~n27158 & n27159 ) ;
  assign n27161 = n10998 | n18396 ;
  assign n27162 = n27161 ^ n6119 ^ 1'b0 ;
  assign n27163 = n26474 ^ n3944 ^ n2607 ;
  assign n27164 = n27163 ^ n2222 ^ 1'b0 ;
  assign n27165 = n26583 | n27164 ;
  assign n27166 = ( n9471 & ~n20697 ) | ( n9471 & n23108 ) | ( ~n20697 & n23108 ) ;
  assign n27167 = n22766 ^ n8759 ^ 1'b0 ;
  assign n27168 = ~n17885 & n27167 ;
  assign n27169 = n27168 ^ n18282 ^ 1'b0 ;
  assign n27170 = ( n18130 & ~n27166 ) | ( n18130 & n27169 ) | ( ~n27166 & n27169 ) ;
  assign n27171 = n15192 ^ n1492 ^ 1'b0 ;
  assign n27174 = n15484 ^ n5177 ^ n535 ;
  assign n27172 = ~n5865 & n8559 ;
  assign n27173 = ( ~n3735 & n22067 ) | ( ~n3735 & n27172 ) | ( n22067 & n27172 ) ;
  assign n27175 = n27174 ^ n27173 ^ 1'b0 ;
  assign n27176 = ( n12487 & n27171 ) | ( n12487 & n27175 ) | ( n27171 & n27175 ) ;
  assign n27177 = n27176 ^ n12580 ^ n8293 ;
  assign n27178 = ( n8962 & ~n10567 ) | ( n8962 & n20699 ) | ( ~n10567 & n20699 ) ;
  assign n27181 = n9333 ^ n5932 ^ n3257 ;
  assign n27179 = ~n23656 & n24831 ;
  assign n27180 = n7587 & n27179 ;
  assign n27182 = n27181 ^ n27180 ^ 1'b0 ;
  assign n27183 = n19164 ^ n12899 ^ n2806 ;
  assign n27184 = ( n2098 & n9962 ) | ( n2098 & ~n27183 ) | ( n9962 & ~n27183 ) ;
  assign n27185 = n1787 | n27184 ;
  assign n27186 = n25410 ^ n17663 ^ n5747 ;
  assign n27187 = n11773 ^ n5233 ^ n4768 ;
  assign n27188 = ( n7059 & ~n8750 ) | ( n7059 & n27187 ) | ( ~n8750 & n27187 ) ;
  assign n27189 = n27188 ^ n27145 ^ n17255 ;
  assign n27190 = n12512 | n21961 ;
  assign n27191 = n8932 ^ n6482 ^ n5070 ;
  assign n27192 = n20887 ^ n16357 ^ n12075 ;
  assign n27193 = n26441 ^ n8548 ^ n5659 ;
  assign n27194 = ( n3144 & ~n10115 ) | ( n3144 & n12702 ) | ( ~n10115 & n12702 ) ;
  assign n27195 = n27194 ^ n16999 ^ n15881 ;
  assign n27196 = n26555 ^ n10775 ^ n6269 ;
  assign n27197 = ( n1725 & n5885 ) | ( n1725 & n8496 ) | ( n5885 & n8496 ) ;
  assign n27198 = ( ~n5902 & n25319 ) | ( ~n5902 & n27197 ) | ( n25319 & n27197 ) ;
  assign n27199 = n12097 & ~n14541 ;
  assign n27200 = n12889 & n27199 ;
  assign n27201 = n14553 ^ n13307 ^ n5822 ;
  assign n27202 = n27201 ^ n6001 ^ 1'b0 ;
  assign n27203 = n17132 ^ n16902 ^ n480 ;
  assign n27204 = n15880 ^ n2361 ^ n656 ;
  assign n27205 = ( ~n8425 & n27203 ) | ( ~n8425 & n27204 ) | ( n27203 & n27204 ) ;
  assign n27206 = ( n15396 & n23769 ) | ( n15396 & n27205 ) | ( n23769 & n27205 ) ;
  assign n27207 = ( n1848 & n4289 ) | ( n1848 & n16135 ) | ( n4289 & n16135 ) ;
  assign n27208 = n7827 ^ n5114 ^ n1204 ;
  assign n27209 = n10416 ^ n9202 ^ n1625 ;
  assign n27210 = ( n826 & n7152 ) | ( n826 & ~n18871 ) | ( n7152 & ~n18871 ) ;
  assign n27211 = ( n10264 & n11123 ) | ( n10264 & n13834 ) | ( n11123 & n13834 ) ;
  assign n27212 = n27211 ^ n15575 ^ n373 ;
  assign n27215 = ( ~n10047 & n12676 ) | ( ~n10047 & n25513 ) | ( n12676 & n25513 ) ;
  assign n27213 = ( n1430 & n12092 ) | ( n1430 & n23597 ) | ( n12092 & n23597 ) ;
  assign n27214 = ( ~n3468 & n7065 ) | ( ~n3468 & n27213 ) | ( n7065 & n27213 ) ;
  assign n27216 = n27215 ^ n27214 ^ n3113 ;
  assign n27217 = ( n16758 & ~n19275 ) | ( n16758 & n21188 ) | ( ~n19275 & n21188 ) ;
  assign n27218 = n7598 & n27217 ;
  assign n27219 = n27218 ^ n3107 ^ 1'b0 ;
  assign n27220 = n7714 & n22590 ;
  assign n27221 = n27220 ^ n14258 ^ 1'b0 ;
  assign n27222 = ( n8096 & ~n10558 ) | ( n8096 & n25141 ) | ( ~n10558 & n25141 ) ;
  assign n27223 = ( n9020 & ~n10894 ) | ( n9020 & n15518 ) | ( ~n10894 & n15518 ) ;
  assign n27224 = n24726 ^ n12994 ^ 1'b0 ;
  assign n27225 = ( n2055 & n8612 ) | ( n2055 & ~n27224 ) | ( n8612 & ~n27224 ) ;
  assign n27226 = n8503 ^ n1712 ^ 1'b0 ;
  assign n27227 = n1158 & n25018 ;
  assign n27228 = n7003 & n27227 ;
  assign n27229 = ( ~n9967 & n27039 ) | ( ~n9967 & n27228 ) | ( n27039 & n27228 ) ;
  assign n27230 = ( n3207 & n18580 ) | ( n3207 & ~n21739 ) | ( n18580 & ~n21739 ) ;
  assign n27231 = ( n21828 & n21955 ) | ( n21828 & n27230 ) | ( n21955 & n27230 ) ;
  assign n27232 = ( n2304 & n11337 ) | ( n2304 & ~n27231 ) | ( n11337 & ~n27231 ) ;
  assign n27233 = n9892 ^ n9837 ^ 1'b0 ;
  assign n27234 = n27233 ^ n17189 ^ n13653 ;
  assign n27235 = n12533 ^ n7333 ^ n3351 ;
  assign n27236 = ( ~n13279 & n15251 ) | ( ~n13279 & n27235 ) | ( n15251 & n27235 ) ;
  assign n27237 = ~n1270 & n2091 ;
  assign n27238 = ~n13667 & n27237 ;
  assign n27239 = n5559 ^ n4712 ^ n394 ;
  assign n27240 = n27239 ^ n1760 ^ n1440 ;
  assign n27241 = n15142 ^ n9212 ^ n3892 ;
  assign n27246 = n3652 & n16222 ;
  assign n27247 = ~n6891 & n27246 ;
  assign n27248 = ( ~n2941 & n11494 ) | ( ~n2941 & n27247 ) | ( n11494 & n27247 ) ;
  assign n27245 = n22427 ^ n16893 ^ n3364 ;
  assign n27242 = ~n216 & n13377 ;
  assign n27243 = ~n4693 & n27242 ;
  assign n27244 = n27243 ^ n22968 ^ n19289 ;
  assign n27249 = n27248 ^ n27245 ^ n27244 ;
  assign n27250 = n4907 & ~n15400 ;
  assign n27251 = n27250 ^ n9570 ^ n3716 ;
  assign n27252 = n25855 ^ n9529 ^ n5087 ;
  assign n27253 = ( ~n8609 & n17052 ) | ( ~n8609 & n24474 ) | ( n17052 & n24474 ) ;
  assign n27254 = n16134 ^ n2381 ^ n542 ;
  assign n27255 = n27254 ^ n12915 ^ n7638 ;
  assign n27256 = n26882 ^ n5550 ^ x25 ;
  assign n27257 = ( n2717 & n4134 ) | ( n2717 & n4990 ) | ( n4134 & n4990 ) ;
  assign n27258 = n9864 | n13925 ;
  assign n27259 = n7088 & n7865 ;
  assign n27260 = ( n4856 & n4998 ) | ( n4856 & n27259 ) | ( n4998 & n27259 ) ;
  assign n27261 = n15962 ^ n9752 ^ 1'b0 ;
  assign n27262 = ( n2019 & n7056 ) | ( n2019 & n16717 ) | ( n7056 & n16717 ) ;
  assign n27263 = ( n24154 & n26171 ) | ( n24154 & ~n27262 ) | ( n26171 & ~n27262 ) ;
  assign n27264 = n20614 ^ n4755 ^ n3375 ;
  assign n27265 = ( n19750 & ~n26008 ) | ( n19750 & n27264 ) | ( ~n26008 & n27264 ) ;
  assign n27266 = n6180 & ~n16911 ;
  assign n27267 = n27266 ^ n2348 ^ 1'b0 ;
  assign n27268 = n22996 ^ n21081 ^ n13170 ;
  assign n27269 = ( n5378 & ~n8509 ) | ( n5378 & n10382 ) | ( ~n8509 & n10382 ) ;
  assign n27270 = ( n2131 & n26353 ) | ( n2131 & ~n27269 ) | ( n26353 & ~n27269 ) ;
  assign n27271 = ( n527 & n19815 ) | ( n527 & n27270 ) | ( n19815 & n27270 ) ;
  assign n27272 = ( ~n4762 & n27268 ) | ( ~n4762 & n27271 ) | ( n27268 & n27271 ) ;
  assign n27273 = ( n10689 & ~n27267 ) | ( n10689 & n27272 ) | ( ~n27267 & n27272 ) ;
  assign n27274 = n21227 ^ n14799 ^ n6157 ;
  assign n27275 = ( n268 & n2059 ) | ( n268 & n7409 ) | ( n2059 & n7409 ) ;
  assign n27276 = n9035 & ~n20209 ;
  assign n27277 = n27275 & n27276 ;
  assign n27282 = n8681 ^ n4408 ^ n573 ;
  assign n27280 = n18001 ^ n12066 ^ n11715 ;
  assign n27281 = n27280 ^ n5568 ^ n2179 ;
  assign n27278 = n12789 ^ n10534 ^ n5079 ;
  assign n27279 = ( n2877 & ~n15474 ) | ( n2877 & n27278 ) | ( ~n15474 & n27278 ) ;
  assign n27283 = n27282 ^ n27281 ^ n27279 ;
  assign n27284 = ( n1339 & n8375 ) | ( n1339 & ~n12342 ) | ( n8375 & ~n12342 ) ;
  assign n27285 = n3251 | n27284 ;
  assign n27286 = ( n2410 & n16968 ) | ( n2410 & ~n27285 ) | ( n16968 & ~n27285 ) ;
  assign n27287 = ( n3637 & ~n9603 ) | ( n3637 & n16244 ) | ( ~n9603 & n16244 ) ;
  assign n27288 = n26059 ^ n24910 ^ n17966 ;
  assign n27289 = n20196 ^ n4956 ^ n3770 ;
  assign n27291 = ( n1556 & ~n4676 ) | ( n1556 & n5828 ) | ( ~n4676 & n5828 ) ;
  assign n27292 = n27291 ^ n8487 ^ n7748 ;
  assign n27290 = ( n9407 & n10685 ) | ( n9407 & ~n12610 ) | ( n10685 & ~n12610 ) ;
  assign n27293 = n27292 ^ n27290 ^ n16404 ;
  assign n27294 = ( n3158 & n3474 ) | ( n3158 & n3839 ) | ( n3474 & n3839 ) ;
  assign n27295 = ~n1696 & n11720 ;
  assign n27296 = ~n20520 & n27295 ;
  assign n27297 = ( ~n14129 & n18443 ) | ( ~n14129 & n27296 ) | ( n18443 & n27296 ) ;
  assign n27298 = ( n17847 & n27294 ) | ( n17847 & n27297 ) | ( n27294 & n27297 ) ;
  assign n27299 = ( n545 & ~n13748 ) | ( n545 & n27298 ) | ( ~n13748 & n27298 ) ;
  assign n27300 = n5931 ^ n4758 ^ 1'b0 ;
  assign n27301 = n12920 & ~n27300 ;
  assign n27302 = n27083 ^ n22270 ^ n6521 ;
  assign n27303 = n8252 ^ n4167 ^ n914 ;
  assign n27304 = n13307 ^ n5922 ^ n5655 ;
  assign n27305 = ( n16082 & ~n17096 ) | ( n16082 & n22217 ) | ( ~n17096 & n22217 ) ;
  assign n27306 = ( n27303 & n27304 ) | ( n27303 & ~n27305 ) | ( n27304 & ~n27305 ) ;
  assign n27307 = x100 & n9754 ;
  assign n27308 = n12240 & n27307 ;
  assign n27309 = n27308 ^ n16190 ^ n13902 ;
  assign n27310 = n2840 & n9499 ;
  assign n27311 = n27310 ^ n20604 ^ n8844 ;
  assign n27312 = n15080 ^ n9143 ^ n326 ;
  assign n27313 = n27312 ^ n26070 ^ n14707 ;
  assign n27314 = n7256 ^ n6704 ^ 1'b0 ;
  assign n27315 = ~n19915 & n27314 ;
  assign n27316 = ( n1451 & ~n25586 ) | ( n1451 & n27315 ) | ( ~n25586 & n27315 ) ;
  assign n27317 = n19007 ^ n5290 ^ n4836 ;
  assign n27318 = n12928 & ~n27317 ;
  assign n27319 = ~n9673 & n15468 ;
  assign n27320 = n27319 ^ n22833 ^ n5947 ;
  assign n27321 = n27320 ^ n23119 ^ n21157 ;
  assign n27322 = n27321 ^ n788 ^ 1'b0 ;
  assign n27323 = n21085 | n27322 ;
  assign n27324 = n21442 ^ n15473 ^ n4313 ;
  assign n27325 = n27324 ^ n22752 ^ n22504 ;
  assign n27326 = n25290 ^ n7311 ^ n4048 ;
  assign n27327 = n19266 ^ n9591 ^ 1'b0 ;
  assign n27328 = ( n2697 & n11130 ) | ( n2697 & ~n27327 ) | ( n11130 & ~n27327 ) ;
  assign n27330 = n3056 & n25263 ;
  assign n27331 = n21677 & n27330 ;
  assign n27332 = ( ~n9477 & n12850 ) | ( ~n9477 & n27331 ) | ( n12850 & n27331 ) ;
  assign n27329 = ~n11556 & n19228 ;
  assign n27333 = n27332 ^ n27329 ^ 1'b0 ;
  assign n27334 = n16916 ^ n4032 ^ n1957 ;
  assign n27335 = n27334 ^ n25572 ^ n22869 ;
  assign n27336 = n5183 ^ n4830 ^ n1717 ;
  assign n27337 = ( n7860 & n26162 ) | ( n7860 & n27336 ) | ( n26162 & n27336 ) ;
  assign n27338 = n26791 ^ n10103 ^ 1'b0 ;
  assign n27339 = ( n1027 & ~n27337 ) | ( n1027 & n27338 ) | ( ~n27337 & n27338 ) ;
  assign n27340 = ( ~n1386 & n4468 ) | ( ~n1386 & n27339 ) | ( n4468 & n27339 ) ;
  assign n27341 = n8047 ^ n4870 ^ n4799 ;
  assign n27342 = n16655 & ~n27341 ;
  assign n27343 = n27342 ^ n11299 ^ n2953 ;
  assign n27344 = n20353 ^ n2207 ^ n915 ;
  assign n27345 = n19459 ^ n594 ^ 1'b0 ;
  assign n27346 = n24158 & ~n27345 ;
  assign n27347 = ( n10099 & n10199 ) | ( n10099 & ~n27346 ) | ( n10199 & ~n27346 ) ;
  assign n27348 = ( n20009 & ~n27344 ) | ( n20009 & n27347 ) | ( ~n27344 & n27347 ) ;
  assign n27349 = n2063 & n2253 ;
  assign n27350 = n27349 ^ n14121 ^ 1'b0 ;
  assign n27351 = ( n934 & ~n10334 ) | ( n934 & n22831 ) | ( ~n10334 & n22831 ) ;
  assign n27352 = n27351 ^ n16423 ^ 1'b0 ;
  assign n27353 = n13170 ^ n12633 ^ n6685 ;
  assign n27360 = n19063 ^ n18404 ^ n2572 ;
  assign n27361 = n27360 ^ n23922 ^ n18405 ;
  assign n27354 = ( n3860 & ~n8162 ) | ( n3860 & n23449 ) | ( ~n8162 & n23449 ) ;
  assign n27355 = n27354 ^ n11202 ^ n3282 ;
  assign n27356 = n21338 ^ n3407 ^ n1791 ;
  assign n27357 = n27356 ^ n16987 ^ n5409 ;
  assign n27358 = n27357 ^ n13026 ^ n3071 ;
  assign n27359 = ( n8982 & ~n27355 ) | ( n8982 & n27358 ) | ( ~n27355 & n27358 ) ;
  assign n27362 = n27361 ^ n27359 ^ n314 ;
  assign n27363 = ( n14089 & n18735 ) | ( n14089 & ~n20130 ) | ( n18735 & ~n20130 ) ;
  assign n27364 = n27363 ^ n19442 ^ n17726 ;
  assign n27365 = ( n9223 & n11546 ) | ( n9223 & ~n13327 ) | ( n11546 & ~n13327 ) ;
  assign n27366 = n15585 ^ n13607 ^ n7852 ;
  assign n27367 = n27366 ^ n24699 ^ n4727 ;
  assign n27368 = ( n4781 & n19825 ) | ( n4781 & ~n24745 ) | ( n19825 & ~n24745 ) ;
  assign n27369 = ( n2471 & n5318 ) | ( n2471 & n18320 ) | ( n5318 & n18320 ) ;
  assign n27370 = n27369 ^ n24273 ^ 1'b0 ;
  assign n27371 = ~n199 & n1459 ;
  assign n27372 = n1363 | n6959 ;
  assign n27373 = n27372 ^ n8943 ^ 1'b0 ;
  assign n27374 = n13400 ^ n8248 ^ 1'b0 ;
  assign n27375 = ( ~x72 & n4969 ) | ( ~x72 & n27374 ) | ( n4969 & n27374 ) ;
  assign n27376 = ( ~n12113 & n23091 ) | ( ~n12113 & n27375 ) | ( n23091 & n27375 ) ;
  assign n27377 = ( n2699 & n6366 ) | ( n2699 & n19806 ) | ( n6366 & n19806 ) ;
  assign n27378 = ( n7130 & n19645 ) | ( n7130 & ~n27377 ) | ( n19645 & ~n27377 ) ;
  assign n27379 = ( n2246 & n2976 ) | ( n2246 & ~n17920 ) | ( n2976 & ~n17920 ) ;
  assign n27380 = ( n6477 & n7328 ) | ( n6477 & n12466 ) | ( n7328 & n12466 ) ;
  assign n27381 = ( n9355 & ~n15799 ) | ( n9355 & n27380 ) | ( ~n15799 & n27380 ) ;
  assign n27382 = ( ~n15719 & n27379 ) | ( ~n15719 & n27381 ) | ( n27379 & n27381 ) ;
  assign n27383 = ~n7644 & n16028 ;
  assign n27384 = ~n2737 & n27383 ;
  assign n27385 = ( ~n11096 & n12402 ) | ( ~n11096 & n27384 ) | ( n12402 & n27384 ) ;
  assign n27386 = ( ~n8798 & n16346 ) | ( ~n8798 & n20732 ) | ( n16346 & n20732 ) ;
  assign n27387 = n27386 ^ n1838 ^ n765 ;
  assign n27388 = n16536 ^ n9683 ^ n4248 ;
  assign n27389 = n27388 ^ n10228 ^ n7535 ;
  assign n27392 = n12308 ^ n2018 ^ n855 ;
  assign n27390 = ( n951 & ~n3713 ) | ( n951 & n5782 ) | ( ~n3713 & n5782 ) ;
  assign n27391 = n17791 & ~n27390 ;
  assign n27393 = n27392 ^ n27391 ^ n25860 ;
  assign n27394 = ~n4090 & n27030 ;
  assign n27395 = n27394 ^ n17649 ^ 1'b0 ;
  assign n27396 = n8932 | n14289 ;
  assign n27397 = n27396 ^ n10425 ^ 1'b0 ;
  assign n27399 = ( n2446 & n8729 ) | ( n2446 & ~n10070 ) | ( n8729 & ~n10070 ) ;
  assign n27398 = n22069 ^ n15623 ^ n814 ;
  assign n27400 = n27399 ^ n27398 ^ n1793 ;
  assign n27401 = ~n4703 & n7140 ;
  assign n27405 = ( n4648 & ~n4867 ) | ( n4648 & n15382 ) | ( ~n4867 & n15382 ) ;
  assign n27402 = n15404 ^ n11471 ^ 1'b0 ;
  assign n27403 = n10928 & ~n27402 ;
  assign n27404 = n27403 ^ n20863 ^ 1'b0 ;
  assign n27406 = n27405 ^ n27404 ^ n6060 ;
  assign n27407 = n19201 ^ n10495 ^ n7740 ;
  assign n27408 = ( n2315 & n10191 ) | ( n2315 & n17176 ) | ( n10191 & n17176 ) ;
  assign n27409 = n1158 & n26074 ;
  assign n27410 = n12261 ^ n1726 ^ 1'b0 ;
  assign n27411 = ~n8448 & n27410 ;
  assign n27412 = n7013 & n21301 ;
  assign n27413 = n27412 ^ n4132 ^ 1'b0 ;
  assign n27414 = n1534 | n1668 ;
  assign n27415 = n9884 & ~n9891 ;
  assign n27416 = n27415 ^ n21274 ^ 1'b0 ;
  assign n27417 = n502 & n27416 ;
  assign n27418 = ( n9860 & ~n11552 ) | ( n9860 & n11763 ) | ( ~n11552 & n11763 ) ;
  assign n27421 = ( n1854 & n4052 ) | ( n1854 & ~n6005 ) | ( n4052 & ~n6005 ) ;
  assign n27419 = n13821 ^ n5885 ^ x113 ;
  assign n27420 = n27419 ^ n19837 ^ n5660 ;
  assign n27422 = n27421 ^ n27420 ^ n13836 ;
  assign n27423 = ( ~n11983 & n27418 ) | ( ~n11983 & n27422 ) | ( n27418 & n27422 ) ;
  assign n27424 = n13272 ^ n4106 ^ 1'b0 ;
  assign n27425 = ( n16237 & n26814 ) | ( n16237 & ~n27424 ) | ( n26814 & ~n27424 ) ;
  assign n27426 = ( n1940 & n7834 ) | ( n1940 & ~n27425 ) | ( n7834 & ~n27425 ) ;
  assign n27427 = ~n14133 & n27426 ;
  assign n27428 = n22110 & n27427 ;
  assign n27429 = n21333 ^ n15528 ^ n14166 ;
  assign n27430 = n22598 ^ n20058 ^ n11702 ;
  assign n27431 = ( x49 & n960 ) | ( x49 & n27430 ) | ( n960 & n27430 ) ;
  assign n27432 = n3284 & ~n5432 ;
  assign n27433 = n1130 | n6087 ;
  assign n27434 = n27433 ^ n14715 ^ 1'b0 ;
  assign n27435 = ( n2311 & n6364 ) | ( n2311 & ~n7428 ) | ( n6364 & ~n7428 ) ;
  assign n27436 = n6200 & ~n27435 ;
  assign n27437 = ( n3444 & n8120 ) | ( n3444 & n8311 ) | ( n8120 & n8311 ) ;
  assign n27442 = n24708 ^ n17266 ^ n17243 ;
  assign n27440 = n16976 ^ n12537 ^ n588 ;
  assign n27438 = ( n4629 & n9396 ) | ( n4629 & n10287 ) | ( n9396 & n10287 ) ;
  assign n27439 = n27438 ^ n6306 ^ 1'b0 ;
  assign n27441 = n27440 ^ n27439 ^ n14680 ;
  assign n27443 = n27442 ^ n27441 ^ n12709 ;
  assign n27444 = ~n6482 & n21663 ;
  assign n27445 = n27425 ^ n19693 ^ n18288 ;
  assign n27446 = ( n1348 & n9642 ) | ( n1348 & n27374 ) | ( n9642 & n27374 ) ;
  assign n27447 = n27446 ^ n7568 ^ x68 ;
  assign n27448 = n19712 ^ n14604 ^ n7462 ;
  assign n27449 = n6676 | n27448 ;
  assign n27450 = n6650 | n27449 ;
  assign n27451 = ~n18111 & n27450 ;
  assign n27452 = n27451 ^ n19082 ^ 1'b0 ;
  assign n27453 = n18747 ^ n7651 ^ 1'b0 ;
  assign n27454 = ( ~n8934 & n18683 ) | ( ~n8934 & n27453 ) | ( n18683 & n27453 ) ;
  assign n27455 = n17308 ^ n11438 ^ n1263 ;
  assign n27458 = ( n1770 & n12506 ) | ( n1770 & ~n15898 ) | ( n12506 & ~n15898 ) ;
  assign n27456 = n8191 ^ n5358 ^ n1287 ;
  assign n27457 = ( n6782 & n7126 ) | ( n6782 & n27456 ) | ( n7126 & n27456 ) ;
  assign n27459 = n27458 ^ n27457 ^ n5566 ;
  assign n27460 = n26956 ^ n18933 ^ n1408 ;
  assign n27461 = n17590 ^ n11868 ^ n9857 ;
  assign n27464 = n848 | n8035 ;
  assign n27465 = n27464 ^ n22895 ^ 1'b0 ;
  assign n27462 = n25571 ^ n18963 ^ 1'b0 ;
  assign n27463 = n27462 ^ n19423 ^ 1'b0 ;
  assign n27466 = n27465 ^ n27463 ^ 1'b0 ;
  assign n27467 = ( n7985 & n13415 ) | ( n7985 & ~n21535 ) | ( n13415 & ~n21535 ) ;
  assign n27468 = n4231 & n27467 ;
  assign n27475 = n19154 ^ n242 ^ 1'b0 ;
  assign n27476 = n27475 ^ n24026 ^ n6606 ;
  assign n27477 = n27476 ^ n20564 ^ n2973 ;
  assign n27470 = n4916 ^ n167 ^ 1'b0 ;
  assign n27471 = n22110 | n27470 ;
  assign n27472 = n27471 ^ n22410 ^ n18571 ;
  assign n27473 = n4652 & ~n27472 ;
  assign n27474 = n27473 ^ n15734 ^ 1'b0 ;
  assign n27469 = ( n3716 & n8374 ) | ( n3716 & n27359 ) | ( n8374 & n27359 ) ;
  assign n27478 = n27477 ^ n27474 ^ n27469 ;
  assign n27479 = n12284 | n21447 ;
  assign n27480 = n27479 ^ n2843 ^ 1'b0 ;
  assign n27486 = n10421 | n12519 ;
  assign n27487 = n27475 & ~n27486 ;
  assign n27488 = n27487 ^ n2247 ^ 1'b0 ;
  assign n27485 = n19722 ^ n18807 ^ n4241 ;
  assign n27481 = n19287 ^ n5827 ^ n4530 ;
  assign n27482 = n16317 ^ n9594 ^ 1'b0 ;
  assign n27483 = ~n27481 & n27482 ;
  assign n27484 = ( n307 & n22530 ) | ( n307 & n27483 ) | ( n22530 & n27483 ) ;
  assign n27489 = n27488 ^ n27485 ^ n27484 ;
  assign n27490 = n24889 ^ n4704 ^ 1'b0 ;
  assign n27491 = n27490 ^ n7243 ^ n907 ;
  assign n27492 = n27491 ^ n21070 ^ 1'b0 ;
  assign n27493 = n24744 ^ n23736 ^ n9017 ;
  assign n27494 = n2408 & ~n19422 ;
  assign n27495 = n27494 ^ n5504 ^ 1'b0 ;
  assign n27496 = ( ~n10020 & n25795 ) | ( ~n10020 & n27495 ) | ( n25795 & n27495 ) ;
  assign n27497 = n9959 & n12617 ;
  assign n27498 = ( n5933 & ~n20291 ) | ( n5933 & n20317 ) | ( ~n20291 & n20317 ) ;
  assign n27499 = n27498 ^ n23172 ^ n4388 ;
  assign n27501 = n18412 ^ n14929 ^ n5656 ;
  assign n27500 = n27158 ^ n8273 ^ n5982 ;
  assign n27502 = n27501 ^ n27500 ^ n918 ;
  assign n27503 = ( ~n1102 & n14178 ) | ( ~n1102 & n22427 ) | ( n14178 & n22427 ) ;
  assign n27504 = ( n280 & n15110 ) | ( n280 & n16109 ) | ( n15110 & n16109 ) ;
  assign n27505 = n27504 ^ n2051 ^ 1'b0 ;
  assign n27506 = n7186 & n27505 ;
  assign n27507 = n27506 ^ n16483 ^ 1'b0 ;
  assign n27508 = ( n1179 & n5878 ) | ( n1179 & n18640 ) | ( n5878 & n18640 ) ;
  assign n27509 = n27508 ^ n13433 ^ n2541 ;
  assign n27510 = ( n1679 & n21784 ) | ( n1679 & n24291 ) | ( n21784 & n24291 ) ;
  assign n27511 = ( n22305 & n27509 ) | ( n22305 & n27510 ) | ( n27509 & n27510 ) ;
  assign n27512 = ( n1480 & n8359 ) | ( n1480 & n27197 ) | ( n8359 & n27197 ) ;
  assign n27513 = ( n1821 & n2425 ) | ( n1821 & ~n3431 ) | ( n2425 & ~n3431 ) ;
  assign n27514 = n17795 & ~n27513 ;
  assign n27515 = ( n5615 & n8938 ) | ( n5615 & ~n27514 ) | ( n8938 & ~n27514 ) ;
  assign n27516 = ( n24905 & n27512 ) | ( n24905 & ~n27515 ) | ( n27512 & ~n27515 ) ;
  assign n27517 = n23990 ^ n12886 ^ n824 ;
  assign n27518 = ( n3171 & n7991 ) | ( n3171 & n27517 ) | ( n7991 & n27517 ) ;
  assign n27519 = ( n18302 & ~n19986 ) | ( n18302 & n27518 ) | ( ~n19986 & n27518 ) ;
  assign n27520 = n2026 & n5260 ;
  assign n27521 = ~n13975 & n27520 ;
  assign n27522 = n12901 ^ n5855 ^ 1'b0 ;
  assign n27523 = n8748 | n27522 ;
  assign n27524 = ( n24658 & ~n25238 ) | ( n24658 & n27166 ) | ( ~n25238 & n27166 ) ;
  assign n27525 = n5703 ^ n5210 ^ n4477 ;
  assign n27526 = ( n9939 & n21746 ) | ( n9939 & ~n27525 ) | ( n21746 & ~n27525 ) ;
  assign n27527 = ( n10276 & n21455 ) | ( n10276 & n27526 ) | ( n21455 & n27526 ) ;
  assign n27530 = ( n357 & n7525 ) | ( n357 & n9630 ) | ( n7525 & n9630 ) ;
  assign n27531 = n27530 ^ n9431 ^ 1'b0 ;
  assign n27528 = ( ~n494 & n12385 ) | ( ~n494 & n21387 ) | ( n12385 & n21387 ) ;
  assign n27529 = n27087 & ~n27528 ;
  assign n27532 = n27531 ^ n27529 ^ 1'b0 ;
  assign n27533 = n27532 ^ n19838 ^ 1'b0 ;
  assign n27534 = ( n1701 & n10842 ) | ( n1701 & ~n27533 ) | ( n10842 & ~n27533 ) ;
  assign n27535 = n27534 ^ n19115 ^ n13391 ;
  assign n27536 = n17403 ^ n12113 ^ n6006 ;
  assign n27537 = n27536 ^ n9972 ^ n2895 ;
  assign n27540 = n5040 ^ n4045 ^ n2010 ;
  assign n27538 = ( n5931 & n15713 ) | ( n5931 & n15838 ) | ( n15713 & n15838 ) ;
  assign n27539 = n27538 ^ n25371 ^ n16471 ;
  assign n27541 = n27540 ^ n27539 ^ n5768 ;
  assign n27542 = n27405 ^ n11063 ^ n229 ;
  assign n27543 = n15692 ^ n6042 ^ n3984 ;
  assign n27544 = n27543 ^ n21992 ^ n1955 ;
  assign n27546 = n24770 ^ n22217 ^ 1'b0 ;
  assign n27547 = n27546 ^ n12276 ^ n7539 ;
  assign n27545 = ( n1928 & ~n4203 ) | ( n1928 & n4559 ) | ( ~n4203 & n4559 ) ;
  assign n27548 = n27547 ^ n27545 ^ 1'b0 ;
  assign n27549 = n5498 & n20062 ;
  assign n27550 = n27549 ^ n17781 ^ 1'b0 ;
  assign n27551 = n10523 ^ n1465 ^ n634 ;
  assign n27552 = ~n10460 & n27551 ;
  assign n27553 = n27552 ^ n6586 ^ 1'b0 ;
  assign n27554 = ( n8570 & ~n17885 ) | ( n8570 & n25087 ) | ( ~n17885 & n25087 ) ;
  assign n27555 = n20313 ^ n14611 ^ n10309 ;
  assign n27556 = ( ~x111 & n2390 ) | ( ~x111 & n7194 ) | ( n2390 & n7194 ) ;
  assign n27557 = ( ~n4297 & n9184 ) | ( ~n4297 & n27556 ) | ( n9184 & n27556 ) ;
  assign n27558 = ( n18576 & n23691 ) | ( n18576 & n27557 ) | ( n23691 & n27557 ) ;
  assign n27559 = n6982 ^ n2501 ^ n503 ;
  assign n27560 = n16284 ^ n15814 ^ n228 ;
  assign n27561 = ( n22526 & n27559 ) | ( n22526 & ~n27560 ) | ( n27559 & ~n27560 ) ;
  assign n27562 = ( n26670 & n27558 ) | ( n26670 & ~n27561 ) | ( n27558 & ~n27561 ) ;
  assign n27563 = ( n5644 & n17816 ) | ( n5644 & ~n19753 ) | ( n17816 & ~n19753 ) ;
  assign n27564 = n27563 ^ n14632 ^ 1'b0 ;
  assign n27565 = n6176 ^ n2218 ^ n646 ;
  assign n27566 = n27565 ^ n23413 ^ n5522 ;
  assign n27567 = ( ~n10954 & n13876 ) | ( ~n10954 & n14896 ) | ( n13876 & n14896 ) ;
  assign n27568 = ~n1474 & n10465 ;
  assign n27569 = ( ~n3827 & n3999 ) | ( ~n3827 & n18922 ) | ( n3999 & n18922 ) ;
  assign n27570 = ( ~n16996 & n27568 ) | ( ~n16996 & n27569 ) | ( n27568 & n27569 ) ;
  assign n27571 = ( n7361 & n27567 ) | ( n7361 & n27570 ) | ( n27567 & n27570 ) ;
  assign n27572 = n15296 ^ n8787 ^ n6214 ;
  assign n27573 = n27572 ^ n9966 ^ n3213 ;
  assign n27574 = ( n3740 & n5136 ) | ( n3740 & n21695 ) | ( n5136 & n21695 ) ;
  assign n27575 = n27574 ^ n21556 ^ n19139 ;
  assign n27576 = n27575 ^ n19920 ^ n5546 ;
  assign n27577 = n15960 & n16428 ;
  assign n27578 = n27576 & n27577 ;
  assign n27579 = n8405 ^ n7949 ^ n5454 ;
  assign n27580 = ( n11333 & n17006 ) | ( n11333 & n22520 ) | ( n17006 & n22520 ) ;
  assign n27581 = ( n20415 & n27579 ) | ( n20415 & n27580 ) | ( n27579 & n27580 ) ;
  assign n27582 = n15675 ^ n2566 ^ 1'b0 ;
  assign n27583 = n27581 & ~n27582 ;
  assign n27584 = n13421 ^ n10704 ^ n1919 ;
  assign n27585 = n11003 & n22642 ;
  assign n27586 = ~n27176 & n27585 ;
  assign n27588 = n8634 ^ n5029 ^ n3758 ;
  assign n27589 = n27588 ^ n17729 ^ n12172 ;
  assign n27587 = ( n404 & ~n5533 ) | ( n404 & n25781 ) | ( ~n5533 & n25781 ) ;
  assign n27590 = n27589 ^ n27587 ^ n942 ;
  assign n27591 = n14478 ^ n6352 ^ n2434 ;
  assign n27592 = n23840 ^ n17625 ^ n454 ;
  assign n27594 = n18436 ^ n6553 ^ n2568 ;
  assign n27593 = ( n2167 & n4060 ) | ( n2167 & n25134 ) | ( n4060 & n25134 ) ;
  assign n27595 = n27594 ^ n27593 ^ n16741 ;
  assign n27596 = ( ~n4045 & n19757 ) | ( ~n4045 & n27595 ) | ( n19757 & n27595 ) ;
  assign n27598 = n8497 ^ n6430 ^ n4711 ;
  assign n27597 = n17543 | n18897 ;
  assign n27599 = n27598 ^ n27597 ^ n22444 ;
  assign n27600 = ( n4146 & ~n5037 ) | ( n4146 & n21340 ) | ( ~n5037 & n21340 ) ;
  assign n27601 = n12696 ^ n11014 ^ n8881 ;
  assign n27602 = n27601 ^ n3684 ^ 1'b0 ;
  assign n27603 = n4775 & ~n27602 ;
  assign n27604 = ( n13192 & n16681 ) | ( n13192 & ~n27603 ) | ( n16681 & ~n27603 ) ;
  assign n27605 = ( n10658 & n13003 ) | ( n10658 & n21075 ) | ( n13003 & n21075 ) ;
  assign n27606 = n8099 & n24887 ;
  assign n27607 = n27605 & n27606 ;
  assign n27608 = n13971 ^ n10297 ^ n10098 ;
  assign n27609 = n27608 ^ n5016 ^ n1240 ;
  assign n27610 = n27609 ^ n10029 ^ n2942 ;
  assign n27611 = n27458 ^ n16369 ^ n3466 ;
  assign n27612 = n13518 & n27611 ;
  assign n27613 = ( n8309 & n9585 ) | ( n8309 & n24145 ) | ( n9585 & n24145 ) ;
  assign n27615 = n2924 & ~n11298 ;
  assign n27616 = n27615 ^ n23331 ^ 1'b0 ;
  assign n27614 = ( n1269 & n10012 ) | ( n1269 & ~n11890 ) | ( n10012 & ~n11890 ) ;
  assign n27617 = n27616 ^ n27614 ^ n14136 ;
  assign n27618 = n27617 ^ n3244 ^ n694 ;
  assign n27624 = n3183 & ~n3817 ;
  assign n27625 = n18931 & n27624 ;
  assign n27619 = n4759 ^ n3214 ^ n985 ;
  assign n27620 = n357 & ~n27619 ;
  assign n27621 = ~n9307 & n27620 ;
  assign n27622 = n27621 ^ n19026 ^ n13080 ;
  assign n27623 = n27622 ^ n19198 ^ 1'b0 ;
  assign n27626 = n27625 ^ n27623 ^ n12607 ;
  assign n27627 = n17197 ^ n13125 ^ n8858 ;
  assign n27628 = ( ~n3961 & n23999 ) | ( ~n3961 & n27627 ) | ( n23999 & n27627 ) ;
  assign n27629 = n26027 ^ n16492 ^ n5579 ;
  assign n27630 = ( n6541 & n14769 ) | ( n6541 & n27629 ) | ( n14769 & n27629 ) ;
  assign n27631 = n11768 ^ n264 ^ 1'b0 ;
  assign n27632 = n24348 & n27631 ;
  assign n27633 = n14745 ^ n1032 ^ 1'b0 ;
  assign n27634 = ( n12938 & n21491 ) | ( n12938 & n27633 ) | ( n21491 & n27633 ) ;
  assign n27635 = ( ~n4760 & n15709 ) | ( ~n4760 & n27634 ) | ( n15709 & n27634 ) ;
  assign n27636 = n17433 ^ n9477 ^ 1'b0 ;
  assign n27637 = n27211 ^ n15837 ^ n10372 ;
  assign n27638 = n13428 ^ n13187 ^ n3161 ;
  assign n27639 = n9744 | n27638 ;
  assign n27640 = n27639 ^ n21332 ^ n20047 ;
  assign n27643 = n24891 ^ n23182 ^ n4667 ;
  assign n27641 = ( ~n681 & n2808 ) | ( ~n681 & n12258 ) | ( n2808 & n12258 ) ;
  assign n27642 = n27641 ^ n4651 ^ 1'b0 ;
  assign n27644 = n27643 ^ n27642 ^ n3484 ;
  assign n27645 = n22240 ^ n15110 ^ n439 ;
  assign n27646 = ( n12954 & n14532 ) | ( n12954 & n25087 ) | ( n14532 & n25087 ) ;
  assign n27647 = ( n4711 & ~n20250 ) | ( n4711 & n24569 ) | ( ~n20250 & n24569 ) ;
  assign n27648 = ( n9062 & ~n11253 ) | ( n9062 & n27647 ) | ( ~n11253 & n27647 ) ;
  assign n27649 = ( x14 & ~n8624 ) | ( x14 & n27281 ) | ( ~n8624 & n27281 ) ;
  assign n27650 = ( n6694 & n21556 ) | ( n6694 & n27649 ) | ( n21556 & n27649 ) ;
  assign n27651 = ( n14810 & ~n20868 ) | ( n14810 & n27650 ) | ( ~n20868 & n27650 ) ;
  assign n27652 = ( n9591 & n27648 ) | ( n9591 & n27651 ) | ( n27648 & n27651 ) ;
  assign n27655 = ( ~n3697 & n11480 ) | ( ~n3697 & n19282 ) | ( n11480 & n19282 ) ;
  assign n27654 = ( ~n3102 & n18745 ) | ( ~n3102 & n21152 ) | ( n18745 & n21152 ) ;
  assign n27653 = ( n18989 & n26418 ) | ( n18989 & ~n26463 ) | ( n26418 & ~n26463 ) ;
  assign n27656 = n27655 ^ n27654 ^ n27653 ;
  assign n27657 = ( n230 & n5699 ) | ( n230 & ~n16342 ) | ( n5699 & ~n16342 ) ;
  assign n27658 = ( n3926 & n8125 ) | ( n3926 & n19313 ) | ( n8125 & n19313 ) ;
  assign n27659 = n11493 ^ n10203 ^ n1624 ;
  assign n27660 = n27659 ^ n21387 ^ 1'b0 ;
  assign n27661 = n27660 ^ n26577 ^ n18481 ;
  assign n27662 = n2486 & ~n16967 ;
  assign n27663 = n5369 & n27662 ;
  assign n27664 = ( ~x118 & n1166 ) | ( ~x118 & n27663 ) | ( n1166 & n27663 ) ;
  assign n27665 = n27664 ^ n22436 ^ n17996 ;
  assign n27666 = n20363 ^ n3870 ^ n1261 ;
  assign n27667 = ( n16147 & n23045 ) | ( n16147 & ~n27666 ) | ( n23045 & ~n27666 ) ;
  assign n27668 = ( n1192 & n4499 ) | ( n1192 & ~n9107 ) | ( n4499 & ~n9107 ) ;
  assign n27669 = ( n23034 & ~n25040 ) | ( n23034 & n27668 ) | ( ~n25040 & n27668 ) ;
  assign n27670 = ( n3574 & n9370 ) | ( n3574 & ~n13900 ) | ( n9370 & ~n13900 ) ;
  assign n27671 = ( n2288 & n5019 ) | ( n2288 & n27670 ) | ( n5019 & n27670 ) ;
  assign n27672 = ( ~n897 & n27669 ) | ( ~n897 & n27671 ) | ( n27669 & n27671 ) ;
  assign n27673 = ( n5333 & n19323 ) | ( n5333 & n20465 ) | ( n19323 & n20465 ) ;
  assign n27674 = ( ~n7717 & n14001 ) | ( ~n7717 & n27673 ) | ( n14001 & n27673 ) ;
  assign n27675 = n12178 ^ n4447 ^ n1146 ;
  assign n27676 = n27675 ^ n12865 ^ 1'b0 ;
  assign n27677 = ( ~n4396 & n7387 ) | ( ~n4396 & n9333 ) | ( n7387 & n9333 ) ;
  assign n27678 = n3583 ^ n2047 ^ 1'b0 ;
  assign n27679 = n27677 & ~n27678 ;
  assign n27680 = n27679 ^ n25724 ^ n15625 ;
  assign n27681 = ( ~n1176 & n2765 ) | ( ~n1176 & n4562 ) | ( n2765 & n4562 ) ;
  assign n27682 = n27681 ^ n5820 ^ x27 ;
  assign n27683 = n19492 ^ n168 ^ 1'b0 ;
  assign n27684 = n1676 & n27683 ;
  assign n27685 = ~n16196 & n27684 ;
  assign n27686 = ( n3741 & n7491 ) | ( n3741 & ~n26343 ) | ( n7491 & ~n26343 ) ;
  assign n27687 = n10246 ^ n5059 ^ 1'b0 ;
  assign n27688 = n4044 & n27687 ;
  assign n27689 = n7143 ^ n5773 ^ n2776 ;
  assign n27690 = n27689 ^ n15560 ^ n13561 ;
  assign n27691 = ( n4964 & n14417 ) | ( n4964 & ~n27690 ) | ( n14417 & ~n27690 ) ;
  assign n27695 = ( n2235 & n2929 ) | ( n2235 & n15565 ) | ( n2929 & n15565 ) ;
  assign n27692 = ( ~x85 & n9670 ) | ( ~x85 & n14648 ) | ( n9670 & n14648 ) ;
  assign n27693 = n27692 ^ n12094 ^ n4368 ;
  assign n27694 = n27693 ^ n19089 ^ 1'b0 ;
  assign n27696 = n27695 ^ n27694 ^ n19758 ;
  assign n27697 = ( n6612 & n7816 ) | ( n6612 & n27696 ) | ( n7816 & n27696 ) ;
  assign n27698 = ( n575 & n10688 ) | ( n575 & ~n15911 ) | ( n10688 & ~n15911 ) ;
  assign n27699 = ~n11535 & n27698 ;
  assign n27700 = ( n13964 & n18368 ) | ( n13964 & ~n27699 ) | ( n18368 & ~n27699 ) ;
  assign n27701 = ( n2716 & ~n6947 ) | ( n2716 & n27700 ) | ( ~n6947 & n27700 ) ;
  assign n27702 = ( n2848 & n19064 ) | ( n2848 & ~n19816 ) | ( n19064 & ~n19816 ) ;
  assign n27703 = n22640 ^ n15518 ^ n10065 ;
  assign n27704 = n27702 & ~n27703 ;
  assign n27705 = n15494 ^ n12787 ^ n4668 ;
  assign n27706 = ( ~n4167 & n15929 ) | ( ~n4167 & n23662 ) | ( n15929 & n23662 ) ;
  assign n27707 = n10642 ^ n4854 ^ 1'b0 ;
  assign n27708 = n12850 | n27707 ;
  assign n27709 = n27708 ^ n19265 ^ n8302 ;
  assign n27710 = n1555 & ~n11143 ;
  assign n27711 = n17887 & ~n27710 ;
  assign n27712 = n27709 & n27711 ;
  assign n27713 = ( ~n2877 & n4892 ) | ( ~n2877 & n11252 ) | ( n4892 & n11252 ) ;
  assign n27714 = n27713 ^ n2981 ^ 1'b0 ;
  assign n27715 = ( ~n7817 & n15446 ) | ( ~n7817 & n27714 ) | ( n15446 & n27714 ) ;
  assign n27716 = ~n5725 & n19366 ;
  assign n27717 = n27627 ^ n11121 ^ n9246 ;
  assign n27718 = n17609 ^ n15130 ^ n12000 ;
  assign n27719 = ( n3415 & n10524 ) | ( n3415 & ~n24206 ) | ( n10524 & ~n24206 ) ;
  assign n27720 = n21614 ^ n16344 ^ n8089 ;
  assign n27721 = n18575 ^ n5680 ^ 1'b0 ;
  assign n27722 = ( n6102 & n15371 ) | ( n6102 & ~n27425 ) | ( n15371 & ~n27425 ) ;
  assign n27723 = ( n12704 & ~n27721 ) | ( n12704 & n27722 ) | ( ~n27721 & n27722 ) ;
  assign n27724 = n27723 ^ n22457 ^ n6396 ;
  assign n27725 = n3709 & n6901 ;
  assign n27726 = n27725 ^ n20191 ^ 1'b0 ;
  assign n27727 = n15247 & ~n27381 ;
  assign n27728 = ~n14468 & n27727 ;
  assign n27729 = ( ~n9836 & n13882 ) | ( ~n9836 & n19986 ) | ( n13882 & n19986 ) ;
  assign n27730 = n17797 ^ n16223 ^ n10831 ;
  assign n27731 = ( n5936 & ~n27729 ) | ( n5936 & n27730 ) | ( ~n27729 & n27730 ) ;
  assign n27732 = n27731 ^ n19874 ^ n6880 ;
  assign n27733 = n12317 ^ n7796 ^ n6280 ;
  assign n27734 = n27733 ^ n10178 ^ 1'b0 ;
  assign n27735 = n17885 ^ n11321 ^ n9980 ;
  assign n27736 = n27735 ^ n10076 ^ n5359 ;
  assign n27737 = n15363 ^ n10680 ^ n4566 ;
  assign n27739 = n6240 | n23656 ;
  assign n27740 = n27739 ^ n1037 ^ 1'b0 ;
  assign n27738 = n25887 ^ n13920 ^ n11584 ;
  assign n27741 = n27740 ^ n27738 ^ n14786 ;
  assign n27742 = ( n251 & ~n1640 ) | ( n251 & n3871 ) | ( ~n1640 & n3871 ) ;
  assign n27743 = ( n313 & n18801 ) | ( n313 & n27742 ) | ( n18801 & n27742 ) ;
  assign n27744 = ( n948 & n9431 ) | ( n948 & n14588 ) | ( n9431 & n14588 ) ;
  assign n27745 = n27744 ^ n26615 ^ n20183 ;
  assign n27746 = ( n18636 & ~n27743 ) | ( n18636 & n27745 ) | ( ~n27743 & n27745 ) ;
  assign n27747 = ( n3687 & n8122 ) | ( n3687 & ~n13579 ) | ( n8122 & ~n13579 ) ;
  assign n27748 = ( n24113 & n25169 ) | ( n24113 & n27747 ) | ( n25169 & n27747 ) ;
  assign n27749 = n11595 ^ n8762 ^ n7917 ;
  assign n27750 = ( n15081 & ~n21519 ) | ( n15081 & n23932 ) | ( ~n21519 & n23932 ) ;
  assign n27751 = ( n7165 & n27749 ) | ( n7165 & ~n27750 ) | ( n27749 & ~n27750 ) ;
  assign n27752 = n19211 & n27751 ;
  assign n27753 = ~n13551 & n27752 ;
  assign n27754 = ( ~n8661 & n11195 ) | ( ~n8661 & n24701 ) | ( n11195 & n24701 ) ;
  assign n27755 = ( n9381 & n9874 ) | ( n9381 & ~n14209 ) | ( n9874 & ~n14209 ) ;
  assign n27756 = ( n1375 & ~n1447 ) | ( n1375 & n27755 ) | ( ~n1447 & n27755 ) ;
  assign n27757 = ( n4639 & n8869 ) | ( n4639 & ~n9035 ) | ( n8869 & ~n9035 ) ;
  assign n27758 = n27757 ^ n20392 ^ n9584 ;
  assign n27759 = ~n15220 & n18459 ;
  assign n27760 = ( n5400 & n21724 ) | ( n5400 & n27759 ) | ( n21724 & n27759 ) ;
  assign n27761 = ( n10939 & n23190 ) | ( n10939 & ~n27760 ) | ( n23190 & ~n27760 ) ;
  assign n27763 = n3197 & ~n25563 ;
  assign n27762 = n25727 ^ n25295 ^ n7676 ;
  assign n27764 = n27763 ^ n27762 ^ n7738 ;
  assign n27765 = n22780 ^ n11096 ^ n2115 ;
  assign n27766 = n20449 | n27765 ;
  assign n27769 = n9967 ^ n8094 ^ n833 ;
  assign n27770 = n27769 ^ n9821 ^ n9661 ;
  assign n27771 = ( ~n12236 & n23366 ) | ( ~n12236 & n27770 ) | ( n23366 & n27770 ) ;
  assign n27767 = n8991 ^ n3371 ^ 1'b0 ;
  assign n27768 = n27767 ^ n25757 ^ n22144 ;
  assign n27772 = n27771 ^ n27768 ^ n2811 ;
  assign n27773 = n7808 ^ n2401 ^ 1'b0 ;
  assign n27774 = ( n7581 & n10186 ) | ( n7581 & n26222 ) | ( n10186 & n26222 ) ;
  assign n27775 = n7505 ^ n4056 ^ n2106 ;
  assign n27776 = n21063 ^ n15864 ^ n15623 ;
  assign n27777 = n6243 ^ n4365 ^ n3222 ;
  assign n27778 = n18740 ^ n1438 ^ 1'b0 ;
  assign n27779 = n9386 & ~n27778 ;
  assign n27780 = n13404 ^ n12030 ^ n178 ;
  assign n27781 = n26070 ^ n16719 ^ n12890 ;
  assign n27782 = n27781 ^ n5970 ^ n2217 ;
  assign n27783 = ( ~n10194 & n11901 ) | ( ~n10194 & n18006 ) | ( n11901 & n18006 ) ;
  assign n27785 = n8380 ^ n6229 ^ n347 ;
  assign n27784 = n13185 | n27651 ;
  assign n27786 = n27785 ^ n27784 ^ 1'b0 ;
  assign n27787 = ( n15439 & ~n25593 ) | ( n15439 & n27786 ) | ( ~n25593 & n27786 ) ;
  assign n27789 = n16462 ^ n9933 ^ n5989 ;
  assign n27788 = n23576 ^ n21788 ^ n21601 ;
  assign n27790 = n27789 ^ n27788 ^ n20279 ;
  assign n27791 = ( ~n4779 & n14062 ) | ( ~n4779 & n18497 ) | ( n14062 & n18497 ) ;
  assign n27792 = ( n785 & n3444 ) | ( n785 & n11768 ) | ( n3444 & n11768 ) ;
  assign n27793 = ~n486 & n9851 ;
  assign n27794 = ~n27792 & n27793 ;
  assign n27795 = n27794 ^ n25035 ^ n2107 ;
  assign n27796 = ( n6484 & n7605 ) | ( n6484 & ~n14942 ) | ( n7605 & ~n14942 ) ;
  assign n27801 = n12163 ^ n4787 ^ n592 ;
  assign n27797 = n13571 & n15755 ;
  assign n27798 = n27797 ^ n5757 ^ 1'b0 ;
  assign n27799 = n10808 ^ n10102 ^ n6116 ;
  assign n27800 = ( n14570 & n27798 ) | ( n14570 & ~n27799 ) | ( n27798 & ~n27799 ) ;
  assign n27802 = n27801 ^ n27800 ^ n24128 ;
  assign n27803 = n23149 ^ n3504 ^ n1630 ;
  assign n27804 = n21655 ^ n6407 ^ 1'b0 ;
  assign n27805 = n25319 ^ n23078 ^ n2552 ;
  assign n27806 = n27805 ^ n23911 ^ n21507 ;
  assign n27807 = n11696 ^ n3090 ^ n2352 ;
  assign n27808 = ( ~n15379 & n25226 ) | ( ~n15379 & n27807 ) | ( n25226 & n27807 ) ;
  assign n27809 = ( ~n3199 & n5033 ) | ( ~n3199 & n13459 ) | ( n5033 & n13459 ) ;
  assign n27810 = ( n8666 & ~n13910 ) | ( n8666 & n27809 ) | ( ~n13910 & n27809 ) ;
  assign n27811 = n27810 ^ n4313 ^ x24 ;
  assign n27812 = n7764 ^ n5762 ^ 1'b0 ;
  assign n27813 = n11894 & n27812 ;
  assign n27814 = n21096 ^ n10671 ^ 1'b0 ;
  assign n27815 = n6668 & n27814 ;
  assign n27816 = ( n4163 & n4288 ) | ( n4163 & ~n20196 ) | ( n4288 & ~n20196 ) ;
  assign n27817 = n27816 ^ n636 ^ 1'b0 ;
  assign n27818 = n14061 ^ n12816 ^ n10815 ;
  assign n27819 = ( n12604 & n14072 ) | ( n12604 & ~n27818 ) | ( n14072 & ~n27818 ) ;
  assign n27820 = ( n12524 & n14159 ) | ( n12524 & n27819 ) | ( n14159 & n27819 ) ;
  assign n27821 = n17460 ^ n8646 ^ n6328 ;
  assign n27822 = n27821 ^ n14895 ^ n11187 ;
  assign n27823 = n826 | n18982 ;
  assign n27824 = ( n16711 & n27822 ) | ( n16711 & n27823 ) | ( n27822 & n27823 ) ;
  assign n27825 = ( n4301 & n13121 ) | ( n4301 & n17821 ) | ( n13121 & n17821 ) ;
  assign n27826 = n12612 ^ n6796 ^ n1032 ;
  assign n27827 = ( n1809 & ~n21484 ) | ( n1809 & n27826 ) | ( ~n21484 & n27826 ) ;
  assign n27828 = ( n949 & n7340 ) | ( n949 & ~n25427 ) | ( n7340 & ~n25427 ) ;
  assign n27829 = n3815 ^ n2021 ^ n248 ;
  assign n27830 = ( n13355 & n16290 ) | ( n13355 & n27829 ) | ( n16290 & n27829 ) ;
  assign n27831 = ( n2680 & ~n27828 ) | ( n2680 & n27830 ) | ( ~n27828 & n27830 ) ;
  assign n27832 = ( ~n2714 & n10485 ) | ( ~n2714 & n10626 ) | ( n10485 & n10626 ) ;
  assign n27833 = n20066 ^ n8735 ^ n543 ;
  assign n27834 = ( ~n12432 & n27832 ) | ( ~n12432 & n27833 ) | ( n27832 & n27833 ) ;
  assign n27835 = ~n6843 & n24469 ;
  assign n27836 = ~n14042 & n27835 ;
  assign n27837 = n15979 ^ n10219 ^ n2804 ;
  assign n27842 = n20036 ^ n16817 ^ n11422 ;
  assign n27839 = n2853 ^ n859 ^ n527 ;
  assign n27838 = ( ~n14280 & n21256 ) | ( ~n14280 & n27821 ) | ( n21256 & n27821 ) ;
  assign n27840 = n27839 ^ n27838 ^ n10708 ;
  assign n27841 = n27840 ^ n20524 ^ 1'b0 ;
  assign n27843 = n27842 ^ n27841 ^ n20812 ;
  assign n27844 = n27442 ^ n27384 ^ n1447 ;
  assign n27845 = ( n3407 & n4248 ) | ( n3407 & ~n6601 ) | ( n4248 & ~n6601 ) ;
  assign n27846 = n1148 | n14714 ;
  assign n27847 = n27846 ^ n2569 ^ 1'b0 ;
  assign n27851 = n17094 & ~n20584 ;
  assign n27852 = n27851 ^ n9265 ^ 1'b0 ;
  assign n27848 = n1104 & ~n1557 ;
  assign n27849 = n17178 ^ n12668 ^ n11500 ;
  assign n27850 = ( n4566 & n27848 ) | ( n4566 & ~n27849 ) | ( n27848 & ~n27849 ) ;
  assign n27853 = n27852 ^ n27850 ^ 1'b0 ;
  assign n27854 = n25871 ^ n23489 ^ n6077 ;
  assign n27855 = ( n843 & n11910 ) | ( n843 & n12760 ) | ( n11910 & n12760 ) ;
  assign n27856 = ( n17503 & ~n27854 ) | ( n17503 & n27855 ) | ( ~n27854 & n27855 ) ;
  assign n27857 = n11018 ^ n2768 ^ 1'b0 ;
  assign n27858 = n22811 ^ n9917 ^ n8768 ;
  assign n27859 = n11307 ^ n10527 ^ 1'b0 ;
  assign n27860 = n27858 & n27859 ;
  assign n27861 = ( n1299 & ~n17720 ) | ( n1299 & n19554 ) | ( ~n17720 & n19554 ) ;
  assign n27862 = n11456 & n27861 ;
  assign n27863 = n27664 & n27862 ;
  assign n27864 = ( n4334 & n10006 ) | ( n4334 & ~n27863 ) | ( n10006 & ~n27863 ) ;
  assign n27865 = n14788 & n16622 ;
  assign n27866 = ( n9349 & ~n17559 ) | ( n9349 & n21095 ) | ( ~n17559 & n21095 ) ;
  assign n27867 = n27866 ^ n19776 ^ n4289 ;
  assign n27868 = ( n27864 & n27865 ) | ( n27864 & ~n27867 ) | ( n27865 & ~n27867 ) ;
  assign n27874 = ( n3389 & n7658 ) | ( n3389 & n26254 ) | ( n7658 & n26254 ) ;
  assign n27871 = ( n8081 & n8437 ) | ( n8081 & ~n9975 ) | ( n8437 & ~n9975 ) ;
  assign n27872 = n19726 ^ n8382 ^ n5131 ;
  assign n27873 = ( ~n12402 & n27871 ) | ( ~n12402 & n27872 ) | ( n27871 & n27872 ) ;
  assign n27869 = n11407 ^ n4788 ^ 1'b0 ;
  assign n27870 = ~n12041 & n27869 ;
  assign n27875 = n27874 ^ n27873 ^ n27870 ;
  assign n27876 = ( n7654 & n11291 ) | ( n7654 & n15677 ) | ( n11291 & n15677 ) ;
  assign n27877 = n10125 ^ n3220 ^ n982 ;
  assign n27878 = ( n3202 & n8529 ) | ( n3202 & n27877 ) | ( n8529 & n27877 ) ;
  assign n27879 = ( ~n3118 & n7190 ) | ( ~n3118 & n27878 ) | ( n7190 & n27878 ) ;
  assign n27880 = ( ~n8537 & n21804 ) | ( ~n8537 & n26534 ) | ( n21804 & n26534 ) ;
  assign n27881 = n1135 | n2947 ;
  assign n27882 = n27668 ^ n2198 ^ 1'b0 ;
  assign n27883 = n3825 | n27882 ;
  assign n27884 = n13582 ^ n9688 ^ n3693 ;
  assign n27885 = n18989 | n27884 ;
  assign n27886 = n22030 & ~n27885 ;
  assign n27887 = ( n15872 & n20652 ) | ( n15872 & ~n24272 ) | ( n20652 & ~n24272 ) ;
  assign n27888 = ~n12142 & n13428 ;
  assign n27889 = n17407 & n27888 ;
  assign n27890 = ( n2493 & n12182 ) | ( n2493 & ~n27889 ) | ( n12182 & ~n27889 ) ;
  assign n27891 = n2188 | n5351 ;
  assign n27892 = n6991 & ~n27891 ;
  assign n27893 = ( n1768 & n9374 ) | ( n1768 & ~n27892 ) | ( n9374 & ~n27892 ) ;
  assign n27894 = ~n2606 & n2646 ;
  assign n27895 = ( n10954 & n11068 ) | ( n10954 & n27894 ) | ( n11068 & n27894 ) ;
  assign n27896 = ( n17619 & n27893 ) | ( n17619 & ~n27895 ) | ( n27893 & ~n27895 ) ;
  assign n27898 = n23437 ^ n11257 ^ n10788 ;
  assign n27897 = ( n1061 & ~n8295 ) | ( n1061 & n18292 ) | ( ~n8295 & n18292 ) ;
  assign n27899 = n27898 ^ n27897 ^ n1824 ;
  assign n27900 = n9307 ^ n4891 ^ n2740 ;
  assign n27901 = ( ~n3668 & n6403 ) | ( ~n3668 & n8509 ) | ( n6403 & n8509 ) ;
  assign n27902 = n27901 ^ n20960 ^ n277 ;
  assign n27903 = ( n4116 & n5792 ) | ( n4116 & n25255 ) | ( n5792 & n25255 ) ;
  assign n27904 = ~n19649 & n27903 ;
  assign n27905 = ~n26713 & n27904 ;
  assign n27906 = ( ~n18911 & n20289 ) | ( ~n18911 & n27905 ) | ( n20289 & n27905 ) ;
  assign n27907 = n27392 ^ n19504 ^ n7065 ;
  assign n27913 = ~n19542 & n21594 ;
  assign n27910 = n3083 & n15287 ;
  assign n27911 = n27910 ^ n1733 ^ 1'b0 ;
  assign n27912 = n27911 ^ n18736 ^ n597 ;
  assign n27908 = n17690 ^ n16278 ^ n5878 ;
  assign n27909 = ( n2924 & n25753 ) | ( n2924 & n27908 ) | ( n25753 & n27908 ) ;
  assign n27914 = n27913 ^ n27912 ^ n27909 ;
  assign n27915 = n27914 ^ n21272 ^ n20359 ;
  assign n27916 = ( ~n10077 & n27907 ) | ( ~n10077 & n27915 ) | ( n27907 & n27915 ) ;
  assign n27917 = n18170 ^ n11546 ^ 1'b0 ;
  assign n27918 = n8768 & ~n27917 ;
  assign n27919 = ( ~n12976 & n16448 ) | ( ~n12976 & n18147 ) | ( n16448 & n18147 ) ;
  assign n27920 = n5500 ^ n3502 ^ n1061 ;
  assign n27921 = n14612 ^ n10774 ^ n7148 ;
  assign n27922 = ( ~x55 & n8578 ) | ( ~x55 & n14000 ) | ( n8578 & n14000 ) ;
  assign n27923 = n27922 ^ n24155 ^ n23612 ;
  assign n27924 = n27923 ^ n21792 ^ n7961 ;
  assign n27925 = n26607 ^ n25149 ^ n15667 ;
  assign n27926 = n3092 & ~n12440 ;
  assign n27927 = n27926 ^ n26714 ^ 1'b0 ;
  assign n27928 = ~n3687 & n18556 ;
  assign n27929 = n27928 ^ n3300 ^ 1'b0 ;
  assign n27930 = ( n2624 & ~n7134 ) | ( n2624 & n21292 ) | ( ~n7134 & n21292 ) ;
  assign n27931 = n21067 ^ n18008 ^ n12024 ;
  assign n27932 = n17532 ^ n1759 ^ 1'b0 ;
  assign n27933 = n4488 & n27932 ;
  assign n27934 = ( ~n2176 & n4468 ) | ( ~n2176 & n27933 ) | ( n4468 & n27933 ) ;
  assign n27935 = ( n7539 & n19802 ) | ( n7539 & ~n27934 ) | ( n19802 & ~n27934 ) ;
  assign n27936 = n27442 ^ n16264 ^ n7680 ;
  assign n27937 = n26765 ^ n21798 ^ n17700 ;
  assign n27938 = n27937 ^ n3324 ^ n3086 ;
  assign n27941 = n611 & n17029 ;
  assign n27942 = ( ~n18593 & n22010 ) | ( ~n18593 & n27941 ) | ( n22010 & n27941 ) ;
  assign n27939 = n23106 ^ n22312 ^ n8229 ;
  assign n27940 = ( n3172 & n24992 ) | ( n3172 & ~n27939 ) | ( n24992 & ~n27939 ) ;
  assign n27943 = n27942 ^ n27940 ^ n8450 ;
  assign n27944 = n18813 ^ n10619 ^ n6961 ;
  assign n27945 = ( ~n3054 & n8606 ) | ( ~n3054 & n27944 ) | ( n8606 & n27944 ) ;
  assign n27946 = ( n8890 & n9239 ) | ( n8890 & ~n15776 ) | ( n9239 & ~n15776 ) ;
  assign n27948 = ( n11692 & ~n13472 ) | ( n11692 & n21787 ) | ( ~n13472 & n21787 ) ;
  assign n27947 = ( ~n1012 & n7800 ) | ( ~n1012 & n10403 ) | ( n7800 & n10403 ) ;
  assign n27949 = n27948 ^ n27947 ^ n7439 ;
  assign n27950 = n27949 ^ n27634 ^ n9222 ;
  assign n27952 = n15952 ^ n6034 ^ 1'b0 ;
  assign n27953 = ( n14818 & n19946 ) | ( n14818 & n27952 ) | ( n19946 & n27952 ) ;
  assign n27951 = ( n3531 & ~n15851 ) | ( n3531 & n22218 ) | ( ~n15851 & n22218 ) ;
  assign n27954 = n27953 ^ n27951 ^ n13895 ;
  assign n27955 = ( n5653 & ~n15667 ) | ( n5653 & n27954 ) | ( ~n15667 & n27954 ) ;
  assign n27956 = ( n4496 & n14604 ) | ( n4496 & n27955 ) | ( n14604 & n27955 ) ;
  assign n27957 = n22841 ^ n13983 ^ n604 ;
  assign n27958 = ( n756 & ~n11673 ) | ( n756 & n12624 ) | ( ~n11673 & n12624 ) ;
  assign n27959 = n25491 ^ n19643 ^ n16264 ;
  assign n27961 = ( n4062 & ~n6675 ) | ( n4062 & n18953 ) | ( ~n6675 & n18953 ) ;
  assign n27962 = n27961 ^ n19266 ^ n5828 ;
  assign n27960 = ~n6351 & n10328 ;
  assign n27963 = n27962 ^ n27960 ^ n7526 ;
  assign n27964 = ( n686 & n12386 ) | ( n686 & n12885 ) | ( n12386 & n12885 ) ;
  assign n27965 = n27964 ^ n10644 ^ 1'b0 ;
  assign n27966 = ( n6158 & n14682 ) | ( n6158 & ~n19428 ) | ( n14682 & ~n19428 ) ;
  assign n27967 = n27966 ^ n11412 ^ 1'b0 ;
  assign n27968 = n4036 & ~n10262 ;
  assign n27969 = n27968 ^ n13045 ^ 1'b0 ;
  assign n27970 = n24267 ^ n18935 ^ n5962 ;
  assign n27971 = ( n15584 & n27969 ) | ( n15584 & n27970 ) | ( n27969 & n27970 ) ;
  assign n27972 = ( ~n6395 & n6875 ) | ( ~n6395 & n14077 ) | ( n6875 & n14077 ) ;
  assign n27973 = ( n21844 & n23641 ) | ( n21844 & n27972 ) | ( n23641 & n27972 ) ;
  assign n27974 = n27973 ^ n26619 ^ n13629 ;
  assign n27975 = n17229 ^ n9173 ^ n8666 ;
  assign n27976 = n18612 ^ n18273 ^ n15494 ;
  assign n27977 = n27976 ^ n17227 ^ n5408 ;
  assign n27978 = ( n6031 & ~n7253 ) | ( n6031 & n9495 ) | ( ~n7253 & n9495 ) ;
  assign n27979 = n27978 ^ n12205 ^ n5135 ;
  assign n27980 = n27979 ^ n6288 ^ n4853 ;
  assign n27981 = n22010 ^ n20147 ^ n6357 ;
  assign n27982 = n7401 ^ n3025 ^ n2026 ;
  assign n27983 = ( n767 & n1845 ) | ( n767 & n3467 ) | ( n1845 & n3467 ) ;
  assign n27984 = n27983 ^ n17105 ^ n5136 ;
  assign n27985 = ( n19142 & n27982 ) | ( n19142 & n27984 ) | ( n27982 & n27984 ) ;
  assign n27986 = n27985 ^ n23529 ^ n152 ;
  assign n27987 = n18437 ^ n6211 ^ n5132 ;
  assign n27988 = n18499 ^ n17584 ^ n13966 ;
  assign n27989 = n1436 & n5000 ;
  assign n27990 = ~n11093 & n27989 ;
  assign n27991 = n17250 ^ n8354 ^ 1'b0 ;
  assign n27992 = n19816 ^ n14860 ^ 1'b0 ;
  assign n27993 = n14902 ^ n6453 ^ n2745 ;
  assign n27994 = ( n5957 & n10168 ) | ( n5957 & ~n18886 ) | ( n10168 & ~n18886 ) ;
  assign n27995 = n25246 ^ n14848 ^ n4571 ;
  assign n27996 = ( n2436 & n3120 ) | ( n2436 & n14048 ) | ( n3120 & n14048 ) ;
  assign n28000 = n9843 ^ n7571 ^ n3535 ;
  assign n27997 = n2527 | n5747 ;
  assign n27998 = n270 | n27997 ;
  assign n27999 = n27998 ^ n16333 ^ n8577 ;
  assign n28001 = n28000 ^ n27999 ^ n7796 ;
  assign n28002 = n7033 ^ n4479 ^ 1'b0 ;
  assign n28003 = ( n5645 & n21977 ) | ( n5645 & ~n28002 ) | ( n21977 & ~n28002 ) ;
  assign n28004 = n9674 ^ n4064 ^ n2570 ;
  assign n28005 = ( n9845 & ~n15358 ) | ( n9845 & n28004 ) | ( ~n15358 & n28004 ) ;
  assign n28006 = ( n3253 & n27203 ) | ( n3253 & ~n28005 ) | ( n27203 & ~n28005 ) ;
  assign n28007 = n20279 ^ n18173 ^ 1'b0 ;
  assign n28008 = ~n12027 & n28007 ;
  assign n28009 = ( n1730 & ~n8728 ) | ( n1730 & n10870 ) | ( ~n8728 & n10870 ) ;
  assign n28010 = ( n13656 & n21422 ) | ( n13656 & ~n23610 ) | ( n21422 & ~n23610 ) ;
  assign n28011 = n28010 ^ n5618 ^ n5070 ;
  assign n28012 = n21055 ^ n7785 ^ n717 ;
  assign n28013 = ( n6099 & n7504 ) | ( n6099 & n17511 ) | ( n7504 & n17511 ) ;
  assign n28014 = n25519 ^ n22245 ^ n3165 ;
  assign n28015 = n18224 ^ n3016 ^ n1936 ;
  assign n28016 = n9629 & n9954 ;
  assign n28017 = ( n4354 & ~n9294 ) | ( n4354 & n10644 ) | ( ~n9294 & n10644 ) ;
  assign n28018 = n28017 ^ n4571 ^ n1545 ;
  assign n28019 = ( n23481 & n28016 ) | ( n23481 & n28018 ) | ( n28016 & n28018 ) ;
  assign n28020 = n28019 ^ n23954 ^ n15209 ;
  assign n28021 = n1707 & ~n10375 ;
  assign n28022 = ~n20224 & n28021 ;
  assign n28023 = ( ~n8330 & n15726 ) | ( ~n8330 & n28022 ) | ( n15726 & n28022 ) ;
  assign n28024 = n4235 & n20676 ;
  assign n28025 = n28024 ^ n247 ^ 1'b0 ;
  assign n28026 = ( n2946 & ~n11992 ) | ( n2946 & n28025 ) | ( ~n11992 & n28025 ) ;
  assign n28027 = n28026 ^ n13397 ^ n3408 ;
  assign n28028 = ( n19162 & n28023 ) | ( n19162 & n28027 ) | ( n28023 & n28027 ) ;
  assign n28029 = n17869 ^ n12454 ^ 1'b0 ;
  assign n28030 = n11629 | n28029 ;
  assign n28031 = ( ~n6064 & n8015 ) | ( ~n6064 & n9416 ) | ( n8015 & n9416 ) ;
  assign n28032 = n28031 ^ n14765 ^ n10699 ;
  assign n28033 = n17535 & ~n20151 ;
  assign n28034 = n28032 & n28033 ;
  assign n28035 = n17271 ^ n16934 ^ 1'b0 ;
  assign n28036 = ( n3715 & n12722 ) | ( n3715 & n27878 ) | ( n12722 & n27878 ) ;
  assign n28037 = n18898 ^ n4420 ^ 1'b0 ;
  assign n28038 = ( ~n2560 & n3072 ) | ( ~n2560 & n21095 ) | ( n3072 & n21095 ) ;
  assign n28039 = ( n3383 & ~n15598 ) | ( n3383 & n28038 ) | ( ~n15598 & n28038 ) ;
  assign n28040 = ( ~n2044 & n9698 ) | ( ~n2044 & n14222 ) | ( n9698 & n14222 ) ;
  assign n28041 = n18576 ^ n10769 ^ n954 ;
  assign n28042 = n28041 ^ n21594 ^ n1593 ;
  assign n28043 = ( n2330 & ~n23097 ) | ( n2330 & n28042 ) | ( ~n23097 & n28042 ) ;
  assign n28044 = ( n7731 & n14792 ) | ( n7731 & n14901 ) | ( n14792 & n14901 ) ;
  assign n28045 = ( n3327 & n10753 ) | ( n3327 & n23738 ) | ( n10753 & n23738 ) ;
  assign n28048 = n10131 ^ n6764 ^ 1'b0 ;
  assign n28049 = n2669 & n28048 ;
  assign n28050 = n28049 ^ n25713 ^ n7468 ;
  assign n28046 = ( n2263 & ~n6874 ) | ( n2263 & n18802 ) | ( ~n6874 & n18802 ) ;
  assign n28047 = ( n5116 & n14193 ) | ( n5116 & ~n28046 ) | ( n14193 & ~n28046 ) ;
  assign n28051 = n28050 ^ n28047 ^ 1'b0 ;
  assign n28052 = n10783 | n28051 ;
  assign n28053 = ( ~n27324 & n28045 ) | ( ~n27324 & n28052 ) | ( n28045 & n28052 ) ;
  assign n28054 = ( ~n27669 & n28044 ) | ( ~n27669 & n28053 ) | ( n28044 & n28053 ) ;
  assign n28055 = n25799 ^ n17453 ^ n4650 ;
  assign n28056 = ( n7393 & n11610 ) | ( n7393 & n11910 ) | ( n11610 & n11910 ) ;
  assign n28057 = n28056 ^ n3366 ^ 1'b0 ;
  assign n28058 = n1693 & ~n28057 ;
  assign n28059 = n6558 ^ n4747 ^ n3389 ;
  assign n28060 = ( n11679 & n24721 ) | ( n11679 & n28059 ) | ( n24721 & n28059 ) ;
  assign n28061 = ( n7890 & n8387 ) | ( n7890 & ~n9870 ) | ( n8387 & ~n9870 ) ;
  assign n28062 = n12747 ^ n3729 ^ 1'b0 ;
  assign n28063 = n28062 ^ n22667 ^ n4006 ;
  assign n28064 = ( n4285 & n28061 ) | ( n4285 & ~n28063 ) | ( n28061 & ~n28063 ) ;
  assign n28065 = n14412 ^ n13552 ^ 1'b0 ;
  assign n28070 = ( n2932 & n8872 ) | ( n2932 & ~n9360 ) | ( n8872 & ~n9360 ) ;
  assign n28066 = n3617 & ~n16355 ;
  assign n28067 = n10841 & n28066 ;
  assign n28068 = ( n1701 & n10964 ) | ( n1701 & ~n22952 ) | ( n10964 & ~n22952 ) ;
  assign n28069 = ( n20317 & n28067 ) | ( n20317 & n28068 ) | ( n28067 & n28068 ) ;
  assign n28071 = n28070 ^ n28069 ^ n22931 ;
  assign n28072 = n19426 ^ n4444 ^ n1889 ;
  assign n28073 = ( ~n1650 & n19417 ) | ( ~n1650 & n28072 ) | ( n19417 & n28072 ) ;
  assign n28074 = ( n9206 & n22611 ) | ( n9206 & ~n27483 ) | ( n22611 & ~n27483 ) ;
  assign n28075 = n326 | n16393 ;
  assign n28076 = n28074 & ~n28075 ;
  assign n28077 = n28076 ^ n11343 ^ n1600 ;
  assign n28078 = ( n3656 & n13792 ) | ( n3656 & ~n18632 ) | ( n13792 & ~n18632 ) ;
  assign n28079 = n14121 ^ n11720 ^ 1'b0 ;
  assign n28080 = ( ~n9994 & n27176 ) | ( ~n9994 & n28079 ) | ( n27176 & n28079 ) ;
  assign n28083 = ( ~n2147 & n3091 ) | ( ~n2147 & n18725 ) | ( n3091 & n18725 ) ;
  assign n28084 = n28083 ^ n18457 ^ n12147 ;
  assign n28081 = n19624 ^ n5599 ^ 1'b0 ;
  assign n28082 = n8948 & ~n28081 ;
  assign n28085 = n28084 ^ n28082 ^ n792 ;
  assign n28086 = n17289 ^ n11897 ^ n5692 ;
  assign n28087 = ( n2369 & n8438 ) | ( n2369 & n10861 ) | ( n8438 & n10861 ) ;
  assign n28088 = ( n1995 & n2054 ) | ( n1995 & n6931 ) | ( n2054 & n6931 ) ;
  assign n28089 = n28088 ^ n9495 ^ n3441 ;
  assign n28090 = n20675 ^ n15272 ^ n10223 ;
  assign n28092 = ( ~n3731 & n11374 ) | ( ~n3731 & n15424 ) | ( n11374 & n15424 ) ;
  assign n28091 = ( ~n157 & n424 ) | ( ~n157 & n8212 ) | ( n424 & n8212 ) ;
  assign n28093 = n28092 ^ n28091 ^ 1'b0 ;
  assign n28094 = ( ~n460 & n7920 ) | ( ~n460 & n9070 ) | ( n7920 & n9070 ) ;
  assign n28095 = n28094 ^ n6631 ^ n2141 ;
  assign n28096 = n28095 ^ n4933 ^ n1902 ;
  assign n28097 = n28096 ^ n6386 ^ n5381 ;
  assign n28098 = n21476 ^ n9283 ^ n464 ;
  assign n28099 = n9145 ^ n3438 ^ 1'b0 ;
  assign n28100 = n9555 & ~n28099 ;
  assign n28101 = n28100 ^ n26441 ^ 1'b0 ;
  assign n28102 = n4219 & n23530 ;
  assign n28103 = n24332 & n28102 ;
  assign n28104 = n3529 ^ n2534 ^ 1'b0 ;
  assign n28105 = n11271 | n28104 ;
  assign n28106 = n16002 ^ n10065 ^ x107 ;
  assign n28107 = n19027 & n28106 ;
  assign n28108 = ( n10573 & ~n19460 ) | ( n10573 & n28107 ) | ( ~n19460 & n28107 ) ;
  assign n28109 = n21472 ^ n13591 ^ n738 ;
  assign n28110 = ( n5701 & n12524 ) | ( n5701 & ~n27243 ) | ( n12524 & ~n27243 ) ;
  assign n28111 = ( n6923 & ~n18953 ) | ( n6923 & n23197 ) | ( ~n18953 & n23197 ) ;
  assign n28112 = ( n7594 & n15964 ) | ( n7594 & ~n28111 ) | ( n15964 & ~n28111 ) ;
  assign n28113 = n26128 ^ n25124 ^ n8015 ;
  assign n28116 = ~n2215 & n4436 ;
  assign n28117 = n28116 ^ n1499 ^ 1'b0 ;
  assign n28118 = ( n3332 & n7850 ) | ( n3332 & n28117 ) | ( n7850 & n28117 ) ;
  assign n28114 = n14378 ^ n3208 ^ 1'b0 ;
  assign n28115 = n28114 ^ n23589 ^ n3390 ;
  assign n28119 = n28118 ^ n28115 ^ n24289 ;
  assign n28120 = ( n14118 & ~n16288 ) | ( n14118 & n28096 ) | ( ~n16288 & n28096 ) ;
  assign n28121 = n4501 ^ n4046 ^ n995 ;
  assign n28122 = ( ~n1881 & n6312 ) | ( ~n1881 & n8380 ) | ( n6312 & n8380 ) ;
  assign n28123 = ( n6230 & ~n28121 ) | ( n6230 & n28122 ) | ( ~n28121 & n28122 ) ;
  assign n28124 = n28123 ^ n23288 ^ n18539 ;
  assign n28125 = n20483 ^ n16874 ^ 1'b0 ;
  assign n28126 = n10392 | n28125 ;
  assign n28127 = ~n5161 & n15755 ;
  assign n28128 = n28127 ^ n10947 ^ 1'b0 ;
  assign n28129 = n22499 & n28128 ;
  assign n28130 = ( n354 & n2937 ) | ( n354 & n9951 ) | ( n2937 & n9951 ) ;
  assign n28131 = ( n6410 & ~n7137 ) | ( n6410 & n8953 ) | ( ~n7137 & n8953 ) ;
  assign n28132 = n16530 ^ n14655 ^ n1632 ;
  assign n28133 = ( n28130 & n28131 ) | ( n28130 & ~n28132 ) | ( n28131 & ~n28132 ) ;
  assign n28134 = ( n4319 & ~n6561 ) | ( n4319 & n10971 ) | ( ~n6561 & n10971 ) ;
  assign n28135 = n28134 ^ n24701 ^ n4924 ;
  assign n28136 = ( ~n5971 & n14853 ) | ( ~n5971 & n27134 ) | ( n14853 & n27134 ) ;
  assign n28137 = ( n12337 & n28135 ) | ( n12337 & ~n28136 ) | ( n28135 & ~n28136 ) ;
  assign n28138 = n28137 ^ n23908 ^ 1'b0 ;
  assign n28139 = n3802 | n22096 ;
  assign n28140 = n21491 ^ n14383 ^ n11810 ;
  assign n28141 = ( n10704 & n20657 ) | ( n10704 & n28140 ) | ( n20657 & n28140 ) ;
  assign n28142 = n28141 ^ n15069 ^ n10968 ;
  assign n28143 = n4884 | n21505 ;
  assign n28144 = ( n216 & n14013 ) | ( n216 & ~n24203 ) | ( n14013 & ~n24203 ) ;
  assign n28145 = n5337 ^ n3765 ^ n491 ;
  assign n28146 = n28145 ^ n9484 ^ n670 ;
  assign n28147 = ( ~n3373 & n14378 ) | ( ~n3373 & n26146 ) | ( n14378 & n26146 ) ;
  assign n28148 = n16734 ^ n8129 ^ n7919 ;
  assign n28149 = n9889 & n25429 ;
  assign n28150 = n20156 ^ n16315 ^ 1'b0 ;
  assign n28151 = n27933 & ~n28150 ;
  assign n28152 = n26567 & ~n28151 ;
  assign n28153 = n28152 ^ n26110 ^ n18736 ;
  assign n28154 = n24444 ^ n19174 ^ n7926 ;
  assign n28155 = ( ~n19139 & n26606 ) | ( ~n19139 & n28154 ) | ( n26606 & n28154 ) ;
  assign n28156 = n19315 ^ n18316 ^ n1291 ;
  assign n28158 = ( ~n7334 & n18638 ) | ( ~n7334 & n22382 ) | ( n18638 & n22382 ) ;
  assign n28159 = ( n4100 & ~n4637 ) | ( n4100 & n28158 ) | ( ~n4637 & n28158 ) ;
  assign n28157 = ( ~n9558 & n14760 ) | ( ~n9558 & n18745 ) | ( n14760 & n18745 ) ;
  assign n28160 = n28159 ^ n28157 ^ n12486 ;
  assign n28161 = ( n13299 & ~n18650 ) | ( n13299 & n22960 ) | ( ~n18650 & n22960 ) ;
  assign n28162 = n14716 ^ n6493 ^ n582 ;
  assign n28163 = n5930 ^ n3222 ^ n499 ;
  assign n28164 = n5903 & ~n22626 ;
  assign n28165 = n23675 | n28164 ;
  assign n28166 = ( n28162 & n28163 ) | ( n28162 & n28165 ) | ( n28163 & n28165 ) ;
  assign n28167 = ( n1472 & n13169 ) | ( n1472 & ~n13778 ) | ( n13169 & ~n13778 ) ;
  assign n28168 = n11414 & ~n28167 ;
  assign n28169 = ~n3710 & n28168 ;
  assign n28170 = ~n1888 & n27638 ;
  assign n28171 = n1352 & n28170 ;
  assign n28172 = n10884 & ~n13658 ;
  assign n28173 = ( n783 & n14818 ) | ( n783 & n18439 ) | ( n14818 & n18439 ) ;
  assign n28174 = n20492 ^ n15370 ^ n1745 ;
  assign n28175 = n8286 & n11696 ;
  assign n28176 = n28175 ^ n23754 ^ n936 ;
  assign n28177 = ( n9577 & n28174 ) | ( n9577 & ~n28176 ) | ( n28174 & ~n28176 ) ;
  assign n28178 = ( ~n26071 & n28173 ) | ( ~n26071 & n28177 ) | ( n28173 & n28177 ) ;
  assign n28179 = n17090 ^ n15541 ^ n14844 ;
  assign n28180 = ( ~n5052 & n5195 ) | ( ~n5052 & n19162 ) | ( n5195 & n19162 ) ;
  assign n28181 = ( n13827 & n22126 ) | ( n13827 & n28180 ) | ( n22126 & n28180 ) ;
  assign n28182 = ( n6889 & n10785 ) | ( n6889 & n27183 ) | ( n10785 & n27183 ) ;
  assign n28183 = ( ~n2274 & n3333 ) | ( ~n2274 & n9335 ) | ( n3333 & n9335 ) ;
  assign n28184 = n16500 ^ n3503 ^ n2019 ;
  assign n28185 = n24228 ^ n15655 ^ n13915 ;
  assign n28186 = ( n28183 & n28184 ) | ( n28183 & n28185 ) | ( n28184 & n28185 ) ;
  assign n28187 = n13062 ^ n9432 ^ 1'b0 ;
  assign n28188 = ~n15128 & n28187 ;
  assign n28189 = ( ~n6519 & n11335 ) | ( ~n6519 & n11699 ) | ( n11335 & n11699 ) ;
  assign n28191 = n8091 ^ n7623 ^ n7370 ;
  assign n28192 = ( n5112 & n11735 ) | ( n5112 & ~n28191 ) | ( n11735 & ~n28191 ) ;
  assign n28190 = n10814 ^ n10752 ^ n4527 ;
  assign n28193 = n28192 ^ n28190 ^ 1'b0 ;
  assign n28194 = n28189 & ~n28193 ;
  assign n28195 = n12459 ^ n8072 ^ n906 ;
  assign n28196 = n28195 ^ n12986 ^ n676 ;
  assign n28197 = n28196 ^ n11193 ^ n3824 ;
  assign n28198 = ( ~n4633 & n28194 ) | ( ~n4633 & n28197 ) | ( n28194 & n28197 ) ;
  assign n28199 = n28198 ^ n27915 ^ 1'b0 ;
  assign n28200 = n14061 & ~n28199 ;
  assign n28201 = n7545 & ~n23909 ;
  assign n28202 = n28201 ^ n11199 ^ 1'b0 ;
  assign n28203 = n2735 & ~n28202 ;
  assign n28204 = ( ~n6890 & n12327 ) | ( ~n6890 & n27346 ) | ( n12327 & n27346 ) ;
  assign n28207 = ( ~n454 & n1663 ) | ( ~n454 & n10039 ) | ( n1663 & n10039 ) ;
  assign n28205 = ~n17988 & n20647 ;
  assign n28206 = ( n1792 & n22136 ) | ( n1792 & n28205 ) | ( n22136 & n28205 ) ;
  assign n28208 = n28207 ^ n28206 ^ n9679 ;
  assign n28209 = n10686 & ~n27113 ;
  assign n28210 = n28209 ^ n16582 ^ n12314 ;
  assign n28211 = ( n134 & n21978 ) | ( n134 & ~n24455 ) | ( n21978 & ~n24455 ) ;
  assign n28212 = ( ~n6673 & n11631 ) | ( ~n6673 & n19944 ) | ( n11631 & n19944 ) ;
  assign n28214 = ~n15742 & n16342 ;
  assign n28215 = n28214 ^ n12154 ^ 1'b0 ;
  assign n28213 = ~n2658 & n9431 ;
  assign n28216 = n28215 ^ n28213 ^ 1'b0 ;
  assign n28217 = ( n8851 & n10121 ) | ( n8851 & n28216 ) | ( n10121 & n28216 ) ;
  assign n28218 = n28217 ^ n11731 ^ n2393 ;
  assign n28219 = n3914 | n13860 ;
  assign n28220 = ( n10586 & ~n14103 ) | ( n10586 & n28219 ) | ( ~n14103 & n28219 ) ;
  assign n28221 = n28220 ^ n13574 ^ n10344 ;
  assign n28222 = n10039 & n10049 ;
  assign n28223 = n28222 ^ n22233 ^ 1'b0 ;
  assign n28224 = n22283 ^ n12213 ^ n10406 ;
  assign n28225 = ( ~n4558 & n19371 ) | ( ~n4558 & n28224 ) | ( n19371 & n28224 ) ;
  assign n28226 = ( n1635 & n6789 ) | ( n1635 & n28225 ) | ( n6789 & n28225 ) ;
  assign n28230 = n7815 ^ n2360 ^ n503 ;
  assign n28229 = n14313 ^ n11571 ^ n401 ;
  assign n28227 = ( ~n1673 & n7660 ) | ( ~n1673 & n25426 ) | ( n7660 & n25426 ) ;
  assign n28228 = n28227 ^ n7560 ^ n5614 ;
  assign n28231 = n28230 ^ n28229 ^ n28228 ;
  assign n28232 = n20289 ^ n16049 ^ n12024 ;
  assign n28233 = ( n3721 & n20663 ) | ( n3721 & ~n28232 ) | ( n20663 & ~n28232 ) ;
  assign n28234 = n15283 & ~n28233 ;
  assign n28235 = ~n17440 & n21343 ;
  assign n28236 = ( ~n14227 & n26880 ) | ( ~n14227 & n28235 ) | ( n26880 & n28235 ) ;
  assign n28237 = n24752 ^ n18775 ^ n10443 ;
  assign n28238 = ( n8221 & n9356 ) | ( n8221 & n10148 ) | ( n9356 & n10148 ) ;
  assign n28239 = n28238 ^ n4898 ^ n3170 ;
  assign n28240 = ~n133 & n28239 ;
  assign n28241 = n28240 ^ n18201 ^ 1'b0 ;
  assign n28242 = ( n1048 & n10315 ) | ( n1048 & n28241 ) | ( n10315 & n28241 ) ;
  assign n28243 = n20518 ^ n8029 ^ n7408 ;
  assign n28244 = n28243 ^ n17890 ^ n8694 ;
  assign n28245 = ( n569 & n10934 ) | ( n569 & ~n28244 ) | ( n10934 & ~n28244 ) ;
  assign n28246 = n28245 ^ n18339 ^ 1'b0 ;
  assign n28247 = n27675 ^ n19809 ^ n10510 ;
  assign n28248 = ( ~n13461 & n18260 ) | ( ~n13461 & n27095 ) | ( n18260 & n27095 ) ;
  assign n28249 = ( n9551 & n28247 ) | ( n9551 & ~n28248 ) | ( n28247 & ~n28248 ) ;
  assign n28250 = ( n1752 & ~n3942 ) | ( n1752 & n7243 ) | ( ~n3942 & n7243 ) ;
  assign n28251 = ( n14837 & ~n24070 ) | ( n14837 & n28250 ) | ( ~n24070 & n28250 ) ;
  assign n28252 = n18014 & ~n28251 ;
  assign n28253 = n3203 & ~n7642 ;
  assign n28254 = n28253 ^ n4321 ^ 1'b0 ;
  assign n28255 = n11931 ^ n9610 ^ n8083 ;
  assign n28256 = ( ~n969 & n20732 ) | ( ~n969 & n28255 ) | ( n20732 & n28255 ) ;
  assign n28257 = ( n6222 & n28254 ) | ( n6222 & n28256 ) | ( n28254 & n28256 ) ;
  assign n28258 = ( n8331 & ~n9334 ) | ( n8331 & n28257 ) | ( ~n9334 & n28257 ) ;
  assign n28259 = n25863 ^ n10196 ^ n5174 ;
  assign n28260 = ( n3307 & ~n3452 ) | ( n3307 & n6051 ) | ( ~n3452 & n6051 ) ;
  assign n28261 = ( n1535 & n8933 ) | ( n1535 & n12036 ) | ( n8933 & n12036 ) ;
  assign n28262 = ( ~n4614 & n12348 ) | ( ~n4614 & n28261 ) | ( n12348 & n28261 ) ;
  assign n28266 = ( ~n6979 & n13274 ) | ( ~n6979 & n22755 ) | ( n13274 & n22755 ) ;
  assign n28264 = n3530 ^ n1961 ^ 1'b0 ;
  assign n28265 = ( n9637 & n14207 ) | ( n9637 & n28264 ) | ( n14207 & n28264 ) ;
  assign n28263 = ( n6407 & n15881 ) | ( n6407 & n17291 ) | ( n15881 & n17291 ) ;
  assign n28267 = n28266 ^ n28265 ^ n28263 ;
  assign n28268 = ( n10481 & n16921 ) | ( n10481 & ~n27947 ) | ( n16921 & ~n27947 ) ;
  assign n28269 = n5400 & n10613 ;
  assign n28270 = n28269 ^ n20953 ^ 1'b0 ;
  assign n28273 = ( n5448 & n5780 ) | ( n5448 & ~n12120 ) | ( n5780 & ~n12120 ) ;
  assign n28271 = n19056 ^ n3468 ^ n888 ;
  assign n28272 = n28271 ^ n20946 ^ n12763 ;
  assign n28274 = n28273 ^ n28272 ^ n16650 ;
  assign n28276 = n24634 ^ n19244 ^ 1'b0 ;
  assign n28275 = n21297 ^ n18801 ^ n11893 ;
  assign n28277 = n28276 ^ n28275 ^ 1'b0 ;
  assign n28281 = n9534 ^ n7826 ^ n7216 ;
  assign n28282 = ( n3255 & n22258 ) | ( n3255 & n28281 ) | ( n22258 & n28281 ) ;
  assign n28278 = n12950 ^ n8081 ^ n930 ;
  assign n28279 = n28278 ^ n380 ^ x40 ;
  assign n28280 = ( n12113 & n12305 ) | ( n12113 & ~n28279 ) | ( n12305 & ~n28279 ) ;
  assign n28283 = n28282 ^ n28280 ^ n7476 ;
  assign n28284 = ( ~n7818 & n15474 ) | ( ~n7818 & n19577 ) | ( n15474 & n19577 ) ;
  assign n28285 = n28284 ^ n15557 ^ n12686 ;
  assign n28286 = ( ~n2386 & n6220 ) | ( ~n2386 & n11688 ) | ( n6220 & n11688 ) ;
  assign n28287 = n28286 ^ n8115 ^ n1422 ;
  assign n28288 = ( n8076 & n12524 ) | ( n8076 & n16068 ) | ( n12524 & n16068 ) ;
  assign n28289 = n28288 ^ n8540 ^ n373 ;
  assign n28290 = ( n3357 & n20877 ) | ( n3357 & ~n28289 ) | ( n20877 & ~n28289 ) ;
  assign n28291 = ( n15614 & n28287 ) | ( n15614 & ~n28290 ) | ( n28287 & ~n28290 ) ;
  assign n28292 = n3587 ^ n3085 ^ 1'b0 ;
  assign n28293 = ~n3897 & n28292 ;
  assign n28294 = ( n1823 & n9300 ) | ( n1823 & ~n28293 ) | ( n9300 & ~n28293 ) ;
  assign n28295 = ( ~n18304 & n18500 ) | ( ~n18304 & n20532 ) | ( n18500 & n20532 ) ;
  assign n28296 = ( ~n6338 & n21341 ) | ( ~n6338 & n28295 ) | ( n21341 & n28295 ) ;
  assign n28297 = n7905 ^ n2109 ^ x93 ;
  assign n28298 = n3936 | n18933 ;
  assign n28299 = ( ~n14657 & n16353 ) | ( ~n14657 & n17245 ) | ( n16353 & n17245 ) ;
  assign n28300 = ( n5063 & ~n10134 ) | ( n5063 & n20821 ) | ( ~n10134 & n20821 ) ;
  assign n28304 = n27964 ^ n9960 ^ 1'b0 ;
  assign n28305 = ~n4886 & n28304 ;
  assign n28306 = ( n14564 & n15812 ) | ( n14564 & ~n28305 ) | ( n15812 & ~n28305 ) ;
  assign n28301 = ~n3194 & n6284 ;
  assign n28302 = ~n3786 & n28301 ;
  assign n28303 = n28302 ^ n610 ^ 1'b0 ;
  assign n28307 = n28306 ^ n28303 ^ n15087 ;
  assign n28308 = ( n2752 & n9349 ) | ( n2752 & n17992 ) | ( n9349 & n17992 ) ;
  assign n28309 = n4993 & ~n28308 ;
  assign n28310 = n15862 ^ n7932 ^ n731 ;
  assign n28311 = ( n12311 & n14304 ) | ( n12311 & ~n14976 ) | ( n14304 & ~n14976 ) ;
  assign n28312 = n12739 ^ n8271 ^ n8225 ;
  assign n28313 = n28312 ^ n14030 ^ n1072 ;
  assign n28315 = n19798 ^ n11839 ^ n5327 ;
  assign n28314 = n25683 ^ n17130 ^ n3829 ;
  assign n28316 = n28315 ^ n28314 ^ n3480 ;
  assign n28317 = n7535 & n9366 ;
  assign n28319 = ( ~n1246 & n3573 ) | ( ~n1246 & n27278 ) | ( n3573 & n27278 ) ;
  assign n28320 = n23882 & n28319 ;
  assign n28318 = n17227 & n26749 ;
  assign n28321 = n28320 ^ n28318 ^ 1'b0 ;
  assign n28322 = n10717 ^ n7777 ^ n3853 ;
  assign n28323 = ( n2820 & n22415 ) | ( n2820 & ~n28322 ) | ( n22415 & ~n28322 ) ;
  assign n28324 = n28323 ^ n25425 ^ n7592 ;
  assign n28325 = n15704 & ~n25493 ;
  assign n28326 = n28325 ^ n14168 ^ 1'b0 ;
  assign n28327 = ( n1594 & n8585 ) | ( n1594 & n28326 ) | ( n8585 & n28326 ) ;
  assign n28328 = n4448 & ~n7698 ;
  assign n28329 = ( n884 & ~n2600 ) | ( n884 & n27292 ) | ( ~n2600 & n27292 ) ;
  assign n28330 = ( n2557 & n10225 ) | ( n2557 & ~n28329 ) | ( n10225 & ~n28329 ) ;
  assign n28331 = n14966 ^ n9062 ^ n4550 ;
  assign n28332 = ( n3567 & ~n4785 ) | ( n3567 & n28331 ) | ( ~n4785 & n28331 ) ;
  assign n28333 = ( n4543 & ~n6286 ) | ( n4543 & n23613 ) | ( ~n6286 & n23613 ) ;
  assign n28334 = n670 | n11391 ;
  assign n28335 = n11148 | n28334 ;
  assign n28336 = n17946 ^ n14054 ^ 1'b0 ;
  assign n28337 = n28335 & n28336 ;
  assign n28338 = ( n14174 & n14646 ) | ( n14174 & ~n27327 ) | ( n14646 & ~n27327 ) ;
  assign n28339 = n12872 | n22694 ;
  assign n28340 = n18667 ^ n10393 ^ n7912 ;
  assign n28341 = ( n1727 & n11377 ) | ( n1727 & ~n19221 ) | ( n11377 & ~n19221 ) ;
  assign n28342 = ( n3813 & ~n5783 ) | ( n3813 & n16224 ) | ( ~n5783 & n16224 ) ;
  assign n28343 = ( ~n6468 & n28341 ) | ( ~n6468 & n28342 ) | ( n28341 & n28342 ) ;
  assign n28344 = ( n4733 & n6581 ) | ( n4733 & n28343 ) | ( n6581 & n28343 ) ;
  assign n28347 = ( n1711 & ~n5002 ) | ( n1711 & n7366 ) | ( ~n5002 & n7366 ) ;
  assign n28345 = n14708 ^ n6812 ^ n1036 ;
  assign n28346 = n28345 ^ n14790 ^ n3731 ;
  assign n28348 = n28347 ^ n28346 ^ n16361 ;
  assign n28349 = n15551 ^ n6486 ^ n1219 ;
  assign n28350 = ( n4201 & n17061 ) | ( n4201 & n28349 ) | ( n17061 & n28349 ) ;
  assign n28351 = n8285 & ~n14253 ;
  assign n28352 = n28351 ^ n15307 ^ 1'b0 ;
  assign n28353 = n3154 | n26354 ;
  assign n28354 = n28353 ^ n6915 ^ 1'b0 ;
  assign n28355 = ( ~n20281 & n28352 ) | ( ~n20281 & n28354 ) | ( n28352 & n28354 ) ;
  assign n28356 = n3994 | n27581 ;
  assign n28357 = ( n3550 & n10194 ) | ( n3550 & n13683 ) | ( n10194 & n13683 ) ;
  assign n28358 = n8540 & ~n28357 ;
  assign n28359 = n24518 ^ n5566 ^ n4562 ;
  assign n28360 = n28359 ^ n7394 ^ 1'b0 ;
  assign n28361 = n28358 & n28360 ;
  assign n28362 = n9647 ^ n6965 ^ n6405 ;
  assign n28363 = n5457 & n28362 ;
  assign n28364 = ~n27083 & n28363 ;
  assign n28369 = n15336 ^ n8221 ^ n1754 ;
  assign n28365 = n8363 & n23129 ;
  assign n28366 = n28365 ^ n12932 ^ 1'b0 ;
  assign n28367 = n28366 ^ n15103 ^ n5164 ;
  assign n28368 = n28367 ^ n7660 ^ n2562 ;
  assign n28370 = n28369 ^ n28368 ^ n9456 ;
  assign n28371 = ( n6863 & n13217 ) | ( n6863 & n13460 ) | ( n13217 & n13460 ) ;
  assign n28372 = n28371 ^ n23249 ^ n7318 ;
  assign n28374 = ( n5144 & ~n11896 ) | ( n5144 & n12247 ) | ( ~n11896 & n12247 ) ;
  assign n28373 = ( n4379 & ~n23248 ) | ( n4379 & n23533 ) | ( ~n23248 & n23533 ) ;
  assign n28375 = n28374 ^ n28373 ^ n2589 ;
  assign n28381 = n12066 ^ n1863 ^ 1'b0 ;
  assign n28379 = n15119 ^ n13885 ^ n12706 ;
  assign n28376 = n12436 & ~n15630 ;
  assign n28377 = ~n5541 & n28376 ;
  assign n28378 = n28377 ^ n18074 ^ n13748 ;
  assign n28380 = n28379 ^ n28378 ^ n1901 ;
  assign n28382 = n28381 ^ n28380 ^ n24513 ;
  assign n28383 = n27023 ^ n26438 ^ n22939 ;
  assign n28384 = ( n6402 & n20216 ) | ( n6402 & ~n25388 ) | ( n20216 & ~n25388 ) ;
  assign n28385 = n965 & n1669 ;
  assign n28386 = ~n25138 & n28385 ;
  assign n28387 = ( ~n2196 & n9646 ) | ( ~n2196 & n20723 ) | ( n9646 & n20723 ) ;
  assign n28388 = n25777 ^ n20888 ^ n19692 ;
  assign n28389 = ( n3519 & n5150 ) | ( n3519 & ~n12835 ) | ( n5150 & ~n12835 ) ;
  assign n28390 = ~n7105 & n7762 ;
  assign n28391 = ~n4371 & n28390 ;
  assign n28392 = ( n18604 & n27420 ) | ( n18604 & ~n28391 ) | ( n27420 & ~n28391 ) ;
  assign n28393 = n7985 & n15831 ;
  assign n28394 = n28393 ^ n10249 ^ 1'b0 ;
  assign n28395 = n8412 | n27146 ;
  assign n28397 = n8663 ^ n6136 ^ 1'b0 ;
  assign n28396 = ( n5570 & n16142 ) | ( n5570 & ~n28235 ) | ( n16142 & ~n28235 ) ;
  assign n28398 = n28397 ^ n28396 ^ n18066 ;
  assign n28399 = n20431 ^ n1757 ^ n1568 ;
  assign n28400 = n28399 ^ n16824 ^ n13185 ;
  assign n28401 = ( n1634 & n4570 ) | ( n1634 & n5361 ) | ( n4570 & n5361 ) ;
  assign n28402 = n28401 ^ n23592 ^ n19990 ;
  assign n28403 = n5505 & n17709 ;
  assign n28404 = n5164 ^ n2826 ^ 1'b0 ;
  assign n28405 = ( n15905 & n18781 ) | ( n15905 & n28404 ) | ( n18781 & n28404 ) ;
  assign n28406 = n22394 ^ n6694 ^ n4151 ;
  assign n28407 = ( ~n3294 & n28405 ) | ( ~n3294 & n28406 ) | ( n28405 & n28406 ) ;
  assign n28408 = n28407 ^ n18921 ^ n513 ;
  assign n28409 = n7577 ^ n6887 ^ n2565 ;
  assign n28410 = ( n524 & n2747 ) | ( n524 & ~n28409 ) | ( n2747 & ~n28409 ) ;
  assign n28411 = n5067 & n8531 ;
  assign n28412 = n25937 & n28411 ;
  assign n28413 = ( n1612 & n4975 ) | ( n1612 & ~n12488 ) | ( n4975 & ~n12488 ) ;
  assign n28414 = ( n11466 & n20147 ) | ( n11466 & n28413 ) | ( n20147 & n28413 ) ;
  assign n28415 = n11611 ^ n10699 ^ n8778 ;
  assign n28416 = ( ~n3630 & n26086 ) | ( ~n3630 & n28415 ) | ( n26086 & n28415 ) ;
  assign n28417 = n28416 ^ n13139 ^ n2008 ;
  assign n28418 = n19896 ^ n16312 ^ 1'b0 ;
  assign n28419 = n4804 & ~n28418 ;
  assign n28420 = ( ~n19876 & n28417 ) | ( ~n19876 & n28419 ) | ( n28417 & n28419 ) ;
  assign n28421 = ( n579 & ~n2347 ) | ( n579 & n4566 ) | ( ~n2347 & n4566 ) ;
  assign n28422 = n28421 ^ n12076 ^ n10051 ;
  assign n28423 = ( ~n14755 & n20105 ) | ( ~n14755 & n21426 ) | ( n20105 & n21426 ) ;
  assign n28424 = n17652 ^ n2479 ^ n718 ;
  assign n28428 = ( n6436 & n8279 ) | ( n6436 & ~n14964 ) | ( n8279 & ~n14964 ) ;
  assign n28425 = ( n2917 & ~n3268 ) | ( n2917 & n3337 ) | ( ~n3268 & n3337 ) ;
  assign n28426 = n28425 ^ n1824 ^ n160 ;
  assign n28427 = n1573 | n28426 ;
  assign n28429 = n28428 ^ n28427 ^ 1'b0 ;
  assign n28430 = n28429 ^ n22263 ^ n14028 ;
  assign n28431 = ( n1397 & n24342 ) | ( n1397 & ~n28430 ) | ( n24342 & ~n28430 ) ;
  assign n28432 = n22100 ^ n4696 ^ 1'b0 ;
  assign n28433 = ( ~n4841 & n18766 ) | ( ~n4841 & n28432 ) | ( n18766 & n28432 ) ;
  assign n28434 = ( n3817 & ~n13384 ) | ( n3817 & n21158 ) | ( ~n13384 & n21158 ) ;
  assign n28435 = ( n5880 & n11399 ) | ( n5880 & n19683 ) | ( n11399 & n19683 ) ;
  assign n28436 = n10482 ^ n6317 ^ n3635 ;
  assign n28437 = n28436 ^ n21806 ^ n6883 ;
  assign n28438 = ( n5216 & n28435 ) | ( n5216 & ~n28437 ) | ( n28435 & ~n28437 ) ;
  assign n28439 = n15414 ^ n11735 ^ n7262 ;
  assign n28440 = ( n7596 & n16805 ) | ( n7596 & n28439 ) | ( n16805 & n28439 ) ;
  assign n28441 = ( ~n6465 & n12120 ) | ( ~n6465 & n22364 ) | ( n12120 & n22364 ) ;
  assign n28442 = n12439 ^ n7760 ^ 1'b0 ;
  assign n28443 = ( n5869 & ~n10389 ) | ( n5869 & n28442 ) | ( ~n10389 & n28442 ) ;
  assign n28444 = ( ~n3129 & n14366 ) | ( ~n3129 & n28443 ) | ( n14366 & n28443 ) ;
  assign n28445 = n20421 ^ n4014 ^ n2287 ;
  assign n28446 = ( n2586 & n15300 ) | ( n2586 & ~n24824 ) | ( n15300 & ~n24824 ) ;
  assign n28447 = ( n5701 & n7021 ) | ( n5701 & n7879 ) | ( n7021 & n7879 ) ;
  assign n28448 = n28447 ^ n2530 ^ n1125 ;
  assign n28449 = n2014 | n28448 ;
  assign n28450 = n28449 ^ n10351 ^ 1'b0 ;
  assign n28451 = n28450 ^ n9524 ^ n530 ;
  assign n28452 = ~n906 & n9973 ;
  assign n28453 = n17826 & n28452 ;
  assign n28454 = n1097 & ~n11250 ;
  assign n28455 = n28454 ^ n3182 ^ 1'b0 ;
  assign n28456 = ( n1575 & ~n2285 ) | ( n1575 & n28455 ) | ( ~n2285 & n28455 ) ;
  assign n28457 = n25321 ^ n16431 ^ n16402 ;
  assign n28458 = n28457 ^ n26662 ^ n444 ;
  assign n28459 = ( ~n7715 & n20688 ) | ( ~n7715 & n22070 ) | ( n20688 & n22070 ) ;
  assign n28460 = ( n1329 & ~n3212 ) | ( n1329 & n5145 ) | ( ~n3212 & n5145 ) ;
  assign n28461 = ( n16905 & n25920 ) | ( n16905 & n28460 ) | ( n25920 & n28460 ) ;
  assign n28462 = n28461 ^ n14109 ^ n1629 ;
  assign n28463 = ( n12442 & n15004 ) | ( n12442 & ~n28462 ) | ( n15004 & ~n28462 ) ;
  assign n28464 = ( n2015 & n12166 ) | ( n2015 & ~n22315 ) | ( n12166 & ~n22315 ) ;
  assign n28465 = ( ~n1487 & n3191 ) | ( ~n1487 & n20804 ) | ( n3191 & n20804 ) ;
  assign n28466 = ( n15288 & ~n19092 ) | ( n15288 & n28465 ) | ( ~n19092 & n28465 ) ;
  assign n28467 = ( ~n19937 & n28464 ) | ( ~n19937 & n28466 ) | ( n28464 & n28466 ) ;
  assign n28468 = n25102 ^ n22780 ^ 1'b0 ;
  assign n28469 = n16353 ^ n5430 ^ n4578 ;
  assign n28470 = n14932 ^ n5224 ^ n1717 ;
  assign n28471 = ( ~n20023 & n28469 ) | ( ~n20023 & n28470 ) | ( n28469 & n28470 ) ;
  assign n28472 = ( n8823 & n10356 ) | ( n8823 & ~n28471 ) | ( n10356 & ~n28471 ) ;
  assign n28473 = n5769 ^ n4562 ^ 1'b0 ;
  assign n28474 = ~n18092 & n28473 ;
  assign n28475 = ( n8730 & ~n14237 ) | ( n8730 & n18065 ) | ( ~n14237 & n18065 ) ;
  assign n28476 = ( ~n4836 & n23358 ) | ( ~n4836 & n27002 ) | ( n23358 & n27002 ) ;
  assign n28477 = ( n3257 & ~n3723 ) | ( n3257 & n4120 ) | ( ~n3723 & n4120 ) ;
  assign n28478 = n6867 & ~n28477 ;
  assign n28479 = n28476 & n28478 ;
  assign n28480 = ( n15404 & n28475 ) | ( n15404 & n28479 ) | ( n28475 & n28479 ) ;
  assign n28483 = ~n12189 & n15820 ;
  assign n28484 = n28483 ^ n12467 ^ n1765 ;
  assign n28485 = ( n4390 & ~n17776 ) | ( n4390 & n28484 ) | ( ~n17776 & n28484 ) ;
  assign n28481 = n13298 ^ n11076 ^ n9860 ;
  assign n28482 = n28481 ^ n24586 ^ n13878 ;
  assign n28486 = n28485 ^ n28482 ^ n586 ;
  assign n28487 = ( n12026 & n28480 ) | ( n12026 & n28486 ) | ( n28480 & n28486 ) ;
  assign n28488 = ( n2138 & n6229 ) | ( n2138 & n7603 ) | ( n6229 & n7603 ) ;
  assign n28489 = n28488 ^ n25183 ^ n8448 ;
  assign n28491 = n971 & n2583 ;
  assign n28492 = n7898 & n28491 ;
  assign n28490 = n18593 ^ n4471 ^ n888 ;
  assign n28493 = n28492 ^ n28490 ^ n26139 ;
  assign n28494 = ( n5659 & n21754 ) | ( n5659 & n25134 ) | ( n21754 & n25134 ) ;
  assign n28495 = n16278 ^ n12460 ^ n4204 ;
  assign n28496 = ( n1781 & ~n7210 ) | ( n1781 & n28495 ) | ( ~n7210 & n28495 ) ;
  assign n28497 = n18996 | n22759 ;
  assign n28498 = ( ~n6534 & n14158 ) | ( ~n6534 & n26102 ) | ( n14158 & n26102 ) ;
  assign n28499 = n28498 ^ n11728 ^ x54 ;
  assign n28500 = ( n8006 & n28429 ) | ( n8006 & n28499 ) | ( n28429 & n28499 ) ;
  assign n28501 = n11240 | n12071 ;
  assign n28502 = n11741 | n28501 ;
  assign n28503 = n28502 ^ n5191 ^ 1'b0 ;
  assign n28504 = n23966 ^ n17620 ^ n5254 ;
  assign n28505 = n28504 ^ n26191 ^ 1'b0 ;
  assign n28506 = ( n10746 & n12739 ) | ( n10746 & n25784 ) | ( n12739 & n25784 ) ;
  assign n28507 = ( ~n18951 & n27169 ) | ( ~n18951 & n28506 ) | ( n27169 & n28506 ) ;
  assign n28508 = n26477 ^ n21363 ^ n16081 ;
  assign n28509 = n28508 ^ n24412 ^ n20049 ;
  assign n28510 = ~n13543 & n19495 ;
  assign n28511 = ( n12095 & n14062 ) | ( n12095 & ~n17128 ) | ( n14062 & ~n17128 ) ;
  assign n28512 = n12660 ^ n10551 ^ n7525 ;
  assign n28513 = n28512 ^ n9030 ^ n6889 ;
  assign n28514 = ( n9795 & ~n28511 ) | ( n9795 & n28513 ) | ( ~n28511 & n28513 ) ;
  assign n28517 = ( n3533 & n8497 ) | ( n3533 & ~n10176 ) | ( n8497 & ~n10176 ) ;
  assign n28515 = n14356 ^ n8002 ^ n6227 ;
  assign n28516 = ( n6926 & n8974 ) | ( n6926 & ~n28515 ) | ( n8974 & ~n28515 ) ;
  assign n28518 = n28517 ^ n28516 ^ n27305 ;
  assign n28519 = n22944 ^ n14421 ^ n13194 ;
  assign n28520 = n19414 & ~n20947 ;
  assign n28521 = ~n28519 & n28520 ;
  assign n28522 = n28521 ^ n8897 ^ n6665 ;
  assign n28523 = n22833 ^ n15344 ^ n6613 ;
  assign n28524 = n18740 ^ n11651 ^ n2383 ;
  assign n28525 = ~n4878 & n9729 ;
  assign n28526 = ~n787 & n28525 ;
  assign n28527 = ( n2471 & n8648 ) | ( n2471 & ~n18589 ) | ( n8648 & ~n18589 ) ;
  assign n28528 = n4073 | n28527 ;
  assign n28529 = n28528 ^ n23691 ^ 1'b0 ;
  assign n28530 = n20611 ^ n12161 ^ n11601 ;
  assign n28531 = ( n6697 & n8854 ) | ( n6697 & n28530 ) | ( n8854 & n28530 ) ;
  assign n28532 = n15576 ^ n14776 ^ n6109 ;
  assign n28533 = n25289 ^ n14166 ^ n8365 ;
  assign n28534 = ( n19447 & n28532 ) | ( n19447 & n28533 ) | ( n28532 & n28533 ) ;
  assign n28535 = n28534 ^ n13340 ^ n779 ;
  assign n28536 = n23659 ^ n17302 ^ n9381 ;
  assign n28537 = n25710 ^ n18087 ^ n10798 ;
  assign n28538 = n1598 | n5066 ;
  assign n28539 = n7541 & ~n28538 ;
  assign n28540 = ( ~n12906 & n28537 ) | ( ~n12906 & n28539 ) | ( n28537 & n28539 ) ;
  assign n28541 = ( n5312 & ~n12643 ) | ( n5312 & n18276 ) | ( ~n12643 & n18276 ) ;
  assign n28542 = ( ~n17463 & n23907 ) | ( ~n17463 & n28541 ) | ( n23907 & n28541 ) ;
  assign n28543 = n19109 ^ n13193 ^ n12305 ;
  assign n28544 = ( n4527 & n10097 ) | ( n4527 & ~n28543 ) | ( n10097 & ~n28543 ) ;
  assign n28547 = ( n6220 & ~n15905 ) | ( n6220 & n24752 ) | ( ~n15905 & n24752 ) ;
  assign n28545 = n3775 & n12199 ;
  assign n28546 = n28545 ^ n9495 ^ 1'b0 ;
  assign n28548 = n28547 ^ n28546 ^ n5773 ;
  assign n28549 = n15771 ^ n12086 ^ 1'b0 ;
  assign n28550 = n28549 ^ n21816 ^ n9461 ;
  assign n28551 = ( ~n15195 & n28548 ) | ( ~n15195 & n28550 ) | ( n28548 & n28550 ) ;
  assign n28552 = n11863 ^ n4003 ^ 1'b0 ;
  assign n28553 = ~n3565 & n28552 ;
  assign n28554 = n28553 ^ n18447 ^ n11108 ;
  assign n28555 = n18005 ^ n11782 ^ n6387 ;
  assign n28556 = ( n1204 & ~n18514 ) | ( n1204 & n20808 ) | ( ~n18514 & n20808 ) ;
  assign n28557 = n28556 ^ n27398 ^ n16229 ;
  assign n28558 = ( ~n3530 & n9558 ) | ( ~n3530 & n26781 ) | ( n9558 & n26781 ) ;
  assign n28559 = n28558 ^ n24306 ^ n8298 ;
  assign n28560 = n6242 ^ n4575 ^ n1283 ;
  assign n28561 = n22747 ^ n18077 ^ n9884 ;
  assign n28562 = n25383 ^ n9554 ^ n4807 ;
  assign n28563 = n16999 ^ n8727 ^ n1533 ;
  assign n28564 = ( n5318 & n13518 ) | ( n5318 & ~n21362 ) | ( n13518 & ~n21362 ) ;
  assign n28565 = n20310 ^ n2948 ^ 1'b0 ;
  assign n28566 = n27996 & n28565 ;
  assign n28567 = n28564 & n28566 ;
  assign n28568 = x37 & n16553 ;
  assign n28569 = n28568 ^ n20442 ^ 1'b0 ;
  assign n28570 = ( n9671 & n10264 ) | ( n9671 & ~n28569 ) | ( n10264 & ~n28569 ) ;
  assign n28571 = n15540 ^ n14832 ^ n6946 ;
  assign n28572 = n1716 & ~n16784 ;
  assign n28573 = ~n3698 & n28572 ;
  assign n28574 = n28573 ^ n22170 ^ n7661 ;
  assign n28576 = ( n7249 & n23528 ) | ( n7249 & n27075 ) | ( n23528 & n27075 ) ;
  assign n28575 = ( n13571 & n15104 ) | ( n13571 & n22061 ) | ( n15104 & n22061 ) ;
  assign n28577 = n28576 ^ n28575 ^ n24344 ;
  assign n28578 = n3444 ^ n2380 ^ n2198 ;
  assign n28580 = ( n8400 & n11842 ) | ( n8400 & n12789 ) | ( n11842 & n12789 ) ;
  assign n28579 = n13694 ^ n12121 ^ n7118 ;
  assign n28581 = n28580 ^ n28579 ^ n11511 ;
  assign n28582 = ( n8274 & n28578 ) | ( n8274 & ~n28581 ) | ( n28578 & ~n28581 ) ;
  assign n28583 = n28235 ^ n13649 ^ 1'b0 ;
  assign n28584 = n703 & ~n3879 ;
  assign n28585 = ~n5910 & n28584 ;
  assign n28586 = n10315 & n23458 ;
  assign n28587 = n8902 & n28586 ;
  assign n28588 = ( ~n4461 & n11408 ) | ( ~n4461 & n24740 ) | ( n11408 & n24740 ) ;
  assign n28589 = ( n28585 & ~n28587 ) | ( n28585 & n28588 ) | ( ~n28587 & n28588 ) ;
  assign n28590 = ~n17619 & n19260 ;
  assign n28591 = ( n9013 & n12096 ) | ( n9013 & ~n17514 ) | ( n12096 & ~n17514 ) ;
  assign n28592 = ( n21324 & ~n27560 ) | ( n21324 & n28591 ) | ( ~n27560 & n28591 ) ;
  assign n28593 = ( n20760 & ~n28590 ) | ( n20760 & n28592 ) | ( ~n28590 & n28592 ) ;
  assign n28594 = n28593 ^ n24594 ^ n3570 ;
  assign n28595 = n20443 ^ n16317 ^ n8506 ;
  assign n28596 = n13790 & n23411 ;
  assign n28597 = n28596 ^ n9414 ^ 1'b0 ;
  assign n28598 = n14068 ^ n13486 ^ n10452 ;
  assign n28599 = ( n8103 & n15221 ) | ( n8103 & n28598 ) | ( n15221 & n28598 ) ;
  assign n28600 = ( n6307 & n7005 ) | ( n6307 & ~n14259 ) | ( n7005 & ~n14259 ) ;
  assign n28601 = n28600 ^ n2629 ^ 1'b0 ;
  assign n28602 = n28599 & n28601 ;
  assign n28606 = n6955 | n8374 ;
  assign n28607 = n21658 & ~n28606 ;
  assign n28603 = ( n12537 & ~n14237 ) | ( n12537 & n14754 ) | ( ~n14237 & n14754 ) ;
  assign n28604 = n5771 | n28603 ;
  assign n28605 = n1022 | n28604 ;
  assign n28608 = n28607 ^ n28605 ^ 1'b0 ;
  assign n28609 = n21549 ^ n11414 ^ 1'b0 ;
  assign n28610 = ( n26389 & n28608 ) | ( n26389 & ~n28609 ) | ( n28608 & ~n28609 ) ;
  assign n28611 = n18781 ^ n4104 ^ n827 ;
  assign n28612 = ( ~n4721 & n5882 ) | ( ~n4721 & n18345 ) | ( n5882 & n18345 ) ;
  assign n28613 = ( n5290 & ~n5382 ) | ( n5290 & n19766 ) | ( ~n5382 & n19766 ) ;
  assign n28614 = n1778 | n13923 ;
  assign n28615 = n15547 ^ n5861 ^ 1'b0 ;
  assign n28616 = ( ~n212 & n21009 ) | ( ~n212 & n28615 ) | ( n21009 & n28615 ) ;
  assign n28617 = ( ~n21216 & n28614 ) | ( ~n21216 & n28616 ) | ( n28614 & n28616 ) ;
  assign n28618 = ( ~n22934 & n28613 ) | ( ~n22934 & n28617 ) | ( n28613 & n28617 ) ;
  assign n28619 = ( ~n2171 & n5505 ) | ( ~n2171 & n7553 ) | ( n5505 & n7553 ) ;
  assign n28620 = ( ~n7980 & n21447 ) | ( ~n7980 & n21768 ) | ( n21447 & n21768 ) ;
  assign n28621 = n21449 ^ n15779 ^ n1725 ;
  assign n28622 = n28366 ^ n27450 ^ n9686 ;
  assign n28623 = ( ~n1047 & n1410 ) | ( ~n1047 & n13509 ) | ( n1410 & n13509 ) ;
  assign n28624 = n28623 ^ n19446 ^ n12691 ;
  assign n28625 = ( n567 & n20051 ) | ( n567 & ~n28624 ) | ( n20051 & ~n28624 ) ;
  assign n28626 = n21948 ^ n5077 ^ n506 ;
  assign n28632 = ( n507 & n1477 ) | ( n507 & ~n13362 ) | ( n1477 & ~n13362 ) ;
  assign n28630 = n7383 & ~n16725 ;
  assign n28631 = n12683 & n28630 ;
  assign n28627 = n16040 ^ n13542 ^ n2273 ;
  assign n28628 = n301 & n28627 ;
  assign n28629 = ~n19900 & n28628 ;
  assign n28633 = n28632 ^ n28631 ^ n28629 ;
  assign n28634 = ( ~n3232 & n5775 ) | ( ~n3232 & n13111 ) | ( n5775 & n13111 ) ;
  assign n28635 = ( n5851 & n15228 ) | ( n5851 & n28634 ) | ( n15228 & n28634 ) ;
  assign n28636 = n28635 ^ n26614 ^ n23504 ;
  assign n28639 = ( ~n3656 & n3675 ) | ( ~n3656 & n7665 ) | ( n3675 & n7665 ) ;
  assign n28637 = ( n10825 & n11901 ) | ( n10825 & n17061 ) | ( n11901 & n17061 ) ;
  assign n28638 = ( n16951 & n19620 ) | ( n16951 & n28637 ) | ( n19620 & n28637 ) ;
  assign n28640 = n28639 ^ n28638 ^ n11193 ;
  assign n28641 = ( n13479 & n15265 ) | ( n13479 & ~n28640 ) | ( n15265 & ~n28640 ) ;
  assign n28642 = n5602 ^ n1198 ^ 1'b0 ;
  assign n28643 = n16223 ^ n6516 ^ 1'b0 ;
  assign n28644 = n432 & n28643 ;
  assign n28645 = n17282 ^ n13473 ^ n5671 ;
  assign n28646 = n16836 & ~n28645 ;
  assign n28647 = n9171 ^ n5675 ^ n1637 ;
  assign n28648 = ( n10310 & n10844 ) | ( n10310 & ~n25905 ) | ( n10844 & ~n25905 ) ;
  assign n28649 = ( n5015 & ~n7564 ) | ( n5015 & n27594 ) | ( ~n7564 & n27594 ) ;
  assign n28650 = n22626 ^ n19043 ^ n5782 ;
  assign n28651 = ( ~n9775 & n11241 ) | ( ~n9775 & n26570 ) | ( n11241 & n26570 ) ;
  assign n28652 = ( n7096 & n8279 ) | ( n7096 & n11853 ) | ( n8279 & n11853 ) ;
  assign n28653 = ~n1835 & n4771 ;
  assign n28654 = n28653 ^ n1210 ^ 1'b0 ;
  assign n28655 = ( ~n18654 & n28652 ) | ( ~n18654 & n28654 ) | ( n28652 & n28654 ) ;
  assign n28662 = n9114 & ~n22822 ;
  assign n28663 = ~n9445 & n28662 ;
  assign n28664 = n28663 ^ n8021 ^ 1'b0 ;
  assign n28661 = ( ~n8519 & n17288 ) | ( ~n8519 & n27733 ) | ( n17288 & n27733 ) ;
  assign n28657 = ( n1438 & n1841 ) | ( n1438 & ~n5430 ) | ( n1841 & ~n5430 ) ;
  assign n28656 = n14208 ^ n10616 ^ n3657 ;
  assign n28658 = n28657 ^ n28656 ^ n12359 ;
  assign n28659 = ( ~n1323 & n11217 ) | ( ~n1323 & n16687 ) | ( n11217 & n16687 ) ;
  assign n28660 = ( n13514 & n28658 ) | ( n13514 & n28659 ) | ( n28658 & n28659 ) ;
  assign n28665 = n28664 ^ n28661 ^ n28660 ;
  assign n28666 = n23550 ^ n4301 ^ 1'b0 ;
  assign n28667 = n10021 ^ n9035 ^ n6148 ;
  assign n28668 = n22535 ^ n3851 ^ 1'b0 ;
  assign n28669 = n28667 & n28668 ;
  assign n28670 = n28669 ^ n20201 ^ n745 ;
  assign n28671 = n27351 ^ n7182 ^ 1'b0 ;
  assign n28672 = ( ~n5599 & n18933 ) | ( ~n5599 & n28415 ) | ( n18933 & n28415 ) ;
  assign n28673 = ( n12314 & ~n12578 ) | ( n12314 & n28159 ) | ( ~n12578 & n28159 ) ;
  assign n28674 = n20018 ^ n9780 ^ n2138 ;
  assign n28675 = n6086 & n8323 ;
  assign n28676 = n20214 & n28675 ;
  assign n28677 = ( ~n20820 & n28674 ) | ( ~n20820 & n28676 ) | ( n28674 & n28676 ) ;
  assign n28679 = n25263 ^ n10682 ^ n1935 ;
  assign n28678 = n9365 ^ n6275 ^ 1'b0 ;
  assign n28680 = n28679 ^ n28678 ^ n24483 ;
  assign n28681 = n1379 & n13292 ;
  assign n28682 = n28681 ^ n4149 ^ 1'b0 ;
  assign n28683 = n3735 & n6601 ;
  assign n28684 = n28683 ^ n22609 ^ 1'b0 ;
  assign n28685 = n18239 & ~n26418 ;
  assign n28686 = ~n2530 & n11088 ;
  assign n28687 = n27966 ^ n17261 ^ n1692 ;
  assign n28688 = ( ~n204 & n12422 ) | ( ~n204 & n17085 ) | ( n12422 & n17085 ) ;
  assign n28689 = n28688 ^ n18881 ^ n11926 ;
  assign n28690 = ( n26199 & ~n28687 ) | ( n26199 & n28689 ) | ( ~n28687 & n28689 ) ;
  assign n28691 = ( n3218 & n11222 ) | ( n3218 & n28107 ) | ( n11222 & n28107 ) ;
  assign n28692 = ~n6894 & n25190 ;
  assign n28693 = ~n16266 & n28692 ;
  assign n28694 = n28693 ^ n25922 ^ n9517 ;
  assign n28695 = n3047 & ~n9321 ;
  assign n28696 = n28695 ^ n6727 ^ 1'b0 ;
  assign n28697 = ~n21662 & n28696 ;
  assign n28698 = ( n2953 & n3124 ) | ( n2953 & n7769 ) | ( n3124 & n7769 ) ;
  assign n28699 = n26690 ^ n21446 ^ n4723 ;
  assign n28700 = n27418 ^ n7467 ^ n2717 ;
  assign n28701 = ( n28698 & n28699 ) | ( n28698 & ~n28700 ) | ( n28699 & ~n28700 ) ;
  assign n28702 = n12643 ^ n5998 ^ n1478 ;
  assign n28703 = n28702 ^ n16529 ^ n1208 ;
  assign n28704 = n28703 ^ n14710 ^ n3141 ;
  assign n28705 = n9629 ^ n3303 ^ 1'b0 ;
  assign n28706 = n23935 ^ n17500 ^ n8360 ;
  assign n28707 = ( ~n442 & n2981 ) | ( ~n442 & n21752 ) | ( n2981 & n21752 ) ;
  assign n28708 = ( n12348 & n19765 ) | ( n12348 & n28707 ) | ( n19765 & n28707 ) ;
  assign n28709 = n13676 ^ n1583 ^ n576 ;
  assign n28710 = n24807 ^ n9942 ^ 1'b0 ;
  assign n28711 = n27500 ^ n11636 ^ n5217 ;
  assign n28712 = ~n2475 & n21503 ;
  assign n28713 = ( ~n1881 & n11716 ) | ( ~n1881 & n19728 ) | ( n11716 & n19728 ) ;
  assign n28714 = ( n12744 & ~n16585 ) | ( n12744 & n28654 ) | ( ~n16585 & n28654 ) ;
  assign n28715 = ~n6496 & n13590 ;
  assign n28716 = n24864 ^ n15621 ^ n3951 ;
  assign n28717 = n28716 ^ n23337 ^ 1'b0 ;
  assign n28718 = n28715 & ~n28717 ;
  assign n28719 = n10066 ^ n3519 ^ 1'b0 ;
  assign n28720 = ~n9302 & n28719 ;
  assign n28721 = ( n3574 & n6762 ) | ( n3574 & ~n11672 ) | ( n6762 & ~n11672 ) ;
  assign n28722 = n9569 ^ n6475 ^ n2413 ;
  assign n28723 = n28722 ^ n9042 ^ n2770 ;
  assign n28724 = ( n1339 & ~n28721 ) | ( n1339 & n28723 ) | ( ~n28721 & n28723 ) ;
  assign n28725 = ( n460 & ~n5287 ) | ( n460 & n28724 ) | ( ~n5287 & n28724 ) ;
  assign n28726 = n28725 ^ n22427 ^ 1'b0 ;
  assign n28727 = n20538 ^ n4633 ^ n2193 ;
  assign n28728 = ( n1083 & n1537 ) | ( n1083 & n16568 ) | ( n1537 & n16568 ) ;
  assign n28729 = ( ~n28284 & n28727 ) | ( ~n28284 & n28728 ) | ( n28727 & n28728 ) ;
  assign n28730 = n25286 ^ n12112 ^ n10531 ;
  assign n28731 = n28730 ^ n10371 ^ 1'b0 ;
  assign n28732 = ( n3514 & ~n9479 ) | ( n3514 & n10418 ) | ( ~n9479 & n10418 ) ;
  assign n28733 = ( n793 & n1892 ) | ( n793 & ~n5387 ) | ( n1892 & ~n5387 ) ;
  assign n28734 = n28733 ^ n12128 ^ n3366 ;
  assign n28735 = ( n5425 & n28732 ) | ( n5425 & ~n28734 ) | ( n28732 & ~n28734 ) ;
  assign n28736 = ( n2235 & ~n14609 ) | ( n2235 & n21260 ) | ( ~n14609 & n21260 ) ;
  assign n28737 = ( n3942 & n25924 ) | ( n3942 & n26298 ) | ( n25924 & n26298 ) ;
  assign n28738 = n26514 ^ n23805 ^ 1'b0 ;
  assign n28739 = n21415 ^ n7851 ^ 1'b0 ;
  assign n28740 = n23292 ^ n14876 ^ n8057 ;
  assign n28741 = n28740 ^ n4556 ^ x93 ;
  assign n28749 = ( n5860 & ~n7783 ) | ( n5860 & n12077 ) | ( ~n7783 & n12077 ) ;
  assign n28742 = n18493 ^ n17402 ^ n6609 ;
  assign n28743 = ( ~n8260 & n12251 ) | ( ~n8260 & n17056 ) | ( n12251 & n17056 ) ;
  assign n28744 = ( n19561 & n28742 ) | ( n19561 & n28743 ) | ( n28742 & n28743 ) ;
  assign n28745 = ( n9897 & n11048 ) | ( n9897 & ~n19315 ) | ( n11048 & ~n19315 ) ;
  assign n28746 = ( n19658 & n28744 ) | ( n19658 & ~n28745 ) | ( n28744 & ~n28745 ) ;
  assign n28747 = n28746 ^ n1941 ^ 1'b0 ;
  assign n28748 = n26868 & n28747 ;
  assign n28750 = n28749 ^ n28748 ^ n26670 ;
  assign n28751 = n11097 ^ n2062 ^ n841 ;
  assign n28752 = ( ~n5304 & n21025 ) | ( ~n5304 & n28751 ) | ( n21025 & n28751 ) ;
  assign n28754 = ( ~n7187 & n13619 ) | ( ~n7187 & n23951 ) | ( n13619 & n23951 ) ;
  assign n28755 = ~n7189 & n28754 ;
  assign n28753 = ( n10749 & n23175 ) | ( n10749 & n27483 ) | ( n23175 & n27483 ) ;
  assign n28756 = n28755 ^ n28753 ^ n7533 ;
  assign n28757 = n6849 ^ n6360 ^ n3538 ;
  assign n28758 = n22740 ^ n16913 ^ n11484 ;
  assign n28759 = ~n22447 & n28758 ;
  assign n28760 = ~n4737 & n13992 ;
  assign n28761 = ( n3628 & n6922 ) | ( n3628 & n20373 ) | ( n6922 & n20373 ) ;
  assign n28762 = ( n9349 & n20798 ) | ( n9349 & n28761 ) | ( n20798 & n28761 ) ;
  assign n28763 = ( ~n16204 & n23933 ) | ( ~n16204 & n25007 ) | ( n23933 & n25007 ) ;
  assign n28764 = n5087 | n9134 ;
  assign n28765 = n28764 ^ n9325 ^ 1'b0 ;
  assign n28766 = n12725 ^ n11061 ^ n7890 ;
  assign n28767 = ( n508 & ~n11412 ) | ( n508 & n15225 ) | ( ~n11412 & n15225 ) ;
  assign n28768 = ( n7460 & ~n12119 ) | ( n7460 & n28767 ) | ( ~n12119 & n28767 ) ;
  assign n28769 = ( n2728 & ~n28549 ) | ( n2728 & n28768 ) | ( ~n28549 & n28768 ) ;
  assign n28770 = ( n4270 & ~n11146 ) | ( n4270 & n25651 ) | ( ~n11146 & n25651 ) ;
  assign n28771 = n21011 ^ n7373 ^ n2970 ;
  assign n28772 = ( n2105 & n9493 ) | ( n2105 & n28771 ) | ( n9493 & n28771 ) ;
  assign n28773 = n12457 & n28772 ;
  assign n28774 = ( n1376 & n2276 ) | ( n1376 & n7614 ) | ( n2276 & n7614 ) ;
  assign n28775 = n20231 ^ n16605 ^ 1'b0 ;
  assign n28776 = n28774 & ~n28775 ;
  assign n28778 = n10723 ^ n7658 ^ n1448 ;
  assign n28777 = n8905 ^ n7963 ^ n3746 ;
  assign n28779 = n28778 ^ n28777 ^ 1'b0 ;
  assign n28781 = n12907 ^ n4403 ^ n1792 ;
  assign n28780 = n20746 ^ n15751 ^ n11493 ;
  assign n28782 = n28781 ^ n28780 ^ n17630 ;
  assign n28783 = ( n7281 & ~n8412 ) | ( n7281 & n14374 ) | ( ~n8412 & n14374 ) ;
  assign n28784 = ( n4993 & n7997 ) | ( n4993 & ~n28783 ) | ( n7997 & ~n28783 ) ;
  assign n28785 = ( ~n7622 & n15948 ) | ( ~n7622 & n28784 ) | ( n15948 & n28784 ) ;
  assign n28786 = ( n1363 & n16094 ) | ( n1363 & n24262 ) | ( n16094 & n24262 ) ;
  assign n28787 = ( n7912 & ~n25331 ) | ( n7912 & n25765 ) | ( ~n25331 & n25765 ) ;
  assign n28788 = ( n13137 & n28786 ) | ( n13137 & ~n28787 ) | ( n28786 & ~n28787 ) ;
  assign n28789 = n28788 ^ n15246 ^ n13990 ;
  assign n28790 = ( ~n134 & n5836 ) | ( ~n134 & n8220 ) | ( n5836 & n8220 ) ;
  assign n28791 = ( n1552 & ~n11218 ) | ( n1552 & n11862 ) | ( ~n11218 & n11862 ) ;
  assign n28792 = ( n2558 & ~n28790 ) | ( n2558 & n28791 ) | ( ~n28790 & n28791 ) ;
  assign n28793 = n28792 ^ n12019 ^ n10376 ;
  assign n28794 = ( n7307 & n17801 ) | ( n7307 & ~n28793 ) | ( n17801 & ~n28793 ) ;
  assign n28795 = ( n14066 & ~n15301 ) | ( n14066 & n23828 ) | ( ~n15301 & n23828 ) ;
  assign n28796 = ( n14174 & n25600 ) | ( n14174 & ~n28795 ) | ( n25600 & ~n28795 ) ;
  assign n28797 = n23529 ^ n10961 ^ 1'b0 ;
  assign n28798 = n16422 & n25760 ;
  assign n28799 = n28798 ^ n3590 ^ 1'b0 ;
  assign n28800 = ( n5261 & n24114 ) | ( n5261 & n25470 ) | ( n24114 & n25470 ) ;
  assign n28801 = ( n11847 & ~n28799 ) | ( n11847 & n28800 ) | ( ~n28799 & n28800 ) ;
  assign n28802 = n16423 ^ n6430 ^ 1'b0 ;
  assign n28803 = n14061 & n28802 ;
  assign n28804 = ~n3401 & n28803 ;
  assign n28805 = n28804 ^ n16657 ^ 1'b0 ;
  assign n28806 = ( n11776 & n12261 ) | ( n11776 & n19216 ) | ( n12261 & n19216 ) ;
  assign n28807 = ~n4106 & n28806 ;
  assign n28808 = n28807 ^ n15570 ^ 1'b0 ;
  assign n28809 = ( ~n363 & n1459 ) | ( ~n363 & n7558 ) | ( n1459 & n7558 ) ;
  assign n28810 = ( n13927 & n14688 ) | ( n13927 & n20912 ) | ( n14688 & n20912 ) ;
  assign n28811 = ( n2437 & n15635 ) | ( n2437 & ~n28810 ) | ( n15635 & ~n28810 ) ;
  assign n28812 = ( n23884 & ~n28809 ) | ( n23884 & n28811 ) | ( ~n28809 & n28811 ) ;
  assign n28813 = ( n7963 & ~n25861 ) | ( n7963 & n27231 ) | ( ~n25861 & n27231 ) ;
  assign n28814 = ( n1173 & ~n4621 ) | ( n1173 & n5818 ) | ( ~n4621 & n5818 ) ;
  assign n28818 = n19164 ^ n7539 ^ n1548 ;
  assign n28819 = n28818 ^ n7064 ^ n5519 ;
  assign n28820 = n28819 ^ n10239 ^ n5025 ;
  assign n28816 = n6984 ^ n4975 ^ n543 ;
  assign n28815 = n18379 ^ n9495 ^ n8849 ;
  assign n28817 = n28816 ^ n28815 ^ n2756 ;
  assign n28821 = n28820 ^ n28817 ^ n24250 ;
  assign n28822 = n27863 ^ n13870 ^ n8932 ;
  assign n28823 = n28822 ^ n19105 ^ n6570 ;
  assign n28824 = n28823 ^ n20920 ^ n7087 ;
  assign n28825 = n19495 ^ n19454 ^ n3544 ;
  assign n28827 = ( ~n9064 & n12521 ) | ( ~n9064 & n16153 ) | ( n12521 & n16153 ) ;
  assign n28826 = ( n8060 & n17162 ) | ( n8060 & ~n24506 ) | ( n17162 & ~n24506 ) ;
  assign n28828 = n28827 ^ n28826 ^ n24359 ;
  assign n28829 = ( ~n1608 & n27655 ) | ( ~n1608 & n28828 ) | ( n27655 & n28828 ) ;
  assign n28830 = n6896 ^ n4391 ^ 1'b0 ;
  assign n28831 = n28830 ^ n13091 ^ n9438 ;
  assign n28832 = ~n11046 & n11250 ;
  assign n28833 = ( n1804 & n26622 ) | ( n1804 & n28832 ) | ( n26622 & n28832 ) ;
  assign n28834 = n28833 ^ n1692 ^ 1'b0 ;
  assign n28835 = n7303 & n28834 ;
  assign n28836 = ( n8100 & ~n16492 ) | ( n8100 & n18747 ) | ( ~n16492 & n18747 ) ;
  assign n28837 = ( n4703 & ~n12115 ) | ( n4703 & n23766 ) | ( ~n12115 & n23766 ) ;
  assign n28838 = ( n1839 & n10456 ) | ( n1839 & n12436 ) | ( n10456 & n12436 ) ;
  assign n28839 = ( n7355 & ~n17501 ) | ( n7355 & n23942 ) | ( ~n17501 & n23942 ) ;
  assign n28840 = ( ~n14200 & n15049 ) | ( ~n14200 & n24007 ) | ( n15049 & n24007 ) ;
  assign n28841 = ( n16851 & n16902 ) | ( n16851 & n18109 ) | ( n16902 & n18109 ) ;
  assign n28842 = ( n8041 & n10052 ) | ( n8041 & ~n28841 ) | ( n10052 & ~n28841 ) ;
  assign n28844 = ( n8550 & n11878 ) | ( n8550 & n20285 ) | ( n11878 & n20285 ) ;
  assign n28843 = n18580 ^ n6348 ^ 1'b0 ;
  assign n28845 = n28844 ^ n28843 ^ n22461 ;
  assign n28846 = n6313 ^ n4666 ^ n1163 ;
  assign n28847 = ( ~n13849 & n16079 ) | ( ~n13849 & n28846 ) | ( n16079 & n28846 ) ;
  assign n28848 = n9717 ^ n6567 ^ n5622 ;
  assign n28849 = n18243 ^ n6726 ^ x101 ;
  assign n28850 = n28849 ^ n23964 ^ n5225 ;
  assign n28851 = n28850 ^ n25516 ^ n23600 ;
  assign n28852 = n19270 ^ n2332 ^ 1'b0 ;
  assign n28853 = n1639 & ~n28852 ;
  assign n28854 = n28853 ^ n17776 ^ n13145 ;
  assign n28855 = n16455 ^ n15016 ^ n2927 ;
  assign n28856 = n24169 ^ n7885 ^ 1'b0 ;
  assign n28857 = ( n761 & n3382 ) | ( n761 & ~n11768 ) | ( n3382 & ~n11768 ) ;
  assign n28858 = n22760 ^ n10386 ^ n5033 ;
  assign n28859 = ( n591 & ~n15845 ) | ( n591 & n28858 ) | ( ~n15845 & n28858 ) ;
  assign n28860 = n28859 ^ n14683 ^ n6863 ;
  assign n28861 = n23222 ^ n20003 ^ n1354 ;
  assign n28862 = ( x68 & ~n28860 ) | ( x68 & n28861 ) | ( ~n28860 & n28861 ) ;
  assign n28863 = ( n7956 & n28857 ) | ( n7956 & ~n28862 ) | ( n28857 & ~n28862 ) ;
  assign n28864 = n25275 ^ n9526 ^ n2112 ;
  assign n28865 = n2741 | n15209 ;
  assign n28866 = n28865 ^ n12097 ^ 1'b0 ;
  assign n28867 = ( n1095 & n11804 ) | ( n1095 & n28866 ) | ( n11804 & n28866 ) ;
  assign n28868 = ( ~n2609 & n12276 ) | ( ~n2609 & n19854 ) | ( n12276 & n19854 ) ;
  assign n28869 = n4390 & ~n28868 ;
  assign n28870 = ~n28867 & n28869 ;
  assign n28874 = ( n3499 & ~n7468 ) | ( n3499 & n10749 ) | ( ~n7468 & n10749 ) ;
  assign n28873 = ( n2924 & n4550 ) | ( n2924 & ~n11580 ) | ( n4550 & ~n11580 ) ;
  assign n28871 = n9250 ^ n1271 ^ 1'b0 ;
  assign n28872 = n19731 & ~n28871 ;
  assign n28875 = n28874 ^ n28873 ^ n28872 ;
  assign n28876 = ( ~n971 & n1024 ) | ( ~n971 & n12421 ) | ( n1024 & n12421 ) ;
  assign n28877 = ( n4685 & ~n10124 ) | ( n4685 & n28876 ) | ( ~n10124 & n28876 ) ;
  assign n28878 = ( n10095 & n22137 ) | ( n10095 & ~n28877 ) | ( n22137 & ~n28877 ) ;
  assign n28879 = n6959 | n28878 ;
  assign n28880 = n28875 & ~n28879 ;
  assign n28881 = ( n13136 & n15793 ) | ( n13136 & ~n25489 ) | ( n15793 & ~n25489 ) ;
  assign n28882 = ( n3340 & n22064 ) | ( n3340 & ~n28151 ) | ( n22064 & ~n28151 ) ;
  assign n28883 = ~n3281 & n27467 ;
  assign n28884 = ( n4338 & ~n26492 ) | ( n4338 & n28883 ) | ( ~n26492 & n28883 ) ;
  assign n28885 = n14904 ^ n4589 ^ 1'b0 ;
  assign n28886 = n13478 & ~n28885 ;
  assign n28887 = ( ~n10390 & n10817 ) | ( ~n10390 & n25381 ) | ( n10817 & n25381 ) ;
  assign n28888 = ( ~n12816 & n12833 ) | ( ~n12816 & n28887 ) | ( n12833 & n28887 ) ;
  assign n28889 = ( n3261 & n28886 ) | ( n3261 & ~n28888 ) | ( n28886 & ~n28888 ) ;
  assign n28890 = ( ~n5625 & n13215 ) | ( ~n5625 & n21580 ) | ( n13215 & n21580 ) ;
  assign n28891 = n28890 ^ n22113 ^ n9229 ;
  assign n28892 = n16714 ^ n1140 ^ 1'b0 ;
  assign n28893 = ( ~n9451 & n14952 ) | ( ~n9451 & n28892 ) | ( n14952 & n28892 ) ;
  assign n28894 = n28893 ^ n1679 ^ 1'b0 ;
  assign n28895 = n16726 ^ n10957 ^ n3432 ;
  assign n28896 = n28895 ^ n27952 ^ n3997 ;
  assign n28897 = ( n3975 & ~n10412 ) | ( n3975 & n13986 ) | ( ~n10412 & n13986 ) ;
  assign n28898 = n22893 ^ n19623 ^ 1'b0 ;
  assign n28899 = n18702 & n28898 ;
  assign n28902 = ( n4155 & n4602 ) | ( n4155 & n7981 ) | ( n4602 & n7981 ) ;
  assign n28903 = n28902 ^ n24122 ^ n4134 ;
  assign n28900 = n16486 ^ n14449 ^ n9204 ;
  assign n28901 = n13151 | n28900 ;
  assign n28904 = n28903 ^ n28901 ^ 1'b0 ;
  assign n28905 = ( n767 & ~n13325 ) | ( n767 & n25302 ) | ( ~n13325 & n25302 ) ;
  assign n28906 = ( ~n2877 & n7248 ) | ( ~n2877 & n16861 ) | ( n7248 & n16861 ) ;
  assign n28907 = ( ~n3351 & n6640 ) | ( ~n3351 & n13686 ) | ( n6640 & n13686 ) ;
  assign n28908 = ( n6493 & n14609 ) | ( n6493 & n18378 ) | ( n14609 & n18378 ) ;
  assign n28909 = ( n13311 & n28907 ) | ( n13311 & n28908 ) | ( n28907 & n28908 ) ;
  assign n28910 = n9934 ^ n3929 ^ n183 ;
  assign n28911 = n28910 ^ n19641 ^ n18931 ;
  assign n28912 = n28121 ^ n3158 ^ n2885 ;
  assign n28913 = n28912 ^ n22625 ^ n17326 ;
  assign n28914 = n28913 ^ n2375 ^ 1'b0 ;
  assign n28915 = n5313 | n28914 ;
  assign n28916 = n28915 ^ n15959 ^ n3652 ;
  assign n28917 = n16210 ^ n6880 ^ 1'b0 ;
  assign n28918 = ( ~n13918 & n15804 ) | ( ~n13918 & n22859 ) | ( n15804 & n22859 ) ;
  assign n28919 = n15060 ^ n10303 ^ n4447 ;
  assign n28920 = ( n853 & ~n3772 ) | ( n853 & n25905 ) | ( ~n3772 & n25905 ) ;
  assign n28921 = ( n5987 & ~n26578 ) | ( n5987 & n28920 ) | ( ~n26578 & n28920 ) ;
  assign n28922 = n5092 & ~n28921 ;
  assign n28923 = n14153 ^ n8301 ^ n7194 ;
  assign n28924 = ( n7315 & n14388 ) | ( n7315 & ~n28923 ) | ( n14388 & ~n28923 ) ;
  assign n28925 = n11503 ^ n8162 ^ n965 ;
  assign n28926 = n18828 & ~n28925 ;
  assign n28927 = ~n28924 & n28926 ;
  assign n28928 = n15557 ^ n11139 ^ n3226 ;
  assign n28929 = ( n15631 & ~n23862 ) | ( n15631 & n28928 ) | ( ~n23862 & n28928 ) ;
  assign n28930 = ~n4828 & n28929 ;
  assign n28931 = ~n25864 & n28930 ;
  assign n28932 = n22035 ^ n5442 ^ n1126 ;
  assign n28933 = n28932 ^ n23560 ^ n14993 ;
  assign n28934 = n17218 ^ n15286 ^ n11489 ;
  assign n28935 = n28934 ^ n16349 ^ n312 ;
  assign n28936 = ( n4252 & ~n20337 ) | ( n4252 & n28935 ) | ( ~n20337 & n28935 ) ;
  assign n28937 = ( ~n539 & n5482 ) | ( ~n539 & n24707 ) | ( n5482 & n24707 ) ;
  assign n28938 = n28937 ^ n16911 ^ n6282 ;
  assign n28939 = ( n734 & n9036 ) | ( n734 & n17778 ) | ( n9036 & n17778 ) ;
  assign n28940 = ( n15347 & ~n24813 ) | ( n15347 & n28939 ) | ( ~n24813 & n28939 ) ;
  assign n28941 = n28940 ^ n7217 ^ n1719 ;
  assign n28942 = n23195 ^ n7903 ^ n7512 ;
  assign n28943 = ( n8430 & n20240 ) | ( n8430 & ~n20353 ) | ( n20240 & ~n20353 ) ;
  assign n28947 = n1377 | n5014 ;
  assign n28944 = n10569 ^ n3574 ^ n293 ;
  assign n28945 = n28944 ^ n20163 ^ n14995 ;
  assign n28946 = ( n11454 & ~n14661 ) | ( n11454 & n28945 ) | ( ~n14661 & n28945 ) ;
  assign n28948 = n28947 ^ n28946 ^ n8393 ;
  assign n28949 = ( n11064 & n22520 ) | ( n11064 & ~n22708 ) | ( n22520 & ~n22708 ) ;
  assign n28950 = ~n1403 & n8617 ;
  assign n28951 = n3907 & n28950 ;
  assign n28952 = n9114 ^ n8491 ^ 1'b0 ;
  assign n28953 = n3898 | n28952 ;
  assign n28954 = n28953 ^ n16118 ^ n1354 ;
  assign n28955 = ( ~n3865 & n12893 ) | ( ~n3865 & n28954 ) | ( n12893 & n28954 ) ;
  assign n28956 = n28955 ^ n15246 ^ n753 ;
  assign n28957 = n19253 ^ n8749 ^ 1'b0 ;
  assign n28958 = ( ~n721 & n14421 ) | ( ~n721 & n28957 ) | ( n14421 & n28957 ) ;
  assign n28959 = ( n1852 & ~n7033 ) | ( n1852 & n28958 ) | ( ~n7033 & n28958 ) ;
  assign n28960 = n28959 ^ n28849 ^ n20027 ;
  assign n28969 = ( n2527 & n5603 ) | ( n2527 & ~n8138 ) | ( n5603 & ~n8138 ) ;
  assign n28970 = n28969 ^ n16535 ^ n8099 ;
  assign n28971 = n28970 ^ n16429 ^ n2046 ;
  assign n28966 = n19283 ^ n9728 ^ n2839 ;
  assign n28967 = n28966 ^ n19575 ^ n13710 ;
  assign n28968 = ( n7756 & ~n21054 ) | ( n7756 & n28967 ) | ( ~n21054 & n28967 ) ;
  assign n28961 = ( ~n2591 & n20343 ) | ( ~n2591 & n22998 ) | ( n20343 & n22998 ) ;
  assign n28962 = n28961 ^ n2775 ^ 1'b0 ;
  assign n28963 = n28962 ^ n5002 ^ 1'b0 ;
  assign n28964 = n25987 & n28963 ;
  assign n28965 = n28964 ^ n18492 ^ 1'b0 ;
  assign n28972 = n28971 ^ n28968 ^ n28965 ;
  assign n28973 = n9364 ^ n1674 ^ 1'b0 ;
  assign n28974 = n19489 ^ n6175 ^ 1'b0 ;
  assign n28975 = n6050 & n28974 ;
  assign n28976 = n9005 ^ n8259 ^ n2367 ;
  assign n28977 = ( n6616 & ~n28975 ) | ( n6616 & n28976 ) | ( ~n28975 & n28976 ) ;
  assign n28978 = n21055 ^ n12371 ^ n1315 ;
  assign n28979 = n26736 ^ n21461 ^ n2803 ;
  assign n28980 = ( n2410 & n15232 ) | ( n2410 & n17895 ) | ( n15232 & n17895 ) ;
  assign n28981 = ( n4657 & n18432 ) | ( n4657 & n28980 ) | ( n18432 & n28980 ) ;
  assign n28982 = ~n20575 & n26874 ;
  assign n28983 = n28982 ^ n7721 ^ 1'b0 ;
  assign n28984 = ( n2188 & ~n2243 ) | ( n2188 & n5194 ) | ( ~n2243 & n5194 ) ;
  assign n28985 = n28984 ^ n28656 ^ 1'b0 ;
  assign n28986 = ( ~n15752 & n23665 ) | ( ~n15752 & n28985 ) | ( n23665 & n28985 ) ;
  assign n28987 = n27324 ^ n19250 ^ n10159 ;
  assign n28988 = ( n2549 & n5322 ) | ( n2549 & ~n12154 ) | ( n5322 & ~n12154 ) ;
  assign n28989 = n28988 ^ n28100 ^ n24440 ;
  assign n28990 = n22430 ^ n15153 ^ n1461 ;
  assign n28991 = n28990 ^ n21489 ^ n9167 ;
  assign n28992 = n21985 ^ n2686 ^ n282 ;
  assign n28993 = ( n3074 & n11880 ) | ( n3074 & n28992 ) | ( n11880 & n28992 ) ;
  assign n28994 = ( x67 & n24607 ) | ( x67 & n28993 ) | ( n24607 & n28993 ) ;
  assign n28995 = n28994 ^ n24959 ^ n22939 ;
  assign n28996 = n17400 ^ n12256 ^ n4447 ;
  assign n28997 = n28996 ^ n19361 ^ 1'b0 ;
  assign n28998 = n25302 ^ n9999 ^ n7051 ;
  assign n28999 = n17065 ^ n4483 ^ 1'b0 ;
  assign n29000 = n10104 & n28999 ;
  assign n29001 = ( ~n13808 & n28998 ) | ( ~n13808 & n29000 ) | ( n28998 & n29000 ) ;
  assign n29002 = ( ~n14013 & n17296 ) | ( ~n14013 & n22721 ) | ( n17296 & n22721 ) ;
  assign n29003 = n20229 ^ n17252 ^ n11306 ;
  assign n29004 = ~n12426 & n19817 ;
  assign n29005 = ( n14718 & ~n15636 ) | ( n14718 & n28053 ) | ( ~n15636 & n28053 ) ;
  assign n29006 = n18967 ^ n13836 ^ n11454 ;
  assign n29007 = ( n1942 & n12365 ) | ( n1942 & ~n21074 ) | ( n12365 & ~n21074 ) ;
  assign n29008 = n21793 ^ n19338 ^ n9816 ;
  assign n29009 = n29008 ^ n16352 ^ n8408 ;
  assign n29011 = n210 | n12899 ;
  assign n29012 = n29011 ^ n12967 ^ n5757 ;
  assign n29010 = ( n746 & n2425 ) | ( n746 & ~n28290 ) | ( n2425 & ~n28290 ) ;
  assign n29013 = n29012 ^ n29010 ^ n14931 ;
  assign n29014 = n7129 ^ n6812 ^ n2373 ;
  assign n29015 = ( n8609 & ~n10613 ) | ( n8609 & n10968 ) | ( ~n10613 & n10968 ) ;
  assign n29017 = n4137 ^ n230 ^ 1'b0 ;
  assign n29016 = n26670 ^ n21917 ^ n6422 ;
  assign n29018 = n29017 ^ n29016 ^ n28939 ;
  assign n29019 = n15466 ^ n6038 ^ 1'b0 ;
  assign n29020 = ( n277 & n3203 ) | ( n277 & n12935 ) | ( n3203 & n12935 ) ;
  assign n29021 = n23610 ^ n4612 ^ n3628 ;
  assign n29022 = n2236 | n29021 ;
  assign n29023 = ( ~n1739 & n12643 ) | ( ~n1739 & n29022 ) | ( n12643 & n29022 ) ;
  assign n29024 = ( n12264 & ~n15151 ) | ( n12264 & n23570 ) | ( ~n15151 & n23570 ) ;
  assign n29025 = n29024 ^ n16470 ^ n13514 ;
  assign n29026 = ( n21984 & n29023 ) | ( n21984 & n29025 ) | ( n29023 & n29025 ) ;
  assign n29027 = n4358 & n29026 ;
  assign n29028 = ~n29020 & n29027 ;
  assign n29029 = n1328 & ~n2466 ;
  assign n29030 = n29029 ^ n19770 ^ n1207 ;
  assign n29031 = ( n642 & n1589 ) | ( n642 & ~n22649 ) | ( n1589 & ~n22649 ) ;
  assign n29032 = n29031 ^ n23024 ^ n20214 ;
  assign n29033 = n18169 ^ n9603 ^ n5452 ;
  assign n29034 = ( n8864 & n12626 ) | ( n8864 & ~n16923 ) | ( n12626 & ~n16923 ) ;
  assign n29036 = n17101 ^ n7622 ^ 1'b0 ;
  assign n29037 = ~n2048 & n29036 ;
  assign n29035 = n14464 ^ n14009 ^ n11909 ;
  assign n29038 = n29037 ^ n29035 ^ n12255 ;
  assign n29039 = ( n1845 & n29034 ) | ( n1845 & ~n29038 ) | ( n29034 & ~n29038 ) ;
  assign n29040 = ( n5771 & n15530 ) | ( n5771 & n21820 ) | ( n15530 & n21820 ) ;
  assign n29041 = n29040 ^ n28044 ^ n16066 ;
  assign n29042 = n18578 ^ n13590 ^ 1'b0 ;
  assign n29043 = n27678 ^ n18619 ^ 1'b0 ;
  assign n29044 = ( n5556 & n20872 ) | ( n5556 & ~n24494 ) | ( n20872 & ~n24494 ) ;
  assign n29045 = ( n7688 & n13523 ) | ( n7688 & ~n13804 ) | ( n13523 & ~n13804 ) ;
  assign n29046 = n2203 | n8533 ;
  assign n29047 = n3342 | n7119 ;
  assign n29048 = n10928 | n29047 ;
  assign n29049 = ( n4559 & ~n18581 ) | ( n4559 & n20061 ) | ( ~n18581 & n20061 ) ;
  assign n29050 = ( n11216 & n24848 ) | ( n11216 & ~n29049 ) | ( n24848 & ~n29049 ) ;
  assign n29051 = n29050 ^ n12396 ^ n5266 ;
  assign n29052 = n2111 | n9355 ;
  assign n29053 = n10060 | n29052 ;
  assign n29054 = n29053 ^ n19603 ^ n17760 ;
  assign n29055 = n26694 ^ n16905 ^ n10898 ;
  assign n29056 = n29055 ^ n26191 ^ 1'b0 ;
  assign n29057 = ( n2691 & n7263 ) | ( n2691 & n9855 ) | ( n7263 & n9855 ) ;
  assign n29058 = ( n8410 & ~n17459 ) | ( n8410 & n29057 ) | ( ~n17459 & n29057 ) ;
  assign n29059 = n12070 ^ n10166 ^ n2352 ;
  assign n29060 = n29059 ^ n24975 ^ n17815 ;
  assign n29061 = ( ~n15437 & n18729 ) | ( ~n15437 & n22350 ) | ( n18729 & n22350 ) ;
  assign n29062 = ( n284 & ~n3154 ) | ( n284 & n7661 ) | ( ~n3154 & n7661 ) ;
  assign n29063 = ( ~n1960 & n3094 ) | ( ~n1960 & n29062 ) | ( n3094 & n29062 ) ;
  assign n29064 = n7498 & n10890 ;
  assign n29065 = n19040 & n29064 ;
  assign n29066 = n22798 ^ n17605 ^ n5410 ;
  assign n29067 = ( n22548 & n29065 ) | ( n22548 & n29066 ) | ( n29065 & n29066 ) ;
  assign n29068 = n29067 ^ n13331 ^ n4285 ;
  assign n29070 = ( ~x5 & n2450 ) | ( ~x5 & n8341 ) | ( n2450 & n8341 ) ;
  assign n29069 = n19481 ^ n1681 ^ 1'b0 ;
  assign n29071 = n29070 ^ n29069 ^ n6300 ;
  assign n29072 = n29071 ^ n18883 ^ n12006 ;
  assign n29073 = ( n16576 & n21540 ) | ( n16576 & ~n29072 ) | ( n21540 & ~n29072 ) ;
  assign n29074 = n11467 | n28664 ;
  assign n29075 = n15458 ^ n3825 ^ 1'b0 ;
  assign n29076 = n29074 & n29075 ;
  assign n29077 = ( n4842 & ~n10398 ) | ( n4842 & n15451 ) | ( ~n10398 & n15451 ) ;
  assign n29078 = n12154 ^ n9249 ^ n5470 ;
  assign n29079 = ~n8416 & n29078 ;
  assign n29080 = ( n14643 & n15666 ) | ( n14643 & ~n29079 ) | ( n15666 & ~n29079 ) ;
  assign n29081 = n19826 ^ n10177 ^ 1'b0 ;
  assign n29082 = n29081 ^ n6624 ^ n6251 ;
  assign n29086 = n27052 ^ n20599 ^ 1'b0 ;
  assign n29085 = n16448 ^ n7309 ^ n414 ;
  assign n29083 = n6300 & n14445 ;
  assign n29084 = n29083 ^ n21980 ^ 1'b0 ;
  assign n29087 = n29086 ^ n29085 ^ n29084 ;
  assign n29088 = n12957 | n14198 ;
  assign n29089 = n9279 ^ n1422 ^ x16 ;
  assign n29090 = n14038 ^ n801 ^ x107 ;
  assign n29091 = ( ~n7408 & n12965 ) | ( ~n7408 & n29090 ) | ( n12965 & n29090 ) ;
  assign n29092 = ( ~n15076 & n17481 ) | ( ~n15076 & n18139 ) | ( n17481 & n18139 ) ;
  assign n29093 = ( n1569 & n4895 ) | ( n1569 & n16686 ) | ( n4895 & n16686 ) ;
  assign n29094 = n15966 ^ n15584 ^ 1'b0 ;
  assign n29095 = n7069 | n29094 ;
  assign n29096 = ( ~n20345 & n26929 ) | ( ~n20345 & n29095 ) | ( n26929 & n29095 ) ;
  assign n29097 = n29096 ^ n8577 ^ n5619 ;
  assign n29098 = ( ~n450 & n4234 ) | ( ~n450 & n4245 ) | ( n4234 & n4245 ) ;
  assign n29099 = n27568 ^ n12803 ^ n7423 ;
  assign n29100 = ( ~n17991 & n29098 ) | ( ~n17991 & n29099 ) | ( n29098 & n29099 ) ;
  assign n29101 = ( n8268 & ~n8889 ) | ( n8268 & n11157 ) | ( ~n8889 & n11157 ) ;
  assign n29102 = n10645 ^ n9837 ^ n3673 ;
  assign n29103 = ( n13730 & n14384 ) | ( n13730 & ~n29040 ) | ( n14384 & ~n29040 ) ;
  assign n29104 = n10089 ^ n6229 ^ n3909 ;
  assign n29105 = n6785 | n9140 ;
  assign n29106 = n1770 & ~n29105 ;
  assign n29107 = ( ~n12058 & n16529 ) | ( ~n12058 & n29106 ) | ( n16529 & n29106 ) ;
  assign n29108 = ( ~n5239 & n29104 ) | ( ~n5239 & n29107 ) | ( n29104 & n29107 ) ;
  assign n29109 = ( n7749 & n21493 ) | ( n7749 & n29108 ) | ( n21493 & n29108 ) ;
  assign n29110 = n18280 ^ n736 ^ 1'b0 ;
  assign n29111 = n29110 ^ n7157 ^ n2257 ;
  assign n29112 = n29111 ^ n26853 ^ n932 ;
  assign n29113 = n20441 ^ n4959 ^ 1'b0 ;
  assign n29114 = n25896 & n29113 ;
  assign n29115 = n16101 & ~n27709 ;
  assign n29116 = ( ~n16212 & n24217 ) | ( ~n16212 & n29115 ) | ( n24217 & n29115 ) ;
  assign n29117 = ( n26240 & n29114 ) | ( n26240 & n29116 ) | ( n29114 & n29116 ) ;
  assign n29118 = n29117 ^ n27280 ^ 1'b0 ;
  assign n29119 = n8657 & ~n9143 ;
  assign n29120 = n29119 ^ n1775 ^ 1'b0 ;
  assign n29121 = n8071 & ~n9028 ;
  assign n29122 = n14806 ^ n6987 ^ n6021 ;
  assign n29123 = n4314 & ~n29122 ;
  assign n29124 = n29121 & n29123 ;
  assign n29125 = ( n13650 & n16775 ) | ( n13650 & n29124 ) | ( n16775 & n29124 ) ;
  assign n29126 = ~n3860 & n21198 ;
  assign n29127 = ~n29125 & n29126 ;
  assign n29128 = x81 & ~n25429 ;
  assign n29129 = n29128 ^ n17286 ^ 1'b0 ;
  assign n29130 = ( n19071 & n22774 ) | ( n19071 & ~n29129 ) | ( n22774 & ~n29129 ) ;
  assign n29131 = ( n5139 & n9973 ) | ( n5139 & ~n19964 ) | ( n9973 & ~n19964 ) ;
  assign n29133 = n26557 ^ n9924 ^ n4972 ;
  assign n29132 = ( n1429 & ~n2516 ) | ( n1429 & n17214 ) | ( ~n2516 & n17214 ) ;
  assign n29134 = n29133 ^ n29132 ^ n27952 ;
  assign n29135 = n24686 ^ n19865 ^ n1718 ;
  assign n29136 = n25593 ^ n23033 ^ 1'b0 ;
  assign n29137 = n20315 ^ n3602 ^ n1977 ;
  assign n29138 = n29137 ^ n22903 ^ n3931 ;
  assign n29139 = n23046 ^ n18191 ^ n16529 ;
  assign n29140 = n29139 ^ n1403 ^ 1'b0 ;
  assign n29141 = n28290 ^ n14905 ^ n12039 ;
  assign n29142 = n20667 ^ n13776 ^ 1'b0 ;
  assign n29143 = n14211 & ~n29034 ;
  assign n29144 = n29143 ^ n28118 ^ 1'b0 ;
  assign n29145 = n27693 ^ n13212 ^ 1'b0 ;
  assign n29146 = n25524 ^ n14209 ^ n4814 ;
  assign n29147 = ( n15684 & n19655 ) | ( n15684 & ~n25344 ) | ( n19655 & ~n25344 ) ;
  assign n29148 = n29147 ^ n21006 ^ n16747 ;
  assign n29149 = n29148 ^ n24893 ^ n18659 ;
  assign n29150 = n22580 ^ n14141 ^ n8381 ;
  assign n29151 = n29150 ^ n17850 ^ n1692 ;
  assign n29152 = n28435 ^ n24986 ^ 1'b0 ;
  assign n29153 = ( n1281 & n9686 ) | ( n1281 & n29152 ) | ( n9686 & n29152 ) ;
  assign n29154 = n237 | n20711 ;
  assign n29155 = n19946 & ~n29154 ;
  assign n29156 = ( ~n5391 & n29153 ) | ( ~n5391 & n29155 ) | ( n29153 & n29155 ) ;
  assign n29157 = ( ~n7195 & n27530 ) | ( ~n7195 & n28174 ) | ( n27530 & n28174 ) ;
  assign n29158 = ( ~n6440 & n27159 ) | ( ~n6440 & n29157 ) | ( n27159 & n29157 ) ;
  assign n29159 = n4758 | n11835 ;
  assign n29160 = n29159 ^ n10569 ^ 1'b0 ;
  assign n29161 = ( n3372 & n6449 ) | ( n3372 & n29160 ) | ( n6449 & n29160 ) ;
  assign n29162 = n29161 ^ n28658 ^ 1'b0 ;
  assign n29163 = ( n5484 & ~n12419 ) | ( n5484 & n21555 ) | ( ~n12419 & n21555 ) ;
  assign n29164 = n3428 & n14542 ;
  assign n29165 = n8985 & n29164 ;
  assign n29166 = n29165 ^ n8584 ^ 1'b0 ;
  assign n29167 = n22861 ^ n7907 ^ 1'b0 ;
  assign n29168 = n26399 & ~n29167 ;
  assign n29169 = n11017 ^ n10783 ^ n6551 ;
  assign n29170 = ( ~n868 & n1998 ) | ( ~n868 & n21821 ) | ( n1998 & n21821 ) ;
  assign n29171 = ( n6665 & n20305 ) | ( n6665 & n29170 ) | ( n20305 & n29170 ) ;
  assign n29174 = n11099 | n16581 ;
  assign n29175 = n25695 & ~n29174 ;
  assign n29173 = ( n11385 & n13679 ) | ( n11385 & n16650 ) | ( n13679 & n16650 ) ;
  assign n29172 = n17432 ^ n11882 ^ n2721 ;
  assign n29176 = n29175 ^ n29173 ^ n29172 ;
  assign n29177 = ( ~n551 & n9261 ) | ( ~n551 & n29176 ) | ( n9261 & n29176 ) ;
  assign n29178 = x54 & n27792 ;
  assign n29179 = n29178 ^ n24678 ^ n8520 ;
  assign n29180 = n29179 ^ n16199 ^ n572 ;
  assign n29181 = ( n8693 & ~n12011 ) | ( n8693 & n13235 ) | ( ~n12011 & n13235 ) ;
  assign n29182 = ( n3984 & n20605 ) | ( n3984 & n22713 ) | ( n20605 & n22713 ) ;
  assign n29183 = n16805 ^ n6361 ^ n3802 ;
  assign n29184 = n29183 ^ n18857 ^ n13800 ;
  assign n29185 = n23189 ^ n11080 ^ n9662 ;
  assign n29186 = ( n9623 & n10828 ) | ( n9623 & ~n29185 ) | ( n10828 & ~n29185 ) ;
  assign n29187 = n29186 ^ n25724 ^ n2686 ;
  assign n29192 = ( n4770 & n12393 ) | ( n4770 & ~n16049 ) | ( n12393 & ~n16049 ) ;
  assign n29193 = ( n936 & n2590 ) | ( n936 & n29192 ) | ( n2590 & n29192 ) ;
  assign n29194 = n1462 | n6177 ;
  assign n29195 = n29194 ^ n9503 ^ 1'b0 ;
  assign n29196 = n29193 & ~n29195 ;
  assign n29191 = n13836 ^ n7229 ^ n1048 ;
  assign n29197 = n29196 ^ n29191 ^ n19855 ;
  assign n29188 = ( ~n3826 & n4343 ) | ( ~n3826 & n5622 ) | ( n4343 & n5622 ) ;
  assign n29189 = n29188 ^ n14723 ^ n11723 ;
  assign n29190 = ~n13204 & n29189 ;
  assign n29198 = n29197 ^ n29190 ^ 1'b0 ;
  assign n29199 = n28162 ^ n26126 ^ n1507 ;
  assign n29200 = ( n7435 & n9237 ) | ( n7435 & ~n9319 ) | ( n9237 & ~n9319 ) ;
  assign n29201 = n29200 ^ n16045 ^ 1'b0 ;
  assign n29202 = ( n1331 & n10318 ) | ( n1331 & ~n18563 ) | ( n10318 & ~n18563 ) ;
  assign n29203 = n29202 ^ n23404 ^ n13491 ;
  assign n29204 = ( n28484 & n29201 ) | ( n28484 & n29203 ) | ( n29201 & n29203 ) ;
  assign n29206 = n18967 ^ n2063 ^ n572 ;
  assign n29207 = ( n7640 & n22654 ) | ( n7640 & ~n29206 ) | ( n22654 & ~n29206 ) ;
  assign n29208 = n13789 & n29207 ;
  assign n29205 = ( n11118 & n19381 ) | ( n11118 & ~n22818 ) | ( n19381 & ~n22818 ) ;
  assign n29209 = n29208 ^ n29205 ^ n29125 ;
  assign n29210 = n6422 | n20451 ;
  assign n29211 = n5466 ^ n5348 ^ n4888 ;
  assign n29212 = ( n28660 & n29210 ) | ( n28660 & ~n29211 ) | ( n29210 & ~n29211 ) ;
  assign n29213 = n468 | n15510 ;
  assign n29214 = n29213 ^ n14118 ^ n5367 ;
  assign n29215 = ( ~n2441 & n2893 ) | ( ~n2441 & n16374 ) | ( n2893 & n16374 ) ;
  assign n29216 = ( n2478 & n10442 ) | ( n2478 & n12084 ) | ( n10442 & n12084 ) ;
  assign n29217 = n196 & n25861 ;
  assign n29218 = ~n3716 & n29217 ;
  assign n29219 = n29216 | n29218 ;
  assign n29220 = ( ~n2632 & n19351 ) | ( ~n2632 & n22683 ) | ( n19351 & n22683 ) ;
  assign n29221 = n10688 ^ n3007 ^ 1'b0 ;
  assign n29222 = ~n11364 & n29221 ;
  assign n29223 = n4433 & n24848 ;
  assign n29224 = n29223 ^ n1768 ^ 1'b0 ;
  assign n29225 = ~n4499 & n8998 ;
  assign n29226 = ( ~n10112 & n15640 ) | ( ~n10112 & n29225 ) | ( n15640 & n29225 ) ;
  assign n29227 = n29226 ^ n4077 ^ n1366 ;
  assign n29228 = ( n12168 & n21491 ) | ( n12168 & n29227 ) | ( n21491 & n29227 ) ;
  assign n29229 = n8771 & ~n22190 ;
  assign n29230 = n29229 ^ n21216 ^ n17484 ;
  assign n29231 = ( n10331 & n11707 ) | ( n10331 & ~n13695 ) | ( n11707 & ~n13695 ) ;
  assign n29232 = n29231 ^ n8932 ^ n5331 ;
  assign n29233 = n13782 | n27694 ;
  assign n29234 = n21836 & ~n29233 ;
  assign n29235 = ( n18924 & n21961 ) | ( n18924 & ~n29234 ) | ( n21961 & ~n29234 ) ;
  assign n29236 = ( n10395 & ~n16755 ) | ( n10395 & n18563 ) | ( ~n16755 & n18563 ) ;
  assign n29237 = ( n6539 & ~n9883 ) | ( n6539 & n12115 ) | ( ~n9883 & n12115 ) ;
  assign n29238 = ( ~n1715 & n1872 ) | ( ~n1715 & n25868 ) | ( n1872 & n25868 ) ;
  assign n29239 = x83 & n5716 ;
  assign n29240 = ~n345 & n29239 ;
  assign n29241 = n29240 ^ n12480 ^ n455 ;
  assign n29242 = n29241 ^ n21017 ^ n670 ;
  assign n29243 = ( n13996 & ~n17047 ) | ( n13996 & n29242 ) | ( ~n17047 & n29242 ) ;
  assign n29244 = n5069 | n29243 ;
  assign n29245 = n29244 ^ n26352 ^ 1'b0 ;
  assign n29246 = n29238 & ~n29245 ;
  assign n29247 = n29246 ^ n5353 ^ 1'b0 ;
  assign n29248 = n24312 ^ n11099 ^ 1'b0 ;
  assign n29249 = n8581 ^ n1988 ^ n715 ;
  assign n29250 = ( n8628 & n18572 ) | ( n8628 & ~n29249 ) | ( n18572 & ~n29249 ) ;
  assign n29251 = ( n404 & n799 ) | ( n404 & n29250 ) | ( n799 & n29250 ) ;
  assign n29255 = n3995 & n13077 ;
  assign n29256 = n20043 & n29255 ;
  assign n29252 = n22213 ^ n10569 ^ n346 ;
  assign n29253 = n29252 ^ n9107 ^ n4707 ;
  assign n29254 = ( n456 & ~n21774 ) | ( n456 & n29253 ) | ( ~n21774 & n29253 ) ;
  assign n29257 = n29256 ^ n29254 ^ n4136 ;
  assign n29260 = n23119 ^ n18677 ^ n11135 ;
  assign n29261 = n29260 ^ n5576 ^ n5277 ;
  assign n29262 = ( n3500 & n12674 ) | ( n3500 & ~n29261 ) | ( n12674 & ~n29261 ) ;
  assign n29258 = ~n4270 & n10660 ;
  assign n29259 = n6828 & n29258 ;
  assign n29263 = n29262 ^ n29259 ^ n15311 ;
  assign n29264 = n6835 & ~n11983 ;
  assign n29265 = n29264 ^ n10546 ^ 1'b0 ;
  assign n29266 = n4106 ^ n3976 ^ n178 ;
  assign n29267 = ( n4859 & n20413 ) | ( n4859 & ~n29266 ) | ( n20413 & ~n29266 ) ;
  assign n29268 = n24676 ^ n13532 ^ n5349 ;
  assign n29269 = ( n8386 & n20609 ) | ( n8386 & ~n29268 ) | ( n20609 & ~n29268 ) ;
  assign n29270 = n16732 ^ n13653 ^ n10236 ;
  assign n29271 = ~n3437 & n29270 ;
  assign n29272 = ~n17962 & n29271 ;
  assign n29273 = n29272 ^ n20926 ^ n8479 ;
  assign n29274 = ( ~n1371 & n12296 ) | ( ~n1371 & n17617 ) | ( n12296 & n17617 ) ;
  assign n29275 = n12412 ^ n9256 ^ n3614 ;
  assign n29276 = n29275 ^ n3481 ^ 1'b0 ;
  assign n29277 = n29276 ^ n15031 ^ n9034 ;
  assign n29278 = ( n3582 & ~n24734 ) | ( n3582 & n29277 ) | ( ~n24734 & n29277 ) ;
  assign n29279 = ( n7642 & n10468 ) | ( n7642 & ~n15592 ) | ( n10468 & ~n15592 ) ;
  assign n29290 = ( n1554 & ~n13967 ) | ( n1554 & n14446 ) | ( ~n13967 & n14446 ) ;
  assign n29288 = n7263 & ~n27366 ;
  assign n29285 = n13143 ^ n10397 ^ n8280 ;
  assign n29286 = n26976 ^ n6300 ^ 1'b0 ;
  assign n29287 = n29285 & ~n29286 ;
  assign n29289 = n29288 ^ n29287 ^ n9936 ;
  assign n29280 = ( n7611 & ~n8478 ) | ( n7611 & n15087 ) | ( ~n8478 & n15087 ) ;
  assign n29281 = n29280 ^ n11325 ^ 1'b0 ;
  assign n29282 = ( n14323 & ~n15724 ) | ( n14323 & n29281 ) | ( ~n15724 & n29281 ) ;
  assign n29283 = ( ~n9222 & n28841 ) | ( ~n9222 & n29282 ) | ( n28841 & n29282 ) ;
  assign n29284 = n29283 ^ n296 ^ 1'b0 ;
  assign n29291 = n29290 ^ n29289 ^ n29284 ;
  assign n29292 = n5091 ^ n2852 ^ n526 ;
  assign n29293 = n29292 ^ n23193 ^ n15801 ;
  assign n29297 = ( ~n782 & n21837 ) | ( ~n782 & n26071 ) | ( n21837 & n26071 ) ;
  assign n29294 = ( n1080 & n7301 ) | ( n1080 & n14384 ) | ( n7301 & n14384 ) ;
  assign n29295 = ~n3460 & n29294 ;
  assign n29296 = ~n20020 & n29295 ;
  assign n29298 = n29297 ^ n29296 ^ n6440 ;
  assign n29299 = ~n14953 & n16943 ;
  assign n29300 = n29299 ^ n24773 ^ 1'b0 ;
  assign n29301 = ( n7794 & n28696 ) | ( n7794 & ~n29300 ) | ( n28696 & ~n29300 ) ;
  assign n29302 = ( n2669 & n22738 ) | ( n2669 & n29301 ) | ( n22738 & n29301 ) ;
  assign n29303 = ( ~n17233 & n28537 ) | ( ~n17233 & n29302 ) | ( n28537 & n29302 ) ;
  assign n29304 = ( n3997 & n10461 ) | ( n3997 & n19963 ) | ( n10461 & n19963 ) ;
  assign n29306 = n10281 ^ n6452 ^ n5296 ;
  assign n29305 = n27215 ^ n11466 ^ n7647 ;
  assign n29307 = n29306 ^ n29305 ^ n25190 ;
  assign n29308 = n29307 ^ n25873 ^ n23787 ;
  assign n29309 = n26692 ^ n7848 ^ n4364 ;
  assign n29310 = n29309 ^ n25528 ^ n24462 ;
  assign n29311 = n5303 & ~n25161 ;
  assign n29312 = n27723 ^ n1240 ^ 1'b0 ;
  assign n29313 = n25190 & n29312 ;
  assign n29314 = ( n14137 & n29311 ) | ( n14137 & ~n29313 ) | ( n29311 & ~n29313 ) ;
  assign n29315 = n384 & n24344 ;
  assign n29316 = ~n28541 & n29315 ;
  assign n29317 = n14711 | n24962 ;
  assign n29318 = ( n15755 & n22578 ) | ( n15755 & n29011 ) | ( n22578 & n29011 ) ;
  assign n29319 = ( n8182 & n10695 ) | ( n8182 & ~n29318 ) | ( n10695 & ~n29318 ) ;
  assign n29320 = ( ~n1507 & n3562 ) | ( ~n1507 & n6822 ) | ( n3562 & n6822 ) ;
  assign n29321 = n29320 ^ n18911 ^ n7893 ;
  assign n29322 = ( n16442 & ~n19016 ) | ( n16442 & n21183 ) | ( ~n19016 & n21183 ) ;
  assign n29323 = ( n471 & n3665 ) | ( n471 & n11624 ) | ( n3665 & n11624 ) ;
  assign n29324 = ( n8225 & n8539 ) | ( n8225 & ~n14030 ) | ( n8539 & ~n14030 ) ;
  assign n29325 = ( ~n812 & n5885 ) | ( ~n812 & n29324 ) | ( n5885 & n29324 ) ;
  assign n29326 = ( n5439 & n29323 ) | ( n5439 & ~n29325 ) | ( n29323 & ~n29325 ) ;
  assign n29327 = n24746 ^ n20890 ^ n16298 ;
  assign n29328 = n29327 ^ n22546 ^ n4367 ;
  assign n29329 = ( n4708 & n13965 ) | ( n4708 & n21091 ) | ( n13965 & n21091 ) ;
  assign n29330 = n7206 & ~n10642 ;
  assign n29331 = n3647 & n29330 ;
  assign n29332 = ( n2029 & n7229 ) | ( n2029 & ~n29331 ) | ( n7229 & ~n29331 ) ;
  assign n29333 = n29332 ^ n3248 ^ 1'b0 ;
  assign n29334 = n8232 ^ n3514 ^ n1297 ;
  assign n29335 = ( n9701 & ~n28661 ) | ( n9701 & n29334 ) | ( ~n28661 & n29334 ) ;
  assign n29336 = n20924 ^ n4446 ^ 1'b0 ;
  assign n29337 = ( n2388 & n4562 ) | ( n2388 & ~n16816 ) | ( n4562 & ~n16816 ) ;
  assign n29338 = ( n8536 & ~n10402 ) | ( n8536 & n14980 ) | ( ~n10402 & n14980 ) ;
  assign n29339 = n29338 ^ n28876 ^ n6931 ;
  assign n29340 = ( n11387 & ~n11672 ) | ( n11387 & n19495 ) | ( ~n11672 & n19495 ) ;
  assign n29341 = n29340 ^ n26845 ^ n3441 ;
  assign n29342 = n10773 ^ n7837 ^ n774 ;
  assign n29343 = ( n16288 & n21945 ) | ( n16288 & ~n29342 ) | ( n21945 & ~n29342 ) ;
  assign n29344 = n29343 ^ n3115 ^ n3054 ;
  assign n29345 = ( n16109 & n17403 ) | ( n16109 & ~n29344 ) | ( n17403 & ~n29344 ) ;
  assign n29346 = ( ~n1148 & n7055 ) | ( ~n1148 & n9486 ) | ( n7055 & n9486 ) ;
  assign n29347 = n29346 ^ n21041 ^ n510 ;
  assign n29348 = n3526 ^ n2259 ^ n839 ;
  assign n29349 = n29348 ^ n11511 ^ n8393 ;
  assign n29350 = n29349 ^ n16260 ^ 1'b0 ;
  assign n29351 = ~n3725 & n22968 ;
  assign n29352 = ~n20047 & n29351 ;
  assign n29353 = ( n5953 & n7686 ) | ( n5953 & ~n7870 ) | ( n7686 & ~n7870 ) ;
  assign n29354 = ( ~n2422 & n29352 ) | ( ~n2422 & n29353 ) | ( n29352 & n29353 ) ;
  assign n29355 = ( n8055 & n19759 ) | ( n8055 & ~n29354 ) | ( n19759 & ~n29354 ) ;
  assign n29356 = n29355 ^ n22659 ^ n15898 ;
  assign n29357 = n18605 ^ n8054 ^ 1'b0 ;
  assign n29358 = ~n6589 & n29357 ;
  assign n29359 = n1049 & n6922 ;
  assign n29360 = n29359 ^ n7559 ^ 1'b0 ;
  assign n29361 = ( ~x122 & n8161 ) | ( ~x122 & n12171 ) | ( n8161 & n12171 ) ;
  assign n29362 = n29361 ^ n19260 ^ n8920 ;
  assign n29363 = n24513 ^ n19737 ^ n19064 ;
  assign n29364 = n20916 ^ n18062 ^ n8567 ;
  assign n29365 = ( ~n4628 & n6621 ) | ( ~n4628 & n29364 ) | ( n6621 & n29364 ) ;
  assign n29373 = ( n3750 & n6216 ) | ( n3750 & ~n6484 ) | ( n6216 & ~n6484 ) ;
  assign n29374 = n29373 ^ n14290 ^ n1886 ;
  assign n29372 = n11584 & ~n16572 ;
  assign n29375 = n29374 ^ n29372 ^ 1'b0 ;
  assign n29367 = n16987 & ~n24130 ;
  assign n29368 = n29367 ^ n13976 ^ 1'b0 ;
  assign n29369 = n29368 ^ n20151 ^ n5407 ;
  assign n29370 = ( n4189 & ~n5722 ) | ( n4189 & n29369 ) | ( ~n5722 & n29369 ) ;
  assign n29366 = ( n9140 & n10583 ) | ( n9140 & ~n11396 ) | ( n10583 & ~n11396 ) ;
  assign n29371 = n29370 ^ n29366 ^ n21846 ;
  assign n29376 = n29375 ^ n29371 ^ n22750 ;
  assign n29381 = n6796 ^ n814 ^ 1'b0 ;
  assign n29377 = ~n7364 & n8642 ;
  assign n29378 = n29377 ^ n6738 ^ 1'b0 ;
  assign n29379 = ~n10897 & n23378 ;
  assign n29380 = n29378 & n29379 ;
  assign n29382 = n29381 ^ n29380 ^ n7865 ;
  assign n29383 = ( n17604 & ~n24979 ) | ( n17604 & n26209 ) | ( ~n24979 & n26209 ) ;
  assign n29385 = ( ~n1434 & n4859 ) | ( ~n1434 & n4984 ) | ( n4859 & n4984 ) ;
  assign n29384 = ( n6078 & n14762 ) | ( n6078 & ~n16547 ) | ( n14762 & ~n16547 ) ;
  assign n29386 = n29385 ^ n29384 ^ n9313 ;
  assign n29387 = n17151 ^ n16290 ^ n11004 ;
  assign n29388 = ( ~n8908 & n28964 ) | ( ~n8908 & n29387 ) | ( n28964 & n29387 ) ;
  assign n29389 = ( n2579 & ~n3043 ) | ( n2579 & n10788 ) | ( ~n3043 & n10788 ) ;
  assign n29390 = n29389 ^ n20744 ^ n8228 ;
  assign n29391 = n24002 | n24511 ;
  assign n29392 = n29390 & ~n29391 ;
  assign n29393 = ( n1286 & n1350 ) | ( n1286 & n2250 ) | ( n1350 & n2250 ) ;
  assign n29394 = ( n7727 & ~n27914 ) | ( n7727 & n29393 ) | ( ~n27914 & n29393 ) ;
  assign n29395 = n29394 ^ n8094 ^ 1'b0 ;
  assign n29396 = n20085 & n29395 ;
  assign n29397 = n27565 ^ n23367 ^ n16454 ;
  assign n29398 = ( n2619 & n27171 ) | ( n2619 & ~n29397 ) | ( n27171 & ~n29397 ) ;
  assign n29399 = n24123 ^ n8659 ^ n6160 ;
  assign n29400 = n14891 ^ n5830 ^ n5143 ;
  assign n29401 = ( n1927 & ~n3107 ) | ( n1927 & n29400 ) | ( ~n3107 & n29400 ) ;
  assign n29402 = ( n2360 & n3044 ) | ( n2360 & n11930 ) | ( n3044 & n11930 ) ;
  assign n29403 = n26649 & n29402 ;
  assign n29404 = ( n9038 & n13886 ) | ( n9038 & ~n24992 ) | ( n13886 & ~n24992 ) ;
  assign n29405 = n29404 ^ n27742 ^ n10310 ;
  assign n29406 = n12043 ^ n5628 ^ 1'b0 ;
  assign n29407 = n29406 ^ n12478 ^ n4015 ;
  assign n29408 = n18096 ^ n15034 ^ n5508 ;
  assign n29409 = ( n15407 & n29407 ) | ( n15407 & ~n29408 ) | ( n29407 & ~n29408 ) ;
  assign n29410 = ( n3793 & ~n9617 ) | ( n3793 & n13793 ) | ( ~n9617 & n13793 ) ;
  assign n29411 = n29410 ^ n29115 ^ n20224 ;
  assign n29412 = ( n523 & ~n2157 ) | ( n523 & n9657 ) | ( ~n2157 & n9657 ) ;
  assign n29413 = n29412 ^ n12206 ^ n8396 ;
  assign n29414 = n18066 ^ n7695 ^ n6799 ;
  assign n29415 = n29414 ^ n15434 ^ n1106 ;
  assign n29416 = ( ~n14130 & n20275 ) | ( ~n14130 & n23322 ) | ( n20275 & n23322 ) ;
  assign n29417 = n17972 ^ n10995 ^ 1'b0 ;
  assign n29418 = ~n29416 & n29417 ;
  assign n29419 = ( x59 & n3316 ) | ( x59 & n23207 ) | ( n3316 & n23207 ) ;
  assign n29420 = n13143 ^ n8585 ^ n3028 ;
  assign n29421 = n13119 | n29420 ;
  assign n29422 = n29419 | n29421 ;
  assign n29423 = ~n14358 & n25024 ;
  assign n29424 = n26400 & n29423 ;
  assign n29425 = ( ~n10778 & n23994 ) | ( ~n10778 & n29424 ) | ( n23994 & n29424 ) ;
  assign n29426 = n11411 ^ n7686 ^ n291 ;
  assign n29427 = ( n655 & ~n23070 ) | ( n655 & n29426 ) | ( ~n23070 & n29426 ) ;
  assign n29428 = ( ~n6984 & n16601 ) | ( ~n6984 & n29427 ) | ( n16601 & n29427 ) ;
  assign n29433 = n15024 ^ n7150 ^ n4376 ;
  assign n29434 = n29433 ^ n2652 ^ x91 ;
  assign n29432 = ( n7310 & ~n10393 ) | ( n7310 & n12640 ) | ( ~n10393 & n12640 ) ;
  assign n29435 = n29434 ^ n29432 ^ n8577 ;
  assign n29429 = ( n3496 & ~n9978 ) | ( n3496 & n14832 ) | ( ~n9978 & n14832 ) ;
  assign n29430 = n29429 ^ n12140 ^ n843 ;
  assign n29431 = ( n1134 & n28790 ) | ( n1134 & n29430 ) | ( n28790 & n29430 ) ;
  assign n29436 = n29435 ^ n29431 ^ n24308 ;
  assign n29437 = n5188 & n9069 ;
  assign n29438 = ~n1905 & n29437 ;
  assign n29439 = n2104 & ~n10174 ;
  assign n29440 = n9619 & n29439 ;
  assign n29441 = ( n19150 & n29438 ) | ( n19150 & ~n29440 ) | ( n29438 & ~n29440 ) ;
  assign n29442 = ( n7853 & n11272 ) | ( n7853 & ~n29441 ) | ( n11272 & ~n29441 ) ;
  assign n29443 = n29442 ^ n16836 ^ 1'b0 ;
  assign n29444 = n11155 | n24699 ;
  assign n29445 = ( n14347 & ~n24651 ) | ( n14347 & n29444 ) | ( ~n24651 & n29444 ) ;
  assign n29446 = ( n517 & ~n5762 ) | ( n517 & n9135 ) | ( ~n5762 & n9135 ) ;
  assign n29447 = ( n641 & n18407 ) | ( n641 & n29446 ) | ( n18407 & n29446 ) ;
  assign n29448 = n11689 ^ n1715 ^ n1241 ;
  assign n29449 = ~n6421 & n11291 ;
  assign n29450 = ~n17925 & n29449 ;
  assign n29451 = n29450 ^ n23996 ^ n20568 ;
  assign n29452 = n25864 ^ n6970 ^ n4398 ;
  assign n29453 = n29452 ^ n10784 ^ 1'b0 ;
  assign n29454 = n6173 & n29453 ;
  assign n29455 = n16001 & n24866 ;
  assign n29456 = n29455 ^ n860 ^ 1'b0 ;
  assign n29457 = ( ~n12968 & n21907 ) | ( ~n12968 & n26304 ) | ( n21907 & n26304 ) ;
  assign n29460 = ( n2840 & n5050 ) | ( n2840 & n13676 ) | ( n5050 & n13676 ) ;
  assign n29458 = ~n4167 & n4804 ;
  assign n29459 = ~n19288 & n29458 ;
  assign n29461 = n29460 ^ n29459 ^ n10952 ;
  assign n29462 = ( n282 & n10263 ) | ( n282 & ~n10664 ) | ( n10263 & ~n10664 ) ;
  assign n29463 = n29462 ^ n9121 ^ n7201 ;
  assign n29464 = n21804 ^ n19447 ^ n2510 ;
  assign n29465 = n29464 ^ n18270 ^ n12148 ;
  assign n29466 = n22081 ^ n12961 ^ n7639 ;
  assign n29467 = n29466 ^ n27153 ^ n2908 ;
  assign n29468 = n29467 ^ n2851 ^ n2141 ;
  assign n29469 = ( n6696 & ~n12840 ) | ( n6696 & n20253 ) | ( ~n12840 & n20253 ) ;
  assign n29470 = n7103 | n24490 ;
  assign n29471 = n11213 & ~n29470 ;
  assign n29472 = n22762 ^ n6081 ^ n408 ;
  assign n29474 = n28696 ^ n10360 ^ n9910 ;
  assign n29473 = ( n5674 & n6301 ) | ( n5674 & n22788 ) | ( n6301 & n22788 ) ;
  assign n29475 = n29474 ^ n29473 ^ n10844 ;
  assign n29476 = ( n526 & n9643 ) | ( n526 & ~n10262 ) | ( n9643 & ~n10262 ) ;
  assign n29477 = n29476 ^ n7862 ^ n7688 ;
  assign n29478 = n1904 ^ n699 ^ 1'b0 ;
  assign n29479 = n18791 ^ n14002 ^ 1'b0 ;
  assign n29480 = ~n1496 & n12965 ;
  assign n29481 = ( n7206 & n14950 ) | ( n7206 & ~n29480 ) | ( n14950 & ~n29480 ) ;
  assign n29482 = ( n6702 & n11653 ) | ( n6702 & ~n22681 ) | ( n11653 & ~n22681 ) ;
  assign n29483 = n29481 & n29482 ;
  assign n29485 = ( n741 & ~n2203 ) | ( n741 & n11208 ) | ( ~n2203 & n11208 ) ;
  assign n29484 = ( n7129 & n16273 ) | ( n7129 & ~n17315 ) | ( n16273 & ~n17315 ) ;
  assign n29486 = n29485 ^ n29484 ^ n2465 ;
  assign n29487 = n16185 ^ n2856 ^ 1'b0 ;
  assign n29488 = n29487 ^ n10342 ^ n1251 ;
  assign n29489 = ( n836 & n1739 ) | ( n836 & ~n3002 ) | ( n1739 & ~n3002 ) ;
  assign n29490 = n29489 ^ n26090 ^ n3067 ;
  assign n29491 = n29490 ^ n13646 ^ n10431 ;
  assign n29492 = n23016 ^ n10681 ^ 1'b0 ;
  assign n29493 = n6873 & n29492 ;
  assign n29494 = n19926 | n23199 ;
  assign n29495 = n20600 | n29494 ;
  assign n29496 = ( ~n10601 & n24631 ) | ( ~n10601 & n27487 ) | ( n24631 & n27487 ) ;
  assign n29497 = n2040 & ~n22047 ;
  assign n29498 = n5599 | n29497 ;
  assign n29499 = ( ~n463 & n12014 ) | ( ~n463 & n29498 ) | ( n12014 & n29498 ) ;
  assign n29500 = ( n2205 & n15049 ) | ( n2205 & n25711 ) | ( n15049 & n25711 ) ;
  assign n29501 = n14442 & ~n20130 ;
  assign n29502 = n29501 ^ n13863 ^ 1'b0 ;
  assign n29503 = ( n4212 & n5281 ) | ( n4212 & ~n29502 ) | ( n5281 & ~n29502 ) ;
  assign n29504 = n13918 ^ n13195 ^ n5464 ;
  assign n29505 = ( n6192 & n7635 ) | ( n6192 & ~n14313 ) | ( n7635 & ~n14313 ) ;
  assign n29506 = n29505 ^ n20132 ^ n17262 ;
  assign n29509 = ( n856 & ~n4767 ) | ( n856 & n16374 ) | ( ~n4767 & n16374 ) ;
  assign n29507 = n24529 ^ n11122 ^ n10744 ;
  assign n29508 = ( n22360 & ~n23573 ) | ( n22360 & n29507 ) | ( ~n23573 & n29507 ) ;
  assign n29510 = n29509 ^ n29508 ^ n21743 ;
  assign n29511 = ( n1441 & n4165 ) | ( n1441 & ~n10381 ) | ( n4165 & ~n10381 ) ;
  assign n29512 = ( n8363 & n29502 ) | ( n8363 & ~n29511 ) | ( n29502 & ~n29511 ) ;
  assign n29513 = n13796 ^ n2518 ^ 1'b0 ;
  assign n29514 = ~n22698 & n29513 ;
  assign n29517 = n23128 ^ n9583 ^ n4083 ;
  assign n29518 = n29517 ^ n4853 ^ n3259 ;
  assign n29515 = ( n3793 & ~n4024 ) | ( n3793 & n9976 ) | ( ~n4024 & n9976 ) ;
  assign n29516 = n29515 ^ n6263 ^ n525 ;
  assign n29519 = n29518 ^ n29516 ^ n27267 ;
  assign n29520 = ( n5489 & ~n23264 ) | ( n5489 & n29519 ) | ( ~n23264 & n29519 ) ;
  assign n29521 = ( n13255 & ~n17976 ) | ( n13255 & n20879 ) | ( ~n17976 & n20879 ) ;
  assign n29522 = ( n2273 & n7727 ) | ( n2273 & n14900 ) | ( n7727 & n14900 ) ;
  assign n29523 = n29522 ^ n21477 ^ n18935 ;
  assign n29524 = n18116 & ~n29523 ;
  assign n29525 = ( ~n771 & n3342 ) | ( ~n771 & n12940 ) | ( n3342 & n12940 ) ;
  assign n29526 = ( n5814 & n22182 ) | ( n5814 & ~n29525 ) | ( n22182 & ~n29525 ) ;
  assign n29527 = n214 | n20342 ;
  assign n29528 = n19336 | n29527 ;
  assign n29529 = n29528 ^ n7140 ^ n5114 ;
  assign n29530 = n27487 ^ n16272 ^ n7988 ;
  assign n29531 = n7536 | n10946 ;
  assign n29532 = n8035 & ~n29531 ;
  assign n29533 = n29532 ^ n19104 ^ n14405 ;
  assign n29534 = n23005 ^ n3479 ^ n1698 ;
  assign n29535 = n29534 ^ n20032 ^ n11617 ;
  assign n29536 = n29535 ^ n20220 ^ n9571 ;
  assign n29537 = n8770 ^ n2240 ^ n358 ;
  assign n29538 = n4658 | n7365 ;
  assign n29539 = n29538 ^ n10358 ^ 1'b0 ;
  assign n29540 = n794 & n29539 ;
  assign n29541 = n29540 ^ n12342 ^ 1'b0 ;
  assign n29542 = ( n12442 & ~n29537 ) | ( n12442 & n29541 ) | ( ~n29537 & n29541 ) ;
  assign n29544 = n13441 ^ n8657 ^ n7324 ;
  assign n29543 = ~n25916 & n27134 ;
  assign n29545 = n29544 ^ n29543 ^ 1'b0 ;
  assign n29546 = n26461 ^ n17020 ^ n6986 ;
  assign n29547 = n21296 ^ n14927 ^ n10189 ;
  assign n29548 = n28573 | n29547 ;
  assign n29549 = n1347 & ~n29548 ;
  assign n29550 = n29549 ^ n16075 ^ n3252 ;
  assign n29551 = ( n487 & n2667 ) | ( n487 & n9183 ) | ( n2667 & n9183 ) ;
  assign n29552 = n17763 ^ n17068 ^ n11888 ;
  assign n29553 = n17859 ^ n7716 ^ n4024 ;
  assign n29554 = n15882 ^ n4636 ^ 1'b0 ;
  assign n29555 = ( n4776 & n12130 ) | ( n4776 & ~n27025 ) | ( n12130 & ~n27025 ) ;
  assign n29556 = ( n8330 & n10391 ) | ( n8330 & ~n23952 ) | ( n10391 & ~n23952 ) ;
  assign n29557 = ( n5475 & ~n5991 ) | ( n5475 & n13607 ) | ( ~n5991 & n13607 ) ;
  assign n29558 = ~n17291 & n21126 ;
  assign n29559 = n10904 ^ n3541 ^ 1'b0 ;
  assign n29560 = ~n29558 & n29559 ;
  assign n29562 = ( n1267 & n2696 ) | ( n1267 & n7486 ) | ( n2696 & n7486 ) ;
  assign n29561 = n5146 & ~n22183 ;
  assign n29563 = n29562 ^ n29561 ^ 1'b0 ;
  assign n29564 = n20244 ^ n19853 ^ n7386 ;
  assign n29565 = ( n20040 & n26619 ) | ( n20040 & ~n29564 ) | ( n26619 & ~n29564 ) ;
  assign n29567 = ( ~n1143 & n16810 ) | ( ~n1143 & n16857 ) | ( n16810 & n16857 ) ;
  assign n29566 = n15942 ^ n8134 ^ n4500 ;
  assign n29568 = n29567 ^ n29566 ^ n3122 ;
  assign n29569 = n11363 ^ n5490 ^ n3611 ;
  assign n29570 = ( n5908 & ~n28428 ) | ( n5908 & n29569 ) | ( ~n28428 & n29569 ) ;
  assign n29571 = ( n859 & ~n10821 ) | ( n859 & n21287 ) | ( ~n10821 & n21287 ) ;
  assign n29572 = n7146 | n9109 ;
  assign n29573 = n29572 ^ n5822 ^ 1'b0 ;
  assign n29574 = n29573 ^ n16868 ^ n14007 ;
  assign n29575 = n29574 ^ n27745 ^ n919 ;
  assign n29576 = n25752 ^ n24565 ^ n17685 ;
  assign n29577 = n16045 ^ n5825 ^ n3753 ;
  assign n29578 = n29577 ^ n7406 ^ n3597 ;
  assign n29579 = n4216 | n17029 ;
  assign n29580 = n29579 ^ n23020 ^ n11012 ;
  assign n29581 = ( n25451 & n25810 ) | ( n25451 & ~n29580 ) | ( n25810 & ~n29580 ) ;
  assign n29582 = n12908 ^ n11323 ^ n2393 ;
  assign n29583 = n29582 ^ n23407 ^ 1'b0 ;
  assign n29584 = n20355 ^ n13676 ^ n1722 ;
  assign n29585 = n29584 ^ n19504 ^ n17460 ;
  assign n29586 = n29585 ^ n6220 ^ n1223 ;
  assign n29587 = n15779 ^ n14627 ^ n4633 ;
  assign n29588 = n25445 ^ n18126 ^ x84 ;
  assign n29589 = n29588 ^ n27915 ^ n6092 ;
  assign n29590 = ~x107 & n220 ;
  assign n29591 = n8018 ^ n373 ^ 1'b0 ;
  assign n29592 = n13428 & ~n29591 ;
  assign n29593 = n29592 ^ n21607 ^ n2465 ;
  assign n29594 = n29593 ^ n18308 ^ n15480 ;
  assign n29595 = ( n3372 & n29590 ) | ( n3372 & n29594 ) | ( n29590 & n29594 ) ;
  assign n29596 = ( n639 & ~n22892 ) | ( n639 & n29595 ) | ( ~n22892 & n29595 ) ;
  assign n29597 = n18171 & n18378 ;
  assign n29598 = n29597 ^ n11057 ^ n1886 ;
  assign n29599 = n2021 | n27832 ;
  assign n29600 = n29599 ^ n6922 ^ 1'b0 ;
  assign n29601 = n29600 ^ n16781 ^ n8328 ;
  assign n29602 = ( n5987 & n6024 ) | ( n5987 & ~n19784 ) | ( n6024 & ~n19784 ) ;
  assign n29603 = ( n2154 & ~n7545 ) | ( n2154 & n29602 ) | ( ~n7545 & n29602 ) ;
  assign n29604 = n11537 ^ n5503 ^ 1'b0 ;
  assign n29605 = n29604 ^ n13320 ^ n9867 ;
  assign n29606 = n27139 & n29605 ;
  assign n29607 = n7671 ^ n265 ^ 1'b0 ;
  assign n29608 = ~n6715 & n29607 ;
  assign n29609 = ( n8396 & ~n16047 ) | ( n8396 & n25261 ) | ( ~n16047 & n25261 ) ;
  assign n29610 = ( n4344 & ~n29608 ) | ( n4344 & n29609 ) | ( ~n29608 & n29609 ) ;
  assign n29611 = n29610 ^ n14366 ^ n10668 ;
  assign n29612 = n29611 ^ n18429 ^ n8243 ;
  assign n29613 = n16976 ^ n13323 ^ n6633 ;
  assign n29614 = n29613 ^ n18672 ^ n4536 ;
  assign n29615 = n23331 ^ n2207 ^ 1'b0 ;
  assign n29616 = n4985 | n16680 ;
  assign n29617 = n29616 ^ n29522 ^ 1'b0 ;
  assign n29618 = ( n3890 & ~n12452 ) | ( n3890 & n29617 ) | ( ~n12452 & n29617 ) ;
  assign n29619 = n15299 ^ n13379 ^ n10206 ;
  assign n29620 = ( n1146 & n22466 ) | ( n1146 & ~n29619 ) | ( n22466 & ~n29619 ) ;
  assign n29621 = n29620 ^ n3456 ^ 1'b0 ;
  assign n29622 = ( ~n22578 & n26078 ) | ( ~n22578 & n29621 ) | ( n26078 & n29621 ) ;
  assign n29623 = ( n7798 & ~n29618 ) | ( n7798 & n29622 ) | ( ~n29618 & n29622 ) ;
  assign n29628 = ( ~n198 & n5822 ) | ( ~n198 & n13111 ) | ( n5822 & n13111 ) ;
  assign n29626 = ( n15560 & ~n18020 ) | ( n15560 & n24207 ) | ( ~n18020 & n24207 ) ;
  assign n29624 = n16423 ^ n6453 ^ n2583 ;
  assign n29625 = n2328 & ~n29624 ;
  assign n29627 = n29626 ^ n29625 ^ 1'b0 ;
  assign n29629 = n29628 ^ n29627 ^ n14161 ;
  assign n29630 = ( n702 & ~n1348 ) | ( n702 & n5062 ) | ( ~n1348 & n5062 ) ;
  assign n29631 = ( ~n6473 & n8341 ) | ( ~n6473 & n29630 ) | ( n8341 & n29630 ) ;
  assign n29632 = ~n12373 & n22082 ;
  assign n29633 = ( ~n9891 & n20603 ) | ( ~n9891 & n25718 ) | ( n20603 & n25718 ) ;
  assign n29634 = n19138 ^ n13205 ^ 1'b0 ;
  assign n29635 = ( n6845 & n14633 ) | ( n6845 & ~n29634 ) | ( n14633 & ~n29634 ) ;
  assign n29636 = n29635 ^ n5783 ^ 1'b0 ;
  assign n29637 = n29633 & n29636 ;
  assign n29638 = ( ~n7035 & n10088 ) | ( ~n7035 & n25513 ) | ( n10088 & n25513 ) ;
  assign n29639 = n8155 | n29638 ;
  assign n29640 = n7735 ^ n6453 ^ n3604 ;
  assign n29641 = ( n11721 & n19802 ) | ( n11721 & ~n29640 ) | ( n19802 & ~n29640 ) ;
  assign n29642 = n19286 ^ n7358 ^ n1822 ;
  assign n29643 = n2877 & ~n20201 ;
  assign n29644 = ( ~n5172 & n29642 ) | ( ~n5172 & n29643 ) | ( n29642 & n29643 ) ;
  assign n29645 = ( n15300 & ~n29641 ) | ( n15300 & n29644 ) | ( ~n29641 & n29644 ) ;
  assign n29646 = n29645 ^ n21805 ^ n14068 ;
  assign n29647 = ( n1130 & n2328 ) | ( n1130 & n26279 ) | ( n2328 & n26279 ) ;
  assign n29648 = n29647 ^ n1750 ^ n1403 ;
  assign n29651 = n2609 & ~n16611 ;
  assign n29649 = ~n6331 & n15800 ;
  assign n29650 = n29649 ^ n2558 ^ 1'b0 ;
  assign n29652 = n29651 ^ n29650 ^ n5150 ;
  assign n29653 = ( ~n2454 & n12329 ) | ( ~n2454 & n16958 ) | ( n12329 & n16958 ) ;
  assign n29654 = ( n13547 & n29652 ) | ( n13547 & ~n29653 ) | ( n29652 & ~n29653 ) ;
  assign n29655 = n29654 ^ n26360 ^ n1983 ;
  assign n29656 = ( n3706 & n6688 ) | ( n3706 & n17071 ) | ( n6688 & n17071 ) ;
  assign n29657 = ( n3563 & n14718 ) | ( n3563 & n29656 ) | ( n14718 & n29656 ) ;
  assign n29658 = n29657 ^ n20887 ^ n8172 ;
  assign n29659 = n16304 ^ n15383 ^ n12336 ;
  assign n29660 = n29659 ^ n28803 ^ n4011 ;
  assign n29661 = n17775 ^ n17694 ^ n4709 ;
  assign n29662 = ( n4618 & n5195 ) | ( n4618 & n8247 ) | ( n5195 & n8247 ) ;
  assign n29663 = n29662 ^ n10140 ^ n757 ;
  assign n29664 = n29663 ^ n4816 ^ 1'b0 ;
  assign n29665 = n24423 ^ n22484 ^ n6170 ;
  assign n29666 = n22499 ^ n10760 ^ n7180 ;
  assign n29667 = ( ~n9146 & n28175 ) | ( ~n9146 & n29666 ) | ( n28175 & n29666 ) ;
  assign n29668 = x118 & ~n7923 ;
  assign n29669 = n29667 & n29668 ;
  assign n29670 = n15026 ^ n6092 ^ n3957 ;
  assign n29671 = ( n7153 & ~n9038 ) | ( n7153 & n29670 ) | ( ~n9038 & n29670 ) ;
  assign n29672 = n10176 ^ n2836 ^ n1662 ;
  assign n29673 = n25709 | n29672 ;
  assign n29674 = n29671 & n29673 ;
  assign n29675 = n16188 & ~n29674 ;
  assign n29676 = n24008 ^ n209 ^ 1'b0 ;
  assign n29677 = n6536 | n10303 ;
  assign n29678 = n29676 & ~n29677 ;
  assign n29679 = n11350 ^ n11013 ^ n761 ;
  assign n29680 = ( n4852 & n18063 ) | ( n4852 & n29679 ) | ( n18063 & n29679 ) ;
  assign n29681 = ( n6978 & n29678 ) | ( n6978 & ~n29680 ) | ( n29678 & ~n29680 ) ;
  assign n29682 = ( n16285 & ~n23809 ) | ( n16285 & n29681 ) | ( ~n23809 & n29681 ) ;
  assign n29683 = n5782 ^ n5263 ^ n161 ;
  assign n29684 = n29683 ^ n16163 ^ n1951 ;
  assign n29685 = n29684 ^ n22907 ^ n10292 ;
  assign n29686 = ( n3658 & n12764 ) | ( n3658 & ~n14554 ) | ( n12764 & ~n14554 ) ;
  assign n29687 = ( n799 & ~n13117 ) | ( n799 & n18372 ) | ( ~n13117 & n18372 ) ;
  assign n29688 = ( ~n8858 & n16395 ) | ( ~n8858 & n23816 ) | ( n16395 & n23816 ) ;
  assign n29689 = n7385 ^ n3613 ^ n2599 ;
  assign n29690 = ( ~n2651 & n10021 ) | ( ~n2651 & n17191 ) | ( n10021 & n17191 ) ;
  assign n29691 = ( n13635 & ~n27448 ) | ( n13635 & n29690 ) | ( ~n27448 & n29690 ) ;
  assign n29692 = n21749 ^ n9709 ^ n8691 ;
  assign n29693 = n29692 ^ n13214 ^ n5022 ;
  assign n29694 = n28656 ^ n25708 ^ n12032 ;
  assign n29695 = ~n3622 & n29694 ;
  assign n29696 = ( n4121 & ~n5819 ) | ( n4121 & n18317 ) | ( ~n5819 & n18317 ) ;
  assign n29697 = ( ~n4117 & n11636 ) | ( ~n4117 & n29696 ) | ( n11636 & n29696 ) ;
  assign n29698 = ( n6417 & n20795 ) | ( n6417 & n21341 ) | ( n20795 & n21341 ) ;
  assign n29702 = n21262 ^ n13106 ^ n7407 ;
  assign n29699 = ( ~n14478 & n19206 ) | ( ~n14478 & n20067 ) | ( n19206 & n20067 ) ;
  assign n29700 = n29699 ^ n13263 ^ n11858 ;
  assign n29701 = n29700 ^ n10211 ^ n9035 ;
  assign n29703 = n29702 ^ n29701 ^ n15183 ;
  assign n29704 = ( n5442 & ~n9046 ) | ( n5442 & n14666 ) | ( ~n9046 & n14666 ) ;
  assign n29705 = n29704 ^ n28929 ^ n9568 ;
  assign n29706 = n14226 ^ n3847 ^ n2664 ;
  assign n29707 = n13887 ^ n1424 ^ n1355 ;
  assign n29708 = n29707 ^ n20151 ^ n788 ;
  assign n29709 = ( n27217 & n29706 ) | ( n27217 & ~n29708 ) | ( n29706 & ~n29708 ) ;
  assign n29710 = n14815 ^ n6087 ^ n2051 ;
  assign n29711 = n29710 ^ n3172 ^ n1570 ;
  assign n29712 = ( n314 & ~n12528 ) | ( n314 & n29160 ) | ( ~n12528 & n29160 ) ;
  assign n29713 = n29712 ^ n8393 ^ n5524 ;
  assign n29714 = n2662 | n12554 ;
  assign n29715 = n7706 & ~n29714 ;
  assign n29716 = n24054 ^ n5653 ^ 1'b0 ;
  assign n29717 = n5023 & ~n8142 ;
  assign n29718 = n29717 ^ n7409 ^ 1'b0 ;
  assign n29719 = ( n7233 & n10557 ) | ( n7233 & ~n17984 ) | ( n10557 & ~n17984 ) ;
  assign n29720 = n29719 ^ n18693 ^ n1610 ;
  assign n29721 = ( ~n3313 & n9538 ) | ( ~n3313 & n25448 ) | ( n9538 & n25448 ) ;
  assign n29722 = ( n7765 & n27158 ) | ( n7765 & n29721 ) | ( n27158 & n29721 ) ;
  assign n29723 = ( ~n29718 & n29720 ) | ( ~n29718 & n29722 ) | ( n29720 & n29722 ) ;
  assign n29724 = n27670 ^ n25811 ^ n7516 ;
  assign n29725 = ~n875 & n26339 ;
  assign n29726 = n22258 | n29725 ;
  assign n29727 = n6002 | n9413 ;
  assign n29728 = ( n20436 & ~n20916 ) | ( n20436 & n29727 ) | ( ~n20916 & n29727 ) ;
  assign n29729 = ( n6326 & n15247 ) | ( n6326 & ~n29728 ) | ( n15247 & ~n29728 ) ;
  assign n29730 = n29729 ^ n28428 ^ n18026 ;
  assign n29731 = n13142 ^ n1045 ^ n945 ;
  assign n29732 = n27474 ^ n14246 ^ n12799 ;
  assign n29733 = ( ~n16817 & n29731 ) | ( ~n16817 & n29732 ) | ( n29731 & n29732 ) ;
  assign n29734 = n6598 ^ n3339 ^ x43 ;
  assign n29737 = n12285 & ~n14272 ;
  assign n29738 = n29737 ^ n26128 ^ 1'b0 ;
  assign n29735 = ~n4258 & n8950 ;
  assign n29736 = n29735 ^ n26555 ^ n12114 ;
  assign n29739 = n29738 ^ n29736 ^ n18576 ;
  assign n29740 = ( n14580 & n23633 ) | ( n14580 & ~n29739 ) | ( n23633 & ~n29739 ) ;
  assign n29741 = n2083 & ~n29740 ;
  assign n29743 = ( ~n1831 & n5722 ) | ( ~n1831 & n7595 ) | ( n5722 & n7595 ) ;
  assign n29742 = n10176 & ~n16572 ;
  assign n29744 = n29743 ^ n29742 ^ 1'b0 ;
  assign n29745 = ( ~n15473 & n29021 ) | ( ~n15473 & n29744 ) | ( n29021 & n29744 ) ;
  assign n29746 = n2875 & n7047 ;
  assign n29747 = n12658 & n29746 ;
  assign n29748 = n29253 ^ n28543 ^ n1827 ;
  assign n29749 = n20525 ^ n10879 ^ n10044 ;
  assign n29750 = ( n8328 & n13994 ) | ( n8328 & ~n15277 ) | ( n13994 & ~n15277 ) ;
  assign n29751 = ( n1872 & n2021 ) | ( n1872 & n11716 ) | ( n2021 & n11716 ) ;
  assign n29752 = n29751 ^ n8243 ^ n6600 ;
  assign n29753 = n29752 ^ n13130 ^ n3409 ;
  assign n29754 = n2050 & ~n10027 ;
  assign n29755 = n29754 ^ n28475 ^ n24697 ;
  assign n29756 = n29755 ^ n21761 ^ n5037 ;
  assign n29757 = n17813 ^ n5546 ^ n3944 ;
  assign n29758 = ( n7567 & ~n15952 ) | ( n7567 & n29757 ) | ( ~n15952 & n29757 ) ;
  assign n29759 = ( n4486 & n13378 ) | ( n4486 & n14583 ) | ( n13378 & n14583 ) ;
  assign n29760 = ~n28185 & n29759 ;
  assign n29761 = ( n343 & n1919 ) | ( n343 & n4317 ) | ( n1919 & n4317 ) ;
  assign n29762 = n29761 ^ n17039 ^ n15515 ;
  assign n29763 = n29762 ^ n23696 ^ n1983 ;
  assign n29764 = n3482 ^ n2694 ^ n2466 ;
  assign n29765 = ( n7609 & ~n18237 ) | ( n7609 & n27528 ) | ( ~n18237 & n27528 ) ;
  assign n29766 = n22402 & ~n29765 ;
  assign n29767 = n1003 & n29766 ;
  assign n29768 = n29767 ^ n14534 ^ n12488 ;
  assign n29769 = n29764 | n29768 ;
  assign n29770 = n29763 & ~n29769 ;
  assign n29771 = ( n1525 & ~n26773 ) | ( n1525 & n29340 ) | ( ~n26773 & n29340 ) ;
  assign n29772 = n17222 & n29771 ;
  assign n29773 = ( n1211 & n1639 ) | ( n1211 & n2326 ) | ( n1639 & n2326 ) ;
  assign n29774 = n26207 ^ n19796 ^ n11241 ;
  assign n29775 = ( n8496 & n19870 ) | ( n8496 & n25069 ) | ( n19870 & n25069 ) ;
  assign n29776 = n10193 ^ n7469 ^ n6659 ;
  assign n29777 = n12660 & ~n29776 ;
  assign n29778 = n29777 ^ n7403 ^ n1920 ;
  assign n29779 = ( n14096 & n16318 ) | ( n14096 & n27842 ) | ( n16318 & n27842 ) ;
  assign n29780 = n18351 ^ n10929 ^ 1'b0 ;
  assign n29781 = ( ~n1844 & n18481 ) | ( ~n1844 & n26272 ) | ( n18481 & n26272 ) ;
  assign n29784 = n18219 ^ n6959 ^ n426 ;
  assign n29782 = n6056 ^ n2184 ^ n2122 ;
  assign n29783 = ( n16485 & n26965 ) | ( n16485 & ~n29782 ) | ( n26965 & ~n29782 ) ;
  assign n29785 = n29784 ^ n29783 ^ n21673 ;
  assign n29786 = n9838 ^ n6762 ^ n1665 ;
  assign n29787 = ( n12685 & ~n19305 ) | ( n12685 & n29786 ) | ( ~n19305 & n29786 ) ;
  assign n29788 = n2003 | n29787 ;
  assign n29789 = n10551 & ~n29788 ;
  assign n29791 = n19414 ^ n14331 ^ n3213 ;
  assign n29790 = n3862 & ~n14623 ;
  assign n29792 = n29791 ^ n29790 ^ 1'b0 ;
  assign n29794 = ( n2206 & n3559 ) | ( n2206 & n24603 ) | ( n3559 & n24603 ) ;
  assign n29793 = ( n906 & n2503 ) | ( n906 & n3962 ) | ( n2503 & n3962 ) ;
  assign n29795 = n29794 ^ n29793 ^ n10321 ;
  assign n29796 = n9620 ^ n1541 ^ x76 ;
  assign n29797 = n16040 ^ n12403 ^ n7994 ;
  assign n29798 = ( ~n15325 & n16662 ) | ( ~n15325 & n20484 ) | ( n16662 & n20484 ) ;
  assign n29799 = n29798 ^ n16344 ^ n11138 ;
  assign n29800 = ( n5800 & n20667 ) | ( n5800 & ~n29799 ) | ( n20667 & ~n29799 ) ;
  assign n29801 = ( n6696 & n11080 ) | ( n6696 & n21354 ) | ( n11080 & n21354 ) ;
  assign n29802 = ( n13842 & ~n29800 ) | ( n13842 & n29801 ) | ( ~n29800 & n29801 ) ;
  assign n29803 = n28151 ^ n28083 ^ n17477 ;
  assign n29804 = n25151 ^ n15249 ^ n9452 ;
  assign n29805 = ( n12413 & n28883 ) | ( n12413 & ~n29804 ) | ( n28883 & ~n29804 ) ;
  assign n29806 = ( n2455 & ~n2503 ) | ( n2455 & n29805 ) | ( ~n2503 & n29805 ) ;
  assign n29807 = n22478 ^ n4667 ^ n528 ;
  assign n29808 = ~n4902 & n8485 ;
  assign n29809 = n29808 ^ n16837 ^ 1'b0 ;
  assign n29810 = n9770 ^ n6581 ^ n3767 ;
  assign n29811 = n29810 ^ n5050 ^ n1270 ;
  assign n29812 = n23143 ^ n15375 ^ n10044 ;
  assign n29813 = n24917 & n29812 ;
  assign n29814 = n29813 ^ n5840 ^ n4658 ;
  assign n29815 = n1690 & ~n14207 ;
  assign n29816 = ( ~n17450 & n21663 ) | ( ~n17450 & n27733 ) | ( n21663 & n27733 ) ;
  assign n29817 = ( n7599 & ~n13820 ) | ( n7599 & n19452 ) | ( ~n13820 & n19452 ) ;
  assign n29818 = n25981 ^ n20112 ^ 1'b0 ;
  assign n29819 = n9310 ^ n9281 ^ 1'b0 ;
  assign n29820 = ~n17682 & n29819 ;
  assign n29821 = n1514 | n24807 ;
  assign n29822 = n29821 ^ n17650 ^ 1'b0 ;
  assign n29824 = n10704 ^ n2230 ^ x15 ;
  assign n29823 = n24684 ^ n17261 ^ n10639 ;
  assign n29825 = n29824 ^ n29823 ^ n3516 ;
  assign n29826 = n27477 ^ n26615 ^ n25012 ;
  assign n29827 = ( n10913 & n13381 ) | ( n10913 & n19770 ) | ( n13381 & n19770 ) ;
  assign n29828 = n13378 | n15432 ;
  assign n29829 = n16911 & ~n29828 ;
  assign n29830 = n20516 | n29829 ;
  assign n29831 = n29830 ^ n16810 ^ n11548 ;
  assign n29832 = ( n1208 & n2980 ) | ( n1208 & n17293 ) | ( n2980 & n17293 ) ;
  assign n29833 = n29832 ^ n13073 ^ n10600 ;
  assign n29834 = ( n29613 & n29831 ) | ( n29613 & n29833 ) | ( n29831 & n29833 ) ;
  assign n29835 = n25709 ^ n16385 ^ x4 ;
  assign n29840 = n11311 ^ n6697 ^ n3179 ;
  assign n29841 = ( n4901 & ~n15265 ) | ( n4901 & n29840 ) | ( ~n15265 & n29840 ) ;
  assign n29836 = ( n2697 & n9445 ) | ( n2697 & n25462 ) | ( n9445 & n25462 ) ;
  assign n29837 = ~n6941 & n9360 ;
  assign n29838 = n11842 & n29837 ;
  assign n29839 = ( n8503 & ~n29836 ) | ( n8503 & n29838 ) | ( ~n29836 & n29838 ) ;
  assign n29842 = n29841 ^ n29839 ^ n6823 ;
  assign n29843 = ( n3112 & n23624 ) | ( n3112 & ~n28984 ) | ( n23624 & ~n28984 ) ;
  assign n29844 = ( ~n5575 & n16851 ) | ( ~n5575 & n29843 ) | ( n16851 & n29843 ) ;
  assign n29845 = n24699 ^ n20201 ^ n5224 ;
  assign n29846 = ~n2560 & n24979 ;
  assign n29847 = n29846 ^ n27601 ^ 1'b0 ;
  assign n29849 = ( n6202 & n8059 ) | ( n6202 & n15241 ) | ( n8059 & n15241 ) ;
  assign n29848 = n5603 & ~n22033 ;
  assign n29850 = n29849 ^ n29848 ^ 1'b0 ;
  assign n29853 = ( n2919 & ~n20663 ) | ( n2919 & n22995 ) | ( ~n20663 & n22995 ) ;
  assign n29851 = ( n2613 & ~n16827 ) | ( n2613 & n29029 ) | ( ~n16827 & n29029 ) ;
  assign n29852 = n29851 ^ n22640 ^ 1'b0 ;
  assign n29854 = n29853 ^ n29852 ^ n16393 ;
  assign n29855 = n29672 ^ n23331 ^ x122 ;
  assign n29856 = n29855 ^ n7726 ^ n5464 ;
  assign n29857 = n29856 ^ n8700 ^ n302 ;
  assign n29858 = n29857 ^ n9208 ^ n8602 ;
  assign n29859 = n29858 ^ n21430 ^ n19667 ;
  assign n29860 = ( n9269 & n14697 ) | ( n9269 & ~n18583 ) | ( n14697 & ~n18583 ) ;
  assign n29861 = n7222 ^ n4919 ^ n3544 ;
  assign n29862 = n29861 ^ n26407 ^ n22768 ;
  assign n29864 = ~n8177 & n12400 ;
  assign n29865 = n19620 & n29864 ;
  assign n29863 = n22378 ^ n17501 ^ n9767 ;
  assign n29866 = n29865 ^ n29863 ^ n12252 ;
  assign n29867 = n29866 ^ n24843 ^ 1'b0 ;
  assign n29868 = n27305 ^ n20720 ^ n4322 ;
  assign n29869 = n21894 ^ n20693 ^ n10003 ;
  assign n29870 = ( n15506 & n17440 ) | ( n15506 & n29869 ) | ( n17440 & n29869 ) ;
  assign n29871 = n3849 | n5987 ;
  assign n29872 = n29871 ^ n14238 ^ 1'b0 ;
  assign n29873 = ( n5168 & ~n6677 ) | ( n5168 & n29872 ) | ( ~n6677 & n29872 ) ;
  assign n29874 = n8743 ^ n7713 ^ n6169 ;
  assign n29875 = ( n3318 & ~n9388 ) | ( n3318 & n29874 ) | ( ~n9388 & n29874 ) ;
  assign n29876 = n29875 ^ n3061 ^ n918 ;
  assign n29877 = n13377 & ~n29876 ;
  assign n29878 = ( n6658 & n24325 ) | ( n6658 & n26287 ) | ( n24325 & n26287 ) ;
  assign n29879 = ( n1872 & n2121 ) | ( n1872 & ~n27308 ) | ( n2121 & ~n27308 ) ;
  assign n29880 = ( ~n19959 & n29878 ) | ( ~n19959 & n29879 ) | ( n29878 & n29879 ) ;
  assign n29881 = n9927 ^ n9096 ^ 1'b0 ;
  assign n29882 = n29881 ^ n13856 ^ n4887 ;
  assign n29883 = n3160 & ~n3920 ;
  assign n29884 = ( n1739 & ~n22154 ) | ( n1739 & n29883 ) | ( ~n22154 & n29883 ) ;
  assign n29885 = n29884 ^ n27647 ^ n23458 ;
  assign n29886 = n17116 ^ n13227 ^ n2837 ;
  assign n29887 = ( n937 & n15680 ) | ( n937 & n29765 ) | ( n15680 & n29765 ) ;
  assign n29888 = n27976 ^ n4257 ^ n364 ;
  assign n29889 = ( ~x122 & n15715 ) | ( ~x122 & n22929 ) | ( n15715 & n22929 ) ;
  assign n29890 = ( n4471 & n6501 ) | ( n4471 & ~n29889 ) | ( n6501 & ~n29889 ) ;
  assign n29891 = n24184 ^ n21172 ^ n21070 ;
  assign n29892 = n29891 ^ n17537 ^ n7577 ;
  assign n29893 = n29892 ^ n10659 ^ n2030 ;
  assign n29894 = ~n202 & n23190 ;
  assign n29895 = n29894 ^ n1713 ^ 1'b0 ;
  assign n29896 = ( n986 & n18403 ) | ( n986 & n28341 ) | ( n18403 & n28341 ) ;
  assign n29897 = n2273 | n29896 ;
  assign n29898 = x0 | n29897 ;
  assign n29899 = ( ~n3250 & n15325 ) | ( ~n3250 & n16347 ) | ( n15325 & n16347 ) ;
  assign n29900 = ( n3435 & n8864 ) | ( n3435 & n16210 ) | ( n8864 & n16210 ) ;
  assign n29901 = ( n3211 & n25826 ) | ( n3211 & ~n29900 ) | ( n25826 & ~n29900 ) ;
  assign n29902 = n15290 & n19732 ;
  assign n29903 = n29902 ^ n21522 ^ n3758 ;
  assign n29904 = n14236 ^ n9362 ^ n2608 ;
  assign n29905 = x2 | n14822 ;
  assign n29906 = ( n5313 & n18816 ) | ( n5313 & ~n29905 ) | ( n18816 & ~n29905 ) ;
  assign n29907 = n13452 & ~n27435 ;
  assign n29908 = n20348 & n29907 ;
  assign n29909 = n29908 ^ n21063 ^ n16151 ;
  assign n29910 = n25133 ^ n5104 ^ n3940 ;
  assign n29911 = n29910 ^ n9012 ^ n4730 ;
  assign n29912 = ( n29547 & ~n29909 ) | ( n29547 & n29911 ) | ( ~n29909 & n29911 ) ;
  assign n29913 = ( n17293 & ~n19232 ) | ( n17293 & n28608 ) | ( ~n19232 & n28608 ) ;
  assign n29914 = n20235 ^ n19062 ^ n9915 ;
  assign n29915 = n16272 & n29914 ;
  assign n29916 = n29915 ^ n17156 ^ 1'b0 ;
  assign n29917 = ( n2547 & n3039 ) | ( n2547 & n29916 ) | ( n3039 & n29916 ) ;
  assign n29918 = ( n8396 & n24008 ) | ( n8396 & ~n29917 ) | ( n24008 & ~n29917 ) ;
  assign n29919 = n28953 | n29597 ;
  assign n29920 = n19286 ^ n16884 ^ 1'b0 ;
  assign n29921 = n13393 & n29920 ;
  assign n29922 = ( n4256 & n8745 ) | ( n4256 & ~n29921 ) | ( n8745 & ~n29921 ) ;
  assign n29923 = ( n6260 & ~n16285 ) | ( n6260 & n26611 ) | ( ~n16285 & n26611 ) ;
  assign n29924 = ( ~n11620 & n11975 ) | ( ~n11620 & n29923 ) | ( n11975 & n29923 ) ;
  assign n29925 = ( ~n8962 & n10739 ) | ( ~n8962 & n15337 ) | ( n10739 & n15337 ) ;
  assign n29926 = ( n29922 & n29924 ) | ( n29922 & ~n29925 ) | ( n29924 & ~n29925 ) ;
  assign n29927 = n19434 ^ n15225 ^ 1'b0 ;
  assign n29928 = ( n10467 & n10556 ) | ( n10467 & ~n29927 ) | ( n10556 & ~n29927 ) ;
  assign n29929 = n14565 ^ n9344 ^ n466 ;
  assign n29930 = n9201 ^ n9112 ^ n4605 ;
  assign n29931 = ( n2993 & n29929 ) | ( n2993 & n29930 ) | ( n29929 & n29930 ) ;
  assign n29932 = ( n1417 & n6619 ) | ( n1417 & n15544 ) | ( n6619 & n15544 ) ;
  assign n29933 = n15049 ^ n9863 ^ n3529 ;
  assign n29934 = n29933 ^ n14099 ^ 1'b0 ;
  assign n29935 = ( n13298 & ~n29932 ) | ( n13298 & n29934 ) | ( ~n29932 & n29934 ) ;
  assign n29936 = n8959 ^ n1364 ^ 1'b0 ;
  assign n29937 = n29936 ^ n29065 ^ n22632 ;
  assign n29938 = n8229 ^ n138 ^ 1'b0 ;
  assign n29939 = n21156 | n29938 ;
  assign n29940 = ( n11310 & ~n29937 ) | ( n11310 & n29939 ) | ( ~n29937 & n29939 ) ;
  assign n29941 = n16004 ^ n10590 ^ n3808 ;
  assign n29942 = n17622 ^ n5162 ^ n2109 ;
  assign n29943 = ( ~n9889 & n13189 ) | ( ~n9889 & n22121 ) | ( n13189 & n22121 ) ;
  assign n29944 = ~n11099 & n29943 ;
  assign n29945 = n28569 ^ n19908 ^ n3227 ;
  assign n29946 = n29945 ^ n14035 ^ n9726 ;
  assign n29947 = n1638 | n29946 ;
  assign n29948 = n29947 ^ n14039 ^ 1'b0 ;
  assign n29951 = n16987 ^ n6479 ^ n5437 ;
  assign n29949 = n17289 ^ n5897 ^ 1'b0 ;
  assign n29950 = n24919 & ~n29949 ;
  assign n29952 = n29951 ^ n29950 ^ 1'b0 ;
  assign n29953 = n15176 & ~n18720 ;
  assign n29954 = n12513 & ~n15792 ;
  assign n29955 = n14954 & n29954 ;
  assign n29956 = n29955 ^ n8659 ^ n5743 ;
  assign n29957 = n18711 ^ n8843 ^ n7781 ;
  assign n29958 = ( n2073 & n8333 ) | ( n2073 & ~n21312 ) | ( n8333 & ~n21312 ) ;
  assign n29959 = ( n12663 & ~n20947 ) | ( n12663 & n25583 ) | ( ~n20947 & n25583 ) ;
  assign n29960 = n13162 | n23670 ;
  assign n29961 = n25243 ^ n13745 ^ n11271 ;
  assign n29962 = n29961 ^ n28878 ^ n2923 ;
  assign n29964 = n5721 ^ n2878 ^ n1148 ;
  assign n29963 = n29234 ^ n15672 ^ n13163 ;
  assign n29965 = n29964 ^ n29963 ^ n28190 ;
  assign n29967 = n14285 ^ n10578 ^ 1'b0 ;
  assign n29968 = n406 & n29967 ;
  assign n29966 = n23007 ^ n22415 ^ n4113 ;
  assign n29969 = n29968 ^ n29966 ^ n24182 ;
  assign n29970 = n24601 ^ n9009 ^ n5526 ;
  assign n29971 = n29970 ^ n18403 ^ n17049 ;
  assign n29972 = n16851 ^ n4172 ^ 1'b0 ;
  assign n29973 = n16058 | n29972 ;
  assign n29974 = ( n15545 & ~n29971 ) | ( n15545 & n29973 ) | ( ~n29971 & n29973 ) ;
  assign n29975 = n22250 ^ n15879 ^ n6010 ;
  assign n29976 = ( n21213 & n22512 ) | ( n21213 & n23097 ) | ( n22512 & n23097 ) ;
  assign n29977 = n13696 ^ n7822 ^ n981 ;
  assign n29978 = ( n13978 & ~n29976 ) | ( n13978 & n29977 ) | ( ~n29976 & n29977 ) ;
  assign n29979 = ( n2097 & n5701 ) | ( n2097 & ~n11038 ) | ( n5701 & ~n11038 ) ;
  assign n29980 = ( n1094 & n11472 ) | ( n1094 & ~n29979 ) | ( n11472 & ~n29979 ) ;
  assign n29981 = ( ~n13872 & n15123 ) | ( ~n13872 & n29980 ) | ( n15123 & n29980 ) ;
  assign n29985 = n15987 ^ n12955 ^ n5804 ;
  assign n29983 = n23425 ^ n5079 ^ n1121 ;
  assign n29984 = n29983 ^ n16249 ^ n3210 ;
  assign n29982 = ( x44 & n8056 ) | ( x44 & ~n13522 ) | ( n8056 & ~n13522 ) ;
  assign n29986 = n29985 ^ n29984 ^ n29982 ;
  assign n29987 = n8240 ^ n2855 ^ 1'b0 ;
  assign n29988 = n10207 & n29987 ;
  assign n29989 = n18459 ^ n10854 ^ 1'b0 ;
  assign n29991 = n14306 ^ n6386 ^ n2337 ;
  assign n29990 = n1934 & ~n23880 ;
  assign n29992 = n29991 ^ n29990 ^ 1'b0 ;
  assign n29993 = ( n29988 & ~n29989 ) | ( n29988 & n29992 ) | ( ~n29989 & n29992 ) ;
  assign n29994 = ( n3236 & ~n6459 ) | ( n3236 & n23452 ) | ( ~n6459 & n23452 ) ;
  assign n29995 = ( n3898 & ~n20926 ) | ( n3898 & n25265 ) | ( ~n20926 & n25265 ) ;
  assign n29996 = ( n6931 & n29994 ) | ( n6931 & n29995 ) | ( n29994 & n29995 ) ;
  assign n29997 = n29996 ^ n24761 ^ n7540 ;
  assign n29998 = n9542 ^ n6858 ^ n2250 ;
  assign n29999 = n5768 & ~n29998 ;
  assign n30000 = ( n10247 & n28873 ) | ( n10247 & n29999 ) | ( n28873 & n29999 ) ;
  assign n30001 = n13974 & ~n19388 ;
  assign n30002 = n30001 ^ n15061 ^ 1'b0 ;
  assign n30003 = ( n5281 & n11987 ) | ( n5281 & n30002 ) | ( n11987 & n30002 ) ;
  assign n30004 = n18552 ^ n12238 ^ n2699 ;
  assign n30005 = n30004 ^ n26755 ^ n5249 ;
  assign n30006 = ( n1219 & ~n17500 ) | ( n1219 & n27338 ) | ( ~n17500 & n27338 ) ;
  assign n30007 = ( n4228 & ~n12719 ) | ( n4228 & n15118 ) | ( ~n12719 & n15118 ) ;
  assign n30008 = n29592 ^ n22382 ^ n5420 ;
  assign n30009 = ( n18504 & n30007 ) | ( n18504 & n30008 ) | ( n30007 & n30008 ) ;
  assign n30010 = ~n8224 & n16522 ;
  assign n30011 = n1075 & n30010 ;
  assign n30012 = n19411 ^ n15536 ^ n14930 ;
  assign n30013 = ( n21634 & ~n30011 ) | ( n21634 & n30012 ) | ( ~n30011 & n30012 ) ;
  assign n30016 = n28421 ^ n9480 ^ n6524 ;
  assign n30014 = n11566 ^ n7635 ^ n5436 ;
  assign n30015 = ( n3414 & n16861 ) | ( n3414 & ~n30014 ) | ( n16861 & ~n30014 ) ;
  assign n30017 = n30016 ^ n30015 ^ n14745 ;
  assign n30020 = n20719 & n22320 ;
  assign n30021 = n2060 & n30020 ;
  assign n30022 = ( n3694 & n16751 ) | ( n3694 & n30021 ) | ( n16751 & n30021 ) ;
  assign n30018 = ~n474 & n3972 ;
  assign n30019 = ~n1368 & n30018 ;
  assign n30023 = n30022 ^ n30019 ^ n3756 ;
  assign n30024 = n16849 ^ n11048 ^ n6320 ;
  assign n30029 = n6702 | n9905 ;
  assign n30030 = n24119 & ~n30029 ;
  assign n30025 = n9617 ^ n7369 ^ n3484 ;
  assign n30026 = ( ~n881 & n7450 ) | ( ~n881 & n26325 ) | ( n7450 & n26325 ) ;
  assign n30027 = n30026 ^ n22529 ^ n18745 ;
  assign n30028 = ( n11566 & n30025 ) | ( n11566 & n30027 ) | ( n30025 & n30027 ) ;
  assign n30031 = n30030 ^ n30028 ^ n12645 ;
  assign n30032 = n7055 & ~n30031 ;
  assign n30036 = n12052 ^ n9853 ^ n3712 ;
  assign n30033 = n1805 | n1953 ;
  assign n30034 = n10425 | n30033 ;
  assign n30035 = ( n4628 & ~n14830 ) | ( n4628 & n30034 ) | ( ~n14830 & n30034 ) ;
  assign n30037 = n30036 ^ n30035 ^ n16755 ;
  assign n30038 = n26667 ^ n22418 ^ 1'b0 ;
  assign n30039 = n25792 & n30038 ;
  assign n30040 = n13624 & ~n27919 ;
  assign n30041 = n30040 ^ n28843 ^ 1'b0 ;
  assign n30046 = ~n588 & n6788 ;
  assign n30047 = n30046 ^ n14587 ^ 1'b0 ;
  assign n30044 = n3227 & n7731 ;
  assign n30042 = n20736 & n28207 ;
  assign n30043 = n3496 & n30042 ;
  assign n30045 = n30044 ^ n30043 ^ n28727 ;
  assign n30048 = n30047 ^ n30045 ^ n11734 ;
  assign n30049 = ( ~n4784 & n15052 ) | ( ~n4784 & n27044 ) | ( n15052 & n27044 ) ;
  assign n30050 = n13304 ^ n9715 ^ n5058 ;
  assign n30051 = ( n1084 & n8878 ) | ( n1084 & ~n10775 ) | ( n8878 & ~n10775 ) ;
  assign n30052 = ( n8430 & n12580 ) | ( n8430 & ~n19582 ) | ( n12580 & ~n19582 ) ;
  assign n30053 = ( n2263 & ~n18226 ) | ( n2263 & n30052 ) | ( ~n18226 & n30052 ) ;
  assign n30055 = ( n367 & n1647 ) | ( n367 & n8895 ) | ( n1647 & n8895 ) ;
  assign n30054 = n7834 & ~n22698 ;
  assign n30056 = n30055 ^ n30054 ^ 1'b0 ;
  assign n30057 = ( ~n3031 & n22619 ) | ( ~n3031 & n30056 ) | ( n22619 & n30056 ) ;
  assign n30058 = n29371 ^ n8047 ^ 1'b0 ;
  assign n30059 = n193 & n12045 ;
  assign n30060 = n30059 ^ n4251 ^ 1'b0 ;
  assign n30061 = n25414 ^ n21916 ^ n226 ;
  assign n30062 = n12137 & ~n21209 ;
  assign n30063 = ( n6563 & ~n8439 ) | ( n6563 & n10447 ) | ( ~n8439 & n10447 ) ;
  assign n30066 = n17673 ^ n13159 ^ n6393 ;
  assign n30064 = n24152 ^ n3349 ^ n822 ;
  assign n30065 = ( ~n3571 & n15183 ) | ( ~n3571 & n30064 ) | ( n15183 & n30064 ) ;
  assign n30067 = n30066 ^ n30065 ^ n1020 ;
  assign n30068 = ( n6948 & n8594 ) | ( n6948 & ~n30067 ) | ( n8594 & ~n30067 ) ;
  assign n30069 = n22413 ^ n7069 ^ 1'b0 ;
  assign n30070 = ( n17233 & n22768 ) | ( n17233 & ~n30069 ) | ( n22768 & ~n30069 ) ;
  assign n30071 = n28481 ^ n10225 ^ n5989 ;
  assign n30072 = ( ~n6998 & n10088 ) | ( ~n6998 & n21228 ) | ( n10088 & n21228 ) ;
  assign n30073 = ( n2840 & ~n5507 ) | ( n2840 & n6702 ) | ( ~n5507 & n6702 ) ;
  assign n30074 = n22096 | n30073 ;
  assign n30075 = ( n13767 & n14183 ) | ( n13767 & ~n15817 ) | ( n14183 & ~n15817 ) ;
  assign n30076 = ( n6943 & n30074 ) | ( n6943 & n30075 ) | ( n30074 & n30075 ) ;
  assign n30077 = n12131 ^ n997 ^ 1'b0 ;
  assign n30078 = ~n23528 & n30077 ;
  assign n30079 = ( ~n9322 & n10599 ) | ( ~n9322 & n21555 ) | ( n10599 & n21555 ) ;
  assign n30080 = n1135 | n14590 ;
  assign n30081 = n15974 | n30080 ;
  assign n30082 = n30081 ^ n20373 ^ n3058 ;
  assign n30085 = n15720 ^ n558 ^ 1'b0 ;
  assign n30086 = ~n15904 & n30085 ;
  assign n30083 = n12661 ^ n8873 ^ n5248 ;
  assign n30084 = ( ~n265 & n21186 ) | ( ~n265 & n30083 ) | ( n21186 & n30083 ) ;
  assign n30087 = n30086 ^ n30084 ^ n4811 ;
  assign n30088 = n8013 ^ n2848 ^ n2730 ;
  assign n30089 = n26943 ^ n25234 ^ n23618 ;
  assign n30090 = ( n2915 & n8694 ) | ( n2915 & ~n19236 ) | ( n8694 & ~n19236 ) ;
  assign n30091 = n30090 ^ n8046 ^ n5256 ;
  assign n30092 = ( n1694 & n16888 ) | ( n1694 & ~n18147 ) | ( n16888 & ~n18147 ) ;
  assign n30093 = ( n6390 & n9364 ) | ( n6390 & ~n12708 ) | ( n9364 & ~n12708 ) ;
  assign n30094 = ( n6775 & ~n18395 ) | ( n6775 & n26294 ) | ( ~n18395 & n26294 ) ;
  assign n30095 = ( ~n3547 & n10017 ) | ( ~n3547 & n19662 ) | ( n10017 & n19662 ) ;
  assign n30096 = n30095 ^ n25106 ^ n1968 ;
  assign n30097 = ~n26787 & n30096 ;
  assign n30098 = n30097 ^ n1251 ^ 1'b0 ;
  assign n30099 = n24119 ^ n18249 ^ n9799 ;
  assign n30100 = n20989 ^ n17213 ^ n13724 ;
  assign n30101 = n6520 ^ n3983 ^ n189 ;
  assign n30102 = ( ~n14742 & n22794 ) | ( ~n14742 & n30101 ) | ( n22794 & n30101 ) ;
  assign n30103 = n10519 ^ n9965 ^ n2710 ;
  assign n30104 = ~n9008 & n28288 ;
  assign n30105 = ~n7850 & n30104 ;
  assign n30106 = n14540 ^ n2587 ^ 1'b0 ;
  assign n30107 = ~n30105 & n30106 ;
  assign n30108 = n30107 ^ n29927 ^ n13665 ;
  assign n30109 = ( n5951 & n18813 ) | ( n5951 & n28241 ) | ( n18813 & n28241 ) ;
  assign n30112 = ( n5949 & n13117 ) | ( n5949 & n17681 ) | ( n13117 & n17681 ) ;
  assign n30110 = n8185 & ~n24994 ;
  assign n30111 = ~n6023 & n30110 ;
  assign n30113 = n30112 ^ n30111 ^ n690 ;
  assign n30114 = n17476 ^ n7786 ^ n7639 ;
  assign n30115 = n29721 ^ n23809 ^ n23612 ;
  assign n30116 = ( ~n11702 & n18752 ) | ( ~n11702 & n24589 ) | ( n18752 & n24589 ) ;
  assign n30117 = ( ~n475 & n4100 ) | ( ~n475 & n5694 ) | ( n4100 & n5694 ) ;
  assign n30118 = ( n1795 & n2552 ) | ( n1795 & ~n2927 ) | ( n2552 & ~n2927 ) ;
  assign n30119 = n30118 ^ n2450 ^ n721 ;
  assign n30120 = n30119 ^ n20853 ^ 1'b0 ;
  assign n30121 = n14076 ^ n10855 ^ n8490 ;
  assign n30122 = ( ~n2183 & n9101 ) | ( ~n2183 & n30121 ) | ( n9101 & n30121 ) ;
  assign n30123 = n29592 ^ n29157 ^ n11052 ;
  assign n30124 = n8282 ^ n1565 ^ n290 ;
  assign n30125 = n30124 ^ n20727 ^ n13568 ;
  assign n30126 = ( ~n4492 & n6452 ) | ( ~n4492 & n18451 ) | ( n6452 & n18451 ) ;
  assign n30127 = n30126 ^ n14676 ^ n2948 ;
  assign n30128 = n30127 ^ n21472 ^ n1513 ;
  assign n30129 = n24986 ^ n11004 ^ n4880 ;
  assign n30130 = n30129 ^ n21689 ^ n10268 ;
  assign n30131 = ( ~n591 & n7335 ) | ( ~n591 & n7513 ) | ( n7335 & n7513 ) ;
  assign n30133 = ( n6800 & n15248 ) | ( n6800 & ~n15459 ) | ( n15248 & ~n15459 ) ;
  assign n30134 = ( n17172 & n21665 ) | ( n17172 & ~n30133 ) | ( n21665 & ~n30133 ) ;
  assign n30132 = n13109 ^ n2485 ^ 1'b0 ;
  assign n30135 = n30134 ^ n30132 ^ n13810 ;
  assign n30136 = n12334 | n19643 ;
  assign n30137 = n30135 | n30136 ;
  assign n30138 = n8599 & ~n17702 ;
  assign n30139 = ~n27551 & n30138 ;
  assign n30140 = n27002 ^ n3406 ^ n726 ;
  assign n30141 = ( ~n1039 & n2188 ) | ( ~n1039 & n12061 ) | ( n2188 & n12061 ) ;
  assign n30142 = ( n5079 & n8059 ) | ( n5079 & ~n15111 ) | ( n8059 & ~n15111 ) ;
  assign n30143 = n15740 ^ n3994 ^ x71 ;
  assign n30144 = ( ~n2525 & n21664 ) | ( ~n2525 & n30143 ) | ( n21664 & n30143 ) ;
  assign n30145 = n4767 & n4959 ;
  assign n30146 = n26639 ^ n22312 ^ 1'b0 ;
  assign n30147 = ( n13037 & n30145 ) | ( n13037 & ~n30146 ) | ( n30145 & ~n30146 ) ;
  assign n30148 = n7087 ^ n2736 ^ 1'b0 ;
  assign n30149 = n30148 ^ n424 ^ 1'b0 ;
  assign n30150 = n4014 | n30149 ;
  assign n30151 = ( n522 & n3424 ) | ( n522 & ~n30150 ) | ( n3424 & ~n30150 ) ;
  assign n30152 = n17049 ^ n15488 ^ n1288 ;
  assign n30153 = ( n944 & n3224 ) | ( n944 & n30152 ) | ( n3224 & n30152 ) ;
  assign n30154 = ( n5623 & n15470 ) | ( n5623 & ~n30153 ) | ( n15470 & ~n30153 ) ;
  assign n30155 = ( n2848 & n6061 ) | ( n2848 & ~n6819 ) | ( n6061 & ~n6819 ) ;
  assign n30156 = n30155 ^ n27912 ^ n2573 ;
  assign n30158 = ( ~n3416 & n6535 ) | ( ~n3416 & n18100 ) | ( n6535 & n18100 ) ;
  assign n30157 = n10722 | n22035 ;
  assign n30159 = n30158 ^ n30157 ^ 1'b0 ;
  assign n30160 = ( ~n18531 & n27966 ) | ( ~n18531 & n30159 ) | ( n27966 & n30159 ) ;
  assign n30161 = n10808 & ~n24986 ;
  assign n30162 = n19826 & n30161 ;
  assign n30163 = n7942 & ~n22692 ;
  assign n30164 = n30163 ^ n2091 ^ 1'b0 ;
  assign n30165 = n25011 ^ n21431 ^ n14587 ;
  assign n30166 = ( n2580 & n10304 ) | ( n2580 & ~n29672 ) | ( n10304 & ~n29672 ) ;
  assign n30167 = ( n4848 & n9738 ) | ( n4848 & n24144 ) | ( n9738 & n24144 ) ;
  assign n30168 = ( n11364 & n24474 ) | ( n11364 & n30167 ) | ( n24474 & n30167 ) ;
  assign n30169 = ( ~n3161 & n6249 ) | ( ~n3161 & n12015 ) | ( n6249 & n12015 ) ;
  assign n30170 = ( n14263 & ~n23356 ) | ( n14263 & n30169 ) | ( ~n23356 & n30169 ) ;
  assign n30172 = n16494 ^ n10774 ^ n9679 ;
  assign n30171 = n2357 | n6910 ;
  assign n30173 = n30172 ^ n30171 ^ n25849 ;
  assign n30174 = ( ~n2186 & n2452 ) | ( ~n2186 & n10083 ) | ( n2452 & n10083 ) ;
  assign n30175 = n30174 ^ n15395 ^ 1'b0 ;
  assign n30176 = n2303 & n10812 ;
  assign n30177 = n30176 ^ n16539 ^ 1'b0 ;
  assign n30178 = ( n6365 & n20130 ) | ( n6365 & n30177 ) | ( n20130 & n30177 ) ;
  assign n30179 = ( n5103 & ~n16491 ) | ( n5103 & n30178 ) | ( ~n16491 & n30178 ) ;
  assign n30180 = n30179 ^ n21388 ^ n11278 ;
  assign n30181 = ( ~n3651 & n6278 ) | ( ~n3651 & n11663 ) | ( n6278 & n11663 ) ;
  assign n30182 = n17195 ^ n7911 ^ n5504 ;
  assign n30183 = ( n8797 & n23599 ) | ( n8797 & n24313 ) | ( n23599 & n24313 ) ;
  assign n30184 = n29664 ^ n25079 ^ 1'b0 ;
  assign n30185 = n30183 | n30184 ;
  assign n30186 = ( n200 & n656 ) | ( n200 & ~n1730 ) | ( n656 & ~n1730 ) ;
  assign n30187 = n24565 ^ n5961 ^ 1'b0 ;
  assign n30188 = ( n10806 & ~n30186 ) | ( n10806 & n30187 ) | ( ~n30186 & n30187 ) ;
  assign n30189 = n11799 ^ n10348 ^ n7246 ;
  assign n30190 = n30189 ^ n18726 ^ n17961 ;
  assign n30191 = n8816 | n10544 ;
  assign n30192 = n4358 | n18650 ;
  assign n30193 = ( n9719 & n30191 ) | ( n9719 & ~n30192 ) | ( n30191 & ~n30192 ) ;
  assign n30194 = n23489 ^ n10945 ^ n2041 ;
  assign n30195 = n10749 | n30194 ;
  assign n30196 = ( n10834 & n12674 ) | ( n10834 & n30195 ) | ( n12674 & n30195 ) ;
  assign n30197 = ~n5969 & n30196 ;
  assign n30198 = n30197 ^ n1006 ^ 1'b0 ;
  assign n30199 = n30198 ^ n18039 ^ n2241 ;
  assign n30200 = n13779 ^ n12276 ^ n8485 ;
  assign n30201 = ( n2408 & n5913 ) | ( n2408 & n30200 ) | ( n5913 & n30200 ) ;
  assign n30203 = ( n1207 & n13416 ) | ( n1207 & n15931 ) | ( n13416 & n15931 ) ;
  assign n30202 = n154 & ~n5464 ;
  assign n30204 = n30203 ^ n30202 ^ n11055 ;
  assign n30205 = n27740 ^ n8750 ^ 1'b0 ;
  assign n30211 = n18300 ^ n5765 ^ n824 ;
  assign n30206 = n7105 ^ n6176 ^ 1'b0 ;
  assign n30207 = n6922 | n30206 ;
  assign n30208 = n30207 ^ n5373 ^ n3615 ;
  assign n30209 = ( n14891 & n22530 ) | ( n14891 & n22577 ) | ( n22530 & n22577 ) ;
  assign n30210 = ( ~n982 & n30208 ) | ( ~n982 & n30209 ) | ( n30208 & n30209 ) ;
  assign n30212 = n30211 ^ n30210 ^ 1'b0 ;
  assign n30213 = ( n14035 & n30205 ) | ( n14035 & ~n30212 ) | ( n30205 & ~n30212 ) ;
  assign n30214 = ( n25350 & n25959 ) | ( n25350 & n30155 ) | ( n25959 & n30155 ) ;
  assign n30215 = ( ~n2076 & n8836 ) | ( ~n2076 & n12327 ) | ( n8836 & n12327 ) ;
  assign n30216 = ( n11574 & n11608 ) | ( n11574 & n11797 ) | ( n11608 & n11797 ) ;
  assign n30217 = n20829 ^ n15386 ^ n678 ;
  assign n30218 = n30217 ^ n15684 ^ n5298 ;
  assign n30221 = n18935 ^ n10010 ^ n6267 ;
  assign n30222 = ( n5448 & ~n8279 ) | ( n5448 & n30221 ) | ( ~n8279 & n30221 ) ;
  assign n30219 = n24125 ^ n19690 ^ n14046 ;
  assign n30220 = n30219 ^ n26239 ^ n14966 ;
  assign n30223 = n30222 ^ n30220 ^ n6913 ;
  assign n30224 = n7608 ^ n3082 ^ n1878 ;
  assign n30225 = n12918 | n30224 ;
  assign n30226 = n19915 & ~n30225 ;
  assign n30227 = ( ~n13245 & n27495 ) | ( ~n13245 & n30226 ) | ( n27495 & n30226 ) ;
  assign n30228 = ( n2396 & n3300 ) | ( n2396 & n4872 ) | ( n3300 & n4872 ) ;
  assign n30229 = n19526 ^ n14000 ^ n10262 ;
  assign n30230 = n23686 | n30229 ;
  assign n30231 = ( n28822 & n30228 ) | ( n28822 & n30230 ) | ( n30228 & n30230 ) ;
  assign n30232 = n21925 ^ n10929 ^ n8408 ;
  assign n30233 = n12451 & n30232 ;
  assign n30234 = ( n8666 & n21840 ) | ( n8666 & ~n26162 ) | ( n21840 & ~n26162 ) ;
  assign n30235 = ( x105 & n17500 ) | ( x105 & ~n30234 ) | ( n17500 & ~n30234 ) ;
  assign n30236 = ( ~n12087 & n18617 ) | ( ~n12087 & n30235 ) | ( n18617 & n30235 ) ;
  assign n30237 = n22550 ^ n8422 ^ 1'b0 ;
  assign n30238 = n4850 & n22515 ;
  assign n30239 = n23923 & n30238 ;
  assign n30240 = n2440 & ~n10556 ;
  assign n30241 = n30240 ^ n12037 ^ 1'b0 ;
  assign n30242 = n10931 ^ n2453 ^ 1'b0 ;
  assign n30243 = ( n4883 & ~n8078 ) | ( n4883 & n9819 ) | ( ~n8078 & n9819 ) ;
  assign n30244 = n30243 ^ n21025 ^ n4183 ;
  assign n30245 = n15004 & ~n30244 ;
  assign n30246 = n4995 & ~n24626 ;
  assign n30247 = n9709 ^ n3020 ^ 1'b0 ;
  assign n30248 = ( n5033 & n5502 ) | ( n5033 & n30247 ) | ( n5502 & n30247 ) ;
  assign n30249 = n17894 ^ n9351 ^ n6425 ;
  assign n30250 = ( n3386 & n23087 ) | ( n3386 & n30249 ) | ( n23087 & n30249 ) ;
  assign n30251 = n30209 ^ n11005 ^ n5132 ;
  assign n30252 = n29633 ^ n17538 ^ n11661 ;
  assign n30253 = n15612 ^ n8952 ^ n5566 ;
  assign n30254 = ( ~n19356 & n20591 ) | ( ~n19356 & n30253 ) | ( n20591 & n30253 ) ;
  assign n30255 = n18615 ^ n12706 ^ 1'b0 ;
  assign n30256 = n16818 & ~n30255 ;
  assign n30258 = n6285 ^ n5411 ^ 1'b0 ;
  assign n30259 = n25964 ^ n13806 ^ 1'b0 ;
  assign n30260 = n30258 & n30259 ;
  assign n30257 = ~n496 & n2196 ;
  assign n30261 = n30260 ^ n30257 ^ n25553 ;
  assign n30262 = n19406 ^ n10937 ^ n7412 ;
  assign n30263 = ( n1818 & ~n3117 ) | ( n1818 & n30262 ) | ( ~n3117 & n30262 ) ;
  assign n30264 = n24874 ^ n13009 ^ n4726 ;
  assign n30265 = ( n403 & n10189 ) | ( n403 & n30264 ) | ( n10189 & n30264 ) ;
  assign n30266 = ( n16207 & n30263 ) | ( n16207 & ~n30265 ) | ( n30263 & ~n30265 ) ;
  assign n30267 = n5697 ^ n2963 ^ 1'b0 ;
  assign n30268 = ( n6205 & ~n15263 ) | ( n6205 & n15652 ) | ( ~n15263 & n15652 ) ;
  assign n30269 = ( n6922 & n13622 ) | ( n6922 & n20347 ) | ( n13622 & n20347 ) ;
  assign n30270 = ( n2637 & n17378 ) | ( n2637 & ~n30269 ) | ( n17378 & ~n30269 ) ;
  assign n30271 = n12240 ^ n12236 ^ n6957 ;
  assign n30272 = ( n14869 & n18332 ) | ( n14869 & ~n24493 ) | ( n18332 & ~n24493 ) ;
  assign n30273 = ~n3360 & n17653 ;
  assign n30274 = n30273 ^ n3764 ^ 1'b0 ;
  assign n30275 = n305 | n15748 ;
  assign n30276 = n16151 & ~n30275 ;
  assign n30278 = ( n5227 & n5884 ) | ( n5227 & n19964 ) | ( n5884 & n19964 ) ;
  assign n30279 = ( n6723 & ~n18935 ) | ( n6723 & n30278 ) | ( ~n18935 & n30278 ) ;
  assign n30277 = ~n12029 & n28731 ;
  assign n30280 = n30279 ^ n30277 ^ 1'b0 ;
  assign n30281 = ~n11278 & n20656 ;
  assign n30282 = ~n10240 & n30281 ;
  assign n30283 = ( n8040 & n11280 ) | ( n8040 & ~n30282 ) | ( n11280 & ~n30282 ) ;
  assign n30284 = n28281 ^ n13627 ^ x85 ;
  assign n30285 = n30283 & ~n30284 ;
  assign n30286 = ( n1600 & ~n3208 ) | ( n1600 & n16499 ) | ( ~n3208 & n16499 ) ;
  assign n30287 = n9885 ^ n7915 ^ n6038 ;
  assign n30288 = ( n7129 & n22829 ) | ( n7129 & ~n30287 ) | ( n22829 & ~n30287 ) ;
  assign n30289 = n6695 ^ n4637 ^ n4425 ;
  assign n30290 = ( n1817 & n16462 ) | ( n1817 & n30289 ) | ( n16462 & n30289 ) ;
  assign n30291 = n30290 ^ n20034 ^ n19964 ;
  assign n30292 = ( ~n4436 & n7293 ) | ( ~n4436 & n8007 ) | ( n7293 & n8007 ) ;
  assign n30293 = ( n294 & ~n6764 ) | ( n294 & n30292 ) | ( ~n6764 & n30292 ) ;
  assign n30294 = ( n12193 & n29062 ) | ( n12193 & n30293 ) | ( n29062 & n30293 ) ;
  assign n30295 = ( n14087 & ~n16195 ) | ( n14087 & n20914 ) | ( ~n16195 & n20914 ) ;
  assign n30296 = ( ~n3133 & n9356 ) | ( ~n3133 & n19668 ) | ( n9356 & n19668 ) ;
  assign n30297 = n30296 ^ n13139 ^ 1'b0 ;
  assign n30298 = n5939 ^ n1328 ^ 1'b0 ;
  assign n30299 = n19946 ^ n19460 ^ 1'b0 ;
  assign n30300 = ( n9625 & n22361 ) | ( n9625 & n30299 ) | ( n22361 & n30299 ) ;
  assign n30301 = ( n2651 & ~n30298 ) | ( n2651 & n30300 ) | ( ~n30298 & n30300 ) ;
  assign n30302 = n399 & ~n24255 ;
  assign n30303 = n30302 ^ n23797 ^ 1'b0 ;
  assign n30305 = n13493 ^ n10333 ^ n8138 ;
  assign n30306 = ( ~n5079 & n28341 ) | ( ~n5079 & n30305 ) | ( n28341 & n30305 ) ;
  assign n30307 = n30306 ^ n17480 ^ x37 ;
  assign n30308 = n30307 ^ n26018 ^ n4074 ;
  assign n30304 = n10724 & ~n19267 ;
  assign n30309 = n30308 ^ n30304 ^ 1'b0 ;
  assign n30310 = ( n5790 & n21068 ) | ( n5790 & ~n25507 ) | ( n21068 & ~n25507 ) ;
  assign n30311 = ( n6100 & n8230 ) | ( n6100 & n30171 ) | ( n8230 & n30171 ) ;
  assign n30312 = n11096 ^ n6855 ^ n3031 ;
  assign n30313 = n28061 ^ n26514 ^ n13216 ;
  assign n30314 = ( ~n8733 & n8783 ) | ( ~n8733 & n17468 ) | ( n8783 & n17468 ) ;
  assign n30315 = ( n15121 & ~n24956 ) | ( n15121 & n25363 ) | ( ~n24956 & n25363 ) ;
  assign n30316 = ( n7110 & n30314 ) | ( n7110 & ~n30315 ) | ( n30314 & ~n30315 ) ;
  assign n30317 = n19869 ^ n18478 ^ n1114 ;
  assign n30318 = n20423 ^ n13976 ^ n11128 ;
  assign n30319 = n28530 ^ n25929 ^ n8129 ;
  assign n30320 = ~n22126 & n30319 ;
  assign n30321 = n9267 ^ n6253 ^ n2812 ;
  assign n30322 = n30321 ^ n3883 ^ 1'b0 ;
  assign n30323 = ~n6593 & n30322 ;
  assign n30327 = n22086 ^ n6809 ^ 1'b0 ;
  assign n30328 = n30327 ^ n6802 ^ n6433 ;
  assign n30326 = ( ~x75 & n2871 ) | ( ~x75 & n5888 ) | ( n2871 & n5888 ) ;
  assign n30324 = ( n8386 & ~n11592 ) | ( n8386 & n28939 ) | ( ~n11592 & n28939 ) ;
  assign n30325 = ( n5937 & n27204 ) | ( n5937 & n30324 ) | ( n27204 & n30324 ) ;
  assign n30329 = n30328 ^ n30326 ^ n30325 ;
  assign n30330 = ( n7211 & n30323 ) | ( n7211 & ~n30329 ) | ( n30323 & ~n30329 ) ;
  assign n30331 = n20460 ^ n7764 ^ 1'b0 ;
  assign n30332 = n10753 & ~n30331 ;
  assign n30333 = n9439 & ~n12787 ;
  assign n30334 = ~n26703 & n30333 ;
  assign n30335 = n21080 ^ n7638 ^ n6260 ;
  assign n30336 = n25955 ^ n2162 ^ 1'b0 ;
  assign n30337 = n30335 | n30336 ;
  assign n30338 = n30337 ^ n4293 ^ n1178 ;
  assign n30339 = ( n3969 & n12368 ) | ( n3969 & ~n12656 ) | ( n12368 & ~n12656 ) ;
  assign n30340 = n22939 ^ n22807 ^ n4329 ;
  assign n30341 = ( n356 & n5623 ) | ( n356 & ~n30340 ) | ( n5623 & ~n30340 ) ;
  assign n30342 = ( n1022 & n13121 ) | ( n1022 & ~n21817 ) | ( n13121 & ~n21817 ) ;
  assign n30343 = n28664 ^ n2165 ^ 1'b0 ;
  assign n30344 = n22048 ^ n11912 ^ n6884 ;
  assign n30345 = ( ~n28215 & n29400 ) | ( ~n28215 & n30344 ) | ( n29400 & n30344 ) ;
  assign n30346 = n30345 ^ n9416 ^ n6909 ;
  assign n30347 = ( n11320 & n18100 ) | ( n11320 & ~n23781 ) | ( n18100 & ~n23781 ) ;
  assign n30348 = ( ~n9435 & n15696 ) | ( ~n9435 & n30347 ) | ( n15696 & n30347 ) ;
  assign n30349 = n30348 ^ n8603 ^ n6667 ;
  assign n30350 = n15747 ^ n11258 ^ n1762 ;
  assign n30351 = n7026 ^ n5828 ^ n4576 ;
  assign n30352 = n30351 ^ n5816 ^ n521 ;
  assign n30353 = ( n12662 & n26766 ) | ( n12662 & ~n30352 ) | ( n26766 & ~n30352 ) ;
  assign n30355 = n26093 ^ n13253 ^ n5884 ;
  assign n30354 = ( n4437 & n10564 ) | ( n4437 & n29287 ) | ( n10564 & n29287 ) ;
  assign n30356 = n30355 ^ n30354 ^ n19603 ;
  assign n30357 = ( ~n7198 & n7345 ) | ( ~n7198 & n30356 ) | ( n7345 & n30356 ) ;
  assign n30358 = ( n1295 & n30353 ) | ( n1295 & ~n30357 ) | ( n30353 & ~n30357 ) ;
  assign n30359 = n17119 ^ n8060 ^ n3768 ;
  assign n30360 = n30359 ^ n9471 ^ n720 ;
  assign n30361 = ( n646 & n2042 ) | ( n646 & n30360 ) | ( n2042 & n30360 ) ;
  assign n30362 = ~n2509 & n30361 ;
  assign n30363 = n19273 & n30362 ;
  assign n30364 = n18520 ^ n3601 ^ 1'b0 ;
  assign n30365 = ~n23497 & n30364 ;
  assign n30366 = ( n17894 & n18554 ) | ( n17894 & n28992 ) | ( n18554 & n28992 ) ;
  assign n30368 = n15637 ^ n1064 ^ 1'b0 ;
  assign n30367 = ( n3340 & n12442 ) | ( n3340 & ~n25709 ) | ( n12442 & ~n25709 ) ;
  assign n30369 = n30368 ^ n30367 ^ n5810 ;
  assign n30370 = n23746 ^ n13754 ^ n8208 ;
  assign n30371 = n4076 & ~n18330 ;
  assign n30372 = ~n1393 & n30371 ;
  assign n30373 = n30372 ^ n6926 ^ n885 ;
  assign n30374 = ( n6413 & n18167 ) | ( n6413 & n30150 ) | ( n18167 & n30150 ) ;
  assign n30375 = ( ~n3566 & n3757 ) | ( ~n3566 & n10910 ) | ( n3757 & n10910 ) ;
  assign n30376 = n15651 ^ n8738 ^ 1'b0 ;
  assign n30377 = ( ~n1098 & n19940 ) | ( ~n1098 & n30376 ) | ( n19940 & n30376 ) ;
  assign n30378 = ( ~n7852 & n23456 ) | ( ~n7852 & n24731 ) | ( n23456 & n24731 ) ;
  assign n30379 = n7633 ^ n7359 ^ n2032 ;
  assign n30380 = n21273 ^ n20520 ^ n1546 ;
  assign n30381 = n30380 ^ n11079 ^ n7731 ;
  assign n30382 = ( n30378 & n30379 ) | ( n30378 & ~n30381 ) | ( n30379 & ~n30381 ) ;
  assign n30383 = n4467 | n18295 ;
  assign n30384 = n26420 | n30383 ;
  assign n30385 = ( n3162 & n28992 ) | ( n3162 & n30384 ) | ( n28992 & n30384 ) ;
  assign n30386 = ( n3550 & n24386 ) | ( n3550 & ~n30385 ) | ( n24386 & ~n30385 ) ;
  assign n30387 = ( n3274 & n7815 ) | ( n3274 & ~n30386 ) | ( n7815 & ~n30386 ) ;
  assign n30388 = ~n10073 & n14433 ;
  assign n30393 = n3641 ^ n1927 ^ n1496 ;
  assign n30394 = ( n1084 & ~n20939 ) | ( n1084 & n30393 ) | ( ~n20939 & n30393 ) ;
  assign n30389 = n13739 ^ n4948 ^ n3788 ;
  assign n30390 = ( ~n12076 & n25499 ) | ( ~n12076 & n30389 ) | ( n25499 & n30389 ) ;
  assign n30391 = n30390 ^ n16069 ^ n1817 ;
  assign n30392 = ( n8569 & n15621 ) | ( n8569 & n30391 ) | ( n15621 & n30391 ) ;
  assign n30395 = n30394 ^ n30392 ^ n2962 ;
  assign n30396 = ( n10287 & ~n12119 ) | ( n10287 & n18548 ) | ( ~n12119 & n18548 ) ;
  assign n30397 = n665 | n20232 ;
  assign n30398 = n30397 ^ n2595 ^ 1'b0 ;
  assign n30399 = ( n19328 & n27800 ) | ( n19328 & ~n30398 ) | ( n27800 & ~n30398 ) ;
  assign n30400 = ( n7891 & n8202 ) | ( n7891 & ~n18619 ) | ( n8202 & ~n18619 ) ;
  assign n30401 = n1682 & n20929 ;
  assign n30402 = n30401 ^ n25284 ^ 1'b0 ;
  assign n30403 = n12186 | n29743 ;
  assign n30404 = n30403 ^ n22906 ^ 1'b0 ;
  assign n30405 = ( n30400 & n30402 ) | ( n30400 & n30404 ) | ( n30402 & n30404 ) ;
  assign n30406 = n10237 ^ n2813 ^ n1785 ;
  assign n30407 = n30406 ^ n16353 ^ n11560 ;
  assign n30408 = n5092 & ~n21836 ;
  assign n30409 = ( ~n2582 & n3483 ) | ( ~n2582 & n8412 ) | ( n3483 & n8412 ) ;
  assign n30410 = ( n318 & n9343 ) | ( n318 & ~n14045 ) | ( n9343 & ~n14045 ) ;
  assign n30411 = n30410 ^ n15609 ^ 1'b0 ;
  assign n30412 = n15185 | n30411 ;
  assign n30413 = n1803 | n8426 ;
  assign n30414 = ( n5948 & n22688 ) | ( n5948 & n27239 ) | ( n22688 & n27239 ) ;
  assign n30415 = n22088 ^ n20794 ^ n14662 ;
  assign n30416 = ( n8425 & ~n11566 ) | ( n8425 & n15277 ) | ( ~n11566 & n15277 ) ;
  assign n30417 = n30172 ^ n25781 ^ n21200 ;
  assign n30418 = n21067 ^ n6760 ^ 1'b0 ;
  assign n30419 = ~n7862 & n30418 ;
  assign n30420 = n10861 & ~n20885 ;
  assign n30421 = n30420 ^ n22283 ^ n7939 ;
  assign n30422 = ( n17172 & ~n30419 ) | ( n17172 & n30421 ) | ( ~n30419 & n30421 ) ;
  assign n30423 = n17235 ^ n3701 ^ n814 ;
  assign n30424 = ( n1181 & n3115 ) | ( n1181 & ~n24069 ) | ( n3115 & ~n24069 ) ;
  assign n30425 = n10063 ^ n735 ^ 1'b0 ;
  assign n30426 = ~n19895 & n30425 ;
  assign n30427 = n24345 ^ n24221 ^ x9 ;
  assign n30428 = ( n1269 & n6342 ) | ( n1269 & n12767 ) | ( n6342 & n12767 ) ;
  assign n30429 = n30428 ^ n3238 ^ n1768 ;
  assign n30430 = ( n16253 & n24887 ) | ( n16253 & n28063 ) | ( n24887 & n28063 ) ;
  assign n30431 = n23884 ^ n17448 ^ n5144 ;
  assign n30432 = n29731 ^ n5338 ^ n1647 ;
  assign n30433 = ( n2735 & ~n28873 ) | ( n2735 & n30432 ) | ( ~n28873 & n30432 ) ;
  assign n30434 = n15424 ^ n15256 ^ n3951 ;
  assign n30435 = n23260 ^ n13393 ^ n1719 ;
  assign n30436 = n26280 ^ n8035 ^ n5501 ;
  assign n30437 = ~n30435 & n30436 ;
  assign n30438 = ( ~n3452 & n20575 ) | ( ~n3452 & n27214 ) | ( n20575 & n27214 ) ;
  assign n30439 = n30438 ^ n16148 ^ n5231 ;
  assign n30440 = n16535 ^ n14677 ^ 1'b0 ;
  assign n30441 = n5260 & n30440 ;
  assign n30442 = n14340 & n30441 ;
  assign n30443 = n20571 ^ n1555 ^ 1'b0 ;
  assign n30444 = ~n10212 & n30443 ;
  assign n30445 = n10052 & n30444 ;
  assign n30446 = ( n1921 & ~n2958 ) | ( n1921 & n5828 ) | ( ~n2958 & n5828 ) ;
  assign n30447 = n30446 ^ n23611 ^ n13947 ;
  assign n30448 = ( n5866 & n13015 ) | ( n5866 & n30447 ) | ( n13015 & n30447 ) ;
  assign n30449 = ( n390 & ~n5273 ) | ( n390 & n28580 ) | ( ~n5273 & n28580 ) ;
  assign n30450 = ( ~n14803 & n15909 ) | ( ~n14803 & n30449 ) | ( n15909 & n30449 ) ;
  assign n30451 = ( n5346 & n9107 ) | ( n5346 & ~n24002 ) | ( n9107 & ~n24002 ) ;
  assign n30452 = ( ~n1414 & n12816 ) | ( ~n1414 & n22736 ) | ( n12816 & n22736 ) ;
  assign n30453 = n22086 ^ n21571 ^ n4149 ;
  assign n30454 = n10612 ^ n4469 ^ n3454 ;
  assign n30455 = n30454 ^ n25664 ^ n8946 ;
  assign n30456 = n18294 ^ n15325 ^ n2895 ;
  assign n30457 = ( ~n3884 & n4382 ) | ( ~n3884 & n30456 ) | ( n4382 & n30456 ) ;
  assign n30458 = ( x37 & n228 ) | ( x37 & ~n7283 ) | ( n228 & ~n7283 ) ;
  assign n30459 = n30458 ^ n21373 ^ n2599 ;
  assign n30460 = n29910 ^ n29132 ^ n26023 ;
  assign n30462 = n26745 ^ n11036 ^ n3288 ;
  assign n30461 = ~n2349 & n7460 ;
  assign n30463 = n30462 ^ n30461 ^ 1'b0 ;
  assign n30464 = n12615 ^ n7335 ^ n1805 ;
  assign n30465 = ( n11415 & n21884 ) | ( n11415 & n30464 ) | ( n21884 & n30464 ) ;
  assign n30466 = ( n5225 & n10102 ) | ( n5225 & n18352 ) | ( n10102 & n18352 ) ;
  assign n30467 = n26580 ^ n13160 ^ n5605 ;
  assign n30468 = n30467 ^ n24703 ^ n20095 ;
  assign n30469 = ( n28623 & ~n30466 ) | ( n28623 & n30468 ) | ( ~n30466 & n30468 ) ;
  assign n30470 = n27101 ^ n22839 ^ n19384 ;
  assign n30471 = ( n21000 & ~n23131 ) | ( n21000 & n23821 ) | ( ~n23131 & n23821 ) ;
  assign n30472 = n30471 ^ n25869 ^ n6378 ;
  assign n30478 = ( n1415 & n4982 ) | ( n1415 & ~n9891 ) | ( n4982 & ~n9891 ) ;
  assign n30473 = n14509 ^ n3092 ^ n2908 ;
  assign n30474 = ( n2141 & n19893 ) | ( n2141 & ~n21172 ) | ( n19893 & ~n21172 ) ;
  assign n30475 = ( n544 & n10182 ) | ( n544 & n30474 ) | ( n10182 & n30474 ) ;
  assign n30476 = n30475 ^ n2943 ^ 1'b0 ;
  assign n30477 = n30473 | n30476 ;
  assign n30479 = n30478 ^ n30477 ^ n26413 ;
  assign n30480 = ( n5720 & n10407 ) | ( n5720 & ~n24809 ) | ( n10407 & ~n24809 ) ;
  assign n30481 = n22190 ^ n10114 ^ x122 ;
  assign n30482 = n13556 ^ n9842 ^ n3779 ;
  assign n30483 = n1572 & n30482 ;
  assign n30484 = n15973 ^ n12873 ^ n8031 ;
  assign n30485 = ( n3636 & ~n17706 ) | ( n3636 & n21717 ) | ( ~n17706 & n21717 ) ;
  assign n30486 = n1551 & n30485 ;
  assign n30487 = n5746 & n30486 ;
  assign n30491 = ~n322 & n3902 ;
  assign n30489 = n21806 ^ n6657 ^ n6370 ;
  assign n30490 = n11333 | n30489 ;
  assign n30492 = n30491 ^ n30490 ^ n19969 ;
  assign n30488 = ~n3005 & n24475 ;
  assign n30493 = n30492 ^ n30488 ^ 1'b0 ;
  assign n30494 = ( n5682 & n9682 ) | ( n5682 & ~n25504 ) | ( n9682 & ~n25504 ) ;
  assign n30495 = ( ~n2157 & n5248 ) | ( ~n2157 & n10400 ) | ( n5248 & n10400 ) ;
  assign n30496 = ( ~n13113 & n21422 ) | ( ~n13113 & n30495 ) | ( n21422 & n30495 ) ;
  assign n30497 = n18826 ^ n4411 ^ n3670 ;
  assign n30498 = n30497 ^ n18927 ^ n17717 ;
  assign n30499 = n30498 ^ n11139 ^ n10636 ;
  assign n30500 = n30499 ^ n5522 ^ n3252 ;
  assign n30501 = ( n160 & ~n14033 ) | ( n160 & n26997 ) | ( ~n14033 & n26997 ) ;
  assign n30502 = n14578 ^ n12094 ^ n11374 ;
  assign n30503 = n27651 | n30502 ;
  assign n30504 = ( n1791 & n18412 ) | ( n1791 & ~n27042 ) | ( n18412 & ~n27042 ) ;
  assign n30505 = n11710 ^ n9837 ^ n340 ;
  assign n30506 = ( n1075 & n7123 ) | ( n1075 & n24021 ) | ( n7123 & n24021 ) ;
  assign n30507 = n23935 ^ n11085 ^ 1'b0 ;
  assign n30509 = n23930 ^ n22621 ^ n1257 ;
  assign n30510 = ( n4112 & n8255 ) | ( n4112 & ~n11355 ) | ( n8255 & ~n11355 ) ;
  assign n30511 = n30510 ^ n15953 ^ n8607 ;
  assign n30512 = ( n3437 & n7948 ) | ( n3437 & ~n10744 ) | ( n7948 & ~n10744 ) ;
  assign n30513 = ( n5064 & ~n30511 ) | ( n5064 & n30512 ) | ( ~n30511 & n30512 ) ;
  assign n30514 = n30509 | n30513 ;
  assign n30508 = n6241 & ~n12168 ;
  assign n30515 = n30514 ^ n30508 ^ 1'b0 ;
  assign n30516 = n11744 ^ n7842 ^ 1'b0 ;
  assign n30517 = n3867 & ~n30516 ;
  assign n30518 = n6623 ^ n401 ^ x13 ;
  assign n30519 = n19020 ^ n8776 ^ n5376 ;
  assign n30520 = n16923 ^ n12686 ^ 1'b0 ;
  assign n30521 = ( ~n12530 & n20072 ) | ( ~n12530 & n23176 ) | ( n20072 & n23176 ) ;
  assign n30522 = n26377 ^ n5678 ^ n5069 ;
  assign n30523 = n3382 & n10237 ;
  assign n30524 = n436 & n30523 ;
  assign n30525 = n30524 ^ n21652 ^ n19174 ;
  assign n30526 = n30525 ^ n21578 ^ n18835 ;
  assign n30527 = n10929 ^ n6181 ^ n3470 ;
  assign n30528 = ( ~n7100 & n24854 ) | ( ~n7100 & n30527 ) | ( n24854 & n30527 ) ;
  assign n30529 = ( n2101 & ~n4410 ) | ( n2101 & n30528 ) | ( ~n4410 & n30528 ) ;
  assign n30530 = n27026 ^ n13382 ^ n226 ;
  assign n30531 = ( ~n172 & n793 ) | ( ~n172 & n27264 ) | ( n793 & n27264 ) ;
  assign n30533 = n13604 | n24687 ;
  assign n30532 = n169 | n19298 ;
  assign n30534 = n30533 ^ n30532 ^ 1'b0 ;
  assign n30535 = n17934 ^ n16485 ^ n5414 ;
  assign n30536 = ~n4385 & n30535 ;
  assign n30537 = ( ~n6860 & n18201 ) | ( ~n6860 & n24257 ) | ( n18201 & n24257 ) ;
  assign n30538 = ( n14267 & n23373 ) | ( n14267 & ~n30537 ) | ( n23373 & ~n30537 ) ;
  assign n30539 = ( n5794 & n16961 ) | ( n5794 & n17045 ) | ( n16961 & n17045 ) ;
  assign n30540 = n30539 ^ n27341 ^ n18114 ;
  assign n30541 = ( n9923 & n27469 ) | ( n9923 & ~n30540 ) | ( n27469 & ~n30540 ) ;
  assign n30542 = ( n6819 & ~n7812 ) | ( n6819 & n15865 ) | ( ~n7812 & n15865 ) ;
  assign n30543 = n25492 ^ n14133 ^ n3506 ;
  assign n30544 = n12115 | n21442 ;
  assign n30545 = n30544 ^ n15558 ^ 1'b0 ;
  assign n30546 = ( n5543 & n8839 ) | ( n5543 & n30545 ) | ( n8839 & n30545 ) ;
  assign n30547 = n15799 ^ n10240 ^ 1'b0 ;
  assign n30548 = n19925 ^ n18812 ^ 1'b0 ;
  assign n30549 = ( n6614 & ~n22677 ) | ( n6614 & n30548 ) | ( ~n22677 & n30548 ) ;
  assign n30552 = n9562 ^ n7455 ^ n7390 ;
  assign n30551 = ( n7064 & n11689 ) | ( n7064 & n18762 ) | ( n11689 & n18762 ) ;
  assign n30550 = n4958 ^ n1217 ^ x18 ;
  assign n30553 = n30552 ^ n30551 ^ n30550 ;
  assign n30554 = n30495 ^ n1814 ^ n972 ;
  assign n30555 = n9890 & ~n20048 ;
  assign n30556 = n30555 ^ n26354 ^ 1'b0 ;
  assign n30557 = n17980 ^ n2636 ^ 1'b0 ;
  assign n30558 = n8646 & ~n30557 ;
  assign n30561 = n5867 ^ n4187 ^ n2814 ;
  assign n30562 = n30561 ^ n16675 ^ n2437 ;
  assign n30559 = ( ~n2959 & n9261 ) | ( ~n2959 & n16124 ) | ( n9261 & n16124 ) ;
  assign n30560 = n30559 ^ n20595 ^ 1'b0 ;
  assign n30563 = n30562 ^ n30560 ^ x49 ;
  assign n30564 = n22530 ^ n15459 ^ n244 ;
  assign n30565 = ( n4271 & n14226 ) | ( n4271 & n30564 ) | ( n14226 & n30564 ) ;
  assign n30566 = ( n1342 & ~n16729 ) | ( n1342 & n30565 ) | ( ~n16729 & n30565 ) ;
  assign n30567 = ( n589 & n4291 ) | ( n589 & n10039 ) | ( n4291 & n10039 ) ;
  assign n30568 = n30567 ^ n7964 ^ 1'b0 ;
  assign n30569 = n14065 ^ n2240 ^ n1422 ;
  assign n30570 = n30569 ^ n21501 ^ n13959 ;
  assign n30571 = n18774 ^ n11928 ^ n1284 ;
  assign n30572 = n3845 ^ n575 ^ 1'b0 ;
  assign n30573 = n25522 & ~n30572 ;
  assign n30574 = n16568 ^ n14738 ^ n7044 ;
  assign n30575 = ( n14674 & n30573 ) | ( n14674 & ~n30574 ) | ( n30573 & ~n30574 ) ;
  assign n30576 = ( n4569 & n5378 ) | ( n4569 & n14775 ) | ( n5378 & n14775 ) ;
  assign n30577 = n14780 ^ n9716 ^ n324 ;
  assign n30578 = n23633 ^ n13326 ^ n3109 ;
  assign n30579 = n601 & ~n28921 ;
  assign n30580 = ~n14099 & n30579 ;
  assign n30581 = ( n8585 & n10411 ) | ( n8585 & ~n26319 ) | ( n10411 & ~n26319 ) ;
  assign n30582 = n27744 ^ n25489 ^ n16597 ;
  assign n30583 = ( n2428 & ~n7826 ) | ( n2428 & n11377 ) | ( ~n7826 & n11377 ) ;
  assign n30584 = n30583 ^ n26337 ^ n1577 ;
  assign n30585 = ( n8575 & n13534 ) | ( n8575 & n24252 ) | ( n13534 & n24252 ) ;
  assign n30586 = n2985 ^ n1052 ^ 1'b0 ;
  assign n30587 = ~n30148 & n30586 ;
  assign n30588 = ( n7733 & ~n19033 ) | ( n7733 & n30587 ) | ( ~n19033 & n30587 ) ;
  assign n30589 = n30588 ^ n11906 ^ n297 ;
  assign n30590 = n8156 ^ n1759 ^ n190 ;
  assign n30591 = n20150 | n30590 ;
  assign n30592 = n20151 ^ n871 ^ 1'b0 ;
  assign n30593 = n12282 ^ n2616 ^ 1'b0 ;
  assign n30594 = n17548 ^ n9153 ^ n1400 ;
  assign n30595 = n14266 & ~n30594 ;
  assign n30596 = n19896 ^ n7837 ^ 1'b0 ;
  assign n30597 = n16327 ^ n1985 ^ 1'b0 ;
  assign n30598 = ~n6998 & n30597 ;
  assign n30599 = n1439 | n13630 ;
  assign n30600 = ( ~n8633 & n18860 ) | ( ~n8633 & n30599 ) | ( n18860 & n30599 ) ;
  assign n30601 = ( n4756 & n23732 ) | ( n4756 & n30600 ) | ( n23732 & n30600 ) ;
  assign n30602 = n11556 ^ n7557 ^ n787 ;
  assign n30603 = ( n1183 & ~n9453 ) | ( n1183 & n22428 ) | ( ~n9453 & n22428 ) ;
  assign n30604 = n21770 ^ n11917 ^ n6845 ;
  assign n30605 = ( n7971 & n13999 ) | ( n7971 & n30604 ) | ( n13999 & n30604 ) ;
  assign n30606 = n29324 ^ n23521 ^ n22180 ;
  assign n30607 = n30449 ^ n8935 ^ n651 ;
  assign n30608 = n30607 ^ n7028 ^ n5640 ;
  assign n30609 = n29782 ^ n14995 ^ n12001 ;
  assign n30610 = ( n6286 & ~n28541 ) | ( n6286 & n30609 ) | ( ~n28541 & n30609 ) ;
  assign n30611 = ( n572 & n9494 ) | ( n572 & n22104 ) | ( n9494 & n22104 ) ;
  assign n30612 = n573 & n25228 ;
  assign n30613 = ~n14073 & n30612 ;
  assign n30614 = n437 & n12151 ;
  assign n30615 = ~n9573 & n30614 ;
  assign n30616 = n21405 ^ n11080 ^ 1'b0 ;
  assign n30617 = ~n30615 & n30616 ;
  assign n30618 = ( n2661 & ~n8350 ) | ( n2661 & n16395 ) | ( ~n8350 & n16395 ) ;
  assign n30619 = ( n7665 & n29368 ) | ( n7665 & ~n30618 ) | ( n29368 & ~n30618 ) ;
  assign n30620 = n4223 | n22825 ;
  assign n30621 = n30620 ^ n6900 ^ 1'b0 ;
  assign n30622 = ( n9149 & ~n17787 ) | ( n9149 & n30621 ) | ( ~n17787 & n30621 ) ;
  assign n30623 = ( n15036 & n26404 ) | ( n15036 & n30622 ) | ( n26404 & n30622 ) ;
  assign n30624 = ( ~n1321 & n10676 ) | ( ~n1321 & n19788 ) | ( n10676 & n19788 ) ;
  assign n30625 = ( n6048 & n18667 ) | ( n6048 & ~n26526 ) | ( n18667 & ~n26526 ) ;
  assign n30626 = ( n7557 & n16903 ) | ( n7557 & ~n27679 ) | ( n16903 & ~n27679 ) ;
  assign n30627 = ( n10305 & n24480 ) | ( n10305 & ~n30626 ) | ( n24480 & ~n30626 ) ;
  assign n30628 = n219 & n8398 ;
  assign n30629 = n30628 ^ n746 ^ 1'b0 ;
  assign n30630 = n30629 ^ n22512 ^ n15557 ;
  assign n30632 = n25535 ^ n10538 ^ 1'b0 ;
  assign n30633 = n30632 ^ n19952 ^ n6660 ;
  assign n30631 = ( n2094 & n8873 ) | ( n2094 & ~n30604 ) | ( n8873 & ~n30604 ) ;
  assign n30634 = n30633 ^ n30631 ^ n22245 ;
  assign n30642 = n4406 ^ n3693 ^ 1'b0 ;
  assign n30643 = ( n910 & n9456 ) | ( n910 & n30642 ) | ( n9456 & n30642 ) ;
  assign n30639 = ( n3973 & ~n15602 ) | ( n3973 & n22146 ) | ( ~n15602 & n22146 ) ;
  assign n30640 = n30639 ^ n10299 ^ n9891 ;
  assign n30636 = n24497 ^ n8603 ^ n2002 ;
  assign n30637 = n3474 & ~n30636 ;
  assign n30638 = ~n13235 & n30637 ;
  assign n30635 = n13654 ^ n11704 ^ n4851 ;
  assign n30641 = n30640 ^ n30638 ^ n30635 ;
  assign n30644 = n30643 ^ n30641 ^ n25985 ;
  assign n30645 = ( ~n11983 & n21454 ) | ( ~n11983 & n28184 ) | ( n21454 & n28184 ) ;
  assign n30646 = n8745 ^ n7544 ^ n1411 ;
  assign n30647 = n30646 ^ n7285 ^ n4342 ;
  assign n30648 = n13082 ^ n8914 ^ n6274 ;
  assign n30649 = n25947 ^ n23517 ^ n22489 ;
  assign n30650 = ( ~n1346 & n15272 ) | ( ~n1346 & n21573 ) | ( n15272 & n21573 ) ;
  assign n30651 = n27543 ^ n18649 ^ n8269 ;
  assign n30652 = ( n3415 & n30650 ) | ( n3415 & n30651 ) | ( n30650 & n30651 ) ;
  assign n30653 = n30652 ^ n9512 ^ n705 ;
  assign n30654 = ( n3500 & n21407 ) | ( n3500 & n30653 ) | ( n21407 & n30653 ) ;
  assign n30655 = n30069 ^ n18158 ^ n15880 ;
  assign n30656 = n30655 ^ n13383 ^ n6275 ;
  assign n30657 = n29277 ^ n23256 ^ n2221 ;
  assign n30658 = ( ~n10925 & n18416 ) | ( ~n10925 & n23016 ) | ( n18416 & n23016 ) ;
  assign n30659 = n30658 ^ n13128 ^ n10240 ;
  assign n30660 = n18099 ^ n15390 ^ 1'b0 ;
  assign n30661 = n718 | n5808 ;
  assign n30662 = n8736 & ~n30661 ;
  assign n30663 = n5533 ^ n3605 ^ 1'b0 ;
  assign n30664 = ( n8831 & ~n15515 ) | ( n8831 & n24976 ) | ( ~n15515 & n24976 ) ;
  assign n30665 = ( n14587 & n19810 ) | ( n14587 & ~n30664 ) | ( n19810 & ~n30664 ) ;
  assign n30666 = n23730 ^ n11592 ^ n4454 ;
  assign n30667 = ( ~n5133 & n16691 ) | ( ~n5133 & n28374 ) | ( n16691 & n28374 ) ;
  assign n30668 = n17041 | n30667 ;
  assign n30669 = ( n23114 & n28725 ) | ( n23114 & n30668 ) | ( n28725 & n30668 ) ;
  assign n30670 = n606 & n1336 ;
  assign n30671 = n30670 ^ n6075 ^ 1'b0 ;
  assign n30672 = n30671 ^ n27017 ^ n10879 ;
  assign n30673 = n14673 ^ n8509 ^ n347 ;
  assign n30674 = ( n523 & ~n3943 ) | ( n523 & n30673 ) | ( ~n3943 & n30673 ) ;
  assign n30675 = n30674 ^ n17831 ^ n11749 ;
  assign n30676 = ~n6355 & n20917 ;
  assign n30677 = ( n6016 & n20538 ) | ( n6016 & n30676 ) | ( n20538 & n30676 ) ;
  assign n30678 = ( n12176 & n16992 ) | ( n12176 & ~n22063 ) | ( n16992 & ~n22063 ) ;
  assign n30679 = ( n26663 & n30677 ) | ( n26663 & n30678 ) | ( n30677 & n30678 ) ;
  assign n30680 = ( ~n888 & n10156 ) | ( ~n888 & n18299 ) | ( n10156 & n18299 ) ;
  assign n30681 = ~n4027 & n8470 ;
  assign n30682 = n30680 & n30681 ;
  assign n30684 = ( n3892 & n15005 ) | ( n3892 & n17684 ) | ( n15005 & n17684 ) ;
  assign n30685 = n30684 ^ n12683 ^ n4595 ;
  assign n30683 = n22812 ^ n9009 ^ n6606 ;
  assign n30686 = n30685 ^ n30683 ^ n30389 ;
  assign n30687 = ( n9355 & n11501 ) | ( n9355 & n13099 ) | ( n11501 & n13099 ) ;
  assign n30690 = ( n1212 & n16835 ) | ( n1212 & ~n25937 ) | ( n16835 & ~n25937 ) ;
  assign n30691 = ( n2508 & n16810 ) | ( n2508 & ~n30690 ) | ( n16810 & ~n30690 ) ;
  assign n30688 = n12895 ^ n8702 ^ n4594 ;
  assign n30689 = n30688 ^ n15780 ^ 1'b0 ;
  assign n30692 = n30691 ^ n30689 ^ n3238 ;
  assign n30693 = n8380 ^ n7991 ^ 1'b0 ;
  assign n30694 = n2980 | n30693 ;
  assign n30695 = n30694 ^ n4824 ^ n1689 ;
  assign n30696 = n30695 ^ n12818 ^ 1'b0 ;
  assign n30697 = ( n2228 & n28969 ) | ( n2228 & n30696 ) | ( n28969 & n30696 ) ;
  assign n30698 = ( n2436 & ~n20352 ) | ( n2436 & n23322 ) | ( ~n20352 & n23322 ) ;
  assign n30699 = ( n6736 & n17024 ) | ( n6736 & n30698 ) | ( n17024 & n30698 ) ;
  assign n30700 = ( n7911 & n12275 ) | ( n7911 & n30699 ) | ( n12275 & n30699 ) ;
  assign n30701 = n9194 ^ n2736 ^ 1'b0 ;
  assign n30702 = ( n1531 & ~n10134 ) | ( n1531 & n14401 ) | ( ~n10134 & n14401 ) ;
  assign n30703 = ( n4554 & n6181 ) | ( n4554 & ~n9933 ) | ( n6181 & ~n9933 ) ;
  assign n30704 = n30703 ^ n24148 ^ n12768 ;
  assign n30705 = n30704 ^ n17875 ^ n6224 ;
  assign n30706 = ( n3032 & ~n10272 ) | ( n3032 & n19394 ) | ( ~n10272 & n19394 ) ;
  assign n30707 = n30706 ^ n18356 ^ n12578 ;
  assign n30708 = n6920 | n30707 ;
  assign n30709 = n30705 | n30708 ;
  assign n30710 = ( n19632 & ~n30702 ) | ( n19632 & n30709 ) | ( ~n30702 & n30709 ) ;
  assign n30711 = n5682 & ~n8622 ;
  assign n30712 = n30711 ^ n5779 ^ n1208 ;
  assign n30713 = ( n2690 & n4883 ) | ( n2690 & n13231 ) | ( n4883 & n13231 ) ;
  assign n30714 = ( ~n14200 & n21041 ) | ( ~n14200 & n30713 ) | ( n21041 & n30713 ) ;
  assign n30715 = ( n1660 & n30712 ) | ( n1660 & ~n30714 ) | ( n30712 & ~n30714 ) ;
  assign n30716 = ( ~n7406 & n11298 ) | ( ~n7406 & n17560 ) | ( n11298 & n17560 ) ;
  assign n30717 = n30716 ^ n10834 ^ n7855 ;
  assign n30718 = ( n14583 & n20694 ) | ( n14583 & ~n30717 ) | ( n20694 & ~n30717 ) ;
  assign n30719 = ~n678 & n10947 ;
  assign n30720 = n2290 & n30719 ;
  assign n30721 = n2453 & ~n3778 ;
  assign n30722 = n30721 ^ n16134 ^ 1'b0 ;
  assign n30723 = n28508 ^ n6202 ^ n4539 ;
  assign n30724 = n30723 ^ n27086 ^ n14655 ;
  assign n30725 = n7491 & ~n12039 ;
  assign n30726 = n15823 & ~n30725 ;
  assign n30727 = ( n12261 & ~n23190 ) | ( n12261 & n27147 ) | ( ~n23190 & n27147 ) ;
  assign n30728 = ( n4051 & n30726 ) | ( n4051 & n30727 ) | ( n30726 & n30727 ) ;
  assign n30729 = ( n8059 & n9848 ) | ( n8059 & ~n17385 ) | ( n9848 & ~n17385 ) ;
  assign n30730 = n17695 ^ n8648 ^ n4532 ;
  assign n30731 = ( n3655 & n3950 ) | ( n3655 & ~n27601 ) | ( n3950 & ~n27601 ) ;
  assign n30732 = n19782 ^ n6310 ^ 1'b0 ;
  assign n30733 = n30732 ^ n29810 ^ n19978 ;
  assign n30734 = ( n757 & n13337 ) | ( n757 & n30733 ) | ( n13337 & n30733 ) ;
  assign n30735 = n15036 ^ n13414 ^ n7392 ;
  assign n30736 = n30735 ^ n23291 ^ n4672 ;
  assign n30737 = ~n13765 & n18630 ;
  assign n30738 = ~n10929 & n30737 ;
  assign n30739 = n30738 ^ n27708 ^ n4877 ;
  assign n30740 = ~n3007 & n4135 ;
  assign n30741 = n30740 ^ n8081 ^ 1'b0 ;
  assign n30742 = ( n3184 & ~n6519 ) | ( n3184 & n19388 ) | ( ~n6519 & n19388 ) ;
  assign n30743 = n30742 ^ n12251 ^ 1'b0 ;
  assign n30744 = ( ~n2912 & n4387 ) | ( ~n2912 & n11906 ) | ( n4387 & n11906 ) ;
  assign n30745 = n30744 ^ n3408 ^ 1'b0 ;
  assign n30746 = n30745 ^ n22013 ^ n11595 ;
  assign n30749 = x53 & ~n8962 ;
  assign n30750 = n30749 ^ n9709 ^ 1'b0 ;
  assign n30747 = n12264 ^ n8247 ^ n8080 ;
  assign n30748 = n30747 ^ n26342 ^ n13494 ;
  assign n30751 = n30750 ^ n30748 ^ n8529 ;
  assign n30752 = n13421 | n13633 ;
  assign n30753 = n30752 ^ n29764 ^ n13064 ;
  assign n30754 = n20190 ^ n16923 ^ n2195 ;
  assign n30755 = ( ~n5747 & n10792 ) | ( ~n5747 & n30754 ) | ( n10792 & n30754 ) ;
  assign n30760 = n9695 ^ n6443 ^ n1069 ;
  assign n30761 = ( n8395 & n11069 ) | ( n8395 & n30760 ) | ( n11069 & n30760 ) ;
  assign n30762 = n30761 ^ n20265 ^ n19419 ;
  assign n30763 = n30762 ^ n29865 ^ n9297 ;
  assign n30756 = ~n8748 & n28910 ;
  assign n30757 = n30756 ^ n11896 ^ 1'b0 ;
  assign n30758 = n9744 ^ n3830 ^ 1'b0 ;
  assign n30759 = ~n30757 & n30758 ;
  assign n30764 = n30763 ^ n30759 ^ n6484 ;
  assign n30765 = n10407 ^ n6818 ^ n5159 ;
  assign n30766 = ( n3818 & n20353 ) | ( n3818 & ~n30765 ) | ( n20353 & ~n30765 ) ;
  assign n30767 = ( ~n6809 & n13544 ) | ( ~n6809 & n30766 ) | ( n13544 & n30766 ) ;
  assign n30768 = ( n133 & ~n4356 ) | ( n133 & n9512 ) | ( ~n4356 & n9512 ) ;
  assign n30769 = ( n5429 & ~n23269 ) | ( n5429 & n30768 ) | ( ~n23269 & n30768 ) ;
  assign n30770 = ( n11688 & ~n13134 ) | ( n11688 & n30769 ) | ( ~n13134 & n30769 ) ;
  assign n30771 = ( ~n6667 & n20762 ) | ( ~n6667 & n29735 ) | ( n20762 & n29735 ) ;
  assign n30772 = ( n10298 & ~n14418 ) | ( n10298 & n14955 ) | ( ~n14418 & n14955 ) ;
  assign n30773 = n30772 ^ n5154 ^ 1'b0 ;
  assign n30776 = n9025 | n9397 ;
  assign n30777 = n27810 ^ n13134 ^ n1059 ;
  assign n30778 = ( n2115 & n30776 ) | ( n2115 & n30777 ) | ( n30776 & n30777 ) ;
  assign n30774 = n30367 ^ n15445 ^ n2901 ;
  assign n30775 = n2031 | n30774 ;
  assign n30779 = n30778 ^ n30775 ^ 1'b0 ;
  assign n30780 = n12308 ^ n9593 ^ 1'b0 ;
  assign n30781 = n30780 ^ n19354 ^ n14267 ;
  assign n30782 = n6592 | n11115 ;
  assign n30783 = n22453 & ~n30782 ;
  assign n30784 = ( n12110 & n23893 ) | ( n12110 & ~n27567 ) | ( n23893 & ~n27567 ) ;
  assign n30785 = ( n4633 & ~n30783 ) | ( n4633 & n30784 ) | ( ~n30783 & n30784 ) ;
  assign n30786 = ( x69 & n7274 ) | ( x69 & ~n14473 ) | ( n7274 & ~n14473 ) ;
  assign n30789 = ( n2932 & n10371 ) | ( n2932 & ~n10808 ) | ( n10371 & ~n10808 ) ;
  assign n30787 = n20447 ^ n384 ^ 1'b0 ;
  assign n30788 = n30787 ^ n18462 ^ n12852 ;
  assign n30790 = n30789 ^ n30788 ^ n9200 ;
  assign n30792 = ( ~n1755 & n13418 ) | ( ~n1755 & n14884 ) | ( n13418 & n14884 ) ;
  assign n30791 = ( n7203 & n24465 ) | ( n7203 & ~n27514 ) | ( n24465 & ~n27514 ) ;
  assign n30793 = n30792 ^ n30791 ^ n10956 ;
  assign n30794 = n30793 ^ n19174 ^ n13364 ;
  assign n30795 = n17619 ^ n8096 ^ 1'b0 ;
  assign n30796 = n25456 ^ n9810 ^ n1824 ;
  assign n30797 = n28177 ^ n6710 ^ 1'b0 ;
  assign n30798 = n1847 & n16403 ;
  assign n30799 = ( n9883 & n27700 ) | ( n9883 & ~n30798 ) | ( n27700 & ~n30798 ) ;
  assign n30800 = n8843 ^ n2129 ^ 1'b0 ;
  assign n30801 = n6241 & ~n30800 ;
  assign n30802 = n16967 ^ n7162 ^ 1'b0 ;
  assign n30803 = ~n20477 & n30802 ;
  assign n30804 = ( n12052 & n12975 ) | ( n12052 & ~n17404 ) | ( n12975 & ~n17404 ) ;
  assign n30805 = n12197 ^ n6299 ^ n4494 ;
  assign n30806 = n30805 ^ n10745 ^ n1187 ;
  assign n30807 = n28616 ^ n17830 ^ n1889 ;
  assign n30808 = n15913 ^ n1417 ^ n665 ;
  assign n30809 = n10664 ^ n6179 ^ n1340 ;
  assign n30810 = n14969 ^ n3395 ^ 1'b0 ;
  assign n30811 = n14096 & n30810 ;
  assign n30812 = ( n6026 & ~n30809 ) | ( n6026 & n30811 ) | ( ~n30809 & n30811 ) ;
  assign n30813 = ( n14959 & n28965 ) | ( n14959 & n30812 ) | ( n28965 & n30812 ) ;
  assign n30814 = n6200 ^ n2729 ^ 1'b0 ;
  assign n30815 = n7404 & ~n30814 ;
  assign n30816 = n30815 ^ n19057 ^ n7187 ;
  assign n30817 = n20406 ^ n17047 ^ n1842 ;
  assign n30818 = ( n9857 & ~n21167 ) | ( n9857 & n25428 ) | ( ~n21167 & n25428 ) ;
  assign n30819 = n21110 ^ n17092 ^ n9259 ;
  assign n30820 = n6629 ^ n4935 ^ 1'b0 ;
  assign n30821 = ~n7744 & n30820 ;
  assign n30822 = n30821 ^ n19178 ^ n6160 ;
  assign n30823 = n22245 & n30822 ;
  assign n30824 = n30823 ^ n19303 ^ 1'b0 ;
  assign n30825 = n7718 ^ n267 ^ 1'b0 ;
  assign n30826 = n11041 & n30825 ;
  assign n30827 = n30826 ^ n18320 ^ n898 ;
  assign n30828 = ( n10655 & ~n15461 ) | ( n10655 & n30827 ) | ( ~n15461 & n30827 ) ;
  assign n30834 = n8458 | n17262 ;
  assign n30835 = n5173 | n30834 ;
  assign n30831 = n14031 ^ n4905 ^ n3527 ;
  assign n30832 = n30831 ^ n8327 ^ n7260 ;
  assign n30829 = n1619 & ~n26776 ;
  assign n30830 = ~n6863 & n30829 ;
  assign n30833 = n30832 ^ n30830 ^ n21731 ;
  assign n30836 = n30835 ^ n30833 ^ n21096 ;
  assign n30837 = ( n4112 & ~n21789 ) | ( n4112 & n28447 ) | ( ~n21789 & n28447 ) ;
  assign n30841 = n20576 ^ n12966 ^ n10177 ;
  assign n30838 = n12190 ^ n1827 ^ x77 ;
  assign n30839 = ~n9350 & n30838 ;
  assign n30840 = n30839 ^ n12825 ^ 1'b0 ;
  assign n30842 = n30841 ^ n30840 ^ n28175 ;
  assign n30843 = n25996 ^ n24765 ^ n15347 ;
  assign n30844 = n14847 ^ n12459 ^ n5921 ;
  assign n30845 = n27937 ^ n3580 ^ 1'b0 ;
  assign n30846 = ( n22011 & n30844 ) | ( n22011 & n30845 ) | ( n30844 & n30845 ) ;
  assign n30847 = ( ~n7934 & n10015 ) | ( ~n7934 & n29305 ) | ( n10015 & n29305 ) ;
  assign n30848 = ( ~n3604 & n11631 ) | ( ~n3604 & n30847 ) | ( n11631 & n30847 ) ;
  assign n30849 = ( ~n5607 & n12645 ) | ( ~n5607 & n16028 ) | ( n12645 & n16028 ) ;
  assign n30850 = n5142 ^ n4932 ^ n4577 ;
  assign n30851 = n30850 ^ n15713 ^ n13546 ;
  assign n30852 = ( n3683 & n28928 ) | ( n3683 & n30851 ) | ( n28928 & n30851 ) ;
  assign n30853 = ( n1595 & n18976 ) | ( n1595 & n30852 ) | ( n18976 & n30852 ) ;
  assign n30854 = ( n2398 & n30849 ) | ( n2398 & n30853 ) | ( n30849 & n30853 ) ;
  assign n30856 = ( n9697 & n9804 ) | ( n9697 & ~n19375 ) | ( n9804 & ~n19375 ) ;
  assign n30855 = n27087 ^ n15069 ^ n5834 ;
  assign n30857 = n30856 ^ n30855 ^ n20333 ;
  assign n30858 = n861 & n24849 ;
  assign n30859 = n30858 ^ n15371 ^ 1'b0 ;
  assign n30860 = n12642 | n19255 ;
  assign n30861 = n14519 | n30860 ;
  assign n30862 = n11254 & ~n15436 ;
  assign n30863 = ~n9166 & n30862 ;
  assign n30864 = ( n8320 & n14826 ) | ( n8320 & n30863 ) | ( n14826 & n30863 ) ;
  assign n30865 = n30069 ^ n11894 ^ n11565 ;
  assign n30866 = n19863 ^ n3138 ^ n2695 ;
  assign n30867 = n30866 ^ n24913 ^ n9766 ;
  assign n30868 = n26659 & ~n28576 ;
  assign n30869 = ( n2733 & n15445 ) | ( n2733 & n19322 ) | ( n15445 & n19322 ) ;
  assign n30870 = n175 & ~n22683 ;
  assign n30871 = n30870 ^ n23229 ^ 1'b0 ;
  assign n30872 = n30871 ^ n16118 ^ n3465 ;
  assign n30873 = ( ~n5395 & n11386 ) | ( ~n5395 & n28910 ) | ( n11386 & n28910 ) ;
  assign n30874 = n30873 ^ n21091 ^ n11830 ;
  assign n30876 = n5977 | n15559 ;
  assign n30877 = n30876 ^ n7686 ^ 1'b0 ;
  assign n30878 = ( ~n578 & n9795 ) | ( ~n578 & n30877 ) | ( n9795 & n30877 ) ;
  assign n30875 = ( n7800 & ~n8743 ) | ( n7800 & n12774 ) | ( ~n8743 & n12774 ) ;
  assign n30879 = n30878 ^ n30875 ^ n15185 ;
  assign n30880 = ( ~n385 & n1516 ) | ( ~n385 & n7543 ) | ( n1516 & n7543 ) ;
  assign n30881 = ( n15035 & n19952 ) | ( n15035 & n30880 ) | ( n19952 & n30880 ) ;
  assign n30882 = n30881 ^ n15594 ^ 1'b0 ;
  assign n30883 = n20468 & n30882 ;
  assign n30884 = ~n1265 & n10692 ;
  assign n30885 = n30884 ^ n1705 ^ 1'b0 ;
  assign n30886 = ( n12913 & ~n13663 ) | ( n12913 & n24875 ) | ( ~n13663 & n24875 ) ;
  assign n30888 = n16020 ^ n14473 ^ n9975 ;
  assign n30889 = n30888 ^ n12523 ^ 1'b0 ;
  assign n30887 = n23376 ^ n18451 ^ n5223 ;
  assign n30890 = n30889 ^ n30887 ^ n22844 ;
  assign n30891 = n21770 ^ n19064 ^ n6339 ;
  assign n30892 = ( n11491 & n23935 ) | ( n11491 & n27547 ) | ( n23935 & n27547 ) ;
  assign n30893 = ( ~n16541 & n30891 ) | ( ~n16541 & n30892 ) | ( n30891 & n30892 ) ;
  assign n30894 = ( ~n926 & n3547 ) | ( ~n926 & n18104 ) | ( n3547 & n18104 ) ;
  assign n30895 = ( n310 & n2934 ) | ( n310 & ~n30894 ) | ( n2934 & ~n30894 ) ;
  assign n30896 = n27268 ^ n25514 ^ n6343 ;
  assign n30897 = ( n13649 & ~n21054 ) | ( n13649 & n30896 ) | ( ~n21054 & n30896 ) ;
  assign n30898 = n3120 & ~n25596 ;
  assign n30899 = n24899 ^ n8244 ^ n5780 ;
  assign n30900 = ( n13657 & n25753 ) | ( n13657 & n30899 ) | ( n25753 & n30899 ) ;
  assign n30901 = ( ~n4174 & n5144 ) | ( ~n4174 & n10878 ) | ( n5144 & n10878 ) ;
  assign n30902 = n6054 | n23980 ;
  assign n30903 = n30902 ^ n13275 ^ n10206 ;
  assign n30904 = ( n3164 & n30901 ) | ( n3164 & n30903 ) | ( n30901 & n30903 ) ;
  assign n30905 = n3917 & n10097 ;
  assign n30906 = n17845 & ~n22578 ;
  assign n30907 = n30906 ^ n297 ^ 1'b0 ;
  assign n30908 = n12280 & ~n19146 ;
  assign n30909 = n30907 & n30908 ;
  assign n30910 = n11762 ^ n3501 ^ 1'b0 ;
  assign n30911 = ( n8476 & n22087 ) | ( n8476 & n30910 ) | ( n22087 & n30910 ) ;
  assign n30912 = n29277 ^ n15621 ^ 1'b0 ;
  assign n30913 = n30912 ^ n11564 ^ n944 ;
  assign n30914 = n10355 ^ n7906 ^ n1677 ;
  assign n30915 = n22014 & n30914 ;
  assign n30916 = n24497 ^ n14363 ^ 1'b0 ;
  assign n30917 = n17087 ^ n10232 ^ n1540 ;
  assign n30918 = n5282 ^ n4327 ^ n3711 ;
  assign n30919 = n12128 ^ n6833 ^ n5811 ;
  assign n30920 = n14145 ^ n11919 ^ n7202 ;
  assign n30921 = ( n21740 & n22431 ) | ( n21740 & n28475 ) | ( n22431 & n28475 ) ;
  assign n30922 = n11232 | n14533 ;
  assign n30923 = n30922 ^ n8030 ^ 1'b0 ;
  assign n30924 = n13746 ^ n12040 ^ 1'b0 ;
  assign n30925 = n10882 & n30924 ;
  assign n30926 = n25261 ^ n19399 ^ n1574 ;
  assign n30928 = n12497 ^ n11939 ^ n8634 ;
  assign n30927 = ( n4325 & n5646 ) | ( n4325 & n28569 ) | ( n5646 & n28569 ) ;
  assign n30929 = n30928 ^ n30927 ^ n983 ;
  assign n30930 = ( n1930 & n15494 ) | ( n1930 & n24887 ) | ( n15494 & n24887 ) ;
  assign n30931 = n30930 ^ n805 ^ 1'b0 ;
  assign n30932 = n30880 ^ n21898 ^ n7365 ;
  assign n30933 = n18807 ^ n749 ^ x56 ;
  assign n30934 = ( ~n18844 & n21006 ) | ( ~n18844 & n30933 ) | ( n21006 & n30933 ) ;
  assign n30935 = ( ~n933 & n4409 ) | ( ~n933 & n27113 ) | ( n4409 & n27113 ) ;
  assign n30936 = n30935 ^ n22633 ^ n15659 ;
  assign n30937 = ( n9998 & ~n27439 ) | ( n9998 & n30936 ) | ( ~n27439 & n30936 ) ;
  assign n30938 = ( n8728 & n14075 ) | ( n8728 & n23610 ) | ( n14075 & n23610 ) ;
  assign n30939 = n30938 ^ n18369 ^ n13652 ;
  assign n30940 = n10942 ^ n10670 ^ n9689 ;
  assign n30941 = ( n2393 & ~n7545 ) | ( n2393 & n28971 ) | ( ~n7545 & n28971 ) ;
  assign n30942 = ~n30940 & n30941 ;
  assign n30943 = ( n3788 & ~n15665 ) | ( n3788 & n29593 ) | ( ~n15665 & n29593 ) ;
  assign n30944 = n30943 ^ n25216 ^ n3949 ;
  assign n30945 = n5500 & ~n19844 ;
  assign n30946 = n30945 ^ n16816 ^ 1'b0 ;
  assign n30947 = ~n6610 & n12836 ;
  assign n30948 = ~n25676 & n30947 ;
  assign n30949 = n9764 & ~n30948 ;
  assign n30950 = n30949 ^ n22206 ^ 1'b0 ;
  assign n30951 = ( n9705 & n11805 ) | ( n9705 & ~n27622 ) | ( n11805 & ~n27622 ) ;
  assign n30952 = n25364 ^ n13997 ^ n9114 ;
  assign n30953 = n30952 ^ n19411 ^ n6180 ;
  assign n30954 = n17503 ^ n4117 ^ n2100 ;
  assign n30955 = n3557 ^ n986 ^ n204 ;
  assign n30956 = n2537 & n30955 ;
  assign n30957 = ( n3456 & n7171 ) | ( n3456 & n22864 ) | ( n7171 & n22864 ) ;
  assign n30958 = ( n18617 & n23286 ) | ( n18617 & n25502 ) | ( n23286 & n25502 ) ;
  assign n30959 = n12855 ^ n8305 ^ n6922 ;
  assign n30960 = ( n2288 & n6643 ) | ( n2288 & n18967 ) | ( n6643 & n18967 ) ;
  assign n30961 = ( n14204 & ~n26909 ) | ( n14204 & n30960 ) | ( ~n26909 & n30960 ) ;
  assign n30962 = n25425 ^ n19420 ^ n8538 ;
  assign n30963 = n4906 & ~n5815 ;
  assign n30964 = n30963 ^ n2449 ^ 1'b0 ;
  assign n30965 = ~n19037 & n23511 ;
  assign n30966 = n30965 ^ n21096 ^ 1'b0 ;
  assign n30967 = ( n6946 & n8520 ) | ( n6946 & ~n30966 ) | ( n8520 & ~n30966 ) ;
  assign n30968 = n30967 ^ n30008 ^ n23022 ;
  assign n30969 = ( ~n2938 & n9016 ) | ( ~n2938 & n19034 ) | ( n9016 & n19034 ) ;
  assign n30970 = ( n4091 & n25965 ) | ( n4091 & n30969 ) | ( n25965 & n30969 ) ;
  assign n30971 = ( n12789 & n18789 ) | ( n12789 & n26745 ) | ( n18789 & n26745 ) ;
  assign n30972 = n9510 ^ n9264 ^ n3258 ;
  assign n30973 = n30972 ^ n19576 ^ n7852 ;
  assign n30974 = n4229 | n20772 ;
  assign n30975 = n30974 ^ n22265 ^ 1'b0 ;
  assign n30976 = ( n10410 & n30973 ) | ( n10410 & ~n30975 ) | ( n30973 & ~n30975 ) ;
  assign n30977 = n11656 ^ n10546 ^ 1'b0 ;
  assign n30978 = ( n1758 & ~n2718 ) | ( n1758 & n4884 ) | ( ~n2718 & n4884 ) ;
  assign n30979 = ( n11446 & n16655 ) | ( n11446 & n30978 ) | ( n16655 & n30978 ) ;
  assign n30980 = n7612 ^ n5306 ^ n1836 ;
  assign n30981 = n30980 ^ n8107 ^ x62 ;
  assign n30982 = ( ~n16529 & n28719 ) | ( ~n16529 & n30981 ) | ( n28719 & n30981 ) ;
  assign n30983 = n1436 & n12657 ;
  assign n30984 = n30983 ^ n28787 ^ n1352 ;
  assign n30985 = n7697 & ~n23376 ;
  assign n30986 = n19904 & ~n21487 ;
  assign n30987 = n23998 & n30986 ;
  assign n30988 = ( n387 & ~n1908 ) | ( n387 & n3330 ) | ( ~n1908 & n3330 ) ;
  assign n30989 = n2884 | n8755 ;
  assign n30990 = n30989 ^ n16875 ^ 1'b0 ;
  assign n30991 = n5021 ^ n2689 ^ 1'b0 ;
  assign n30992 = n30990 & n30991 ;
  assign n30993 = ( n26164 & ~n30988 ) | ( n26164 & n30992 ) | ( ~n30988 & n30992 ) ;
  assign n30994 = n15983 ^ n9857 ^ n4301 ;
  assign n30995 = n30994 ^ n5084 ^ n4086 ;
  assign n30996 = ~n3227 & n5254 ;
  assign n30997 = n6269 & n30996 ;
  assign n30998 = ( ~n6039 & n22670 ) | ( ~n6039 & n30997 ) | ( n22670 & n30997 ) ;
  assign n31000 = ( ~n1225 & n7785 ) | ( ~n1225 & n19295 ) | ( n7785 & n19295 ) ;
  assign n30999 = ( n17101 & n22342 ) | ( n17101 & ~n22872 ) | ( n22342 & ~n22872 ) ;
  assign n31001 = n31000 ^ n30999 ^ n2568 ;
  assign n31002 = n13265 ^ n7887 ^ n4651 ;
  assign n31003 = ( n7956 & n22959 ) | ( n7956 & ~n31002 ) | ( n22959 & ~n31002 ) ;
  assign n31004 = ( n771 & n10039 ) | ( n771 & ~n31003 ) | ( n10039 & ~n31003 ) ;
  assign n31005 = ( n5103 & n13410 ) | ( n5103 & n26830 ) | ( n13410 & n26830 ) ;
  assign n31006 = n31005 ^ n8776 ^ n2388 ;
  assign n31007 = ( n13114 & ~n30667 ) | ( n13114 & n31006 ) | ( ~n30667 & n31006 ) ;
  assign n31008 = n5828 ^ n1483 ^ 1'b0 ;
  assign n31009 = ( ~n171 & n1797 ) | ( ~n171 & n31008 ) | ( n1797 & n31008 ) ;
  assign n31012 = ( n4614 & n5994 ) | ( n4614 & n12134 ) | ( n5994 & n12134 ) ;
  assign n31011 = n13319 ^ n9953 ^ n893 ;
  assign n31010 = ( n12741 & ~n20689 ) | ( n12741 & n21361 ) | ( ~n20689 & n21361 ) ;
  assign n31013 = n31012 ^ n31011 ^ n31010 ;
  assign n31014 = ( n15849 & n24116 ) | ( n15849 & ~n29497 ) | ( n24116 & ~n29497 ) ;
  assign n31015 = ( n374 & n1646 ) | ( n374 & ~n2924 ) | ( n1646 & ~n2924 ) ;
  assign n31016 = n6747 ^ n6534 ^ n5012 ;
  assign n31017 = ( n11264 & ~n31015 ) | ( n11264 & n31016 ) | ( ~n31015 & n31016 ) ;
  assign n31018 = n7125 & ~n31017 ;
  assign n31019 = n31018 ^ n13568 ^ 1'b0 ;
  assign n31020 = ( n4112 & n14640 ) | ( n4112 & n27508 ) | ( n14640 & n27508 ) ;
  assign n31021 = n27510 ^ n10897 ^ n6630 ;
  assign n31022 = ( ~n16592 & n23362 ) | ( ~n16592 & n23729 ) | ( n23362 & n23729 ) ;
  assign n31023 = ( ~n1573 & n9097 ) | ( ~n1573 & n24017 ) | ( n9097 & n24017 ) ;
  assign n31024 = n10235 ^ n9112 ^ n4246 ;
  assign n31025 = ~n3762 & n4764 ;
  assign n31026 = ~n2871 & n31025 ;
  assign n31027 = n31026 ^ n13915 ^ n7498 ;
  assign n31028 = n5494 & ~n18604 ;
  assign n31029 = n31028 ^ n8478 ^ n5724 ;
  assign n31030 = ~n31027 & n31029 ;
  assign n31031 = n29211 ^ n4121 ^ n1208 ;
  assign n31032 = ( n15856 & ~n15907 ) | ( n15856 & n23036 ) | ( ~n15907 & n23036 ) ;
  assign n31033 = ( n3528 & n6154 ) | ( n3528 & n16422 ) | ( n6154 & n16422 ) ;
  assign n31034 = n4325 & ~n18056 ;
  assign n31035 = n31034 ^ n4769 ^ 1'b0 ;
  assign n31036 = ( ~n11907 & n25764 ) | ( ~n11907 & n31035 ) | ( n25764 & n31035 ) ;
  assign n31037 = ( n6057 & n31033 ) | ( n6057 & n31036 ) | ( n31033 & n31036 ) ;
  assign n31038 = ( ~n5745 & n10124 ) | ( ~n5745 & n14965 ) | ( n10124 & n14965 ) ;
  assign n31039 = n31038 ^ n10136 ^ n3711 ;
  assign n31040 = n31039 ^ n13042 ^ n8755 ;
  assign n31041 = ( ~n3986 & n13652 ) | ( ~n3986 & n27217 ) | ( n13652 & n27217 ) ;
  assign n31042 = n31041 ^ n678 ^ 1'b0 ;
  assign n31043 = n31040 & ~n31042 ;
  assign n31044 = n3318 | n6849 ;
  assign n31045 = n31044 ^ n21207 ^ 1'b0 ;
  assign n31046 = ( n3687 & n8788 ) | ( n3687 & ~n16779 ) | ( n8788 & ~n16779 ) ;
  assign n31047 = n31046 ^ n9245 ^ n2653 ;
  assign n31048 = n31047 ^ n12833 ^ x54 ;
  assign n31049 = ( ~n5383 & n8338 ) | ( ~n5383 & n24480 ) | ( n8338 & n24480 ) ;
  assign n31050 = ( n6223 & n19417 ) | ( n6223 & ~n20724 ) | ( n19417 & ~n20724 ) ;
  assign n31051 = ( ~n2069 & n6763 ) | ( ~n2069 & n7122 ) | ( n6763 & n7122 ) ;
  assign n31052 = n31051 ^ n22375 ^ n344 ;
  assign n31053 = n6143 ^ n3558 ^ n2135 ;
  assign n31054 = n31053 ^ n15252 ^ n7363 ;
  assign n31055 = n31054 ^ n28828 ^ n10726 ;
  assign n31056 = n24901 ^ n10232 ^ n5638 ;
  assign n31057 = ( n12363 & n18706 ) | ( n12363 & n31056 ) | ( n18706 & n31056 ) ;
  assign n31061 = ( ~n2471 & n5823 ) | ( ~n2471 & n28861 ) | ( n5823 & n28861 ) ;
  assign n31058 = ( n10539 & n12758 ) | ( n10539 & n23101 ) | ( n12758 & n23101 ) ;
  assign n31059 = ( n6874 & ~n21152 ) | ( n6874 & n31058 ) | ( ~n21152 & n31058 ) ;
  assign n31060 = ( n16484 & ~n25456 ) | ( n16484 & n31059 ) | ( ~n25456 & n31059 ) ;
  assign n31062 = n31061 ^ n31060 ^ 1'b0 ;
  assign n31063 = n17220 ^ n4658 ^ n2701 ;
  assign n31064 = ( n14099 & n15265 ) | ( n14099 & ~n31063 ) | ( n15265 & ~n31063 ) ;
  assign n31065 = n6924 & n15745 ;
  assign n31066 = n30843 ^ n30631 ^ 1'b0 ;
  assign n31067 = n31065 & n31066 ;
  assign n31068 = n7562 & n16875 ;
  assign n31069 = ~n26572 & n31068 ;
  assign n31070 = ( ~n2414 & n10280 ) | ( ~n2414 & n20920 ) | ( n10280 & n20920 ) ;
  assign n31071 = ~n1404 & n6626 ;
  assign n31072 = n17715 & n31071 ;
  assign n31073 = ( n15496 & n24775 ) | ( n15496 & ~n31072 ) | ( n24775 & ~n31072 ) ;
  assign n31074 = ( ~n24905 & n31070 ) | ( ~n24905 & n31073 ) | ( n31070 & n31073 ) ;
  assign n31075 = n21965 ^ n8608 ^ n726 ;
  assign n31076 = n31012 ^ n22560 ^ n5081 ;
  assign n31077 = ( n6855 & ~n31075 ) | ( n6855 & n31076 ) | ( ~n31075 & n31076 ) ;
  assign n31079 = ( n1902 & n2609 ) | ( n1902 & ~n12924 ) | ( n2609 & ~n12924 ) ;
  assign n31078 = n24201 ^ n17977 ^ n9917 ;
  assign n31080 = n31079 ^ n31078 ^ n10045 ;
  assign n31081 = n25792 ^ n18049 ^ n7854 ;
  assign n31082 = ( n15858 & n20229 ) | ( n15858 & n31081 ) | ( n20229 & n31081 ) ;
  assign n31083 = n8875 & ~n31082 ;
  assign n31084 = ( n147 & n11590 ) | ( n147 & n24594 ) | ( n11590 & n24594 ) ;
  assign n31085 = ( n9488 & n13842 ) | ( n9488 & ~n14637 ) | ( n13842 & ~n14637 ) ;
  assign n31086 = n31085 ^ n21041 ^ n7021 ;
  assign n31087 = ( n24366 & n29739 ) | ( n24366 & ~n31086 ) | ( n29739 & ~n31086 ) ;
  assign n31088 = n27404 ^ n24618 ^ n19566 ;
  assign n31090 = ( n5009 & n8657 ) | ( n5009 & ~n23992 ) | ( n8657 & ~n23992 ) ;
  assign n31089 = ( n9613 & ~n10376 ) | ( n9613 & n27188 ) | ( ~n10376 & n27188 ) ;
  assign n31091 = n31090 ^ n31089 ^ n22849 ;
  assign n31092 = n13832 ^ n6253 ^ 1'b0 ;
  assign n31093 = n5709 & n31092 ;
  assign n31094 = ( n17195 & ~n24359 ) | ( n17195 & n31093 ) | ( ~n24359 & n31093 ) ;
  assign n31095 = n310 & n31094 ;
  assign n31096 = ~n14796 & n31095 ;
  assign n31097 = n27648 ^ n11264 ^ n2403 ;
  assign n31098 = n174 & n31097 ;
  assign n31099 = n1461 ^ n1430 ^ 1'b0 ;
  assign n31100 = n3861 & n31099 ;
  assign n31101 = ( n2617 & ~n10121 ) | ( n2617 & n31100 ) | ( ~n10121 & n31100 ) ;
  assign n31102 = ( ~n7386 & n13708 ) | ( ~n7386 & n22398 ) | ( n13708 & n22398 ) ;
  assign n31103 = n29574 ^ n22049 ^ n16111 ;
  assign n31105 = n21966 ^ n9933 ^ n1102 ;
  assign n31106 = ( n16360 & n27052 ) | ( n16360 & n31105 ) | ( n27052 & n31105 ) ;
  assign n31104 = ( n3100 & n10166 ) | ( n3100 & n22685 ) | ( n10166 & n22685 ) ;
  assign n31107 = n31106 ^ n31104 ^ n607 ;
  assign n31108 = n29057 ^ n17791 ^ n17045 ;
  assign n31109 = n17365 ^ n11493 ^ n9149 ;
  assign n31110 = ( n1947 & ~n4317 ) | ( n1947 & n5033 ) | ( ~n4317 & n5033 ) ;
  assign n31111 = n31110 ^ n5724 ^ n2670 ;
  assign n31112 = n24684 ^ n17655 ^ n1316 ;
  assign n31113 = ( ~n4483 & n4553 ) | ( ~n4483 & n9724 ) | ( n4553 & n9724 ) ;
  assign n31114 = ( n17432 & n31112 ) | ( n17432 & ~n31113 ) | ( n31112 & ~n31113 ) ;
  assign n31115 = ( n11311 & n31111 ) | ( n11311 & ~n31114 ) | ( n31111 & ~n31114 ) ;
  assign n31116 = n28512 ^ n18403 ^ n3121 ;
  assign n31117 = ( n14348 & n18682 ) | ( n14348 & ~n21106 ) | ( n18682 & ~n21106 ) ;
  assign n31118 = n31117 ^ n24330 ^ n5566 ;
  assign n31119 = ( n643 & ~n2539 ) | ( n643 & n10671 ) | ( ~n2539 & n10671 ) ;
  assign n31120 = ( ~n18011 & n30973 ) | ( ~n18011 & n31119 ) | ( n30973 & n31119 ) ;
  assign n31121 = n28185 ^ n16617 ^ n16299 ;
  assign n31122 = n25227 ^ n20926 ^ n11441 ;
  assign n31123 = ( n4800 & ~n7357 ) | ( n4800 & n11439 ) | ( ~n7357 & n11439 ) ;
  assign n31124 = n20662 ^ n13108 ^ n3496 ;
  assign n31125 = ( n23703 & n31123 ) | ( n23703 & n31124 ) | ( n31123 & n31124 ) ;
  assign n31126 = ( n5313 & n10776 ) | ( n5313 & ~n17235 ) | ( n10776 & ~n17235 ) ;
  assign n31127 = n17908 ^ n3545 ^ 1'b0 ;
  assign n31128 = ( n5555 & ~n8481 ) | ( n5555 & n31127 ) | ( ~n8481 & n31127 ) ;
  assign n31129 = ( ~n18295 & n24052 ) | ( ~n18295 & n31128 ) | ( n24052 & n31128 ) ;
  assign n31130 = n25612 ^ n6768 ^ n4708 ;
  assign n31131 = n31130 ^ n14440 ^ 1'b0 ;
  assign n31132 = n8309 & ~n8999 ;
  assign n31133 = n31132 ^ n4238 ^ 1'b0 ;
  assign n31134 = n16288 ^ n2146 ^ 1'b0 ;
  assign n31135 = n18247 | n31134 ;
  assign n31136 = n31135 ^ n21455 ^ 1'b0 ;
  assign n31137 = n19780 ^ n13144 ^ n555 ;
  assign n31138 = ( n4143 & n13814 ) | ( n4143 & n29225 ) | ( n13814 & n29225 ) ;
  assign n31139 = ( n30121 & ~n31137 ) | ( n30121 & n31138 ) | ( ~n31137 & n31138 ) ;
  assign n31140 = ( n3959 & ~n4785 ) | ( n3959 & n7224 ) | ( ~n4785 & n7224 ) ;
  assign n31141 = n31140 ^ n4508 ^ 1'b0 ;
  assign n31142 = ~n13355 & n31141 ;
  assign n31143 = n31142 ^ n28958 ^ n25926 ;
  assign n31144 = ( n5469 & n10310 ) | ( n5469 & n15417 ) | ( n10310 & n15417 ) ;
  assign n31145 = n14097 ^ n12533 ^ n3266 ;
  assign n31146 = n31145 ^ n30750 ^ n29855 ;
  assign n31147 = ( n5667 & n15540 ) | ( n5667 & ~n31146 ) | ( n15540 & ~n31146 ) ;
  assign n31148 = ( n10728 & n31144 ) | ( n10728 & n31147 ) | ( n31144 & n31147 ) ;
  assign n31149 = ( n197 & ~n3011 ) | ( n197 & n6077 ) | ( ~n3011 & n6077 ) ;
  assign n31150 = ( n17323 & ~n30952 ) | ( n17323 & n31149 ) | ( ~n30952 & n31149 ) ;
  assign n31151 = ( n10725 & ~n17085 ) | ( n10725 & n30636 ) | ( ~n17085 & n30636 ) ;
  assign n31152 = n24312 ^ n23240 ^ n21227 ;
  assign n31153 = n1861 | n17460 ;
  assign n31154 = n30880 ^ n8656 ^ n1351 ;
  assign n31155 = ( ~n9441 & n9772 ) | ( ~n9441 & n31154 ) | ( n9772 & n31154 ) ;
  assign n31156 = n353 & n30047 ;
  assign n31157 = ( n13121 & ~n26609 ) | ( n13121 & n31156 ) | ( ~n26609 & n31156 ) ;
  assign n31158 = n2793 | n22448 ;
  assign n31159 = n2234 & ~n31158 ;
  assign n31160 = n9699 ^ n6981 ^ n3378 ;
  assign n31161 = ( n10457 & n21256 ) | ( n10457 & n25371 ) | ( n21256 & n25371 ) ;
  assign n31162 = ( n26226 & ~n31160 ) | ( n26226 & n31161 ) | ( ~n31160 & n31161 ) ;
  assign n31164 = ( ~n4034 & n16228 ) | ( ~n4034 & n17726 ) | ( n16228 & n17726 ) ;
  assign n31163 = n22929 ^ n10788 ^ n9818 ;
  assign n31165 = n31164 ^ n31163 ^ n13514 ;
  assign n31166 = n18691 ^ n11099 ^ n1351 ;
  assign n31167 = ( n2106 & n13456 ) | ( n2106 & n16904 ) | ( n13456 & n16904 ) ;
  assign n31168 = ( n9859 & ~n15697 ) | ( n9859 & n31167 ) | ( ~n15697 & n31167 ) ;
  assign n31169 = ( n31165 & n31166 ) | ( n31165 & n31168 ) | ( n31166 & n31168 ) ;
  assign n31170 = n29249 ^ n646 ^ 1'b0 ;
  assign n31177 = n14860 ^ n3590 ^ n764 ;
  assign n31176 = n17184 ^ n13112 ^ 1'b0 ;
  assign n31172 = ( n1532 & ~n5418 ) | ( n1532 & n9098 ) | ( ~n5418 & n9098 ) ;
  assign n31173 = n2318 & ~n31172 ;
  assign n31174 = n31173 ^ n23128 ^ 1'b0 ;
  assign n31171 = n29680 ^ n22889 ^ n5653 ;
  assign n31175 = n31174 ^ n31171 ^ n17619 ;
  assign n31178 = n31177 ^ n31176 ^ n31175 ;
  assign n31179 = n31178 ^ n9498 ^ n3028 ;
  assign n31180 = ( n15596 & n20923 ) | ( n15596 & n26244 ) | ( n20923 & n26244 ) ;
  assign n31181 = ( n7107 & ~n27398 ) | ( n7107 & n31180 ) | ( ~n27398 & n31180 ) ;
  assign n31182 = ( n1954 & n2160 ) | ( n1954 & n10845 ) | ( n2160 & n10845 ) ;
  assign n31183 = ( n4785 & n25998 ) | ( n4785 & ~n31182 ) | ( n25998 & ~n31182 ) ;
  assign n31184 = ( n12275 & ~n15647 ) | ( n12275 & n31183 ) | ( ~n15647 & n31183 ) ;
  assign n31185 = ( ~n213 & n31181 ) | ( ~n213 & n31184 ) | ( n31181 & n31184 ) ;
  assign n31186 = n27874 ^ n14860 ^ n12051 ;
  assign n31187 = n19542 ^ n1707 ^ n1529 ;
  assign n31188 = n31187 ^ n23931 ^ n5705 ;
  assign n31189 = n5414 | n6409 ;
  assign n31190 = n31189 ^ n5276 ^ 1'b0 ;
  assign n31191 = ( n258 & n3456 ) | ( n258 & n15794 ) | ( n3456 & n15794 ) ;
  assign n31192 = ( n4949 & ~n9543 ) | ( n4949 & n31191 ) | ( ~n9543 & n31191 ) ;
  assign n31193 = n5425 | n31192 ;
  assign n31194 = n31193 ^ n10027 ^ 1'b0 ;
  assign n31195 = ( n3402 & ~n31190 ) | ( n3402 & n31194 ) | ( ~n31190 & n31194 ) ;
  assign n31196 = n2157 | n31195 ;
  assign n31197 = n24895 ^ n23499 ^ n13497 ;
  assign n31198 = n21025 ^ n7877 ^ n268 ;
  assign n31199 = n21613 | n31198 ;
  assign n31200 = x29 | n31199 ;
  assign n31201 = n5989 ^ n3204 ^ n881 ;
  assign n31202 = n12845 & ~n31201 ;
  assign n31203 = ( n2105 & n3532 ) | ( n2105 & ~n28656 ) | ( n3532 & ~n28656 ) ;
  assign n31204 = n15371 ^ n8131 ^ n5783 ;
  assign n31205 = ( n302 & ~n16025 ) | ( n302 & n28479 ) | ( ~n16025 & n28479 ) ;
  assign n31206 = ( n16052 & ~n31204 ) | ( n16052 & n31205 ) | ( ~n31204 & n31205 ) ;
  assign n31207 = ( n1422 & ~n13583 ) | ( n1422 & n23526 ) | ( ~n13583 & n23526 ) ;
  assign n31208 = n31207 ^ n4281 ^ n1081 ;
  assign n31209 = n15998 ^ n6751 ^ n6613 ;
  assign n31210 = n12767 ^ n8135 ^ 1'b0 ;
  assign n31211 = n31210 ^ n22272 ^ n6031 ;
  assign n31212 = n31211 ^ n28822 ^ n5653 ;
  assign n31213 = n24918 ^ n11403 ^ 1'b0 ;
  assign n31214 = ( n13520 & n16462 ) | ( n13520 & n31213 ) | ( n16462 & n31213 ) ;
  assign n31215 = n27767 ^ n17848 ^ 1'b0 ;
  assign n31216 = n13203 & ~n31215 ;
  assign n31217 = ( ~n9622 & n21838 ) | ( ~n9622 & n31216 ) | ( n21838 & n31216 ) ;
  assign n31218 = n24199 ^ n21830 ^ n10059 ;
  assign n31219 = n7496 ^ n3042 ^ n923 ;
  assign n31220 = n31219 ^ n7042 ^ n1776 ;
  assign n31221 = n31220 ^ n8054 ^ 1'b0 ;
  assign n31222 = ( n12186 & ~n18104 ) | ( n12186 & n31221 ) | ( ~n18104 & n31221 ) ;
  assign n31223 = n31218 | n31222 ;
  assign n31224 = n26074 ^ n20608 ^ n18609 ;
  assign n31225 = n1072 & ~n1220 ;
  assign n31226 = n31225 ^ n29049 ^ 1'b0 ;
  assign n31227 = n17397 ^ n15872 ^ 1'b0 ;
  assign n31228 = n21117 & ~n31227 ;
  assign n31229 = ( n13087 & n22550 ) | ( n13087 & n30438 ) | ( n22550 & n30438 ) ;
  assign n31230 = n20680 ^ n4887 ^ n446 ;
  assign n31231 = n7568 & n15402 ;
  assign n31232 = n31231 ^ n15534 ^ 1'b0 ;
  assign n31233 = ( n1334 & ~n13910 ) | ( n1334 & n31232 ) | ( ~n13910 & n31232 ) ;
  assign n31237 = n17119 ^ n6965 ^ n2945 ;
  assign n31235 = ( n4294 & n5357 ) | ( n4294 & ~n12000 ) | ( n5357 & ~n12000 ) ;
  assign n31234 = n18126 ^ n9762 ^ 1'b0 ;
  assign n31236 = n31235 ^ n31234 ^ n6633 ;
  assign n31238 = n31237 ^ n31236 ^ n28878 ;
  assign n31239 = ( n19520 & n24084 ) | ( n19520 & ~n28241 ) | ( n24084 & ~n28241 ) ;
  assign n31240 = ( n16127 & ~n26116 ) | ( n16127 & n28878 ) | ( ~n26116 & n28878 ) ;
  assign n31241 = ( n14516 & n26340 ) | ( n14516 & n31240 ) | ( n26340 & n31240 ) ;
  assign n31242 = ( n2221 & n3005 ) | ( n2221 & n4619 ) | ( n3005 & n4619 ) ;
  assign n31243 = n31242 ^ n16561 ^ n13708 ;
  assign n31244 = n16947 & n31243 ;
  assign n31245 = n31244 ^ n14741 ^ n11147 ;
  assign n31249 = n19149 ^ n10404 ^ n8126 ;
  assign n31246 = ( n4395 & n6056 ) | ( n4395 & n11715 ) | ( n6056 & n11715 ) ;
  assign n31247 = ( n7698 & n10066 ) | ( n7698 & n31246 ) | ( n10066 & n31246 ) ;
  assign n31248 = ( n22691 & n25873 ) | ( n22691 & ~n31247 ) | ( n25873 & ~n31247 ) ;
  assign n31250 = n31249 ^ n31248 ^ 1'b0 ;
  assign n31251 = n17018 ^ n11220 ^ 1'b0 ;
  assign n31252 = n9950 ^ n2847 ^ n2028 ;
  assign n31253 = ( n3588 & n13056 ) | ( n3588 & n26099 ) | ( n13056 & n26099 ) ;
  assign n31254 = n7383 ^ n6859 ^ n2403 ;
  assign n31255 = ( n14535 & n23645 ) | ( n14535 & ~n31254 ) | ( n23645 & ~n31254 ) ;
  assign n31256 = ( n31252 & n31253 ) | ( n31252 & ~n31255 ) | ( n31253 & ~n31255 ) ;
  assign n31257 = n15597 ^ n13947 ^ n13369 ;
  assign n31258 = ( n6039 & n8159 ) | ( n6039 & ~n10213 ) | ( n8159 & ~n10213 ) ;
  assign n31259 = n31258 ^ n28964 ^ n11047 ;
  assign n31260 = ( n17942 & ~n22619 ) | ( n17942 & n23561 ) | ( ~n22619 & n23561 ) ;
  assign n31261 = n31260 ^ n14340 ^ n7957 ;
  assign n31262 = n19017 ^ n12733 ^ 1'b0 ;
  assign n31263 = ( n1474 & n20739 ) | ( n1474 & ~n31262 ) | ( n20739 & ~n31262 ) ;
  assign n31264 = n31263 ^ n19477 ^ n6955 ;
  assign n31265 = ( ~n16004 & n18723 ) | ( ~n16004 & n26205 ) | ( n18723 & n26205 ) ;
  assign n31266 = ( n16474 & n26013 ) | ( n16474 & ~n30278 ) | ( n26013 & ~n30278 ) ;
  assign n31267 = ( n15864 & n19929 ) | ( n15864 & ~n31266 ) | ( n19929 & ~n31266 ) ;
  assign n31268 = n31267 ^ n27001 ^ n1594 ;
  assign n31269 = ( n11860 & n24812 ) | ( n11860 & n31268 ) | ( n24812 & n31268 ) ;
  assign n31270 = ( n773 & n29610 ) | ( n773 & ~n31269 ) | ( n29610 & ~n31269 ) ;
  assign n31271 = n23874 ^ n5743 ^ n504 ;
  assign n31272 = x48 & n20884 ;
  assign n31273 = n31272 ^ n10016 ^ 1'b0 ;
  assign n31274 = n31273 ^ n30344 ^ n7242 ;
  assign n31275 = n14616 | n22730 ;
  assign n31276 = n4642 | n31275 ;
  assign n31277 = ( n2999 & ~n13998 ) | ( n2999 & n15733 ) | ( ~n13998 & n15733 ) ;
  assign n31278 = ( ~n5080 & n8138 ) | ( ~n5080 & n13187 ) | ( n8138 & n13187 ) ;
  assign n31279 = n19598 ^ n6806 ^ n3549 ;
  assign n31280 = ( n10519 & n27832 ) | ( n10519 & n30208 ) | ( n27832 & n30208 ) ;
  assign n31281 = n31280 ^ n25383 ^ 1'b0 ;
  assign n31282 = n25657 ^ n22052 ^ n11657 ;
  assign n31283 = n9017 | n28409 ;
  assign n31284 = n31283 ^ n22259 ^ n16147 ;
  assign n31285 = n31284 ^ n19315 ^ n9905 ;
  assign n31286 = ~n7115 & n7515 ;
  assign n31287 = x78 & n31286 ;
  assign n31288 = n9587 & n31287 ;
  assign n31289 = n31288 ^ n18989 ^ n13767 ;
  assign n31290 = n22824 & n29122 ;
  assign n31291 = ( n3215 & ~n11653 ) | ( n3215 & n19301 ) | ( ~n11653 & n19301 ) ;
  assign n31292 = n31291 ^ n20491 ^ 1'b0 ;
  assign n31293 = n31292 ^ n23204 ^ 1'b0 ;
  assign n31294 = ( n1227 & n6171 ) | ( n1227 & n9415 ) | ( n6171 & n9415 ) ;
  assign n31295 = n31294 ^ n14000 ^ n13487 ;
  assign n31296 = n31295 ^ n20388 ^ n14721 ;
  assign n31297 = ( n238 & n24794 ) | ( n238 & ~n31296 ) | ( n24794 & ~n31296 ) ;
  assign n31298 = n16929 & n17912 ;
  assign n31299 = n31298 ^ n20163 ^ 1'b0 ;
  assign n31300 = ( n6310 & ~n13353 ) | ( n6310 & n31299 ) | ( ~n13353 & n31299 ) ;
  assign n31301 = n27272 ^ n20068 ^ 1'b0 ;
  assign n31302 = n19299 ^ n8339 ^ n5090 ;
  assign n31303 = n15277 ^ n5301 ^ n4625 ;
  assign n31304 = n6835 & ~n19908 ;
  assign n31305 = ( ~n10077 & n13272 ) | ( ~n10077 & n15853 ) | ( n13272 & n15853 ) ;
  assign n31306 = ( ~x15 & n4536 ) | ( ~x15 & n31305 ) | ( n4536 & n31305 ) ;
  assign n31307 = n31306 ^ n22711 ^ n6648 ;
  assign n31308 = ( n12610 & n31304 ) | ( n12610 & n31307 ) | ( n31304 & n31307 ) ;
  assign n31309 = ( n10193 & n21514 ) | ( n10193 & ~n29107 ) | ( n21514 & ~n29107 ) ;
  assign n31310 = n31309 ^ n24439 ^ n15694 ;
  assign n31311 = n20789 ^ n6970 ^ x54 ;
  assign n31312 = ( n1836 & n3945 ) | ( n1836 & n6271 ) | ( n3945 & n6271 ) ;
  assign n31313 = n31312 ^ n30421 ^ n25929 ;
  assign n31314 = ( ~n2062 & n19956 ) | ( ~n2062 & n25684 ) | ( n19956 & n25684 ) ;
  assign n31315 = n28696 ^ n3838 ^ 1'b0 ;
  assign n31316 = n31314 & ~n31315 ;
  assign n31317 = n661 & ~n3283 ;
  assign n31318 = n31317 ^ n30198 ^ n23048 ;
  assign n31319 = ( n1377 & n5886 ) | ( n1377 & ~n14920 ) | ( n5886 & ~n14920 ) ;
  assign n31320 = ( n2673 & n4367 ) | ( n2673 & n7390 ) | ( n4367 & n7390 ) ;
  assign n31321 = n17731 ^ n8215 ^ 1'b0 ;
  assign n31322 = n16968 | n31321 ;
  assign n31323 = n12018 & ~n31322 ;
  assign n31324 = n31201 & n31323 ;
  assign n31325 = ( n31319 & ~n31320 ) | ( n31319 & n31324 ) | ( ~n31320 & n31324 ) ;
  assign n31326 = n31325 ^ n14034 ^ n10369 ;
  assign n31327 = n8643 ^ n3605 ^ n2269 ;
  assign n31328 = n31327 ^ n30757 ^ n13009 ;
  assign n31332 = n5134 | n11323 ;
  assign n31329 = ( n2492 & n8155 ) | ( n2492 & ~n13832 ) | ( n8155 & ~n13832 ) ;
  assign n31330 = n31329 ^ n25987 ^ n12087 ;
  assign n31331 = ( n11051 & n16006 ) | ( n11051 & ~n31330 ) | ( n16006 & ~n31330 ) ;
  assign n31333 = n31332 ^ n31331 ^ n8355 ;
  assign n31335 = ( n1669 & n7618 ) | ( n1669 & ~n12134 ) | ( n7618 & ~n12134 ) ;
  assign n31336 = n1410 & n31123 ;
  assign n31337 = ~n31335 & n31336 ;
  assign n31338 = ( n3522 & n9239 ) | ( n3522 & n31337 ) | ( n9239 & n31337 ) ;
  assign n31334 = n30849 ^ n14889 ^ n12459 ;
  assign n31339 = n31338 ^ n31334 ^ 1'b0 ;
  assign n31340 = n4066 ^ n2350 ^ n874 ;
  assign n31341 = ( ~n1467 & n15305 ) | ( ~n1467 & n31340 ) | ( n15305 & n31340 ) ;
  assign n31342 = ( n1237 & n20337 ) | ( n1237 & ~n22932 ) | ( n20337 & ~n22932 ) ;
  assign n31343 = n31342 ^ n27279 ^ x17 ;
  assign n31344 = ( n7580 & n10098 ) | ( n7580 & n21854 ) | ( n10098 & n21854 ) ;
  assign n31345 = ( n2849 & n10356 ) | ( n2849 & ~n31344 ) | ( n10356 & ~n31344 ) ;
  assign n31346 = n26353 ^ n24382 ^ n4851 ;
  assign n31347 = n24462 ^ n7391 ^ 1'b0 ;
  assign n31348 = n2824 & n31347 ;
  assign n31349 = ( n10345 & n11617 ) | ( n10345 & ~n19699 ) | ( n11617 & ~n19699 ) ;
  assign n31350 = n31349 ^ n29245 ^ n28732 ;
  assign n31351 = n5703 ^ n4772 ^ 1'b0 ;
  assign n31352 = ~n29653 & n31351 ;
  assign n31353 = ( ~n8835 & n10931 ) | ( ~n8835 & n31352 ) | ( n10931 & n31352 ) ;
  assign n31354 = n20281 ^ n6020 ^ n2952 ;
  assign n31355 = ( n16413 & n19369 ) | ( n16413 & ~n29884 ) | ( n19369 & ~n29884 ) ;
  assign n31356 = ( n9371 & n14689 ) | ( n9371 & ~n23611 ) | ( n14689 & ~n23611 ) ;
  assign n31357 = n31356 ^ n7337 ^ n4041 ;
  assign n31358 = n5800 ^ n3853 ^ n2005 ;
  assign n31359 = n31358 ^ n1515 ^ 1'b0 ;
  assign n31360 = ( n4828 & n12674 ) | ( n4828 & n20816 ) | ( n12674 & n20816 ) ;
  assign n31361 = n31360 ^ n13671 ^ n5738 ;
  assign n31362 = n31361 ^ n15255 ^ 1'b0 ;
  assign n31363 = ( ~n6494 & n10355 ) | ( ~n6494 & n10828 ) | ( n10355 & n10828 ) ;
  assign n31364 = n18342 ^ n16131 ^ 1'b0 ;
  assign n31365 = n13808 & ~n31364 ;
  assign n31366 = ( n7617 & ~n28362 ) | ( n7617 & n31365 ) | ( ~n28362 & n31365 ) ;
  assign n31367 = ( n7317 & ~n9042 ) | ( n7317 & n31366 ) | ( ~n9042 & n31366 ) ;
  assign n31368 = ( n7563 & n26069 ) | ( n7563 & ~n31367 ) | ( n26069 & ~n31367 ) ;
  assign n31369 = ~n6616 & n15783 ;
  assign n31370 = n1270 & n31369 ;
  assign n31371 = n5599 ^ n4313 ^ 1'b0 ;
  assign n31372 = ( n11684 & n12059 ) | ( n11684 & ~n31371 ) | ( n12059 & ~n31371 ) ;
  assign n31373 = ( ~n6047 & n8217 ) | ( ~n6047 & n31372 ) | ( n8217 & n31372 ) ;
  assign n31374 = n28733 ^ n28352 ^ n25807 ;
  assign n31375 = ( n26307 & ~n29874 ) | ( n26307 & n31374 ) | ( ~n29874 & n31374 ) ;
  assign n31376 = ( n7547 & n24858 ) | ( n7547 & n25122 ) | ( n24858 & n25122 ) ;
  assign n31377 = ( n1778 & n14769 ) | ( n1778 & ~n31376 ) | ( n14769 & ~n31376 ) ;
  assign n31378 = ( n1242 & ~n18312 ) | ( n1242 & n28888 ) | ( ~n18312 & n28888 ) ;
  assign n31379 = n31378 ^ n19580 ^ n1102 ;
  assign n31380 = n28476 ^ n12769 ^ n2293 ;
  assign n31381 = ( n7301 & n14610 ) | ( n7301 & ~n31380 ) | ( n14610 & ~n31380 ) ;
  assign n31382 = ( n12443 & n14502 ) | ( n12443 & ~n26516 ) | ( n14502 & ~n26516 ) ;
  assign n31383 = ~n1206 & n2669 ;
  assign n31384 = ( n2197 & n7595 ) | ( n2197 & ~n31383 ) | ( n7595 & ~n31383 ) ;
  assign n31385 = ( n3545 & ~n15611 ) | ( n3545 & n22619 ) | ( ~n15611 & n22619 ) ;
  assign n31386 = n31385 ^ n27747 ^ n14046 ;
  assign n31387 = ( ~n5986 & n31384 ) | ( ~n5986 & n31386 ) | ( n31384 & n31386 ) ;
  assign n31388 = n31094 ^ n21798 ^ n3002 ;
  assign n31389 = n4325 & n14579 ;
  assign n31390 = n31389 ^ n7746 ^ n5019 ;
  assign n31391 = ~n12538 & n14136 ;
  assign n31392 = n31391 ^ n23227 ^ 1'b0 ;
  assign n31393 = n27630 ^ n9924 ^ 1'b0 ;
  assign n31394 = n29875 & n31393 ;
  assign n31395 = ( n1603 & n2831 ) | ( n1603 & n3989 ) | ( n2831 & n3989 ) ;
  assign n31396 = n31395 ^ n11885 ^ n5806 ;
  assign n31397 = n16364 ^ n11332 ^ 1'b0 ;
  assign n31398 = n8364 ^ n5916 ^ n5604 ;
  assign n31399 = ( ~n2536 & n5946 ) | ( ~n2536 & n7150 ) | ( n5946 & n7150 ) ;
  assign n31400 = n16368 ^ n7718 ^ n835 ;
  assign n31401 = n31400 ^ n9359 ^ n3101 ;
  assign n31402 = ( n31398 & ~n31399 ) | ( n31398 & n31401 ) | ( ~n31399 & n31401 ) ;
  assign n31403 = ( n14366 & n16319 ) | ( n14366 & n31402 ) | ( n16319 & n31402 ) ;
  assign n31404 = ( n3280 & n6415 ) | ( n3280 & ~n11652 ) | ( n6415 & ~n11652 ) ;
  assign n31405 = n29259 ^ n26751 ^ n1602 ;
  assign n31411 = n30146 ^ n14480 ^ n2844 ;
  assign n31409 = n14472 ^ n6216 ^ n3322 ;
  assign n31407 = ( ~n2929 & n3899 ) | ( ~n2929 & n10182 ) | ( n3899 & n10182 ) ;
  assign n31408 = n31407 ^ n23227 ^ n11251 ;
  assign n31406 = ( n3007 & n25750 ) | ( n3007 & n31192 ) | ( n25750 & n31192 ) ;
  assign n31410 = n31409 ^ n31408 ^ n31406 ;
  assign n31412 = n31411 ^ n31410 ^ 1'b0 ;
  assign n31413 = ( ~n8972 & n12962 ) | ( ~n8972 & n19776 ) | ( n12962 & n19776 ) ;
  assign n31414 = n17574 ^ n7490 ^ n447 ;
  assign n31415 = n31414 ^ n6177 ^ n2167 ;
  assign n31416 = ( n11058 & n25019 ) | ( n11058 & ~n31415 ) | ( n25019 & ~n31415 ) ;
  assign n31417 = n3030 & ~n31416 ;
  assign n31418 = n12459 ^ n12120 ^ n5557 ;
  assign n31419 = n31418 ^ n10121 ^ x58 ;
  assign n31420 = n1303 & n12163 ;
  assign n31421 = n2567 & n31420 ;
  assign n31422 = ( n19632 & n31419 ) | ( n19632 & ~n31421 ) | ( n31419 & ~n31421 ) ;
  assign n31423 = ( ~n17172 & n20327 ) | ( ~n17172 & n23931 ) | ( n20327 & n23931 ) ;
  assign n31424 = n3818 ^ n3181 ^ n860 ;
  assign n31425 = n31424 ^ n3376 ^ 1'b0 ;
  assign n31426 = n31423 & n31425 ;
  assign n31427 = ( n1735 & n10211 ) | ( n1735 & n24977 ) | ( n10211 & n24977 ) ;
  assign n31428 = n13055 ^ n12512 ^ n1431 ;
  assign n31429 = n31428 ^ n30548 ^ n3860 ;
  assign n31430 = ( n2053 & n3884 ) | ( n2053 & ~n26422 ) | ( n3884 & ~n26422 ) ;
  assign n31431 = n11776 ^ n7484 ^ 1'b0 ;
  assign n31432 = n31430 & ~n31431 ;
  assign n31433 = n6429 & n9247 ;
  assign n31434 = ( n12751 & n13504 ) | ( n12751 & ~n31433 ) | ( n13504 & ~n31433 ) ;
  assign n31435 = ( n31429 & n31432 ) | ( n31429 & ~n31434 ) | ( n31432 & ~n31434 ) ;
  assign n31436 = n28703 ^ n8759 ^ n3036 ;
  assign n31437 = ( ~n3402 & n16373 ) | ( ~n3402 & n18269 ) | ( n16373 & n18269 ) ;
  assign n31438 = ~n8038 & n24382 ;
  assign n31439 = n31438 ^ n4224 ^ 1'b0 ;
  assign n31440 = n31439 ^ n8492 ^ n2251 ;
  assign n31441 = ( n3875 & ~n7057 ) | ( n3875 & n17779 ) | ( ~n7057 & n17779 ) ;
  assign n31442 = n30379 ^ n21264 ^ n1300 ;
  assign n31443 = n20061 ^ n6674 ^ 1'b0 ;
  assign n31449 = ( ~n5091 & n13827 ) | ( ~n5091 & n17635 ) | ( n13827 & n17635 ) ;
  assign n31444 = n20078 ^ n14130 ^ n11314 ;
  assign n31445 = n31444 ^ n3021 ^ 1'b0 ;
  assign n31446 = n7576 & n31445 ;
  assign n31447 = ( n11594 & ~n29597 ) | ( n11594 & n31446 ) | ( ~n29597 & n31446 ) ;
  assign n31448 = ( n453 & n31219 ) | ( n453 & n31447 ) | ( n31219 & n31447 ) ;
  assign n31450 = n31449 ^ n31448 ^ n22809 ;
  assign n31451 = n1440 & ~n6550 ;
  assign n31452 = ~n18443 & n31451 ;
  assign n31453 = ( ~n5077 & n15582 ) | ( ~n5077 & n18221 ) | ( n15582 & n18221 ) ;
  assign n31454 = n9818 ^ n3978 ^ n2776 ;
  assign n31455 = n10278 & n17101 ;
  assign n31456 = n13140 & n31455 ;
  assign n31457 = n31456 ^ n16419 ^ n15848 ;
  assign n31458 = ( n31453 & ~n31454 ) | ( n31453 & n31457 ) | ( ~n31454 & n31457 ) ;
  assign n31459 = ( n8702 & ~n8816 ) | ( n8702 & n15677 ) | ( ~n8816 & n15677 ) ;
  assign n31460 = n3623 ^ n3389 ^ 1'b0 ;
  assign n31461 = n28667 & ~n31460 ;
  assign n31462 = n29238 ^ n14126 ^ n5845 ;
  assign n31464 = ( ~x110 & n840 ) | ( ~x110 & n2553 ) | ( n840 & n2553 ) ;
  assign n31463 = n15801 ^ n10567 ^ 1'b0 ;
  assign n31465 = n31464 ^ n31463 ^ n7097 ;
  assign n31466 = ( n8659 & ~n9998 ) | ( n8659 & n31465 ) | ( ~n9998 & n31465 ) ;
  assign n31467 = n11243 ^ n8831 ^ 1'b0 ;
  assign n31468 = ( n4104 & n12347 ) | ( n4104 & ~n31467 ) | ( n12347 & ~n31467 ) ;
  assign n31469 = ( n11814 & n30178 ) | ( n11814 & n31468 ) | ( n30178 & n31468 ) ;
  assign n31470 = n15033 ^ n5046 ^ n4310 ;
  assign n31472 = n20945 ^ n10206 ^ n7246 ;
  assign n31471 = n19461 ^ n7373 ^ n6485 ;
  assign n31473 = n31472 ^ n31471 ^ n22631 ;
  assign n31474 = ( ~n879 & n6880 ) | ( ~n879 & n19497 ) | ( n6880 & n19497 ) ;
  assign n31477 = ( n6604 & ~n11394 ) | ( n6604 & n16297 ) | ( ~n11394 & n16297 ) ;
  assign n31475 = n26973 ^ n7908 ^ n7847 ;
  assign n31476 = n26904 & n31475 ;
  assign n31478 = n31477 ^ n31476 ^ 1'b0 ;
  assign n31479 = ( ~n1357 & n16335 ) | ( ~n1357 & n18107 ) | ( n16335 & n18107 ) ;
  assign n31480 = n9024 & n15088 ;
  assign n31481 = ( ~n10834 & n23330 ) | ( ~n10834 & n28993 ) | ( n23330 & n28993 ) ;
  assign n31482 = ( n393 & n11424 ) | ( n393 & n12876 ) | ( n11424 & n12876 ) ;
  assign n31483 = ( ~n4527 & n17840 ) | ( ~n4527 & n31482 ) | ( n17840 & n31482 ) ;
  assign n31484 = n31483 ^ n28131 ^ n19802 ;
  assign n31485 = n9590 ^ n676 ^ 1'b0 ;
  assign n31486 = ~n3719 & n31485 ;
  assign n31487 = ( ~n4354 & n29657 ) | ( ~n4354 & n31486 ) | ( n29657 & n31486 ) ;
  assign n31488 = n3256 & n19510 ;
  assign n31492 = ( n6643 & n9930 ) | ( n6643 & ~n17242 ) | ( n9930 & ~n17242 ) ;
  assign n31489 = ( ~n2694 & n23686 ) | ( ~n2694 & n28492 ) | ( n23686 & n28492 ) ;
  assign n31490 = n31489 ^ n25628 ^ n24856 ;
  assign n31491 = n31490 ^ n24953 ^ n11085 ;
  assign n31493 = n31492 ^ n31491 ^ n2473 ;
  assign n31494 = n31493 ^ n29706 ^ n12523 ;
  assign n31495 = ( ~n398 & n3629 ) | ( ~n398 & n28742 ) | ( n3629 & n28742 ) ;
  assign n31496 = n4367 & ~n8017 ;
  assign n31497 = n5621 | n12630 ;
  assign n31498 = n15933 & ~n31497 ;
  assign n31499 = n24456 ^ n20575 ^ n16183 ;
  assign n31500 = n29199 & ~n31499 ;
  assign n31501 = n31500 ^ n8735 ^ 1'b0 ;
  assign n31502 = ( n2432 & n11116 ) | ( n2432 & ~n16731 ) | ( n11116 & ~n16731 ) ;
  assign n31503 = n329 | n31502 ;
  assign n31504 = n18936 ^ n13667 ^ n2285 ;
  assign n31505 = ( n7309 & ~n10700 ) | ( n7309 & n31504 ) | ( ~n10700 & n31504 ) ;
  assign n31506 = n5275 | n21711 ;
  assign n31507 = n19202 | n31506 ;
  assign n31508 = ( n20872 & n31505 ) | ( n20872 & n31507 ) | ( n31505 & n31507 ) ;
  assign n31509 = n25032 ^ n21147 ^ n7631 ;
  assign n31510 = ( n10961 & ~n15885 ) | ( n10961 & n18219 ) | ( ~n15885 & n18219 ) ;
  assign n31511 = ( n3713 & ~n8591 ) | ( n3713 & n31510 ) | ( ~n8591 & n31510 ) ;
  assign n31512 = ( ~n2116 & n19287 ) | ( ~n2116 & n31511 ) | ( n19287 & n31511 ) ;
  assign n31514 = ( ~n4602 & n5766 ) | ( ~n4602 & n6899 ) | ( n5766 & n6899 ) ;
  assign n31513 = ( n6440 & n8425 ) | ( n6440 & ~n22567 ) | ( n8425 & ~n22567 ) ;
  assign n31515 = n31514 ^ n31513 ^ n14368 ;
  assign n31516 = n31515 ^ n29309 ^ n25784 ;
  assign n31517 = ( n4398 & n19043 ) | ( n4398 & ~n21407 ) | ( n19043 & ~n21407 ) ;
  assign n31518 = n29172 ^ n26013 ^ n14748 ;
  assign n31519 = n31518 ^ n26731 ^ n7958 ;
  assign n31520 = n9995 ^ n4515 ^ n3223 ;
  assign n31521 = n173 | n31520 ;
  assign n31522 = ( ~n17345 & n29114 ) | ( ~n17345 & n31521 ) | ( n29114 & n31521 ) ;
  assign n31523 = n31522 ^ n7515 ^ n621 ;
  assign n31525 = ( n3617 & n5934 ) | ( n3617 & ~n8772 ) | ( n5934 & ~n8772 ) ;
  assign n31524 = ( n12395 & ~n13657 ) | ( n12395 & n25760 ) | ( ~n13657 & n25760 ) ;
  assign n31526 = n31525 ^ n31524 ^ n479 ;
  assign n31527 = n5679 ^ n1687 ^ 1'b0 ;
  assign n31528 = n15139 & ~n31527 ;
  assign n31529 = ~n3560 & n17355 ;
  assign n31530 = n31529 ^ n4766 ^ 1'b0 ;
  assign n31531 = ( n142 & ~n8497 ) | ( n142 & n13180 ) | ( ~n8497 & n13180 ) ;
  assign n31532 = n4680 & n30899 ;
  assign n31533 = n11155 & n15523 ;
  assign n31534 = n1907 | n24426 ;
  assign n31536 = ( n2132 & n10590 ) | ( n2132 & ~n21607 ) | ( n10590 & ~n21607 ) ;
  assign n31535 = n7627 ^ n6476 ^ n5576 ;
  assign n31537 = n31536 ^ n31535 ^ n6184 ;
  assign n31538 = ( n23287 & n31534 ) | ( n23287 & n31537 ) | ( n31534 & n31537 ) ;
  assign n31539 = n21951 ^ n12867 ^ n1815 ;
  assign n31540 = n31539 ^ n23376 ^ n12203 ;
  assign n31541 = n31540 ^ n1985 ^ n329 ;
  assign n31542 = n31541 ^ n30930 ^ n7388 ;
  assign n31543 = n31542 ^ n25093 ^ n24011 ;
  assign n31544 = n31543 ^ n21073 ^ n6973 ;
  assign n31545 = n21727 ^ n20724 ^ n14705 ;
  assign n31546 = ( n7667 & ~n10746 ) | ( n7667 & n31545 ) | ( ~n10746 & n31545 ) ;
  assign n31547 = ( n1870 & ~n31544 ) | ( n1870 & n31546 ) | ( ~n31544 & n31546 ) ;
  assign n31548 = n9261 ^ n7345 ^ n6100 ;
  assign n31549 = n31548 ^ n30118 ^ n18924 ;
  assign n31550 = n15615 ^ n12520 ^ n1355 ;
  assign n31551 = ( n4965 & ~n21843 ) | ( n4965 & n25906 ) | ( ~n21843 & n25906 ) ;
  assign n31552 = n23039 ^ n16184 ^ n4354 ;
  assign n31553 = n25344 ^ n8655 ^ n3888 ;
  assign n31554 = n17897 & ~n31553 ;
  assign n31555 = n31554 ^ n17786 ^ 1'b0 ;
  assign n31556 = n10874 ^ n10833 ^ n5325 ;
  assign n31557 = n23324 ^ n12567 ^ 1'b0 ;
  assign n31558 = n31557 ^ n29878 ^ n14162 ;
  assign n31559 = n30830 ^ n9484 ^ 1'b0 ;
  assign n31560 = ( n6416 & ~n9415 ) | ( n6416 & n31327 ) | ( ~n9415 & n31327 ) ;
  assign n31561 = n10488 ^ n7406 ^ 1'b0 ;
  assign n31562 = n17847 & ~n31561 ;
  assign n31563 = n11323 & ~n13855 ;
  assign n31564 = ( n2930 & n3404 ) | ( n2930 & ~n31563 ) | ( n3404 & ~n31563 ) ;
  assign n31565 = n21899 ^ n12043 ^ n11019 ;
  assign n31566 = n15513 & ~n29294 ;
  assign n31567 = ( n2653 & n6316 ) | ( n2653 & n15926 ) | ( n6316 & n15926 ) ;
  assign n31568 = ( ~n11965 & n31566 ) | ( ~n11965 & n31567 ) | ( n31566 & n31567 ) ;
  assign n31569 = ( ~n8082 & n12607 ) | ( ~n8082 & n17671 ) | ( n12607 & n17671 ) ;
  assign n31570 = ( n12348 & n29400 ) | ( n12348 & ~n31569 ) | ( n29400 & ~n31569 ) ;
  assign n31571 = n4278 & ~n11404 ;
  assign n31572 = n31571 ^ n2091 ^ 1'b0 ;
  assign n31573 = n9168 ^ n7249 ^ n2503 ;
  assign n31574 = n18201 ^ n2923 ^ n1918 ;
  assign n31575 = ( n28430 & ~n29229 ) | ( n28430 & n31574 ) | ( ~n29229 & n31574 ) ;
  assign n31576 = n19859 ^ n7264 ^ n6504 ;
  assign n31577 = n9814 ^ n7508 ^ n3650 ;
  assign n31578 = n28530 ^ n13271 ^ n4062 ;
  assign n31579 = n31578 ^ n20886 ^ 1'b0 ;
  assign n31580 = ( n1902 & ~n18310 ) | ( n1902 & n30026 ) | ( ~n18310 & n30026 ) ;
  assign n31581 = ( n3796 & n15621 ) | ( n3796 & ~n19613 ) | ( n15621 & ~n19613 ) ;
  assign n31582 = ( n3548 & ~n7481 ) | ( n3548 & n8247 ) | ( ~n7481 & n8247 ) ;
  assign n31583 = ( n768 & n17135 ) | ( n768 & ~n24824 ) | ( n17135 & ~n24824 ) ;
  assign n31584 = ~n11438 & n16927 ;
  assign n31585 = n31584 ^ n24676 ^ 1'b0 ;
  assign n31586 = n17533 ^ n9096 ^ n6424 ;
  assign n31587 = ( n416 & n577 ) | ( n416 & n6840 ) | ( n577 & n6840 ) ;
  assign n31588 = ( n1377 & ~n6332 ) | ( n1377 & n23675 ) | ( ~n6332 & n23675 ) ;
  assign n31589 = ( n9670 & ~n31587 ) | ( n9670 & n31588 ) | ( ~n31587 & n31588 ) ;
  assign n31590 = n14721 ^ n10063 ^ n9351 ;
  assign n31591 = ( n13454 & ~n26567 ) | ( n13454 & n31590 ) | ( ~n26567 & n31590 ) ;
  assign n31592 = n17684 ^ n4611 ^ 1'b0 ;
  assign n31593 = ( n6040 & n9141 ) | ( n6040 & n16668 ) | ( n9141 & n16668 ) ;
  assign n31594 = n29594 ^ n18740 ^ n12206 ;
  assign n31595 = ( n26628 & ~n31593 ) | ( n26628 & n31594 ) | ( ~n31593 & n31594 ) ;
  assign n31596 = n18205 ^ n6142 ^ n3708 ;
  assign n31597 = n3527 & n19094 ;
  assign n31598 = n1354 & ~n31597 ;
  assign n31599 = ( n14123 & n16927 ) | ( n14123 & n27757 ) | ( n16927 & n27757 ) ;
  assign n31600 = n1467 & ~n26774 ;
  assign n31601 = ~n29157 & n31600 ;
  assign n31602 = n31601 ^ n1299 ^ 1'b0 ;
  assign n31603 = ~n18000 & n31602 ;
  assign n31604 = ( n2139 & ~n17286 ) | ( n2139 & n31603 ) | ( ~n17286 & n31603 ) ;
  assign n31605 = ( ~n6872 & n13617 ) | ( ~n6872 & n27911 ) | ( n13617 & n27911 ) ;
  assign n31606 = n31605 ^ n3970 ^ n3070 ;
  assign n31607 = n145 | n31606 ;
  assign n31608 = n31607 ^ n4434 ^ 1'b0 ;
  assign n31609 = n3145 & ~n9379 ;
  assign n31610 = n31609 ^ n26568 ^ 1'b0 ;
  assign n31611 = n1967 ^ n1866 ^ n698 ;
  assign n31612 = ( n3535 & n12096 ) | ( n3535 & n23197 ) | ( n12096 & n23197 ) ;
  assign n31613 = n31612 ^ n4575 ^ 1'b0 ;
  assign n31614 = n10992 & ~n15675 ;
  assign n31615 = n29441 & n31614 ;
  assign n31616 = ( n2042 & n4369 ) | ( n2042 & ~n14669 ) | ( n4369 & ~n14669 ) ;
  assign n31617 = ( n4908 & n9190 ) | ( n4908 & ~n31616 ) | ( n9190 & ~n31616 ) ;
  assign n31618 = ( n9211 & ~n13240 ) | ( n9211 & n20503 ) | ( ~n13240 & n20503 ) ;
  assign n31619 = ( n1347 & n6575 ) | ( n1347 & n31618 ) | ( n6575 & n31618 ) ;
  assign n31620 = n31619 ^ n23932 ^ n13930 ;
  assign n31621 = n24302 ^ n6450 ^ n5033 ;
  assign n31622 = n31621 ^ n26543 ^ 1'b0 ;
  assign n31623 = n15364 & ~n31622 ;
  assign n31624 = ( n2349 & ~n27042 ) | ( n2349 & n31623 ) | ( ~n27042 & n31623 ) ;
  assign n31625 = ( n12086 & n12182 ) | ( n12086 & ~n25375 ) | ( n12182 & ~n25375 ) ;
  assign n31626 = ( n775 & n13209 ) | ( n775 & n31625 ) | ( n13209 & n31625 ) ;
  assign n31627 = n13511 ^ n707 ^ 1'b0 ;
  assign n31628 = n13529 ^ n9543 ^ n1974 ;
  assign n31629 = n31628 ^ n7695 ^ 1'b0 ;
  assign n31630 = n10611 & ~n18198 ;
  assign n31631 = ~n3568 & n31630 ;
  assign n31632 = ~n1790 & n6184 ;
  assign n31633 = ( n1147 & ~n10454 ) | ( n1147 & n13482 ) | ( ~n10454 & n13482 ) ;
  assign n31634 = ( n6598 & ~n11148 ) | ( n6598 & n16949 ) | ( ~n11148 & n16949 ) ;
  assign n31635 = n31634 ^ n25182 ^ n11109 ;
  assign n31636 = ( n5686 & n6943 ) | ( n5686 & n25752 ) | ( n6943 & n25752 ) ;
  assign n31637 = n13690 ^ n12276 ^ n5328 ;
  assign n31638 = n16938 ^ n13511 ^ n7081 ;
  assign n31639 = ( ~n742 & n28716 ) | ( ~n742 & n31638 ) | ( n28716 & n31638 ) ;
  assign n31640 = ( n8574 & n10787 ) | ( n8574 & ~n24975 ) | ( n10787 & ~n24975 ) ;
  assign n31641 = ( n1793 & n2188 ) | ( n1793 & n31640 ) | ( n2188 & n31640 ) ;
  assign n31642 = ( n7285 & n10561 ) | ( n7285 & n12139 ) | ( n10561 & n12139 ) ;
  assign n31643 = ( ~n2906 & n23727 ) | ( ~n2906 & n31642 ) | ( n23727 & n31642 ) ;
  assign n31644 = n13377 ^ n5201 ^ 1'b0 ;
  assign n31645 = n31644 ^ n14513 ^ n6435 ;
  assign n31646 = n31645 ^ n19575 ^ n4754 ;
  assign n31647 = ( n2834 & ~n4359 ) | ( n2834 & n5083 ) | ( ~n4359 & n5083 ) ;
  assign n31648 = n7919 & ~n31647 ;
  assign n31649 = ~n289 & n31648 ;
  assign n31650 = ( n5044 & ~n7346 ) | ( n5044 & n11178 ) | ( ~n7346 & n11178 ) ;
  assign n31651 = n6325 ^ n5237 ^ n701 ;
  assign n31652 = n31651 ^ n19187 ^ n5412 ;
  assign n31653 = ( n21982 & ~n31650 ) | ( n21982 & n31652 ) | ( ~n31650 & n31652 ) ;
  assign n31654 = n31653 ^ n11913 ^ n8126 ;
  assign n31655 = ( ~n12518 & n14164 ) | ( ~n12518 & n31654 ) | ( n14164 & n31654 ) ;
  assign n31656 = n30766 ^ n9085 ^ 1'b0 ;
  assign n31657 = ~n21239 & n31656 ;
  assign n31658 = ( n2146 & n31655 ) | ( n2146 & ~n31657 ) | ( n31655 & ~n31657 ) ;
  assign n31659 = ( n12253 & n14401 ) | ( n12253 & n25344 ) | ( n14401 & n25344 ) ;
  assign n31660 = n24040 ^ n20520 ^ n614 ;
  assign n31661 = n23334 ^ n20947 ^ n5121 ;
  assign n31662 = ( n3804 & n4128 ) | ( n3804 & n25804 ) | ( n4128 & n25804 ) ;
  assign n31663 = ( n11854 & ~n18583 ) | ( n11854 & n24787 ) | ( ~n18583 & n24787 ) ;
  assign n31664 = ( ~n4027 & n5418 ) | ( ~n4027 & n31663 ) | ( n5418 & n31663 ) ;
  assign n31665 = n28428 ^ n2128 ^ 1'b0 ;
  assign n31666 = ( n18095 & n31664 ) | ( n18095 & n31665 ) | ( n31664 & n31665 ) ;
  assign n31667 = n23512 ^ n2435 ^ 1'b0 ;
  assign n31668 = ( n7101 & ~n9776 ) | ( n7101 & n22224 ) | ( ~n9776 & n22224 ) ;
  assign n31669 = n31668 ^ n4184 ^ 1'b0 ;
  assign n31670 = n17757 | n29424 ;
  assign n31671 = n4297 & ~n31670 ;
  assign n31672 = n21299 ^ n19457 ^ n5757 ;
  assign n31673 = n31672 ^ n8538 ^ 1'b0 ;
  assign n31674 = n30838 ^ n12172 ^ n3844 ;
  assign n31675 = ( ~n1526 & n29562 ) | ( ~n1526 & n31674 ) | ( n29562 & n31674 ) ;
  assign n31679 = ( n818 & n14452 ) | ( n818 & n16547 ) | ( n14452 & n16547 ) ;
  assign n31677 = n292 | n22754 ;
  assign n31678 = n31677 ^ n2377 ^ 1'b0 ;
  assign n31676 = n27603 ^ n7571 ^ n3828 ;
  assign n31680 = n31679 ^ n31678 ^ n31676 ;
  assign n31681 = ( n2694 & ~n4085 ) | ( n2694 & n22788 ) | ( ~n4085 & n22788 ) ;
  assign n31682 = n31681 ^ n18151 ^ n11565 ;
  assign n31683 = ( n4066 & ~n5299 ) | ( n4066 & n9474 ) | ( ~n5299 & n9474 ) ;
  assign n31684 = n31683 ^ n26203 ^ n24297 ;
  assign n31685 = n15845 ^ n11424 ^ n3601 ;
  assign n31686 = ( ~n15661 & n27095 ) | ( ~n15661 & n31685 ) | ( n27095 & n31685 ) ;
  assign n31687 = ( n7879 & n27281 ) | ( n7879 & ~n31269 ) | ( n27281 & ~n31269 ) ;
  assign n31688 = n6487 ^ n4086 ^ n2274 ;
  assign n31689 = n20157 ^ n12886 ^ n4955 ;
  assign n31690 = ( n5457 & n10829 ) | ( n5457 & ~n31689 ) | ( n10829 & ~n31689 ) ;
  assign n31691 = n5978 & n22772 ;
  assign n31692 = ~n18109 & n31691 ;
  assign n31693 = ( n3997 & n14637 ) | ( n3997 & n18396 ) | ( n14637 & n18396 ) ;
  assign n31694 = n18209 ^ n9030 ^ n8806 ;
  assign n31695 = n28696 ^ n12476 ^ n6986 ;
  assign n31696 = ( n5007 & n16662 ) | ( n5007 & ~n20004 ) | ( n16662 & ~n20004 ) ;
  assign n31697 = n9754 & n10675 ;
  assign n31698 = ( ~n8723 & n12545 ) | ( ~n8723 & n15514 ) | ( n12545 & n15514 ) ;
  assign n31699 = n19077 ^ n4372 ^ 1'b0 ;
  assign n31700 = n31698 & n31699 ;
  assign n31701 = n31700 ^ n15034 ^ n5077 ;
  assign n31702 = n20776 ^ n8682 ^ n1157 ;
  assign n31703 = n29081 ^ n24474 ^ n9388 ;
  assign n31704 = n18458 ^ n16685 ^ n3815 ;
  assign n31705 = n18239 ^ n6850 ^ 1'b0 ;
  assign n31706 = n477 & ~n31705 ;
  assign n31709 = n7327 & ~n13354 ;
  assign n31710 = n31709 ^ n332 ^ 1'b0 ;
  assign n31707 = n287 | n1291 ;
  assign n31708 = n31707 ^ n8392 ^ 1'b0 ;
  assign n31711 = n31710 ^ n31708 ^ n5186 ;
  assign n31712 = n25224 ^ n20864 ^ n17968 ;
  assign n31713 = n16558 ^ n3820 ^ n1617 ;
  assign n31714 = n3359 | n11662 ;
  assign n31715 = n31714 ^ n23658 ^ 1'b0 ;
  assign n31716 = n5804 & ~n7043 ;
  assign n31717 = n31715 & n31716 ;
  assign n31718 = ( n18218 & n31713 ) | ( n18218 & n31717 ) | ( n31713 & n31717 ) ;
  assign n31719 = n31718 ^ n14994 ^ n1883 ;
  assign n31720 = ( n11375 & n14723 ) | ( n11375 & ~n20306 ) | ( n14723 & ~n20306 ) ;
  assign n31721 = n31720 ^ n27848 ^ n1485 ;
  assign n31723 = n25713 ^ n16049 ^ 1'b0 ;
  assign n31722 = n12419 | n27475 ;
  assign n31724 = n31723 ^ n31722 ^ n29932 ;
  assign n31725 = n23665 ^ n23022 ^ n7133 ;
  assign n31726 = n20047 ^ n18557 ^ n8104 ;
  assign n31727 = ( ~n10970 & n12078 ) | ( ~n10970 & n31726 ) | ( n12078 & n31726 ) ;
  assign n31728 = ( n13691 & ~n20902 ) | ( n13691 & n31727 ) | ( ~n20902 & n31727 ) ;
  assign n31729 = ( ~n2564 & n31725 ) | ( ~n2564 & n31728 ) | ( n31725 & n31728 ) ;
  assign n31730 = n16884 ^ n8788 ^ 1'b0 ;
  assign n31731 = ( n6754 & n26634 ) | ( n6754 & ~n31730 ) | ( n26634 & ~n31730 ) ;
  assign n31732 = n16121 ^ n4624 ^ n4150 ;
  assign n31733 = ( ~n1031 & n15604 ) | ( ~n1031 & n18933 ) | ( n15604 & n18933 ) ;
  assign n31734 = n31733 ^ n25233 ^ n13800 ;
  assign n31735 = n7367 & n15474 ;
  assign n31736 = n31734 & n31735 ;
  assign n31737 = ( ~n4956 & n5924 ) | ( ~n4956 & n24876 ) | ( n5924 & n24876 ) ;
  assign n31738 = ( n11256 & n31736 ) | ( n11256 & n31737 ) | ( n31736 & n31737 ) ;
  assign y0 = x6 ;
  assign y1 = x19 ;
  assign y2 = x21 ;
  assign y3 = x33 ;
  assign y4 = x53 ;
  assign y5 = x81 ;
  assign y6 = x83 ;
  assign y7 = x87 ;
  assign y8 = x92 ;
  assign y9 = x100 ;
  assign y10 = x106 ;
  assign y11 = x107 ;
  assign y12 = x113 ;
  assign y13 = x118 ;
  assign y14 = n129 ;
  assign y15 = n130 ;
  assign y16 = n131 ;
  assign y17 = ~n132 ;
  assign y18 = ~n133 ;
  assign y19 = n136 ;
  assign y20 = ~n137 ;
  assign y21 = ~n138 ;
  assign y22 = n140 ;
  assign y23 = ~n143 ;
  assign y24 = ~n144 ;
  assign y25 = ~n145 ;
  assign y26 = n153 ;
  assign y27 = n159 ;
  assign y28 = n168 ;
  assign y29 = n170 ;
  assign y30 = n176 ;
  assign y31 = ~n181 ;
  assign y32 = n193 ;
  assign y33 = n194 ;
  assign y34 = n196 ;
  assign y35 = ~n202 ;
  assign y36 = n207 ;
  assign y37 = n211 ;
  assign y38 = ~n214 ;
  assign y39 = n220 ;
  assign y40 = ~n237 ;
  assign y41 = n250 ;
  assign y42 = n255 ;
  assign y43 = n264 ;
  assign y44 = ~n269 ;
  assign y45 = n270 ;
  assign y46 = n279 ;
  assign y47 = n286 ;
  assign y48 = ~n287 ;
  assign y49 = ~n292 ;
  assign y50 = n301 ;
  assign y51 = n304 ;
  assign y52 = ~n305 ;
  assign y53 = n311 ;
  assign y54 = n330 ;
  assign y55 = n332 ;
  assign y56 = ~n349 ;
  assign y57 = ~n354 ;
  assign y58 = n357 ;
  assign y59 = ~n371 ;
  assign y60 = n382 ;
  assign y61 = n384 ;
  assign y62 = ~n390 ;
  assign y63 = n399 ;
  assign y64 = ~n419 ;
  assign y65 = n427 ;
  assign y66 = ~n436 ;
  assign y67 = n449 ;
  assign y68 = ~n458 ;
  assign y69 = ~1'b0 ;
  assign y70 = n472 ;
  assign y71 = ~n488 ;
  assign y72 = ~n496 ;
  assign y73 = n503 ;
  assign y74 = ~n511 ;
  assign y75 = n540 ;
  assign y76 = n546 ;
  assign y77 = ~n550 ;
  assign y78 = n554 ;
  assign y79 = ~n558 ;
  assign y80 = n573 ;
  assign y81 = ~1'b0 ;
  assign y82 = ~n580 ;
  assign y83 = n583 ;
  assign y84 = n601 ;
  assign y85 = n609 ;
  assign y86 = ~1'b0 ;
  assign y87 = ~n617 ;
  assign y88 = ~n625 ;
  assign y89 = ~1'b0 ;
  assign y90 = n639 ;
  assign y91 = n649 ;
  assign y92 = n657 ;
  assign y93 = ~n661 ;
  assign y94 = ~n668 ;
  assign y95 = ~n678 ;
  assign y96 = ~n681 ;
  assign y97 = ~n700 ;
  assign y98 = ~n702 ;
  assign y99 = ~n706 ;
  assign y100 = ~n708 ;
  assign y101 = ~n730 ;
  assign y102 = ~n735 ;
  assign y103 = ~n746 ;
  assign y104 = n748 ;
  assign y105 = n751 ;
  assign y106 = ~1'b0 ;
  assign y107 = n754 ;
  assign y108 = n758 ;
  assign y109 = ~n781 ;
  assign y110 = n788 ;
  assign y111 = n794 ;
  assign y112 = ~n795 ;
  assign y113 = ~1'b0 ;
  assign y114 = n796 ;
  assign y115 = ~n803 ;
  assign y116 = n836 ;
  assign y117 = ~n848 ;
  assign y118 = ~n851 ;
  assign y119 = n856 ;
  assign y120 = n861 ;
  assign y121 = ~n865 ;
  assign y122 = n883 ;
  assign y123 = n900 ;
  assign y124 = n907 ;
  assign y125 = ~n909 ;
  assign y126 = ~n922 ;
  assign y127 = ~n930 ;
  assign y128 = n940 ;
  assign y129 = n941 ;
  assign y130 = n965 ;
  assign y131 = ~n966 ;
  assign y132 = n978 ;
  assign y133 = n991 ;
  assign y134 = n997 ;
  assign y135 = n1010 ;
  assign y136 = n1023 ;
  assign y137 = ~n1032 ;
  assign y138 = n1049 ;
  assign y139 = ~n1053 ;
  assign y140 = n1060 ;
  assign y141 = n1070 ;
  assign y142 = ~n1076 ;
  assign y143 = ~1'b0 ;
  assign y144 = ~n1086 ;
  assign y145 = ~n1089 ;
  assign y146 = n1097 ;
  assign y147 = ~n1120 ;
  assign y148 = n1122 ;
  assign y149 = ~n1131 ;
  assign y150 = ~n1138 ;
  assign y151 = ~n1144 ;
  assign y152 = n1155 ;
  assign y153 = n1166 ;
  assign y154 = ~n1169 ;
  assign y155 = n1180 ;
  assign y156 = ~n1185 ;
  assign y157 = n1188 ;
  assign y158 = n1193 ;
  assign y159 = n1216 ;
  assign y160 = ~n1220 ;
  assign y161 = ~n1228 ;
  assign y162 = n1231 ;
  assign y163 = n1233 ;
  assign y164 = ~n1235 ;
  assign y165 = n1243 ;
  assign y166 = ~n1258 ;
  assign y167 = ~n1262 ;
  assign y168 = ~n1265 ;
  assign y169 = ~n1267 ;
  assign y170 = ~n1278 ;
  assign y171 = ~n1279 ;
  assign y172 = n1286 ;
  assign y173 = n1289 ;
  assign y174 = ~n1299 ;
  assign y175 = n1303 ;
  assign y176 = ~n1311 ;
  assign y177 = n1314 ;
  assign y178 = n1316 ;
  assign y179 = n1329 ;
  assign y180 = ~1'b0 ;
  assign y181 = n1333 ;
  assign y182 = n1336 ;
  assign y183 = ~n1341 ;
  assign y184 = ~n1347 ;
  assign y185 = ~n1356 ;
  assign y186 = ~1'b0 ;
  assign y187 = ~n1358 ;
  assign y188 = ~n1362 ;
  assign y189 = n1379 ;
  assign y190 = n1388 ;
  assign y191 = n1392 ;
  assign y192 = n1393 ;
  assign y193 = n1419 ;
  assign y194 = ~n1420 ;
  assign y195 = n1427 ;
  assign y196 = n1440 ;
  assign y197 = n1454 ;
  assign y198 = ~n1459 ;
  assign y199 = ~1'b0 ;
  assign y200 = ~n1495 ;
  assign y201 = n1499 ;
  assign y202 = n1502 ;
  assign y203 = n1508 ;
  assign y204 = ~n1514 ;
  assign y205 = ~n1536 ;
  assign y206 = n1551 ;
  assign y207 = ~n1553 ;
  assign y208 = ~n1563 ;
  assign y209 = ~n1568 ;
  assign y210 = n1586 ;
  assign y211 = ~n1599 ;
  assign y212 = ~n1616 ;
  assign y213 = ~n1638 ;
  assign y214 = ~1'b0 ;
  assign y215 = n1640 ;
  assign y216 = n1652 ;
  assign y217 = n1655 ;
  assign y218 = ~n1658 ;
  assign y219 = n1665 ;
  assign y220 = ~1'b0 ;
  assign y221 = n1670 ;
  assign y222 = n1682 ;
  assign y223 = n1687 ;
  assign y224 = ~n1696 ;
  assign y225 = n1702 ;
  assign y226 = ~n1704 ;
  assign y227 = ~n1708 ;
  assign y228 = ~n1711 ;
  assign y229 = n1716 ;
  assign y230 = n1726 ;
  assign y231 = n1734 ;
  assign y232 = n1741 ;
  assign y233 = n1744 ;
  assign y234 = ~n1747 ;
  assign y235 = n1761 ;
  assign y236 = ~n1777 ;
  assign y237 = n1783 ;
  assign y238 = n1800 ;
  assign y239 = ~n1807 ;
  assign y240 = ~n1815 ;
  assign y241 = n1826 ;
  assign y242 = n1829 ;
  assign y243 = ~n1832 ;
  assign y244 = ~n1835 ;
  assign y245 = n1837 ;
  assign y246 = ~n1859 ;
  assign y247 = ~n1877 ;
  assign y248 = ~n1885 ;
  assign y249 = ~n1888 ;
  assign y250 = n1899 ;
  assign y251 = ~n1911 ;
  assign y252 = n1912 ;
  assign y253 = ~n1929 ;
  assign y254 = n1938 ;
  assign y255 = ~n1941 ;
  assign y256 = ~1'b0 ;
  assign y257 = n1943 ;
  assign y258 = n1945 ;
  assign y259 = ~n1953 ;
  assign y260 = ~n1961 ;
  assign y261 = ~n1970 ;
  assign y262 = n1985 ;
  assign y263 = n1992 ;
  assign y264 = ~n2003 ;
  assign y265 = n2007 ;
  assign y266 = ~n2014 ;
  assign y267 = n2026 ;
  assign y268 = ~n2031 ;
  assign y269 = n2046 ;
  assign y270 = n2051 ;
  assign y271 = n2054 ;
  assign y272 = ~n2057 ;
  assign y273 = n2064 ;
  assign y274 = ~n2071 ;
  assign y275 = ~n2078 ;
  assign y276 = n2089 ;
  assign y277 = ~n2123 ;
  assign y278 = ~n2125 ;
  assign y279 = n2128 ;
  assign y280 = n2131 ;
  assign y281 = n2148 ;
  assign y282 = ~1'b0 ;
  assign y283 = n2150 ;
  assign y284 = n2162 ;
  assign y285 = ~n2164 ;
  assign y286 = n2187 ;
  assign y287 = n2191 ;
  assign y288 = n2198 ;
  assign y289 = ~n2215 ;
  assign y290 = n2222 ;
  assign y291 = n2253 ;
  assign y292 = ~n2256 ;
  assign y293 = ~n2270 ;
  assign y294 = ~n2273 ;
  assign y295 = ~n2294 ;
  assign y296 = n2295 ;
  assign y297 = n2300 ;
  assign y298 = ~n2301 ;
  assign y299 = n2318 ;
  assign y300 = n2328 ;
  assign y301 = ~n2332 ;
  assign y302 = ~n2334 ;
  assign y303 = ~n2345 ;
  assign y304 = n2357 ;
  assign y305 = n2361 ;
  assign y306 = n2364 ;
  assign y307 = ~n2372 ;
  assign y308 = n2375 ;
  assign y309 = n2380 ;
  assign y310 = n2400 ;
  assign y311 = n2402 ;
  assign y312 = n2403 ;
  assign y313 = n2404 ;
  assign y314 = n2412 ;
  assign y315 = ~n2422 ;
  assign y316 = ~n2424 ;
  assign y317 = ~n2439 ;
  assign y318 = ~1'b0 ;
  assign y319 = n2444 ;
  assign y320 = ~n2451 ;
  assign y321 = ~n2459 ;
  assign y322 = n2469 ;
  assign y323 = n2501 ;
  assign y324 = n2502 ;
  assign y325 = ~n2504 ;
  assign y326 = ~n2509 ;
  assign y327 = ~n2514 ;
  assign y328 = n2519 ;
  assign y329 = ~n2523 ;
  assign y330 = ~n2533 ;
  assign y331 = ~n2535 ;
  assign y332 = n2542 ;
  assign y333 = n2543 ;
  assign y334 = ~n2545 ;
  assign y335 = ~n2555 ;
  assign y336 = n2566 ;
  assign y337 = ~n2570 ;
  assign y338 = n2577 ;
  assign y339 = ~n2579 ;
  assign y340 = n2592 ;
  assign y341 = n2602 ;
  assign y342 = n2625 ;
  assign y343 = ~n2626 ;
  assign y344 = ~n2627 ;
  assign y345 = ~n2629 ;
  assign y346 = n2630 ;
  assign y347 = ~n2640 ;
  assign y348 = ~n2644 ;
  assign y349 = n2646 ;
  assign y350 = n2648 ;
  assign y351 = ~n2650 ;
  assign y352 = n2671 ;
  assign y353 = n2687 ;
  assign y354 = ~n2690 ;
  assign y355 = ~n2693 ;
  assign y356 = ~n2701 ;
  assign y357 = ~n2704 ;
  assign y358 = ~n2713 ;
  assign y359 = n2714 ;
  assign y360 = n2729 ;
  assign y361 = n2739 ;
  assign y362 = n2755 ;
  assign y363 = n2760 ;
  assign y364 = ~n2763 ;
  assign y365 = n2766 ;
  assign y366 = n2767 ;
  assign y367 = n2777 ;
  assign y368 = ~n2788 ;
  assign y369 = ~n2793 ;
  assign y370 = ~n2794 ;
  assign y371 = n2796 ;
  assign y372 = n2815 ;
  assign y373 = ~n2822 ;
  assign y374 = ~1'b0 ;
  assign y375 = ~n2826 ;
  assign y376 = ~1'b0 ;
  assign y377 = n2836 ;
  assign y378 = n2845 ;
  assign y379 = ~n2855 ;
  assign y380 = ~n2858 ;
  assign y381 = n2863 ;
  assign y382 = ~n2865 ;
  assign y383 = n2871 ;
  assign y384 = ~n2904 ;
  assign y385 = ~n2911 ;
  assign y386 = ~n2928 ;
  assign y387 = n2933 ;
  assign y388 = ~n2936 ;
  assign y389 = ~n2943 ;
  assign y390 = n2954 ;
  assign y391 = n2961 ;
  assign y392 = n2968 ;
  assign y393 = ~n2985 ;
  assign y394 = ~n3003 ;
  assign y395 = ~n3005 ;
  assign y396 = ~1'b0 ;
  assign y397 = ~n3008 ;
  assign y398 = ~n3021 ;
  assign y399 = n3032 ;
  assign y400 = ~n3042 ;
  assign y401 = n3052 ;
  assign y402 = n3061 ;
  assign y403 = ~n3065 ;
  assign y404 = n3069 ;
  assign y405 = ~n3072 ;
  assign y406 = ~n3078 ;
  assign y407 = ~1'b0 ;
  assign y408 = n3089 ;
  assign y409 = n3092 ;
  assign y410 = ~n3099 ;
  assign y411 = n3102 ;
  assign y412 = n3117 ;
  assign y413 = n3123 ;
  assign y414 = n3125 ;
  assign y415 = n3134 ;
  assign y416 = ~n3135 ;
  assign y417 = n3145 ;
  assign y418 = ~n3152 ;
  assign y419 = ~n3174 ;
  assign y420 = ~n3192 ;
  assign y421 = ~n3196 ;
  assign y422 = ~n3200 ;
  assign y423 = n3203 ;
  assign y424 = n3212 ;
  assign y425 = n3219 ;
  assign y426 = ~1'b0 ;
  assign y427 = ~n3227 ;
  assign y428 = n3237 ;
  assign y429 = ~n3246 ;
  assign y430 = ~n3251 ;
  assign y431 = ~n3260 ;
  assign y432 = n3266 ;
  assign y433 = n3270 ;
  assign y434 = n3286 ;
  assign y435 = n3292 ;
  assign y436 = ~n3303 ;
  assign y437 = ~n3317 ;
  assign y438 = n3321 ;
  assign y439 = n3322 ;
  assign y440 = n3328 ;
  assign y441 = n3344 ;
  assign y442 = ~n3347 ;
  assign y443 = ~n3364 ;
  assign y444 = ~n3370 ;
  assign y445 = ~n3376 ;
  assign y446 = n3377 ;
  assign y447 = ~n3384 ;
  assign y448 = ~n3395 ;
  assign y449 = ~n3411 ;
  assign y450 = n3413 ;
  assign y451 = ~n3416 ;
  assign y452 = ~n3420 ;
  assign y453 = n3422 ;
  assign y454 = n3425 ;
  assign y455 = n3426 ;
  assign y456 = ~n3437 ;
  assign y457 = ~n3454 ;
  assign y458 = ~n3457 ;
  assign y459 = ~1'b0 ;
  assign y460 = ~n3460 ;
  assign y461 = n3474 ;
  assign y462 = ~n3485 ;
  assign y463 = n3488 ;
  assign y464 = ~n3490 ;
  assign y465 = n3494 ;
  assign y466 = n3507 ;
  assign y467 = ~n3515 ;
  assign y468 = ~n3529 ;
  assign y469 = ~1'b0 ;
  assign y470 = n3541 ;
  assign y471 = ~n3545 ;
  assign y472 = ~n3552 ;
  assign y473 = ~n3560 ;
  assign y474 = ~n3563 ;
  assign y475 = n3567 ;
  assign y476 = ~n3587 ;
  assign y477 = ~n3591 ;
  assign y478 = n3606 ;
  assign y479 = n3610 ;
  assign y480 = n3612 ;
  assign y481 = n3626 ;
  assign y482 = ~n3632 ;
  assign y483 = n3634 ;
  assign y484 = ~n3643 ;
  assign y485 = ~n3666 ;
  assign y486 = ~n3671 ;
  assign y487 = n3675 ;
  assign y488 = n3678 ;
  assign y489 = ~n3686 ;
  assign y490 = ~n3687 ;
  assign y491 = ~n3690 ;
  assign y492 = n3694 ;
  assign y493 = ~n3696 ;
  assign y494 = ~n3699 ;
  assign y495 = ~n3705 ;
  assign y496 = n3712 ;
  assign y497 = n3728 ;
  assign y498 = n3735 ;
  assign y499 = n3737 ;
  assign y500 = n3739 ;
  assign y501 = ~1'b0 ;
  assign y502 = ~n3745 ;
  assign y503 = ~n3754 ;
  assign y504 = n3767 ;
  assign y505 = n3775 ;
  assign y506 = ~n3778 ;
  assign y507 = ~n3780 ;
  assign y508 = ~n3786 ;
  assign y509 = ~n3801 ;
  assign y510 = ~n3813 ;
  assign y511 = n3818 ;
  assign y512 = ~n3823 ;
  assign y513 = ~n3825 ;
  assign y514 = n3837 ;
  assign y515 = ~n3851 ;
  assign y516 = n3854 ;
  assign y517 = ~n3855 ;
  assign y518 = n3862 ;
  assign y519 = ~n3873 ;
  assign y520 = ~n3879 ;
  assign y521 = n3883 ;
  assign y522 = ~n3886 ;
  assign y523 = n3889 ;
  assign y524 = ~1'b0 ;
  assign y525 = ~n3902 ;
  assign y526 = ~n3932 ;
  assign y527 = n3937 ;
  assign y528 = n3947 ;
  assign y529 = n3958 ;
  assign y530 = ~1'b0 ;
  assign y531 = n3963 ;
  assign y532 = n3972 ;
  assign y533 = ~n3973 ;
  assign y534 = ~n3980 ;
  assign y535 = n3988 ;
  assign y536 = ~n4007 ;
  assign y537 = ~n4012 ;
  assign y538 = n4019 ;
  assign y539 = ~1'b0 ;
  assign y540 = ~n4027 ;
  assign y541 = n4035 ;
  assign y542 = n4040 ;
  assign y543 = ~n4046 ;
  assign y544 = ~n4067 ;
  assign y545 = ~n4073 ;
  assign y546 = ~n4084 ;
  assign y547 = n4088 ;
  assign y548 = ~n4089 ;
  assign y549 = ~1'b0 ;
  assign y550 = ~n4090 ;
  assign y551 = n4095 ;
  assign y552 = n4101 ;
  assign y553 = ~n4106 ;
  assign y554 = ~n4124 ;
  assign y555 = n4135 ;
  assign y556 = ~n4148 ;
  assign y557 = n4159 ;
  assign y558 = n4163 ;
  assign y559 = n4182 ;
  assign y560 = n4193 ;
  assign y561 = ~n4200 ;
  assign y562 = ~n4218 ;
  assign y563 = ~n4223 ;
  assign y564 = ~n4240 ;
  assign y565 = ~n4245 ;
  assign y566 = ~n4254 ;
  assign y567 = ~n4255 ;
  assign y568 = ~n4261 ;
  assign y569 = n4268 ;
  assign y570 = n4280 ;
  assign y571 = ~n4286 ;
  assign y572 = n4292 ;
  assign y573 = n4295 ;
  assign y574 = n4301 ;
  assign y575 = ~1'b0 ;
  assign y576 = ~n4315 ;
  assign y577 = ~n4318 ;
  assign y578 = n4332 ;
  assign y579 = ~n4333 ;
  assign y580 = n4340 ;
  assign y581 = n4358 ;
  assign y582 = ~n4372 ;
  assign y583 = n4375 ;
  assign y584 = n4378 ;
  assign y585 = n4390 ;
  assign y586 = n4412 ;
  assign y587 = n4417 ;
  assign y588 = n4425 ;
  assign y589 = n4427 ;
  assign y590 = n4432 ;
  assign y591 = n4441 ;
  assign y592 = n4442 ;
  assign y593 = ~n4450 ;
  assign y594 = ~n4458 ;
  assign y595 = ~n4467 ;
  assign y596 = n4476 ;
  assign y597 = n4481 ;
  assign y598 = n4484 ;
  assign y599 = ~n4495 ;
  assign y600 = ~n4503 ;
  assign y601 = n4506 ;
  assign y602 = n4508 ;
  assign y603 = n4510 ;
  assign y604 = ~n4524 ;
  assign y605 = ~n4526 ;
  assign y606 = n4529 ;
  assign y607 = ~1'b0 ;
  assign y608 = n4545 ;
  assign y609 = n4547 ;
  assign y610 = n4554 ;
  assign y611 = ~n4565 ;
  assign y612 = n4572 ;
  assign y613 = ~n4573 ;
  assign y614 = ~n4580 ;
  assign y615 = ~n4585 ;
  assign y616 = ~n4600 ;
  assign y617 = n4601 ;
  assign y618 = ~n4615 ;
  assign y619 = n4632 ;
  assign y620 = ~n4642 ;
  assign y621 = n4648 ;
  assign y622 = n4652 ;
  assign y623 = n4675 ;
  assign y624 = ~n4677 ;
  assign y625 = n4681 ;
  assign y626 = n4694 ;
  assign y627 = n4700 ;
  assign y628 = n4710 ;
  assign y629 = n4712 ;
  assign y630 = ~n4715 ;
  assign y631 = ~n4726 ;
  assign y632 = ~n4731 ;
  assign y633 = ~n4732 ;
  assign y634 = ~n4736 ;
  assign y635 = ~n4737 ;
  assign y636 = ~n4752 ;
  assign y637 = ~n4758 ;
  assign y638 = ~n4763 ;
  assign y639 = ~n4765 ;
  assign y640 = n4772 ;
  assign y641 = ~n4773 ;
  assign y642 = n4786 ;
  assign y643 = ~1'b0 ;
  assign y644 = n4788 ;
  assign y645 = ~n4791 ;
  assign y646 = ~n4792 ;
  assign y647 = n4805 ;
  assign y648 = n4806 ;
  assign y649 = ~1'b0 ;
  assign y650 = ~n4819 ;
  assign y651 = ~n4826 ;
  assign y652 = ~n4828 ;
  assign y653 = ~n4832 ;
  assign y654 = ~n4849 ;
  assign y655 = n4854 ;
  assign y656 = n4857 ;
  assign y657 = ~n4862 ;
  assign y658 = n4870 ;
  assign y659 = n4881 ;
  assign y660 = n4893 ;
  assign y661 = ~n4902 ;
  assign y662 = ~1'b0 ;
  assign y663 = n4918 ;
  assign y664 = n4926 ;
  assign y665 = ~n4928 ;
  assign y666 = ~n4935 ;
  assign y667 = ~n4941 ;
  assign y668 = n4946 ;
  assign y669 = n4971 ;
  assign y670 = n4973 ;
  assign y671 = n4976 ;
  assign y672 = n4981 ;
  assign y673 = ~n4982 ;
  assign y674 = ~n4985 ;
  assign y675 = n4989 ;
  assign y676 = n4991 ;
  assign y677 = n4999 ;
  assign y678 = n5000 ;
  assign y679 = n5002 ;
  assign y680 = n5013 ;
  assign y681 = ~n5025 ;
  assign y682 = n5031 ;
  assign y683 = ~n5035 ;
  assign y684 = n5057 ;
  assign y685 = ~n5066 ;
  assign y686 = n5068 ;
  assign y687 = ~1'b0 ;
  assign y688 = n5073 ;
  assign y689 = ~1'b0 ;
  assign y690 = ~n5087 ;
  assign y691 = n5089 ;
  assign y692 = n5097 ;
  assign y693 = n5104 ;
  assign y694 = ~n5107 ;
  assign y695 = ~n5108 ;
  assign y696 = n5109 ;
  assign y697 = ~1'b0 ;
  assign y698 = n5117 ;
  assign y699 = ~n5118 ;
  assign y700 = ~n5123 ;
  assign y701 = n5136 ;
  assign y702 = ~n5141 ;
  assign y703 = n5146 ;
  assign y704 = ~n5148 ;
  assign y705 = ~n5165 ;
  assign y706 = ~n5185 ;
  assign y707 = n5188 ;
  assign y708 = ~n5192 ;
  assign y709 = n5193 ;
  assign y710 = n5199 ;
  assign y711 = n5205 ;
  assign y712 = n5218 ;
  assign y713 = n5229 ;
  assign y714 = n5232 ;
  assign y715 = n5234 ;
  assign y716 = n5244 ;
  assign y717 = ~n5246 ;
  assign y718 = ~n5253 ;
  assign y719 = n5260 ;
  assign y720 = n5265 ;
  assign y721 = ~n5267 ;
  assign y722 = ~n5268 ;
  assign y723 = ~n5275 ;
  assign y724 = n5280 ;
  assign y725 = n5283 ;
  assign y726 = ~n5286 ;
  assign y727 = n5289 ;
  assign y728 = n5291 ;
  assign y729 = n5292 ;
  assign y730 = ~n5302 ;
  assign y731 = n5310 ;
  assign y732 = ~n5321 ;
  assign y733 = n5334 ;
  assign y734 = n5336 ;
  assign y735 = n5345 ;
  assign y736 = ~n5350 ;
  assign y737 = ~n5360 ;
  assign y738 = n5361 ;
  assign y739 = ~n5374 ;
  assign y740 = n5392 ;
  assign y741 = ~n5393 ;
  assign y742 = n5394 ;
  assign y743 = n5397 ;
  assign y744 = n5400 ;
  assign y745 = n5415 ;
  assign y746 = ~n5421 ;
  assign y747 = n5438 ;
  assign y748 = ~n5445 ;
  assign y749 = n5446 ;
  assign y750 = ~n5461 ;
  assign y751 = n5465 ;
  assign y752 = ~n5468 ;
  assign y753 = ~n5471 ;
  assign y754 = n5474 ;
  assign y755 = ~n5477 ;
  assign y756 = ~n5478 ;
  assign y757 = ~n5493 ;
  assign y758 = n5498 ;
  assign y759 = n5500 ;
  assign y760 = n5501 ;
  assign y761 = ~n5510 ;
  assign y762 = ~1'b0 ;
  assign y763 = n5513 ;
  assign y764 = ~1'b0 ;
  assign y765 = n5527 ;
  assign y766 = ~n5528 ;
  assign y767 = n5534 ;
  assign y768 = ~1'b0 ;
  assign y769 = n5541 ;
  assign y770 = n5561 ;
  assign y771 = n5565 ;
  assign y772 = n5571 ;
  assign y773 = ~1'b0 ;
  assign y774 = ~n5574 ;
  assign y775 = n5577 ;
  assign y776 = n5595 ;
  assign y777 = ~n5601 ;
  assign y778 = n5603 ;
  assign y779 = n5609 ;
  assign y780 = n5612 ;
  assign y781 = ~1'b0 ;
  assign y782 = ~n5616 ;
  assign y783 = ~n5621 ;
  assign y784 = ~1'b0 ;
  assign y785 = ~n5624 ;
  assign y786 = n5627 ;
  assign y787 = ~n5633 ;
  assign y788 = ~n5641 ;
  assign y789 = ~n5665 ;
  assign y790 = ~n5688 ;
  assign y791 = ~n5698 ;
  assign y792 = ~n5711 ;
  assign y793 = n5715 ;
  assign y794 = ~1'b0 ;
  assign y795 = ~n5729 ;
  assign y796 = ~n5732 ;
  assign y797 = ~n5753 ;
  assign y798 = ~n5760 ;
  assign y799 = ~n5769 ;
  assign y800 = n5778 ;
  assign y801 = ~n5783 ;
  assign y802 = n5788 ;
  assign y803 = ~n5796 ;
  assign y804 = ~n5797 ;
  assign y805 = ~n5798 ;
  assign y806 = ~n5812 ;
  assign y807 = ~n5815 ;
  assign y808 = ~n5821 ;
  assign y809 = n5832 ;
  assign y810 = ~1'b0 ;
  assign y811 = ~n5833 ;
  assign y812 = ~n5848 ;
  assign y813 = ~1'b0 ;
  assign y814 = ~n5855 ;
  assign y815 = ~n5859 ;
  assign y816 = n5863 ;
  assign y817 = ~n5864 ;
  assign y818 = ~n5868 ;
  assign y819 = n5871 ;
  assign y820 = ~n5872 ;
  assign y821 = n5874 ;
  assign y822 = ~n5876 ;
  assign y823 = ~n5889 ;
  assign y824 = ~n5897 ;
  assign y825 = ~n5927 ;
  assign y826 = n5928 ;
  assign y827 = ~n5938 ;
  assign y828 = ~n5944 ;
  assign y829 = n5955 ;
  assign y830 = ~n5956 ;
  assign y831 = n5963 ;
  assign y832 = n5967 ;
  assign y833 = ~n5973 ;
  assign y834 = ~n5975 ;
  assign y835 = n5978 ;
  assign y836 = n5979 ;
  assign y837 = n5981 ;
  assign y838 = n5984 ;
  assign y839 = ~n5987 ;
  assign y840 = ~n5996 ;
  assign y841 = n6009 ;
  assign y842 = n6015 ;
  assign y843 = ~n6017 ;
  assign y844 = n6024 ;
  assign y845 = ~n6030 ;
  assign y846 = ~n6033 ;
  assign y847 = ~n6038 ;
  assign y848 = n6043 ;
  assign y849 = n6053 ;
  assign y850 = ~n6062 ;
  assign y851 = ~n6071 ;
  assign y852 = ~n6074 ;
  assign y853 = ~n6082 ;
  assign y854 = n6085 ;
  assign y855 = ~n6087 ;
  assign y856 = n6097 ;
  assign y857 = n6102 ;
  assign y858 = n6110 ;
  assign y859 = ~n6124 ;
  assign y860 = n6134 ;
  assign y861 = n6140 ;
  assign y862 = n6144 ;
  assign y863 = n6148 ;
  assign y864 = n6150 ;
  assign y865 = ~n6151 ;
  assign y866 = ~1'b0 ;
  assign y867 = n6167 ;
  assign y868 = ~n6175 ;
  assign y869 = ~1'b0 ;
  assign y870 = ~n6186 ;
  assign y871 = ~n6190 ;
  assign y872 = ~n6191 ;
  assign y873 = n6195 ;
  assign y874 = ~n6196 ;
  assign y875 = ~n6203 ;
  assign y876 = ~1'b0 ;
  assign y877 = n6207 ;
  assign y878 = n6225 ;
  assign y879 = ~n6240 ;
  assign y880 = n6246 ;
  assign y881 = n6262 ;
  assign y882 = n6266 ;
  assign y883 = ~n6281 ;
  assign y884 = ~n6295 ;
  assign y885 = n6319 ;
  assign y886 = ~n6321 ;
  assign y887 = ~n6327 ;
  assign y888 = ~n6334 ;
  assign y889 = n6345 ;
  assign y890 = ~n6349 ;
  assign y891 = n6353 ;
  assign y892 = ~n6355 ;
  assign y893 = ~n6356 ;
  assign y894 = n6360 ;
  assign y895 = ~n6363 ;
  assign y896 = ~1'b0 ;
  assign y897 = ~n6368 ;
  assign y898 = ~n6376 ;
  assign y899 = ~n6379 ;
  assign y900 = ~n6380 ;
  assign y901 = ~n6382 ;
  assign y902 = ~n6385 ;
  assign y903 = n6389 ;
  assign y904 = ~n6397 ;
  assign y905 = ~n6408 ;
  assign y906 = n6414 ;
  assign y907 = n6419 ;
  assign y908 = n6433 ;
  assign y909 = n6445 ;
  assign y910 = n6451 ;
  assign y911 = ~n6464 ;
  assign y912 = ~n6472 ;
  assign y913 = n6481 ;
  assign y914 = ~n6500 ;
  assign y915 = ~1'b0 ;
  assign y916 = n6507 ;
  assign y917 = ~n6516 ;
  assign y918 = n6520 ;
  assign y919 = n6522 ;
  assign y920 = ~n6535 ;
  assign y921 = ~n6549 ;
  assign y922 = n6554 ;
  assign y923 = n6565 ;
  assign y924 = n6569 ;
  assign y925 = ~n6573 ;
  assign y926 = n6576 ;
  assign y927 = n6578 ;
  assign y928 = ~n6582 ;
  assign y929 = ~n6585 ;
  assign y930 = n6595 ;
  assign y931 = n6611 ;
  assign y932 = ~n6617 ;
  assign y933 = ~n6622 ;
  assign y934 = n6626 ;
  assign y935 = n6632 ;
  assign y936 = ~n6634 ;
  assign y937 = ~n6639 ;
  assign y938 = ~n6641 ;
  assign y939 = ~n6652 ;
  assign y940 = ~n6654 ;
  assign y941 = n6661 ;
  assign y942 = ~n6664 ;
  assign y943 = ~n6678 ;
  assign y944 = n6680 ;
  assign y945 = ~n6682 ;
  assign y946 = n6684 ;
  assign y947 = ~n6693 ;
  assign y948 = ~1'b0 ;
  assign y949 = n6699 ;
  assign y950 = n6709 ;
  assign y951 = n6711 ;
  assign y952 = n6714 ;
  assign y953 = ~n6718 ;
  assign y954 = n6721 ;
  assign y955 = n6730 ;
  assign y956 = ~n6734 ;
  assign y957 = ~n6742 ;
  assign y958 = n6744 ;
  assign y959 = n6745 ;
  assign y960 = n6750 ;
  assign y961 = ~n6753 ;
  assign y962 = ~n6759 ;
  assign y963 = n6769 ;
  assign y964 = ~1'b0 ;
  assign y965 = ~n6771 ;
  assign y966 = n6773 ;
  assign y967 = n6778 ;
  assign y968 = n6780 ;
  assign y969 = n6790 ;
  assign y970 = n6797 ;
  assign y971 = ~n6803 ;
  assign y972 = ~n6815 ;
  assign y973 = ~n6825 ;
  assign y974 = ~n6827 ;
  assign y975 = ~n6830 ;
  assign y976 = n6831 ;
  assign y977 = ~n6843 ;
  assign y978 = ~n6844 ;
  assign y979 = ~n6849 ;
  assign y980 = ~n6850 ;
  assign y981 = n6851 ;
  assign y982 = ~n6861 ;
  assign y983 = ~n6865 ;
  assign y984 = n6867 ;
  assign y985 = n6881 ;
  assign y986 = n6887 ;
  assign y987 = n6901 ;
  assign y988 = ~n6908 ;
  assign y989 = ~n6914 ;
  assign y990 = ~n6920 ;
  assign y991 = ~n6929 ;
  assign y992 = n6933 ;
  assign y993 = n1331 ;
  assign y994 = ~1'b0 ;
  assign y995 = n6942 ;
  assign y996 = n6944 ;
  assign y997 = ~n6973 ;
  assign y998 = n6977 ;
  assign y999 = n6980 ;
  assign y1000 = n6983 ;
  assign y1001 = n6987 ;
  assign y1002 = n6990 ;
  assign y1003 = n6997 ;
  assign y1004 = n6999 ;
  assign y1005 = ~n7002 ;
  assign y1006 = ~n7003 ;
  assign y1007 = n7010 ;
  assign y1008 = ~n7018 ;
  assign y1009 = ~n7019 ;
  assign y1010 = ~n7023 ;
  assign y1011 = n7025 ;
  assign y1012 = ~n7031 ;
  assign y1013 = ~n7034 ;
  assign y1014 = n7036 ;
  assign y1015 = ~n7039 ;
  assign y1016 = ~n7043 ;
  assign y1017 = n7047 ;
  assign y1018 = ~n7060 ;
  assign y1019 = ~n7067 ;
  assign y1020 = ~n7070 ;
  assign y1021 = n7076 ;
  assign y1022 = n7077 ;
  assign y1023 = ~n7086 ;
  assign y1024 = n7089 ;
  assign y1025 = ~n7099 ;
  assign y1026 = ~n7103 ;
  assign y1027 = ~n7111 ;
  assign y1028 = n7114 ;
  assign y1029 = ~n7119 ;
  assign y1030 = n7120 ;
  assign y1031 = n7125 ;
  assign y1032 = ~1'b0 ;
  assign y1033 = n7127 ;
  assign y1034 = n7135 ;
  assign y1035 = n7143 ;
  assign y1036 = n7147 ;
  assign y1037 = ~n7154 ;
  assign y1038 = ~n7159 ;
  assign y1039 = ~n7162 ;
  assign y1040 = ~n7177 ;
  assign y1041 = n7179 ;
  assign y1042 = n7188 ;
  assign y1043 = ~n7193 ;
  assign y1044 = n7199 ;
  assign y1045 = n7207 ;
  assign y1046 = n7215 ;
  assign y1047 = n7219 ;
  assign y1048 = ~n7221 ;
  assign y1049 = ~n7231 ;
  assign y1050 = n7235 ;
  assign y1051 = ~n7238 ;
  assign y1052 = n7241 ;
  assign y1053 = ~n7245 ;
  assign y1054 = n7247 ;
  assign y1055 = ~n7256 ;
  assign y1056 = n7259 ;
  assign y1057 = n7261 ;
  assign y1058 = ~n7268 ;
  assign y1059 = ~n7275 ;
  assign y1060 = n7276 ;
  assign y1061 = ~n7277 ;
  assign y1062 = ~n7290 ;
  assign y1063 = n7295 ;
  assign y1064 = n7296 ;
  assign y1065 = ~n1193 ;
  assign y1066 = ~n7306 ;
  assign y1067 = ~n7329 ;
  assign y1068 = n7339 ;
  assign y1069 = n7348 ;
  assign y1070 = n7353 ;
  assign y1071 = n7354 ;
  assign y1072 = n7367 ;
  assign y1073 = n7384 ;
  assign y1074 = ~1'b0 ;
  assign y1075 = ~n7394 ;
  assign y1076 = n7397 ;
  assign y1077 = ~1'b0 ;
  assign y1078 = n7399 ;
  assign y1079 = n7410 ;
  assign y1080 = ~n7417 ;
  assign y1081 = n7424 ;
  assign y1082 = ~n7427 ;
  assign y1083 = n7428 ;
  assign y1084 = n7433 ;
  assign y1085 = n7436 ;
  assign y1086 = ~1'b0 ;
  assign y1087 = ~n7444 ;
  assign y1088 = ~n7446 ;
  assign y1089 = n7448 ;
  assign y1090 = ~n7451 ;
  assign y1091 = ~n7464 ;
  assign y1092 = n7466 ;
  assign y1093 = n7469 ;
  assign y1094 = ~n7473 ;
  assign y1095 = n7483 ;
  assign y1096 = n7484 ;
  assign y1097 = ~1'b0 ;
  assign y1098 = n7492 ;
  assign y1099 = ~n7496 ;
  assign y1100 = n7497 ;
  assign y1101 = ~n7510 ;
  assign y1102 = n7520 ;
  assign y1103 = n7523 ;
  assign y1104 = n7524 ;
  assign y1105 = n7534 ;
  assign y1106 = ~n7549 ;
  assign y1107 = n7551 ;
  assign y1108 = n7552 ;
  assign y1109 = n7562 ;
  assign y1110 = ~n7566 ;
  assign y1111 = ~n7588 ;
  assign y1112 = n7591 ;
  assign y1113 = n7598 ;
  assign y1114 = ~n7610 ;
  assign y1115 = n7613 ;
  assign y1116 = n7624 ;
  assign y1117 = ~n7632 ;
  assign y1118 = n7634 ;
  assign y1119 = n7636 ;
  assign y1120 = ~n7641 ;
  assign y1121 = ~n7644 ;
  assign y1122 = n7646 ;
  assign y1123 = ~n7656 ;
  assign y1124 = ~n7659 ;
  assign y1125 = ~n7662 ;
  assign y1126 = n7674 ;
  assign y1127 = ~n7682 ;
  assign y1128 = n7684 ;
  assign y1129 = ~n7691 ;
  assign y1130 = n7700 ;
  assign y1131 = ~n7701 ;
  assign y1132 = ~n7704 ;
  assign y1133 = n7712 ;
  assign y1134 = n7714 ;
  assign y1135 = ~1'b0 ;
  assign y1136 = n7718 ;
  assign y1137 = ~n7728 ;
  assign y1138 = ~n7732 ;
  assign y1139 = n7736 ;
  assign y1140 = ~n7742 ;
  assign y1141 = n7743 ;
  assign y1142 = n7750 ;
  assign y1143 = ~n7752 ;
  assign y1144 = n7762 ;
  assign y1145 = n7763 ;
  assign y1146 = n7764 ;
  assign y1147 = ~n7768 ;
  assign y1148 = n7776 ;
  assign y1149 = n7788 ;
  assign y1150 = n7791 ;
  assign y1151 = ~n7806 ;
  assign y1152 = n7809 ;
  assign y1153 = n7820 ;
  assign y1154 = n7821 ;
  assign y1155 = ~n7830 ;
  assign y1156 = ~1'b0 ;
  assign y1157 = n7834 ;
  assign y1158 = n7835 ;
  assign y1159 = ~n7840 ;
  assign y1160 = ~n7842 ;
  assign y1161 = ~n7844 ;
  assign y1162 = n7845 ;
  assign y1163 = n7849 ;
  assign y1164 = n7855 ;
  assign y1165 = n7856 ;
  assign y1166 = n7868 ;
  assign y1167 = n7878 ;
  assign y1168 = n7886 ;
  assign y1169 = n7892 ;
  assign y1170 = ~n7894 ;
  assign y1171 = n7896 ;
  assign y1172 = ~n7901 ;
  assign y1173 = ~n7902 ;
  assign y1174 = ~n7907 ;
  assign y1175 = n7919 ;
  assign y1176 = n7928 ;
  assign y1177 = n7936 ;
  assign y1178 = n7941 ;
  assign y1179 = ~n7943 ;
  assign y1180 = ~n7946 ;
  assign y1181 = ~n7954 ;
  assign y1182 = n7960 ;
  assign y1183 = n7962 ;
  assign y1184 = ~n7970 ;
  assign y1185 = ~n7974 ;
  assign y1186 = ~n7977 ;
  assign y1187 = n7984 ;
  assign y1188 = n7986 ;
  assign y1189 = ~n7993 ;
  assign y1190 = n8007 ;
  assign y1191 = ~n8021 ;
  assign y1192 = n8032 ;
  assign y1193 = ~n8037 ;
  assign y1194 = ~n8038 ;
  assign y1195 = ~n8042 ;
  assign y1196 = ~n8045 ;
  assign y1197 = n8051 ;
  assign y1198 = ~n5919 ;
  assign y1199 = ~n8063 ;
  assign y1200 = n8066 ;
  assign y1201 = ~n8067 ;
  assign y1202 = ~n8072 ;
  assign y1203 = n8076 ;
  assign y1204 = ~n8085 ;
  assign y1205 = ~n8094 ;
  assign y1206 = n8099 ;
  assign y1207 = ~1'b0 ;
  assign y1208 = n8110 ;
  assign y1209 = n8113 ;
  assign y1210 = n8123 ;
  assign y1211 = ~n8127 ;
  assign y1212 = n8130 ;
  assign y1213 = ~n8133 ;
  assign y1214 = ~n8137 ;
  assign y1215 = n8141 ;
  assign y1216 = ~n8143 ;
  assign y1217 = n8145 ;
  assign y1218 = n8157 ;
  assign y1219 = n8169 ;
  assign y1220 = ~1'b0 ;
  assign y1221 = n8170 ;
  assign y1222 = n8171 ;
  assign y1223 = n8174 ;
  assign y1224 = ~n8176 ;
  assign y1225 = ~1'b0 ;
  assign y1226 = ~n8177 ;
  assign y1227 = n8183 ;
  assign y1228 = ~n8200 ;
  assign y1229 = ~n8204 ;
  assign y1230 = ~n8210 ;
  assign y1231 = n8213 ;
  assign y1232 = ~1'b0 ;
  assign y1233 = n8215 ;
  assign y1234 = n8218 ;
  assign y1235 = ~n8219 ;
  assign y1236 = n8227 ;
  assign y1237 = n8231 ;
  assign y1238 = ~n8237 ;
  assign y1239 = ~n8242 ;
  assign y1240 = n8252 ;
  assign y1241 = ~n8258 ;
  assign y1242 = ~n8262 ;
  assign y1243 = n8264 ;
  assign y1244 = n8265 ;
  assign y1245 = ~n8276 ;
  assign y1246 = ~n8277 ;
  assign y1247 = ~n8296 ;
  assign y1248 = ~n8304 ;
  assign y1249 = ~n8306 ;
  assign y1250 = n8309 ;
  assign y1251 = n8316 ;
  assign y1252 = n8319 ;
  assign y1253 = n8323 ;
  assign y1254 = n8326 ;
  assign y1255 = ~n8332 ;
  assign y1256 = ~n8335 ;
  assign y1257 = n8336 ;
  assign y1258 = n8342 ;
  assign y1259 = ~n8347 ;
  assign y1260 = n8349 ;
  assign y1261 = ~n8351 ;
  assign y1262 = ~1'b0 ;
  assign y1263 = n8368 ;
  assign y1264 = ~n8373 ;
  assign y1265 = n8388 ;
  assign y1266 = ~n8391 ;
  assign y1267 = n8398 ;
  assign y1268 = ~n8404 ;
  assign y1269 = n8413 ;
  assign y1270 = ~n8414 ;
  assign y1271 = ~n8421 ;
  assign y1272 = n8428 ;
  assign y1273 = n8432 ;
  assign y1274 = ~n8444 ;
  assign y1275 = n8452 ;
  assign y1276 = n8467 ;
  assign y1277 = ~n8494 ;
  assign y1278 = ~n8498 ;
  assign y1279 = n8500 ;
  assign y1280 = ~n8507 ;
  assign y1281 = ~n8508 ;
  assign y1282 = n8511 ;
  assign y1283 = n8513 ;
  assign y1284 = ~n8522 ;
  assign y1285 = n8527 ;
  assign y1286 = n8531 ;
  assign y1287 = n8532 ;
  assign y1288 = ~n8533 ;
  assign y1289 = ~n8547 ;
  assign y1290 = ~n8548 ;
  assign y1291 = n8549 ;
  assign y1292 = ~n8552 ;
  assign y1293 = ~n8554 ;
  assign y1294 = ~n8560 ;
  assign y1295 = ~n8572 ;
  assign y1296 = n8583 ;
  assign y1297 = n8586 ;
  assign y1298 = ~n8590 ;
  assign y1299 = ~n8596 ;
  assign y1300 = n8599 ;
  assign y1301 = n8618 ;
  assign y1302 = ~n8625 ;
  assign y1303 = ~n8631 ;
  assign y1304 = n8636 ;
  assign y1305 = ~n7148 ;
  assign y1306 = ~n8637 ;
  assign y1307 = ~n8649 ;
  assign y1308 = n8657 ;
  assign y1309 = ~n8658 ;
  assign y1310 = n8660 ;
  assign y1311 = ~1'b0 ;
  assign y1312 = ~n8665 ;
  assign y1313 = ~n8668 ;
  assign y1314 = ~n8670 ;
  assign y1315 = ~n8676 ;
  assign y1316 = ~n8699 ;
  assign y1317 = n8708 ;
  assign y1318 = ~n8714 ;
  assign y1319 = ~n8726 ;
  assign y1320 = ~n8732 ;
  assign y1321 = ~n8734 ;
  assign y1322 = n8741 ;
  assign y1323 = ~n8746 ;
  assign y1324 = n8751 ;
  assign y1325 = n8752 ;
  assign y1326 = ~1'b0 ;
  assign y1327 = n8761 ;
  assign y1328 = n8762 ;
  assign y1329 = ~n8763 ;
  assign y1330 = ~n8766 ;
  assign y1331 = ~n8767 ;
  assign y1332 = ~n8769 ;
  assign y1333 = n8780 ;
  assign y1334 = n8789 ;
  assign y1335 = ~n8790 ;
  assign y1336 = ~n8800 ;
  assign y1337 = n8805 ;
  assign y1338 = n8808 ;
  assign y1339 = ~n8812 ;
  assign y1340 = ~n8819 ;
  assign y1341 = ~n8825 ;
  assign y1342 = n8826 ;
  assign y1343 = ~n8837 ;
  assign y1344 = ~1'b0 ;
  assign y1345 = n8843 ;
  assign y1346 = n8855 ;
  assign y1347 = ~n8871 ;
  assign y1348 = ~n8879 ;
  assign y1349 = ~n8882 ;
  assign y1350 = n8888 ;
  assign y1351 = ~n8892 ;
  assign y1352 = n8898 ;
  assign y1353 = n8909 ;
  assign y1354 = n8916 ;
  assign y1355 = n8919 ;
  assign y1356 = ~n8930 ;
  assign y1357 = ~n8937 ;
  assign y1358 = ~n8944 ;
  assign y1359 = n8945 ;
  assign y1360 = n8948 ;
  assign y1361 = ~n8949 ;
  assign y1362 = n8957 ;
  assign y1363 = ~n8964 ;
  assign y1364 = ~n8973 ;
  assign y1365 = ~n8976 ;
  assign y1366 = n8977 ;
  assign y1367 = n8985 ;
  assign y1368 = ~n8994 ;
  assign y1369 = ~n9010 ;
  assign y1370 = n9018 ;
  assign y1371 = n9026 ;
  assign y1372 = n9031 ;
  assign y1373 = ~n9032 ;
  assign y1374 = ~n9033 ;
  assign y1375 = n9039 ;
  assign y1376 = n9041 ;
  assign y1377 = ~n9045 ;
  assign y1378 = ~n9049 ;
  assign y1379 = ~n9053 ;
  assign y1380 = ~1'b0 ;
  assign y1381 = ~n9059 ;
  assign y1382 = ~n9060 ;
  assign y1383 = n9071 ;
  assign y1384 = n9078 ;
  assign y1385 = n9085 ;
  assign y1386 = ~n9100 ;
  assign y1387 = n9104 ;
  assign y1388 = n9106 ;
  assign y1389 = n9108 ;
  assign y1390 = ~n9110 ;
  assign y1391 = ~n9113 ;
  assign y1392 = n9116 ;
  assign y1393 = n9117 ;
  assign y1394 = n9123 ;
  assign y1395 = n9132 ;
  assign y1396 = n9139 ;
  assign y1397 = n9150 ;
  assign y1398 = n9152 ;
  assign y1399 = n9154 ;
  assign y1400 = n9160 ;
  assign y1401 = ~n9163 ;
  assign y1402 = ~n9165 ;
  assign y1403 = n9169 ;
  assign y1404 = n9177 ;
  assign y1405 = n9186 ;
  assign y1406 = ~n9191 ;
  assign y1407 = ~n9199 ;
  assign y1408 = n9201 ;
  assign y1409 = n9207 ;
  assign y1410 = n9213 ;
  assign y1411 = n9214 ;
  assign y1412 = ~n9218 ;
  assign y1413 = n9220 ;
  assign y1414 = n9234 ;
  assign y1415 = n9236 ;
  assign y1416 = n9238 ;
  assign y1417 = n9248 ;
  assign y1418 = ~n9252 ;
  assign y1419 = ~n9262 ;
  assign y1420 = n9263 ;
  assign y1421 = ~n9271 ;
  assign y1422 = ~n9273 ;
  assign y1423 = ~n9282 ;
  assign y1424 = n9287 ;
  assign y1425 = n9289 ;
  assign y1426 = n9296 ;
  assign y1427 = ~n9299 ;
  assign y1428 = n9302 ;
  assign y1429 = ~n9304 ;
  assign y1430 = n9305 ;
  assign y1431 = n9310 ;
  assign y1432 = ~n9323 ;
  assign y1433 = ~n9326 ;
  assign y1434 = n9328 ;
  assign y1435 = n9332 ;
  assign y1436 = ~n9348 ;
  assign y1437 = ~n9350 ;
  assign y1438 = n9363 ;
  assign y1439 = n9366 ;
  assign y1440 = n9368 ;
  assign y1441 = ~n9369 ;
  assign y1442 = ~n9384 ;
  assign y1443 = n9390 ;
  assign y1444 = ~n9393 ;
  assign y1445 = n9401 ;
  assign y1446 = n9405 ;
  assign y1447 = ~n9406 ;
  assign y1448 = n9408 ;
  assign y1449 = ~n9410 ;
  assign y1450 = n9421 ;
  assign y1451 = ~n9428 ;
  assign y1452 = ~n9433 ;
  assign y1453 = n9442 ;
  assign y1454 = ~1'b0 ;
  assign y1455 = n9448 ;
  assign y1456 = ~n9459 ;
  assign y1457 = n9460 ;
  assign y1458 = n9470 ;
  assign y1459 = n9490 ;
  assign y1460 = n9492 ;
  assign y1461 = ~n9503 ;
  assign y1462 = n9509 ;
  assign y1463 = n9515 ;
  assign y1464 = ~n9527 ;
  assign y1465 = n9531 ;
  assign y1466 = n9544 ;
  assign y1467 = n9566 ;
  assign y1468 = n9574 ;
  assign y1469 = ~n9575 ;
  assign y1470 = n9579 ;
  assign y1471 = n9589 ;
  assign y1472 = ~n9594 ;
  assign y1473 = ~1'b0 ;
  assign y1474 = ~n9597 ;
  assign y1475 = n9600 ;
  assign y1476 = ~1'b0 ;
  assign y1477 = ~n9606 ;
  assign y1478 = ~n9615 ;
  assign y1479 = n9621 ;
  assign y1480 = ~n9624 ;
  assign y1481 = n9635 ;
  assign y1482 = n9639 ;
  assign y1483 = ~n9649 ;
  assign y1484 = n9653 ;
  assign y1485 = n9659 ;
  assign y1486 = n9666 ;
  assign y1487 = ~n9668 ;
  assign y1488 = ~n9669 ;
  assign y1489 = ~n9672 ;
  assign y1490 = ~1'b0 ;
  assign y1491 = n9677 ;
  assign y1492 = ~n9678 ;
  assign y1493 = n9691 ;
  assign y1494 = n9702 ;
  assign y1495 = ~n9703 ;
  assign y1496 = n9704 ;
  assign y1497 = n9728 ;
  assign y1498 = n9729 ;
  assign y1499 = ~n9743 ;
  assign y1500 = ~n9744 ;
  assign y1501 = n9751 ;
  assign y1502 = ~n9756 ;
  assign y1503 = ~n9758 ;
  assign y1504 = ~n9763 ;
  assign y1505 = n9764 ;
  assign y1506 = n9771 ;
  assign y1507 = n9779 ;
  assign y1508 = ~n9781 ;
  assign y1509 = n9782 ;
  assign y1510 = ~n9783 ;
  assign y1511 = n9788 ;
  assign y1512 = ~n9796 ;
  assign y1513 = n9798 ;
  assign y1514 = ~n9800 ;
  assign y1515 = n9807 ;
  assign y1516 = ~n9822 ;
  assign y1517 = ~n9823 ;
  assign y1518 = n9835 ;
  assign y1519 = ~n9839 ;
  assign y1520 = n9841 ;
  assign y1521 = n9851 ;
  assign y1522 = n9855 ;
  assign y1523 = n9865 ;
  assign y1524 = n9866 ;
  assign y1525 = n9868 ;
  assign y1526 = n9880 ;
  assign y1527 = n9887 ;
  assign y1528 = n9890 ;
  assign y1529 = n9896 ;
  assign y1530 = ~n9898 ;
  assign y1531 = n9907 ;
  assign y1532 = ~n9912 ;
  assign y1533 = n9916 ;
  assign y1534 = n9919 ;
  assign y1535 = ~n9921 ;
  assign y1536 = n9925 ;
  assign y1537 = ~1'b0 ;
  assign y1538 = ~n9932 ;
  assign y1539 = n9935 ;
  assign y1540 = n9940 ;
  assign y1541 = ~n9944 ;
  assign y1542 = n9950 ;
  assign y1543 = ~n9952 ;
  assign y1544 = ~n9969 ;
  assign y1545 = ~n9971 ;
  assign y1546 = n9974 ;
  assign y1547 = ~n9982 ;
  assign y1548 = n9983 ;
  assign y1549 = n9984 ;
  assign y1550 = n9989 ;
  assign y1551 = n9992 ;
  assign y1552 = n9993 ;
  assign y1553 = n9996 ;
  assign y1554 = ~n10000 ;
  assign y1555 = n10009 ;
  assign y1556 = n10018 ;
  assign y1557 = n10024 ;
  assign y1558 = ~n10027 ;
  assign y1559 = n10028 ;
  assign y1560 = ~1'b0 ;
  assign y1561 = ~1'b0 ;
  assign y1562 = n10030 ;
  assign y1563 = ~n10034 ;
  assign y1564 = ~n10036 ;
  assign y1565 = ~n10043 ;
  assign y1566 = n10049 ;
  assign y1567 = ~n10056 ;
  assign y1568 = n10064 ;
  assign y1569 = ~n10081 ;
  assign y1570 = n10084 ;
  assign y1571 = n10092 ;
  assign y1572 = ~n10100 ;
  assign y1573 = ~n10102 ;
  assign y1574 = ~1'b0 ;
  assign y1575 = n10104 ;
  assign y1576 = ~n10108 ;
  assign y1577 = n10110 ;
  assign y1578 = n10111 ;
  assign y1579 = ~n10116 ;
  assign y1580 = ~n10118 ;
  assign y1581 = ~n10122 ;
  assign y1582 = ~n10128 ;
  assign y1583 = ~n10137 ;
  assign y1584 = n10138 ;
  assign y1585 = n10145 ;
  assign y1586 = ~n10147 ;
  assign y1587 = ~n10151 ;
  assign y1588 = n10155 ;
  assign y1589 = ~1'b0 ;
  assign y1590 = n10161 ;
  assign y1591 = n10167 ;
  assign y1592 = n10171 ;
  assign y1593 = ~1'b0 ;
  assign y1594 = n10173 ;
  assign y1595 = n10185 ;
  assign y1596 = ~1'b0 ;
  assign y1597 = n10188 ;
  assign y1598 = ~n10202 ;
  assign y1599 = ~n10212 ;
  assign y1600 = n10220 ;
  assign y1601 = n10226 ;
  assign y1602 = ~n10229 ;
  assign y1603 = n10241 ;
  assign y1604 = n10246 ;
  assign y1605 = n10248 ;
  assign y1606 = n10250 ;
  assign y1607 = n10253 ;
  assign y1608 = n10255 ;
  assign y1609 = n10256 ;
  assign y1610 = n10259 ;
  assign y1611 = n10266 ;
  assign y1612 = ~n10269 ;
  assign y1613 = ~n10270 ;
  assign y1614 = ~n10283 ;
  assign y1615 = ~n10286 ;
  assign y1616 = ~n10293 ;
  assign y1617 = n10299 ;
  assign y1618 = n10300 ;
  assign y1619 = n4334 ;
  assign y1620 = ~n10312 ;
  assign y1621 = n10316 ;
  assign y1622 = ~n10317 ;
  assign y1623 = n10318 ;
  assign y1624 = n10320 ;
  assign y1625 = n10325 ;
  assign y1626 = n10327 ;
  assign y1627 = n10335 ;
  assign y1628 = ~1'b0 ;
  assign y1629 = ~n10340 ;
  assign y1630 = n10352 ;
  assign y1631 = n10354 ;
  assign y1632 = ~n10368 ;
  assign y1633 = ~1'b0 ;
  assign y1634 = n10374 ;
  assign y1635 = n10377 ;
  assign y1636 = ~n10379 ;
  assign y1637 = n10399 ;
  assign y1638 = ~n10403 ;
  assign y1639 = n10406 ;
  assign y1640 = n10414 ;
  assign y1641 = n10417 ;
  assign y1642 = ~n10421 ;
  assign y1643 = ~n10424 ;
  assign y1644 = ~n10432 ;
  assign y1645 = ~1'b0 ;
  assign y1646 = n10437 ;
  assign y1647 = n10438 ;
  assign y1648 = ~n10440 ;
  assign y1649 = ~1'b0 ;
  assign y1650 = n10450 ;
  assign y1651 = n10451 ;
  assign y1652 = ~n10460 ;
  assign y1653 = n10462 ;
  assign y1654 = n10470 ;
  assign y1655 = n10475 ;
  assign y1656 = n10490 ;
  assign y1657 = n10498 ;
  assign y1658 = ~n10499 ;
  assign y1659 = n10501 ;
  assign y1660 = n10502 ;
  assign y1661 = ~1'b0 ;
  assign y1662 = n10518 ;
  assign y1663 = ~n10525 ;
  assign y1664 = ~n10528 ;
  assign y1665 = n10530 ;
  assign y1666 = ~n10535 ;
  assign y1667 = ~n10542 ;
  assign y1668 = ~n10547 ;
  assign y1669 = ~n10555 ;
  assign y1670 = ~n10556 ;
  assign y1671 = ~n10563 ;
  assign y1672 = n10565 ;
  assign y1673 = ~n10574 ;
  assign y1674 = n10579 ;
  assign y1675 = n10584 ;
  assign y1676 = ~n10594 ;
  assign y1677 = ~n10602 ;
  assign y1678 = n10603 ;
  assign y1679 = ~n10608 ;
  assign y1680 = n10611 ;
  assign y1681 = ~1'b0 ;
  assign y1682 = n10614 ;
  assign y1683 = n10617 ;
  assign y1684 = n10625 ;
  assign y1685 = n10633 ;
  assign y1686 = ~n10634 ;
  assign y1687 = n10637 ;
  assign y1688 = n10651 ;
  assign y1689 = ~n10666 ;
  assign y1690 = ~n10679 ;
  assign y1691 = ~1'b0 ;
  assign y1692 = ~n10684 ;
  assign y1693 = n10693 ;
  assign y1694 = ~n10694 ;
  assign y1695 = ~n10696 ;
  assign y1696 = n10703 ;
  assign y1697 = n10705 ;
  assign y1698 = ~n10707 ;
  assign y1699 = n10719 ;
  assign y1700 = ~n10722 ;
  assign y1701 = ~1'b0 ;
  assign y1702 = n10724 ;
  assign y1703 = ~n10730 ;
  assign y1704 = ~n10732 ;
  assign y1705 = ~1'b0 ;
  assign y1706 = ~n10733 ;
  assign y1707 = n10757 ;
  assign y1708 = n10758 ;
  assign y1709 = ~n10771 ;
  assign y1710 = n10777 ;
  assign y1711 = n10781 ;
  assign y1712 = ~n10782 ;
  assign y1713 = ~n10784 ;
  assign y1714 = n10789 ;
  assign y1715 = n10790 ;
  assign y1716 = n10794 ;
  assign y1717 = ~n10796 ;
  assign y1718 = n10799 ;
  assign y1719 = n10802 ;
  assign y1720 = ~n10803 ;
  assign y1721 = n10808 ;
  assign y1722 = ~n10810 ;
  assign y1723 = ~n10813 ;
  assign y1724 = ~n10827 ;
  assign y1725 = n10832 ;
  assign y1726 = ~n10835 ;
  assign y1727 = ~n10837 ;
  assign y1728 = n10846 ;
  assign y1729 = n10850 ;
  assign y1730 = n10851 ;
  assign y1731 = ~n10853 ;
  assign y1732 = ~n10858 ;
  assign y1733 = n10862 ;
  assign y1734 = ~n10864 ;
  assign y1735 = n10866 ;
  assign y1736 = ~n10869 ;
  assign y1737 = ~n10876 ;
  assign y1738 = n10885 ;
  assign y1739 = n10892 ;
  assign y1740 = ~1'b0 ;
  assign y1741 = n10898 ;
  assign y1742 = ~n10899 ;
  assign y1743 = ~n10907 ;
  assign y1744 = n10914 ;
  assign y1745 = n10915 ;
  assign y1746 = n10920 ;
  assign y1747 = n10933 ;
  assign y1748 = n10935 ;
  assign y1749 = n10941 ;
  assign y1750 = ~n10949 ;
  assign y1751 = ~n10963 ;
  assign y1752 = ~n10965 ;
  assign y1753 = n10967 ;
  assign y1754 = n10972 ;
  assign y1755 = ~n10973 ;
  assign y1756 = ~n10976 ;
  assign y1757 = n10978 ;
  assign y1758 = n10980 ;
  assign y1759 = ~n10986 ;
  assign y1760 = n10987 ;
  assign y1761 = n10989 ;
  assign y1762 = ~n10998 ;
  assign y1763 = n11001 ;
  assign y1764 = ~n11006 ;
  assign y1765 = ~n11009 ;
  assign y1766 = ~n11010 ;
  assign y1767 = ~n11011 ;
  assign y1768 = n11013 ;
  assign y1769 = n11020 ;
  assign y1770 = ~n11021 ;
  assign y1771 = n11022 ;
  assign y1772 = ~n11025 ;
  assign y1773 = n11028 ;
  assign y1774 = ~n11034 ;
  assign y1775 = n11045 ;
  assign y1776 = n11056 ;
  assign y1777 = n11061 ;
  assign y1778 = ~n11075 ;
  assign y1779 = ~n11080 ;
  assign y1780 = ~n11086 ;
  assign y1781 = ~n11089 ;
  assign y1782 = ~n11095 ;
  assign y1783 = ~n11098 ;
  assign y1784 = n11105 ;
  assign y1785 = n11112 ;
  assign y1786 = ~1'b0 ;
  assign y1787 = ~n11113 ;
  assign y1788 = ~n11120 ;
  assign y1789 = n11125 ;
  assign y1790 = n11127 ;
  assign y1791 = n11131 ;
  assign y1792 = ~n11133 ;
  assign y1793 = ~n11142 ;
  assign y1794 = n11160 ;
  assign y1795 = ~n11163 ;
  assign y1796 = n11171 ;
  assign y1797 = n11172 ;
  assign y1798 = ~n11176 ;
  assign y1799 = n11181 ;
  assign y1800 = n11183 ;
  assign y1801 = n11184 ;
  assign y1802 = n11186 ;
  assign y1803 = ~n11190 ;
  assign y1804 = ~n11196 ;
  assign y1805 = n11197 ;
  assign y1806 = ~1'b0 ;
  assign y1807 = n11203 ;
  assign y1808 = ~n11207 ;
  assign y1809 = n11210 ;
  assign y1810 = ~n11212 ;
  assign y1811 = ~n11214 ;
  assign y1812 = ~n11220 ;
  assign y1813 = ~n11232 ;
  assign y1814 = n11239 ;
  assign y1815 = ~n11240 ;
  assign y1816 = n11243 ;
  assign y1817 = n11246 ;
  assign y1818 = ~n11251 ;
  assign y1819 = n11261 ;
  assign y1820 = n11263 ;
  assign y1821 = ~n11265 ;
  assign y1822 = ~n11273 ;
  assign y1823 = ~n11275 ;
  assign y1824 = ~n11276 ;
  assign y1825 = n11282 ;
  assign y1826 = n11283 ;
  assign y1827 = n11288 ;
  assign y1828 = n11294 ;
  assign y1829 = n11295 ;
  assign y1830 = n11302 ;
  assign y1831 = n11303 ;
  assign y1832 = ~n11307 ;
  assign y1833 = ~n11326 ;
  assign y1834 = ~n11328 ;
  assign y1835 = n11331 ;
  assign y1836 = ~n11334 ;
  assign y1837 = n11340 ;
  assign y1838 = n11341 ;
  assign y1839 = ~n11342 ;
  assign y1840 = n11354 ;
  assign y1841 = ~n11358 ;
  assign y1842 = ~1'b0 ;
  assign y1843 = ~n11359 ;
  assign y1844 = n11365 ;
  assign y1845 = ~n11369 ;
  assign y1846 = ~n11378 ;
  assign y1847 = n11379 ;
  assign y1848 = n11384 ;
  assign y1849 = n11396 ;
  assign y1850 = ~n11397 ;
  assign y1851 = n11402 ;
  assign y1852 = ~n11404 ;
  assign y1853 = ~n11405 ;
  assign y1854 = ~n11406 ;
  assign y1855 = n11410 ;
  assign y1856 = n11414 ;
  assign y1857 = n11420 ;
  assign y1858 = n11425 ;
  assign y1859 = n11428 ;
  assign y1860 = n11432 ;
  assign y1861 = ~n11434 ;
  assign y1862 = n11437 ;
  assign y1863 = ~n11438 ;
  assign y1864 = n11456 ;
  assign y1865 = ~n11463 ;
  assign y1866 = ~1'b0 ;
  assign y1867 = ~n11465 ;
  assign y1868 = ~n11469 ;
  assign y1869 = n11476 ;
  assign y1870 = ~n11482 ;
  assign y1871 = ~n11487 ;
  assign y1872 = n11490 ;
  assign y1873 = ~n11497 ;
  assign y1874 = ~n11499 ;
  assign y1875 = n11505 ;
  assign y1876 = ~n11510 ;
  assign y1877 = ~n11512 ;
  assign y1878 = ~n11516 ;
  assign y1879 = n11517 ;
  assign y1880 = n11524 ;
  assign y1881 = n11525 ;
  assign y1882 = ~1'b0 ;
  assign y1883 = n11528 ;
  assign y1884 = n11530 ;
  assign y1885 = n11532 ;
  assign y1886 = ~n11539 ;
  assign y1887 = n11544 ;
  assign y1888 = ~n11546 ;
  assign y1889 = n11549 ;
  assign y1890 = ~n11550 ;
  assign y1891 = ~1'b0 ;
  assign y1892 = ~n11554 ;
  assign y1893 = n11557 ;
  assign y1894 = n11575 ;
  assign y1895 = n11587 ;
  assign y1896 = n11589 ;
  assign y1897 = ~n11593 ;
  assign y1898 = n11596 ;
  assign y1899 = n11600 ;
  assign y1900 = n11606 ;
  assign y1901 = n11613 ;
  assign y1902 = ~n11623 ;
  assign y1903 = n11627 ;
  assign y1904 = n11633 ;
  assign y1905 = ~n11635 ;
  assign y1906 = n11641 ;
  assign y1907 = n11647 ;
  assign y1908 = ~n11654 ;
  assign y1909 = ~n11660 ;
  assign y1910 = ~n11670 ;
  assign y1911 = n11675 ;
  assign y1912 = n11676 ;
  assign y1913 = n11680 ;
  assign y1914 = ~n11697 ;
  assign y1915 = n11698 ;
  assign y1916 = ~n11701 ;
  assign y1917 = n11706 ;
  assign y1918 = n11712 ;
  assign y1919 = n11713 ;
  assign y1920 = ~n11718 ;
  assign y1921 = n11719 ;
  assign y1922 = n11729 ;
  assign y1923 = ~n11732 ;
  assign y1924 = ~n11742 ;
  assign y1925 = ~n11745 ;
  assign y1926 = n11747 ;
  assign y1927 = ~n11751 ;
  assign y1928 = n11753 ;
  assign y1929 = ~n11755 ;
  assign y1930 = ~n11757 ;
  assign y1931 = n11767 ;
  assign y1932 = ~n11778 ;
  assign y1933 = ~n11780 ;
  assign y1934 = n11788 ;
  assign y1935 = n11791 ;
  assign y1936 = ~n11793 ;
  assign y1937 = ~n11795 ;
  assign y1938 = n11796 ;
  assign y1939 = n11801 ;
  assign y1940 = ~n11803 ;
  assign y1941 = ~n11808 ;
  assign y1942 = ~n11813 ;
  assign y1943 = n11816 ;
  assign y1944 = n11817 ;
  assign y1945 = n11818 ;
  assign y1946 = n11819 ;
  assign y1947 = ~n11821 ;
  assign y1948 = ~n11823 ;
  assign y1949 = n11824 ;
  assign y1950 = n11827 ;
  assign y1951 = n11833 ;
  assign y1952 = ~n11845 ;
  assign y1953 = n11846 ;
  assign y1954 = ~n11848 ;
  assign y1955 = n11863 ;
  assign y1956 = n11872 ;
  assign y1957 = n11876 ;
  assign y1958 = n11877 ;
  assign y1959 = ~n11883 ;
  assign y1960 = ~n11884 ;
  assign y1961 = ~n11900 ;
  assign y1962 = n11903 ;
  assign y1963 = n11904 ;
  assign y1964 = ~n11915 ;
  assign y1965 = n11920 ;
  assign y1966 = ~n11921 ;
  assign y1967 = n11922 ;
  assign y1968 = ~n11929 ;
  assign y1969 = n11932 ;
  assign y1970 = n11934 ;
  assign y1971 = ~n11938 ;
  assign y1972 = ~1'b0 ;
  assign y1973 = ~1'b0 ;
  assign y1974 = n11943 ;
  assign y1975 = ~n11946 ;
  assign y1976 = n11947 ;
  assign y1977 = ~1'b0 ;
  assign y1978 = n11949 ;
  assign y1979 = n11954 ;
  assign y1980 = n11957 ;
  assign y1981 = ~n11960 ;
  assign y1982 = n11962 ;
  assign y1983 = ~n11968 ;
  assign y1984 = n11972 ;
  assign y1985 = n11973 ;
  assign y1986 = ~n11977 ;
  assign y1987 = n11978 ;
  assign y1988 = ~n11988 ;
  assign y1989 = ~1'b0 ;
  assign y1990 = ~n11989 ;
  assign y1991 = ~n11993 ;
  assign y1992 = ~n11994 ;
  assign y1993 = ~n11995 ;
  assign y1994 = n11997 ;
  assign y1995 = n12004 ;
  assign y1996 = n12009 ;
  assign y1997 = n12010 ;
  assign y1998 = n12022 ;
  assign y1999 = n12023 ;
  assign y2000 = ~n12028 ;
  assign y2001 = n12034 ;
  assign y2002 = n12040 ;
  assign y2003 = n12056 ;
  assign y2004 = ~n12062 ;
  assign y2005 = ~n12064 ;
  assign y2006 = ~n12069 ;
  assign y2007 = ~n12074 ;
  assign y2008 = ~n12080 ;
  assign y2009 = n12086 ;
  assign y2010 = ~n12098 ;
  assign y2011 = ~n12101 ;
  assign y2012 = n12105 ;
  assign y2013 = ~n12108 ;
  assign y2014 = n12117 ;
  assign y2015 = n12118 ;
  assign y2016 = n12127 ;
  assign y2017 = ~n12131 ;
  assign y2018 = n12144 ;
  assign y2019 = n12151 ;
  assign y2020 = n12153 ;
  assign y2021 = n12162 ;
  assign y2022 = ~n12167 ;
  assign y2023 = n12170 ;
  assign y2024 = n12174 ;
  assign y2025 = ~n12175 ;
  assign y2026 = ~n12179 ;
  assign y2027 = ~n12181 ;
  assign y2028 = ~n12186 ;
  assign y2029 = ~n12187 ;
  assign y2030 = n12196 ;
  assign y2031 = ~n12200 ;
  assign y2032 = n12201 ;
  assign y2033 = n12208 ;
  assign y2034 = ~n12209 ;
  assign y2035 = ~n12210 ;
  assign y2036 = ~n12212 ;
  assign y2037 = ~n12215 ;
  assign y2038 = ~n12217 ;
  assign y2039 = ~n12219 ;
  assign y2040 = n12221 ;
  assign y2041 = n12223 ;
  assign y2042 = n12233 ;
  assign y2043 = n12237 ;
  assign y2044 = n12239 ;
  assign y2045 = n12245 ;
  assign y2046 = ~n12248 ;
  assign y2047 = ~n12249 ;
  assign y2048 = n12250 ;
  assign y2049 = n12254 ;
  assign y2050 = ~n12263 ;
  assign y2051 = ~n12283 ;
  assign y2052 = n12285 ;
  assign y2053 = ~n12288 ;
  assign y2054 = n12289 ;
  assign y2055 = ~n12293 ;
  assign y2056 = ~n12297 ;
  assign y2057 = ~n12298 ;
  assign y2058 = ~n12300 ;
  assign y2059 = ~n12303 ;
  assign y2060 = ~n12306 ;
  assign y2061 = ~n12307 ;
  assign y2062 = ~n12310 ;
  assign y2063 = n12318 ;
  assign y2064 = n12324 ;
  assign y2065 = ~n12330 ;
  assign y2066 = n12332 ;
  assign y2067 = ~n12333 ;
  assign y2068 = ~n12334 ;
  assign y2069 = ~n12339 ;
  assign y2070 = ~1'b0 ;
  assign y2071 = n12341 ;
  assign y2072 = n12345 ;
  assign y2073 = ~n12346 ;
  assign y2074 = ~1'b0 ;
  assign y2075 = ~n12347 ;
  assign y2076 = n12357 ;
  assign y2077 = ~n12360 ;
  assign y2078 = ~n12361 ;
  assign y2079 = ~n12364 ;
  assign y2080 = n12366 ;
  assign y2081 = n12372 ;
  assign y2082 = ~n12380 ;
  assign y2083 = n12383 ;
  assign y2084 = ~n12390 ;
  assign y2085 = n12392 ;
  assign y2086 = ~n12398 ;
  assign y2087 = ~1'b0 ;
  assign y2088 = n12399 ;
  assign y2089 = n12404 ;
  assign y2090 = ~n12408 ;
  assign y2091 = ~n12420 ;
  assign y2092 = n12424 ;
  assign y2093 = n12444 ;
  assign y2094 = n12445 ;
  assign y2095 = n12446 ;
  assign y2096 = n12450 ;
  assign y2097 = n12454 ;
  assign y2098 = n12456 ;
  assign y2099 = ~n12458 ;
  assign y2100 = n12464 ;
  assign y2101 = ~n12470 ;
  assign y2102 = n12477 ;
  assign y2103 = ~n12483 ;
  assign y2104 = n12489 ;
  assign y2105 = ~n12490 ;
  assign y2106 = n12499 ;
  assign y2107 = ~n12500 ;
  assign y2108 = n12501 ;
  assign y2109 = n12508 ;
  assign y2110 = n12522 ;
  assign y2111 = ~n12532 ;
  assign y2112 = ~n12538 ;
  assign y2113 = n12540 ;
  assign y2114 = n12543 ;
  assign y2115 = n12545 ;
  assign y2116 = n12547 ;
  assign y2117 = ~n12549 ;
  assign y2118 = n12550 ;
  assign y2119 = n12551 ;
  assign y2120 = ~n12554 ;
  assign y2121 = n12559 ;
  assign y2122 = n12568 ;
  assign y2123 = n12569 ;
  assign y2124 = ~n12571 ;
  assign y2125 = n12573 ;
  assign y2126 = n12577 ;
  assign y2127 = n12579 ;
  assign y2128 = n12583 ;
  assign y2129 = ~n12585 ;
  assign y2130 = ~n12589 ;
  assign y2131 = n3090 ;
  assign y2132 = n12596 ;
  assign y2133 = n12601 ;
  assign y2134 = ~1'b0 ;
  assign y2135 = ~n12602 ;
  assign y2136 = ~1'b0 ;
  assign y2137 = ~n12609 ;
  assign y2138 = ~n12611 ;
  assign y2139 = n12622 ;
  assign y2140 = ~n12623 ;
  assign y2141 = n12629 ;
  assign y2142 = n12641 ;
  assign y2143 = n12646 ;
  assign y2144 = ~n12649 ;
  assign y2145 = ~n12650 ;
  assign y2146 = n12654 ;
  assign y2147 = ~n12659 ;
  assign y2148 = n12664 ;
  assign y2149 = ~1'b0 ;
  assign y2150 = n12673 ;
  assign y2151 = ~n12675 ;
  assign y2152 = ~n12678 ;
  assign y2153 = ~n12681 ;
  assign y2154 = ~n12684 ;
  assign y2155 = ~n12689 ;
  assign y2156 = ~n12690 ;
  assign y2157 = ~n12693 ;
  assign y2158 = n12694 ;
  assign y2159 = n12698 ;
  assign y2160 = ~n12699 ;
  assign y2161 = ~n12705 ;
  assign y2162 = ~n12714 ;
  assign y2163 = ~n12718 ;
  assign y2164 = n12721 ;
  assign y2165 = ~n12723 ;
  assign y2166 = ~n12724 ;
  assign y2167 = n12728 ;
  assign y2168 = ~n12736 ;
  assign y2169 = n12742 ;
  assign y2170 = ~n12752 ;
  assign y2171 = ~n12753 ;
  assign y2172 = n12754 ;
  assign y2173 = n12762 ;
  assign y2174 = ~n12765 ;
  assign y2175 = ~n12768 ;
  assign y2176 = n12771 ;
  assign y2177 = n12775 ;
  assign y2178 = ~n12777 ;
  assign y2179 = n12778 ;
  assign y2180 = n12783 ;
  assign y2181 = ~n12787 ;
  assign y2182 = ~n12791 ;
  assign y2183 = n12794 ;
  assign y2184 = n12796 ;
  assign y2185 = ~n12798 ;
  assign y2186 = n12806 ;
  assign y2187 = ~1'b0 ;
  assign y2188 = n12810 ;
  assign y2189 = n12813 ;
  assign y2190 = ~1'b0 ;
  assign y2191 = ~n12817 ;
  assign y2192 = n12824 ;
  assign y2193 = n12826 ;
  assign y2194 = n12829 ;
  assign y2195 = n12838 ;
  assign y2196 = n12842 ;
  assign y2197 = n12845 ;
  assign y2198 = n12846 ;
  assign y2199 = ~n12849 ;
  assign y2200 = n12854 ;
  assign y2201 = n12862 ;
  assign y2202 = ~n12870 ;
  assign y2203 = ~1'b0 ;
  assign y2204 = n12871 ;
  assign y2205 = ~n12874 ;
  assign y2206 = n12877 ;
  assign y2207 = n12879 ;
  assign y2208 = n12880 ;
  assign y2209 = ~n12882 ;
  assign y2210 = ~n12884 ;
  assign y2211 = ~n12892 ;
  assign y2212 = n12894 ;
  assign y2213 = n12896 ;
  assign y2214 = n12897 ;
  assign y2215 = ~n12902 ;
  assign y2216 = n12911 ;
  assign y2217 = ~n12914 ;
  assign y2218 = ~n12918 ;
  assign y2219 = n12919 ;
  assign y2220 = ~n12927 ;
  assign y2221 = n12929 ;
  assign y2222 = ~n12931 ;
  assign y2223 = n12933 ;
  assign y2224 = n12934 ;
  assign y2225 = n12936 ;
  assign y2226 = n12937 ;
  assign y2227 = ~n12943 ;
  assign y2228 = n12953 ;
  assign y2229 = ~n12960 ;
  assign y2230 = ~n12973 ;
  assign y2231 = ~1'b0 ;
  assign y2232 = n12980 ;
  assign y2233 = n12987 ;
  assign y2234 = ~n12990 ;
  assign y2235 = ~n12996 ;
  assign y2236 = n12997 ;
  assign y2237 = n12999 ;
  assign y2238 = n13005 ;
  assign y2239 = n13008 ;
  assign y2240 = ~n13013 ;
  assign y2241 = n13019 ;
  assign y2242 = n13020 ;
  assign y2243 = ~n13024 ;
  assign y2244 = ~n13027 ;
  assign y2245 = n13031 ;
  assign y2246 = n13032 ;
  assign y2247 = ~n13033 ;
  assign y2248 = n13040 ;
  assign y2249 = n13041 ;
  assign y2250 = n13043 ;
  assign y2251 = ~n13049 ;
  assign y2252 = ~n13050 ;
  assign y2253 = ~n13053 ;
  assign y2254 = ~n13061 ;
  assign y2255 = ~n13062 ;
  assign y2256 = ~n13063 ;
  assign y2257 = ~n13066 ;
  assign y2258 = ~1'b0 ;
  assign y2259 = n13067 ;
  assign y2260 = ~n13068 ;
  assign y2261 = n13076 ;
  assign y2262 = ~n13084 ;
  assign y2263 = ~n13085 ;
  assign y2264 = n13088 ;
  assign y2265 = ~n13098 ;
  assign y2266 = ~1'b0 ;
  assign y2267 = ~n13100 ;
  assign y2268 = n13101 ;
  assign y2269 = ~n13102 ;
  assign y2270 = n13118 ;
  assign y2271 = ~n13119 ;
  assign y2272 = ~n13123 ;
  assign y2273 = ~n13127 ;
  assign y2274 = ~n13129 ;
  assign y2275 = n13132 ;
  assign y2276 = n13138 ;
  assign y2277 = n13147 ;
  assign y2278 = n13148 ;
  assign y2279 = ~n13150 ;
  assign y2280 = ~n13151 ;
  assign y2281 = ~n13154 ;
  assign y2282 = ~n13156 ;
  assign y2283 = n13165 ;
  assign y2284 = ~n13166 ;
  assign y2285 = n13168 ;
  assign y2286 = ~n13176 ;
  assign y2287 = ~n13179 ;
  assign y2288 = n13181 ;
  assign y2289 = ~n13188 ;
  assign y2290 = ~n13190 ;
  assign y2291 = n13191 ;
  assign y2292 = n13197 ;
  assign y2293 = ~n13204 ;
  assign y2294 = ~n13210 ;
  assign y2295 = ~1'b0 ;
  assign y2296 = ~n13211 ;
  assign y2297 = ~n13217 ;
  assign y2298 = n13218 ;
  assign y2299 = ~n13221 ;
  assign y2300 = n13225 ;
  assign y2301 = ~n13229 ;
  assign y2302 = n13230 ;
  assign y2303 = ~1'b0 ;
  assign y2304 = ~n13232 ;
  assign y2305 = ~n13234 ;
  assign y2306 = n13236 ;
  assign y2307 = ~n13241 ;
  assign y2308 = n13248 ;
  assign y2309 = n13257 ;
  assign y2310 = ~n13258 ;
  assign y2311 = ~n13260 ;
  assign y2312 = n13262 ;
  assign y2313 = ~n13269 ;
  assign y2314 = ~1'b0 ;
  assign y2315 = ~n13280 ;
  assign y2316 = n13288 ;
  assign y2317 = n13293 ;
  assign y2318 = n13295 ;
  assign y2319 = ~n13302 ;
  assign y2320 = ~n13312 ;
  assign y2321 = n13321 ;
  assign y2322 = n13322 ;
  assign y2323 = ~1'b0 ;
  assign y2324 = ~n13328 ;
  assign y2325 = n13330 ;
  assign y2326 = n13336 ;
  assign y2327 = ~n13338 ;
  assign y2328 = n13343 ;
  assign y2329 = n13344 ;
  assign y2330 = ~n13347 ;
  assign y2331 = n13349 ;
  assign y2332 = ~n13359 ;
  assign y2333 = n13372 ;
  assign y2334 = n13373 ;
  assign y2335 = n13375 ;
  assign y2336 = n13386 ;
  assign y2337 = n13388 ;
  assign y2338 = ~n13399 ;
  assign y2339 = n13405 ;
  assign y2340 = ~1'b0 ;
  assign y2341 = n13408 ;
  assign y2342 = ~n13413 ;
  assign y2343 = n13419 ;
  assign y2344 = ~n13422 ;
  assign y2345 = n13427 ;
  assign y2346 = ~n13430 ;
  assign y2347 = n13434 ;
  assign y2348 = n13436 ;
  assign y2349 = n13442 ;
  assign y2350 = n13448 ;
  assign y2351 = ~n13449 ;
  assign y2352 = n13453 ;
  assign y2353 = ~n13462 ;
  assign y2354 = ~n13463 ;
  assign y2355 = ~1'b0 ;
  assign y2356 = ~n13467 ;
  assign y2357 = n13469 ;
  assign y2358 = n13470 ;
  assign y2359 = ~n13477 ;
  assign y2360 = n13490 ;
  assign y2361 = ~n13494 ;
  assign y2362 = n13495 ;
  assign y2363 = ~n13498 ;
  assign y2364 = ~n13500 ;
  assign y2365 = ~n13501 ;
  assign y2366 = ~n13503 ;
  assign y2367 = ~1'b0 ;
  assign y2368 = n13506 ;
  assign y2369 = ~n13508 ;
  assign y2370 = n13510 ;
  assign y2371 = ~n13515 ;
  assign y2372 = n13516 ;
  assign y2373 = ~n13519 ;
  assign y2374 = ~n13521 ;
  assign y2375 = n13524 ;
  assign y2376 = n13530 ;
  assign y2377 = ~n13533 ;
  assign y2378 = ~1'b0 ;
  assign y2379 = ~n13538 ;
  assign y2380 = ~n13540 ;
  assign y2381 = n13550 ;
  assign y2382 = n13557 ;
  assign y2383 = n13565 ;
  assign y2384 = n13570 ;
  assign y2385 = n13572 ;
  assign y2386 = n13576 ;
  assign y2387 = n13588 ;
  assign y2388 = n13589 ;
  assign y2389 = ~1'b0 ;
  assign y2390 = n13594 ;
  assign y2391 = ~n13599 ;
  assign y2392 = ~n13611 ;
  assign y2393 = n13614 ;
  assign y2394 = n13637 ;
  assign y2395 = ~n13641 ;
  assign y2396 = n13647 ;
  assign y2397 = ~n13648 ;
  assign y2398 = n13651 ;
  assign y2399 = ~n13661 ;
  assign y2400 = ~n13664 ;
  assign y2401 = ~1'b0 ;
  assign y2402 = n13670 ;
  assign y2403 = ~n13699 ;
  assign y2404 = n13705 ;
  assign y2405 = ~n13709 ;
  assign y2406 = n13711 ;
  assign y2407 = n13712 ;
  assign y2408 = n13714 ;
  assign y2409 = n13717 ;
  assign y2410 = ~n13719 ;
  assign y2411 = ~n13723 ;
  assign y2412 = ~n13726 ;
  assign y2413 = n13728 ;
  assign y2414 = n13732 ;
  assign y2415 = n13735 ;
  assign y2416 = n13738 ;
  assign y2417 = n13740 ;
  assign y2418 = n13744 ;
  assign y2419 = ~n13749 ;
  assign y2420 = ~n13750 ;
  assign y2421 = ~1'b0 ;
  assign y2422 = ~n13758 ;
  assign y2423 = ~n13764 ;
  assign y2424 = n13768 ;
  assign y2425 = n13769 ;
  assign y2426 = n13772 ;
  assign y2427 = n13773 ;
  assign y2428 = n13778 ;
  assign y2429 = n13781 ;
  assign y2430 = ~n13782 ;
  assign y2431 = n13786 ;
  assign y2432 = ~1'b0 ;
  assign y2433 = n13787 ;
  assign y2434 = ~n13788 ;
  assign y2435 = n13789 ;
  assign y2436 = n13790 ;
  assign y2437 = n13791 ;
  assign y2438 = ~n13796 ;
  assign y2439 = ~n13797 ;
  assign y2440 = n13799 ;
  assign y2441 = ~n13812 ;
  assign y2442 = ~n13813 ;
  assign y2443 = n13815 ;
  assign y2444 = ~n13817 ;
  assign y2445 = ~1'b0 ;
  assign y2446 = ~n13818 ;
  assign y2447 = ~n13819 ;
  assign y2448 = ~n13822 ;
  assign y2449 = n13823 ;
  assign y2450 = ~n13826 ;
  assign y2451 = n13829 ;
  assign y2452 = ~n13838 ;
  assign y2453 = n13850 ;
  assign y2454 = ~n13854 ;
  assign y2455 = n13859 ;
  assign y2456 = n13862 ;
  assign y2457 = ~n13865 ;
  assign y2458 = n13867 ;
  assign y2459 = n13868 ;
  assign y2460 = ~n13874 ;
  assign y2461 = ~n13888 ;
  assign y2462 = n13889 ;
  assign y2463 = n13892 ;
  assign y2464 = n13896 ;
  assign y2465 = ~n13897 ;
  assign y2466 = n13922 ;
  assign y2467 = ~n13924 ;
  assign y2468 = ~n13926 ;
  assign y2469 = n13931 ;
  assign y2470 = n13933 ;
  assign y2471 = n13934 ;
  assign y2472 = ~n13938 ;
  assign y2473 = ~n13942 ;
  assign y2474 = ~n13944 ;
  assign y2475 = n13945 ;
  assign y2476 = n13948 ;
  assign y2477 = n13950 ;
  assign y2478 = ~n13952 ;
  assign y2479 = ~n13955 ;
  assign y2480 = ~n13957 ;
  assign y2481 = n13961 ;
  assign y2482 = ~n13962 ;
  assign y2483 = ~n13968 ;
  assign y2484 = ~1'b0 ;
  assign y2485 = ~n13970 ;
  assign y2486 = n13972 ;
  assign y2487 = ~1'b0 ;
  assign y2488 = ~n13973 ;
  assign y2489 = ~n13980 ;
  assign y2490 = ~1'b0 ;
  assign y2491 = ~n13984 ;
  assign y2492 = ~n13987 ;
  assign y2493 = n13988 ;
  assign y2494 = ~n13989 ;
  assign y2495 = ~n13995 ;
  assign y2496 = ~n14005 ;
  assign y2497 = ~n14014 ;
  assign y2498 = n14016 ;
  assign y2499 = ~n14018 ;
  assign y2500 = ~n14020 ;
  assign y2501 = ~n14023 ;
  assign y2502 = n14036 ;
  assign y2503 = ~n14037 ;
  assign y2504 = n14043 ;
  assign y2505 = ~n14044 ;
  assign y2506 = ~n14050 ;
  assign y2507 = ~n14056 ;
  assign y2508 = n14057 ;
  assign y2509 = n14059 ;
  assign y2510 = n14064 ;
  assign y2511 = ~n14067 ;
  assign y2512 = n14070 ;
  assign y2513 = ~n14074 ;
  assign y2514 = n14079 ;
  assign y2515 = ~n14080 ;
  assign y2516 = ~n14081 ;
  assign y2517 = n14086 ;
  assign y2518 = ~n14093 ;
  assign y2519 = ~n14094 ;
  assign y2520 = n14095 ;
  assign y2521 = n14105 ;
  assign y2522 = ~n14107 ;
  assign y2523 = ~n14108 ;
  assign y2524 = n14109 ;
  assign y2525 = ~n14112 ;
  assign y2526 = ~n14113 ;
  assign y2527 = n14114 ;
  assign y2528 = ~n14117 ;
  assign y2529 = ~1'b0 ;
  assign y2530 = ~n14127 ;
  assign y2531 = ~n14128 ;
  assign y2532 = n14135 ;
  assign y2533 = n14139 ;
  assign y2534 = ~1'b0 ;
  assign y2535 = ~n14146 ;
  assign y2536 = ~n14147 ;
  assign y2537 = n14148 ;
  assign y2538 = n14169 ;
  assign y2539 = n14170 ;
  assign y2540 = n14171 ;
  assign y2541 = ~n14172 ;
  assign y2542 = n14173 ;
  assign y2543 = n14176 ;
  assign y2544 = n14179 ;
  assign y2545 = n14180 ;
  assign y2546 = ~1'b0 ;
  assign y2547 = ~n14181 ;
  assign y2548 = ~n14188 ;
  assign y2549 = n14189 ;
  assign y2550 = ~n14197 ;
  assign y2551 = ~n14199 ;
  assign y2552 = ~1'b0 ;
  assign y2553 = ~n14202 ;
  assign y2554 = n14211 ;
  assign y2555 = n5348 ;
  assign y2556 = ~n14214 ;
  assign y2557 = ~n13667 ;
  assign y2558 = ~n14218 ;
  assign y2559 = ~1'b0 ;
  assign y2560 = ~n14221 ;
  assign y2561 = n14230 ;
  assign y2562 = n14239 ;
  assign y2563 = n14242 ;
  assign y2564 = n14244 ;
  assign y2565 = n14245 ;
  assign y2566 = ~n14251 ;
  assign y2567 = ~n14254 ;
  assign y2568 = n14257 ;
  assign y2569 = ~n14260 ;
  assign y2570 = n14262 ;
  assign y2571 = ~n14265 ;
  assign y2572 = n14268 ;
  assign y2573 = ~n14271 ;
  assign y2574 = ~n14277 ;
  assign y2575 = ~n14279 ;
  assign y2576 = n14281 ;
  assign y2577 = n14296 ;
  assign y2578 = n14300 ;
  assign y2579 = ~n14305 ;
  assign y2580 = n14316 ;
  assign y2581 = n14317 ;
  assign y2582 = n14322 ;
  assign y2583 = ~n14325 ;
  assign y2584 = ~n14328 ;
  assign y2585 = ~1'b0 ;
  assign y2586 = n14330 ;
  assign y2587 = ~n14332 ;
  assign y2588 = n14336 ;
  assign y2589 = ~n14341 ;
  assign y2590 = ~n14343 ;
  assign y2591 = n14345 ;
  assign y2592 = n14352 ;
  assign y2593 = ~n14354 ;
  assign y2594 = ~n14360 ;
  assign y2595 = n14370 ;
  assign y2596 = ~n14372 ;
  assign y2597 = ~n14373 ;
  assign y2598 = ~n14375 ;
  assign y2599 = n14382 ;
  assign y2600 = n14386 ;
  assign y2601 = n14394 ;
  assign y2602 = n14402 ;
  assign y2603 = ~n14408 ;
  assign y2604 = n14411 ;
  assign y2605 = n14415 ;
  assign y2606 = ~n14420 ;
  assign y2607 = ~n14423 ;
  assign y2608 = ~1'b0 ;
  assign y2609 = ~n14425 ;
  assign y2610 = ~n14427 ;
  assign y2611 = ~n190 ;
  assign y2612 = n14429 ;
  assign y2613 = n14437 ;
  assign y2614 = ~n14438 ;
  assign y2615 = n14445 ;
  assign y2616 = ~1'b0 ;
  assign y2617 = n940 ;
  assign y2618 = ~n14447 ;
  assign y2619 = n14451 ;
  assign y2620 = ~n14454 ;
  assign y2621 = n14459 ;
  assign y2622 = ~n14461 ;
  assign y2623 = n14463 ;
  assign y2624 = n14465 ;
  assign y2625 = ~n14471 ;
  assign y2626 = n14479 ;
  assign y2627 = ~n14481 ;
  assign y2628 = n14483 ;
  assign y2629 = ~n14485 ;
  assign y2630 = n14487 ;
  assign y2631 = ~n14495 ;
  assign y2632 = n14496 ;
  assign y2633 = ~n14497 ;
  assign y2634 = ~n14500 ;
  assign y2635 = n14501 ;
  assign y2636 = ~n14504 ;
  assign y2637 = ~n14508 ;
  assign y2638 = n14510 ;
  assign y2639 = ~n14515 ;
  assign y2640 = ~n14517 ;
  assign y2641 = n14524 ;
  assign y2642 = ~1'b0 ;
  assign y2643 = ~n14529 ;
  assign y2644 = n14536 ;
  assign y2645 = ~n14538 ;
  assign y2646 = n5991 ;
  assign y2647 = n14540 ;
  assign y2648 = ~n14541 ;
  assign y2649 = ~n14548 ;
  assign y2650 = ~n14551 ;
  assign y2651 = ~n14555 ;
  assign y2652 = ~n14556 ;
  assign y2653 = n14557 ;
  assign y2654 = ~n14561 ;
  assign y2655 = n14563 ;
  assign y2656 = n14568 ;
  assign y2657 = n14569 ;
  assign y2658 = ~n14574 ;
  assign y2659 = n14577 ;
  assign y2660 = n14585 ;
  assign y2661 = n14595 ;
  assign y2662 = ~n14597 ;
  assign y2663 = ~n14598 ;
  assign y2664 = ~n14601 ;
  assign y2665 = ~n14605 ;
  assign y2666 = ~n14613 ;
  assign y2667 = n14618 ;
  assign y2668 = n14621 ;
  assign y2669 = ~n14626 ;
  assign y2670 = n14634 ;
  assign y2671 = n14636 ;
  assign y2672 = ~n14658 ;
  assign y2673 = ~n14663 ;
  assign y2674 = ~n14667 ;
  assign y2675 = n14671 ;
  assign y2676 = n14675 ;
  assign y2677 = ~n14678 ;
  assign y2678 = ~n14679 ;
  assign y2679 = ~n14681 ;
  assign y2680 = n14686 ;
  assign y2681 = ~n14698 ;
  assign y2682 = ~n14699 ;
  assign y2683 = ~n14701 ;
  assign y2684 = n14704 ;
  assign y2685 = n14706 ;
  assign y2686 = n14712 ;
  assign y2687 = n14719 ;
  assign y2688 = ~n14729 ;
  assign y2689 = n14735 ;
  assign y2690 = ~n14736 ;
  assign y2691 = n14737 ;
  assign y2692 = ~n14743 ;
  assign y2693 = ~n14744 ;
  assign y2694 = ~n14747 ;
  assign y2695 = ~n14756 ;
  assign y2696 = n14758 ;
  assign y2697 = n14763 ;
  assign y2698 = n14766 ;
  assign y2699 = n14768 ;
  assign y2700 = ~n14784 ;
  assign y2701 = ~n14787 ;
  assign y2702 = ~n14794 ;
  assign y2703 = ~n14802 ;
  assign y2704 = ~n14805 ;
  assign y2705 = n14808 ;
  assign y2706 = ~n14814 ;
  assign y2707 = ~n14816 ;
  assign y2708 = ~n14824 ;
  assign y2709 = ~n14829 ;
  assign y2710 = n14835 ;
  assign y2711 = n14836 ;
  assign y2712 = n14846 ;
  assign y2713 = n14850 ;
  assign y2714 = ~1'b0 ;
  assign y2715 = ~n14852 ;
  assign y2716 = n14858 ;
  assign y2717 = ~n14865 ;
  assign y2718 = ~n14866 ;
  assign y2719 = n14871 ;
  assign y2720 = ~1'b0 ;
  assign y2721 = ~n14872 ;
  assign y2722 = n14875 ;
  assign y2723 = ~n14878 ;
  assign y2724 = ~n14882 ;
  assign y2725 = ~n14883 ;
  assign y2726 = ~n14890 ;
  assign y2727 = n14892 ;
  assign y2728 = n14893 ;
  assign y2729 = ~n14906 ;
  assign y2730 = n14910 ;
  assign y2731 = ~n14911 ;
  assign y2732 = n14923 ;
  assign y2733 = ~n14924 ;
  assign y2734 = n14925 ;
  assign y2735 = ~n14934 ;
  assign y2736 = ~n14935 ;
  assign y2737 = ~n14939 ;
  assign y2738 = ~n14941 ;
  assign y2739 = ~n14943 ;
  assign y2740 = n14946 ;
  assign y2741 = ~n14960 ;
  assign y2742 = n14962 ;
  assign y2743 = ~n14974 ;
  assign y2744 = n14975 ;
  assign y2745 = n14979 ;
  assign y2746 = ~n14989 ;
  assign y2747 = n14992 ;
  assign y2748 = ~n14998 ;
  assign y2749 = n15000 ;
  assign y2750 = ~1'b0 ;
  assign y2751 = ~n15003 ;
  assign y2752 = n15009 ;
  assign y2753 = ~n15011 ;
  assign y2754 = ~n15014 ;
  assign y2755 = n15025 ;
  assign y2756 = n15027 ;
  assign y2757 = ~n15029 ;
  assign y2758 = ~n15032 ;
  assign y2759 = ~n15043 ;
  assign y2760 = ~n15045 ;
  assign y2761 = ~n15050 ;
  assign y2762 = n15051 ;
  assign y2763 = n15054 ;
  assign y2764 = ~n15065 ;
  assign y2765 = ~n15068 ;
  assign y2766 = ~n15075 ;
  assign y2767 = n15082 ;
  assign y2768 = ~n15083 ;
  assign y2769 = ~n15084 ;
  assign y2770 = ~n15091 ;
  assign y2771 = n15100 ;
  assign y2772 = n15107 ;
  assign y2773 = n15109 ;
  assign y2774 = n15112 ;
  assign y2775 = ~n15114 ;
  assign y2776 = ~n15117 ;
  assign y2777 = ~1'b0 ;
  assign y2778 = ~n15120 ;
  assign y2779 = n15124 ;
  assign y2780 = n15126 ;
  assign y2781 = ~n15131 ;
  assign y2782 = n15136 ;
  assign y2783 = n15140 ;
  assign y2784 = ~n15141 ;
  assign y2785 = ~n15147 ;
  assign y2786 = ~1'b0 ;
  assign y2787 = n15152 ;
  assign y2788 = n15155 ;
  assign y2789 = ~n15156 ;
  assign y2790 = ~n15158 ;
  assign y2791 = ~n15163 ;
  assign y2792 = ~n15164 ;
  assign y2793 = n15166 ;
  assign y2794 = n15168 ;
  assign y2795 = n15171 ;
  assign y2796 = ~n15172 ;
  assign y2797 = ~n15176 ;
  assign y2798 = n15177 ;
  assign y2799 = n15178 ;
  assign y2800 = ~1'b0 ;
  assign y2801 = ~n15179 ;
  assign y2802 = n15180 ;
  assign y2803 = ~1'b0 ;
  assign y2804 = ~n15190 ;
  assign y2805 = n15194 ;
  assign y2806 = ~n15198 ;
  assign y2807 = ~n15200 ;
  assign y2808 = ~n15204 ;
  assign y2809 = ~n15211 ;
  assign y2810 = ~n15212 ;
  assign y2811 = ~n15217 ;
  assign y2812 = ~n15220 ;
  assign y2813 = ~n15222 ;
  assign y2814 = n15230 ;
  assign y2815 = ~n15234 ;
  assign y2816 = n15236 ;
  assign y2817 = ~1'b0 ;
  assign y2818 = n15237 ;
  assign y2819 = n15238 ;
  assign y2820 = n15243 ;
  assign y2821 = n15246 ;
  assign y2822 = ~1'b0 ;
  assign y2823 = ~n15250 ;
  assign y2824 = n15253 ;
  assign y2825 = ~n15259 ;
  assign y2826 = ~n15262 ;
  assign y2827 = ~n15269 ;
  assign y2828 = n15271 ;
  assign y2829 = n15273 ;
  assign y2830 = ~n15275 ;
  assign y2831 = n15278 ;
  assign y2832 = n15284 ;
  assign y2833 = ~n15289 ;
  assign y2834 = ~n15291 ;
  assign y2835 = n15293 ;
  assign y2836 = n15302 ;
  assign y2837 = ~n15306 ;
  assign y2838 = ~n15310 ;
  assign y2839 = ~n15312 ;
  assign y2840 = ~n15314 ;
  assign y2841 = ~n15316 ;
  assign y2842 = n15320 ;
  assign y2843 = ~n15321 ;
  assign y2844 = n15327 ;
  assign y2845 = ~n15340 ;
  assign y2846 = ~n15341 ;
  assign y2847 = ~n15349 ;
  assign y2848 = n15351 ;
  assign y2849 = n15355 ;
  assign y2850 = ~n15359 ;
  assign y2851 = ~n15361 ;
  assign y2852 = ~n15362 ;
  assign y2853 = n15367 ;
  assign y2854 = ~n15368 ;
  assign y2855 = n15369 ;
  assign y2856 = n15373 ;
  assign y2857 = n15379 ;
  assign y2858 = ~n15384 ;
  assign y2859 = ~n15385 ;
  assign y2860 = n15387 ;
  assign y2861 = n15391 ;
  assign y2862 = ~n15392 ;
  assign y2863 = ~n15400 ;
  assign y2864 = ~1'b0 ;
  assign y2865 = ~n15403 ;
  assign y2866 = ~n15409 ;
  assign y2867 = ~n15410 ;
  assign y2868 = ~1'b0 ;
  assign y2869 = n15411 ;
  assign y2870 = n15412 ;
  assign y2871 = n15413 ;
  assign y2872 = ~n15415 ;
  assign y2873 = n15420 ;
  assign y2874 = n15421 ;
  assign y2875 = ~n15425 ;
  assign y2876 = ~n15433 ;
  assign y2877 = n15438 ;
  assign y2878 = n15440 ;
  assign y2879 = ~1'b0 ;
  assign y2880 = ~n15447 ;
  assign y2881 = ~n15453 ;
  assign y2882 = n15460 ;
  assign y2883 = ~n15462 ;
  assign y2884 = n15467 ;
  assign y2885 = ~n15469 ;
  assign y2886 = ~n15471 ;
  assign y2887 = ~n15481 ;
  assign y2888 = ~n15482 ;
  assign y2889 = n15483 ;
  assign y2890 = ~n15485 ;
  assign y2891 = ~n15487 ;
  assign y2892 = n15489 ;
  assign y2893 = n15490 ;
  assign y2894 = ~n15491 ;
  assign y2895 = ~n15492 ;
  assign y2896 = n15497 ;
  assign y2897 = ~n15499 ;
  assign y2898 = n15501 ;
  assign y2899 = ~n15503 ;
  assign y2900 = ~1'b0 ;
  assign y2901 = n15507 ;
  assign y2902 = n15508 ;
  assign y2903 = n15509 ;
  assign y2904 = ~1'b0 ;
  assign y2905 = ~n15512 ;
  assign y2906 = ~n15527 ;
  assign y2907 = n15532 ;
  assign y2908 = ~n15537 ;
  assign y2909 = ~n15538 ;
  assign y2910 = ~n15543 ;
  assign y2911 = n15546 ;
  assign y2912 = n15550 ;
  assign y2913 = n15562 ;
  assign y2914 = ~1'b0 ;
  assign y2915 = ~n15563 ;
  assign y2916 = n15564 ;
  assign y2917 = n15567 ;
  assign y2918 = ~n15571 ;
  assign y2919 = ~n15572 ;
  assign y2920 = n15573 ;
  assign y2921 = ~n15577 ;
  assign y2922 = ~n15580 ;
  assign y2923 = ~n15586 ;
  assign y2924 = ~n15594 ;
  assign y2925 = ~n15599 ;
  assign y2926 = ~n15600 ;
  assign y2927 = ~n15603 ;
  assign y2928 = ~n15606 ;
  assign y2929 = n15607 ;
  assign y2930 = n15609 ;
  assign y2931 = n15616 ;
  assign y2932 = n15624 ;
  assign y2933 = n15626 ;
  assign y2934 = ~n15639 ;
  assign y2935 = n15644 ;
  assign y2936 = ~n15646 ;
  assign y2937 = n15660 ;
  assign y2938 = ~n15662 ;
  assign y2939 = n15668 ;
  assign y2940 = ~1'b0 ;
  assign y2941 = n15679 ;
  assign y2942 = ~n15685 ;
  assign y2943 = n15686 ;
  assign y2944 = ~n15690 ;
  assign y2945 = ~n15691 ;
  assign y2946 = n15693 ;
  assign y2947 = n15695 ;
  assign y2948 = n15704 ;
  assign y2949 = ~1'b0 ;
  assign y2950 = ~n15712 ;
  assign y2951 = n15716 ;
  assign y2952 = ~n15717 ;
  assign y2953 = n15721 ;
  assign y2954 = n15723 ;
  assign y2955 = ~n15727 ;
  assign y2956 = n15729 ;
  assign y2957 = n15731 ;
  assign y2958 = n15741 ;
  assign y2959 = ~n15754 ;
  assign y2960 = ~n15756 ;
  assign y2961 = n15758 ;
  assign y2962 = ~n15760 ;
  assign y2963 = n15761 ;
  assign y2964 = n15763 ;
  assign y2965 = n15764 ;
  assign y2966 = n15765 ;
  assign y2967 = n15768 ;
  assign y2968 = ~n15774 ;
  assign y2969 = ~n15781 ;
  assign y2970 = ~1'b0 ;
  assign y2971 = ~n15782 ;
  assign y2972 = n15783 ;
  assign y2973 = ~n15786 ;
  assign y2974 = n15787 ;
  assign y2975 = n15788 ;
  assign y2976 = n15789 ;
  assign y2977 = n15790 ;
  assign y2978 = ~n15792 ;
  assign y2979 = n15797 ;
  assign y2980 = ~n15798 ;
  assign y2981 = n15803 ;
  assign y2982 = ~n15805 ;
  assign y2983 = ~n15806 ;
  assign y2984 = n15815 ;
  assign y2985 = n15819 ;
  assign y2986 = ~n15824 ;
  assign y2987 = ~n15826 ;
  assign y2988 = ~n15829 ;
  assign y2989 = ~n15830 ;
  assign y2990 = ~1'b0 ;
  assign y2991 = n15831 ;
  assign y2992 = ~n15833 ;
  assign y2993 = n15844 ;
  assign y2994 = n15854 ;
  assign y2995 = ~n15857 ;
  assign y2996 = ~n15860 ;
  assign y2997 = n15867 ;
  assign y2998 = ~n15869 ;
  assign y2999 = ~n15888 ;
  assign y3000 = n15893 ;
  assign y3001 = n15899 ;
  assign y3002 = n15900 ;
  assign y3003 = ~n15906 ;
  assign y3004 = n15910 ;
  assign y3005 = n15914 ;
  assign y3006 = ~1'b0 ;
  assign y3007 = ~1'b0 ;
  assign y3008 = n15916 ;
  assign y3009 = ~n15917 ;
  assign y3010 = ~n15918 ;
  assign y3011 = n15920 ;
  assign y3012 = n15922 ;
  assign y3013 = n15924 ;
  assign y3014 = n15937 ;
  assign y3015 = n15938 ;
  assign y3016 = ~n15941 ;
  assign y3017 = ~n15945 ;
  assign y3018 = ~1'b0 ;
  assign y3019 = ~n15956 ;
  assign y3020 = ~n15958 ;
  assign y3021 = ~n15961 ;
  assign y3022 = ~n15969 ;
  assign y3023 = ~n15976 ;
  assign y3024 = ~n15978 ;
  assign y3025 = n15981 ;
  assign y3026 = n15984 ;
  assign y3027 = ~n15989 ;
  assign y3028 = ~n15990 ;
  assign y3029 = n15991 ;
  assign y3030 = ~n15995 ;
  assign y3031 = n15996 ;
  assign y3032 = n15999 ;
  assign y3033 = n16001 ;
  assign y3034 = n16003 ;
  assign y3035 = n16005 ;
  assign y3036 = n16011 ;
  assign y3037 = n16017 ;
  assign y3038 = ~n16026 ;
  assign y3039 = ~n16029 ;
  assign y3040 = n16034 ;
  assign y3041 = n16036 ;
  assign y3042 = ~n16038 ;
  assign y3043 = n16039 ;
  assign y3044 = ~n16046 ;
  assign y3045 = n16048 ;
  assign y3046 = ~n16050 ;
  assign y3047 = n16059 ;
  assign y3048 = n16067 ;
  assign y3049 = ~n16076 ;
  assign y3050 = ~n16088 ;
  assign y3051 = n16090 ;
  assign y3052 = ~n16095 ;
  assign y3053 = ~n16096 ;
  assign y3054 = ~n16099 ;
  assign y3055 = ~n16106 ;
  assign y3056 = ~n16108 ;
  assign y3057 = ~1'b0 ;
  assign y3058 = ~n16110 ;
  assign y3059 = ~n16114 ;
  assign y3060 = ~n16116 ;
  assign y3061 = n16117 ;
  assign y3062 = n16119 ;
  assign y3063 = n16122 ;
  assign y3064 = n16123 ;
  assign y3065 = ~n16129 ;
  assign y3066 = ~n16137 ;
  assign y3067 = ~n16141 ;
  assign y3068 = ~n16146 ;
  assign y3069 = ~n16152 ;
  assign y3070 = n16159 ;
  assign y3071 = ~n16164 ;
  assign y3072 = ~n16165 ;
  assign y3073 = n16167 ;
  assign y3074 = ~n16170 ;
  assign y3075 = n16176 ;
  assign y3076 = n16177 ;
  assign y3077 = n16180 ;
  assign y3078 = ~n16187 ;
  assign y3079 = n16191 ;
  assign y3080 = ~n16193 ;
  assign y3081 = n16197 ;
  assign y3082 = ~n16201 ;
  assign y3083 = n16203 ;
  assign y3084 = ~n16206 ;
  assign y3085 = ~n16209 ;
  assign y3086 = n16213 ;
  assign y3087 = n16220 ;
  assign y3088 = n16221 ;
  assign y3089 = ~n16230 ;
  assign y3090 = ~n16239 ;
  assign y3091 = n16241 ;
  assign y3092 = ~n16246 ;
  assign y3093 = ~n16252 ;
  assign y3094 = ~n16254 ;
  assign y3095 = ~n16258 ;
  assign y3096 = n16262 ;
  assign y3097 = n16265 ;
  assign y3098 = ~1'b0 ;
  assign y3099 = ~n16267 ;
  assign y3100 = ~n16274 ;
  assign y3101 = n16281 ;
  assign y3102 = ~n16287 ;
  assign y3103 = ~n16293 ;
  assign y3104 = ~n16303 ;
  assign y3105 = ~n16305 ;
  assign y3106 = ~n16307 ;
  assign y3107 = n16308 ;
  assign y3108 = n16310 ;
  assign y3109 = n16311 ;
  assign y3110 = ~n16312 ;
  assign y3111 = ~n16315 ;
  assign y3112 = ~n16320 ;
  assign y3113 = ~n16321 ;
  assign y3114 = ~n4670 ;
  assign y3115 = ~n16325 ;
  assign y3116 = ~n16328 ;
  assign y3117 = n16330 ;
  assign y3118 = ~n16331 ;
  assign y3119 = n16332 ;
  assign y3120 = ~n16334 ;
  assign y3121 = n16337 ;
  assign y3122 = n16341 ;
  assign y3123 = ~n16343 ;
  assign y3124 = n16350 ;
  assign y3125 = n16358 ;
  assign y3126 = n16359 ;
  assign y3127 = ~n16365 ;
  assign y3128 = ~n16372 ;
  assign y3129 = ~n16377 ;
  assign y3130 = ~1'b0 ;
  assign y3131 = n16382 ;
  assign y3132 = ~n16388 ;
  assign y3133 = n16389 ;
  assign y3134 = n16392 ;
  assign y3135 = ~n16394 ;
  assign y3136 = ~n16397 ;
  assign y3137 = n16399 ;
  assign y3138 = ~1'b0 ;
  assign y3139 = n16406 ;
  assign y3140 = n16407 ;
  assign y3141 = ~n16410 ;
  assign y3142 = ~n16414 ;
  assign y3143 = ~n16416 ;
  assign y3144 = ~n16417 ;
  assign y3145 = ~n16424 ;
  assign y3146 = ~n16425 ;
  assign y3147 = n16428 ;
  assign y3148 = n16434 ;
  assign y3149 = ~n16437 ;
  assign y3150 = n16438 ;
  assign y3151 = n16439 ;
  assign y3152 = ~n16444 ;
  assign y3153 = ~n16446 ;
  assign y3154 = ~n16449 ;
  assign y3155 = ~n16450 ;
  assign y3156 = ~n16453 ;
  assign y3157 = ~n16457 ;
  assign y3158 = n16461 ;
  assign y3159 = n16466 ;
  assign y3160 = n16473 ;
  assign y3161 = n16479 ;
  assign y3162 = ~n16481 ;
  assign y3163 = ~1'b0 ;
  assign y3164 = n16488 ;
  assign y3165 = ~n16489 ;
  assign y3166 = ~n16497 ;
  assign y3167 = ~n16498 ;
  assign y3168 = n16501 ;
  assign y3169 = ~n16502 ;
  assign y3170 = n16505 ;
  assign y3171 = n16507 ;
  assign y3172 = n16510 ;
  assign y3173 = n16512 ;
  assign y3174 = ~n16513 ;
  assign y3175 = ~n16516 ;
  assign y3176 = n16520 ;
  assign y3177 = ~n16523 ;
  assign y3178 = n16532 ;
  assign y3179 = ~n16534 ;
  assign y3180 = ~n16537 ;
  assign y3181 = ~n16540 ;
  assign y3182 = ~n16546 ;
  assign y3183 = n16559 ;
  assign y3184 = n16560 ;
  assign y3185 = ~n16562 ;
  assign y3186 = n16564 ;
  assign y3187 = ~n16565 ;
  assign y3188 = ~n16566 ;
  assign y3189 = ~n16572 ;
  assign y3190 = ~1'b0 ;
  assign y3191 = ~n16575 ;
  assign y3192 = ~n16578 ;
  assign y3193 = ~n16581 ;
  assign y3194 = ~n16584 ;
  assign y3195 = ~n16593 ;
  assign y3196 = ~n16598 ;
  assign y3197 = n16600 ;
  assign y3198 = ~n16604 ;
  assign y3199 = n16605 ;
  assign y3200 = ~n16606 ;
  assign y3201 = n16609 ;
  assign y3202 = ~n16613 ;
  assign y3203 = ~n16619 ;
  assign y3204 = ~n16623 ;
  assign y3205 = n16624 ;
  assign y3206 = n16626 ;
  assign y3207 = n16630 ;
  assign y3208 = n16631 ;
  assign y3209 = n16632 ;
  assign y3210 = n16637 ;
  assign y3211 = n16641 ;
  assign y3212 = ~n16646 ;
  assign y3213 = ~n16648 ;
  assign y3214 = ~n16652 ;
  assign y3215 = n5430 ;
  assign y3216 = n16659 ;
  assign y3217 = ~n16663 ;
  assign y3218 = n16664 ;
  assign y3219 = n16666 ;
  assign y3220 = ~n16669 ;
  assign y3221 = n16670 ;
  assign y3222 = ~n16672 ;
  assign y3223 = n16678 ;
  assign y3224 = ~n16679 ;
  assign y3225 = ~n16682 ;
  assign y3226 = ~n16688 ;
  assign y3227 = n16690 ;
  assign y3228 = ~n16694 ;
  assign y3229 = ~1'b0 ;
  assign y3230 = ~n16696 ;
  assign y3231 = ~n16700 ;
  assign y3232 = ~n16703 ;
  assign y3233 = ~n16704 ;
  assign y3234 = ~n16707 ;
  assign y3235 = ~n16708 ;
  assign y3236 = ~n16709 ;
  assign y3237 = n16712 ;
  assign y3238 = ~n16716 ;
  assign y3239 = ~n16718 ;
  assign y3240 = ~n16720 ;
  assign y3241 = n16728 ;
  assign y3242 = n16733 ;
  assign y3243 = n16737 ;
  assign y3244 = n16740 ;
  assign y3245 = ~n16746 ;
  assign y3246 = n16748 ;
  assign y3247 = ~n16749 ;
  assign y3248 = n16757 ;
  assign y3249 = n16759 ;
  assign y3250 = ~n16761 ;
  assign y3251 = n16762 ;
  assign y3252 = ~n16765 ;
  assign y3253 = ~n16768 ;
  assign y3254 = ~n16769 ;
  assign y3255 = ~n16772 ;
  assign y3256 = n16774 ;
  assign y3257 = n16778 ;
  assign y3258 = n16780 ;
  assign y3259 = ~n16789 ;
  assign y3260 = ~n16792 ;
  assign y3261 = n16793 ;
  assign y3262 = n16795 ;
  assign y3263 = ~n16798 ;
  assign y3264 = ~n16799 ;
  assign y3265 = ~n16800 ;
  assign y3266 = ~n16802 ;
  assign y3267 = ~1'b0 ;
  assign y3268 = ~n16807 ;
  assign y3269 = n16809 ;
  assign y3270 = n16811 ;
  assign y3271 = n16813 ;
  assign y3272 = ~n16815 ;
  assign y3273 = n16819 ;
  assign y3274 = n16820 ;
  assign y3275 = ~n16821 ;
  assign y3276 = ~n16823 ;
  assign y3277 = n16826 ;
  assign y3278 = ~n16830 ;
  assign y3279 = ~n16841 ;
  assign y3280 = ~n16843 ;
  assign y3281 = n16848 ;
  assign y3282 = ~1'b0 ;
  assign y3283 = ~n16852 ;
  assign y3284 = n16856 ;
  assign y3285 = n16867 ;
  assign y3286 = n16873 ;
  assign y3287 = n16874 ;
  assign y3288 = ~n16876 ;
  assign y3289 = n16877 ;
  assign y3290 = n16878 ;
  assign y3291 = ~n16883 ;
  assign y3292 = ~n16890 ;
  assign y3293 = n16892 ;
  assign y3294 = n16894 ;
  assign y3295 = ~n16897 ;
  assign y3296 = n16900 ;
  assign y3297 = n16909 ;
  assign y3298 = ~n16914 ;
  assign y3299 = n16915 ;
  assign y3300 = n16919 ;
  assign y3301 = n16920 ;
  assign y3302 = ~n16924 ;
  assign y3303 = n16929 ;
  assign y3304 = n16935 ;
  assign y3305 = n16936 ;
  assign y3306 = n16940 ;
  assign y3307 = ~1'b0 ;
  assign y3308 = ~n16942 ;
  assign y3309 = n16946 ;
  assign y3310 = n16948 ;
  assign y3311 = n16952 ;
  assign y3312 = n16955 ;
  assign y3313 = n16956 ;
  assign y3314 = ~n16958 ;
  assign y3315 = ~1'b0 ;
  assign y3316 = ~n16960 ;
  assign y3317 = ~n16963 ;
  assign y3318 = ~1'b0 ;
  assign y3319 = ~n16964 ;
  assign y3320 = n16973 ;
  assign y3321 = n16977 ;
  assign y3322 = n16981 ;
  assign y3323 = ~n16984 ;
  assign y3324 = n16986 ;
  assign y3325 = n16991 ;
  assign y3326 = ~n16993 ;
  assign y3327 = n16994 ;
  assign y3328 = ~n16998 ;
  assign y3329 = ~n17002 ;
  assign y3330 = n17004 ;
  assign y3331 = n17007 ;
  assign y3332 = n17013 ;
  assign y3333 = ~n17014 ;
  assign y3334 = ~n17017 ;
  assign y3335 = n17021 ;
  assign y3336 = ~n17023 ;
  assign y3337 = ~n17027 ;
  assign y3338 = n17032 ;
  assign y3339 = ~n17034 ;
  assign y3340 = n17038 ;
  assign y3341 = n17042 ;
  assign y3342 = ~n17043 ;
  assign y3343 = n17046 ;
  assign y3344 = ~n17048 ;
  assign y3345 = ~n17050 ;
  assign y3346 = ~n17053 ;
  assign y3347 = ~n17058 ;
  assign y3348 = ~n17063 ;
  assign y3349 = ~n17067 ;
  assign y3350 = ~n17069 ;
  assign y3351 = n17072 ;
  assign y3352 = ~n17078 ;
  assign y3353 = n17079 ;
  assign y3354 = ~n17080 ;
  assign y3355 = ~n17082 ;
  assign y3356 = ~n17083 ;
  assign y3357 = ~n17089 ;
  assign y3358 = ~n17093 ;
  assign y3359 = n17094 ;
  assign y3360 = n17098 ;
  assign y3361 = n17100 ;
  assign y3362 = ~n17104 ;
  assign y3363 = n17106 ;
  assign y3364 = ~n17109 ;
  assign y3365 = n17111 ;
  assign y3366 = n17114 ;
  assign y3367 = n17115 ;
  assign y3368 = ~n17118 ;
  assign y3369 = ~n17120 ;
  assign y3370 = n17124 ;
  assign y3371 = n17126 ;
  assign y3372 = n17127 ;
  assign y3373 = n17131 ;
  assign y3374 = ~n17136 ;
  assign y3375 = ~n17137 ;
  assign y3376 = n17139 ;
  assign y3377 = ~n17140 ;
  assign y3378 = n17141 ;
  assign y3379 = ~n17144 ;
  assign y3380 = n17146 ;
  assign y3381 = ~n17149 ;
  assign y3382 = ~n17152 ;
  assign y3383 = ~n17157 ;
  assign y3384 = ~n17159 ;
  assign y3385 = n17160 ;
  assign y3386 = n17161 ;
  assign y3387 = n17163 ;
  assign y3388 = ~n17168 ;
  assign y3389 = n17173 ;
  assign y3390 = n17177 ;
  assign y3391 = ~n17179 ;
  assign y3392 = ~n17180 ;
  assign y3393 = ~n17182 ;
  assign y3394 = ~n17186 ;
  assign y3395 = ~n17187 ;
  assign y3396 = n17194 ;
  assign y3397 = n17196 ;
  assign y3398 = n17202 ;
  assign y3399 = ~n17204 ;
  assign y3400 = n17212 ;
  assign y3401 = n17221 ;
  assign y3402 = n17225 ;
  assign y3403 = n17227 ;
  assign y3404 = n11829 ;
  assign y3405 = n17229 ;
  assign y3406 = ~n17231 ;
  assign y3407 = ~n17236 ;
  assign y3408 = ~n17244 ;
  assign y3409 = ~n17246 ;
  assign y3410 = ~n17247 ;
  assign y3411 = n17248 ;
  assign y3412 = n17251 ;
  assign y3413 = n17256 ;
  assign y3414 = n17258 ;
  assign y3415 = ~n17259 ;
  assign y3416 = ~n17260 ;
  assign y3417 = n17264 ;
  assign y3418 = ~n17265 ;
  assign y3419 = n17273 ;
  assign y3420 = n17274 ;
  assign y3421 = n17277 ;
  assign y3422 = ~n17278 ;
  assign y3423 = n17281 ;
  assign y3424 = ~n17283 ;
  assign y3425 = n17299 ;
  assign y3426 = n17305 ;
  assign y3427 = ~n17307 ;
  assign y3428 = n17310 ;
  assign y3429 = ~n17313 ;
  assign y3430 = n17317 ;
  assign y3431 = n17318 ;
  assign y3432 = ~n17322 ;
  assign y3433 = ~n17325 ;
  assign y3434 = ~1'b0 ;
  assign y3435 = ~n17327 ;
  assign y3436 = n17335 ;
  assign y3437 = n17341 ;
  assign y3438 = ~n17342 ;
  assign y3439 = n17343 ;
  assign y3440 = ~n17347 ;
  assign y3441 = ~n17348 ;
  assign y3442 = ~n17352 ;
  assign y3443 = ~n17354 ;
  assign y3444 = ~n17362 ;
  assign y3445 = n17364 ;
  assign y3446 = n17369 ;
  assign y3447 = n17374 ;
  assign y3448 = n17376 ;
  assign y3449 = n17380 ;
  assign y3450 = ~n17388 ;
  assign y3451 = n17390 ;
  assign y3452 = ~n17397 ;
  assign y3453 = n17399 ;
  assign y3454 = ~1'b0 ;
  assign y3455 = ~1'b0 ;
  assign y3456 = n17401 ;
  assign y3457 = ~n17409 ;
  assign y3458 = ~n17413 ;
  assign y3459 = ~n17415 ;
  assign y3460 = ~n17418 ;
  assign y3461 = ~n17419 ;
  assign y3462 = n17422 ;
  assign y3463 = n17426 ;
  assign y3464 = ~n17430 ;
  assign y3465 = ~n17431 ;
  assign y3466 = ~n17437 ;
  assign y3467 = ~n17438 ;
  assign y3468 = n17439 ;
  assign y3469 = n17441 ;
  assign y3470 = n17444 ;
  assign y3471 = n17445 ;
  assign y3472 = n17446 ;
  assign y3473 = n17449 ;
  assign y3474 = ~1'b0 ;
  assign y3475 = ~n17456 ;
  assign y3476 = n17457 ;
  assign y3477 = ~n17464 ;
  assign y3478 = n17465 ;
  assign y3479 = n17466 ;
  assign y3480 = n17471 ;
  assign y3481 = ~n17473 ;
  assign y3482 = n17479 ;
  assign y3483 = n17482 ;
  assign y3484 = n17483 ;
  assign y3485 = n17486 ;
  assign y3486 = ~n17487 ;
  assign y3487 = n17492 ;
  assign y3488 = n17495 ;
  assign y3489 = ~1'b0 ;
  assign y3490 = ~n17498 ;
  assign y3491 = ~n17499 ;
  assign y3492 = n17506 ;
  assign y3493 = ~n17508 ;
  assign y3494 = n17513 ;
  assign y3495 = ~n17515 ;
  assign y3496 = n17516 ;
  assign y3497 = ~n17520 ;
  assign y3498 = ~n17522 ;
  assign y3499 = ~n17524 ;
  assign y3500 = n17525 ;
  assign y3501 = n17526 ;
  assign y3502 = n17531 ;
  assign y3503 = n17535 ;
  assign y3504 = ~n17539 ;
  assign y3505 = n17544 ;
  assign y3506 = n17547 ;
  assign y3507 = ~n17555 ;
  assign y3508 = n17558 ;
  assign y3509 = ~1'b0 ;
  assign y3510 = n17561 ;
  assign y3511 = ~n17562 ;
  assign y3512 = ~n17563 ;
  assign y3513 = n17566 ;
  assign y3514 = n17567 ;
  assign y3515 = ~1'b0 ;
  assign y3516 = n17568 ;
  assign y3517 = n17572 ;
  assign y3518 = n17575 ;
  assign y3519 = n17591 ;
  assign y3520 = ~n17592 ;
  assign y3521 = ~n17595 ;
  assign y3522 = n17596 ;
  assign y3523 = ~n17600 ;
  assign y3524 = n17601 ;
  assign y3525 = ~n17602 ;
  assign y3526 = n17613 ;
  assign y3527 = n17615 ;
  assign y3528 = ~n17629 ;
  assign y3529 = n17631 ;
  assign y3530 = ~n17632 ;
  assign y3531 = n17634 ;
  assign y3532 = n17641 ;
  assign y3533 = n17643 ;
  assign y3534 = ~n17644 ;
  assign y3535 = n17648 ;
  assign y3536 = ~n17651 ;
  assign y3537 = n17671 ;
  assign y3538 = n17672 ;
  assign y3539 = ~n17675 ;
  assign y3540 = n17678 ;
  assign y3541 = n17680 ;
  assign y3542 = n17683 ;
  assign y3543 = n17689 ;
  assign y3544 = ~n17693 ;
  assign y3545 = ~n17697 ;
  assign y3546 = n17699 ;
  assign y3547 = n17704 ;
  assign y3548 = ~1'b0 ;
  assign y3549 = ~1'b0 ;
  assign y3550 = n17707 ;
  assign y3551 = n17710 ;
  assign y3552 = n17714 ;
  assign y3553 = ~n17716 ;
  assign y3554 = n17719 ;
  assign y3555 = ~n17721 ;
  assign y3556 = n17725 ;
  assign y3557 = ~1'b0 ;
  assign y3558 = n17728 ;
  assign y3559 = n17733 ;
  assign y3560 = n17735 ;
  assign y3561 = n17740 ;
  assign y3562 = ~n17741 ;
  assign y3563 = ~n17742 ;
  assign y3564 = n17743 ;
  assign y3565 = n17747 ;
  assign y3566 = ~1'b0 ;
  assign y3567 = ~1'b0 ;
  assign y3568 = ~n17750 ;
  assign y3569 = n17752 ;
  assign y3570 = ~n17754 ;
  assign y3571 = ~n17757 ;
  assign y3572 = ~n17758 ;
  assign y3573 = ~n17761 ;
  assign y3574 = n17768 ;
  assign y3575 = n17769 ;
  assign y3576 = ~n17774 ;
  assign y3577 = n17777 ;
  assign y3578 = n17780 ;
  assign y3579 = ~n17782 ;
  assign y3580 = n17783 ;
  assign y3581 = ~n17785 ;
  assign y3582 = n17789 ;
  assign y3583 = n17790 ;
  assign y3584 = n17798 ;
  assign y3585 = ~n17802 ;
  assign y3586 = ~n17803 ;
  assign y3587 = ~n17810 ;
  assign y3588 = ~1'b0 ;
  assign y3589 = n17812 ;
  assign y3590 = n17819 ;
  assign y3591 = n17823 ;
  assign y3592 = n17825 ;
  assign y3593 = ~n17827 ;
  assign y3594 = ~n17828 ;
  assign y3595 = n17829 ;
  assign y3596 = n17833 ;
  assign y3597 = n17834 ;
  assign y3598 = ~n17835 ;
  assign y3599 = n17842 ;
  assign y3600 = ~n17843 ;
  assign y3601 = n17844 ;
  assign y3602 = ~n17854 ;
  assign y3603 = ~n17856 ;
  assign y3604 = ~n17857 ;
  assign y3605 = ~n17860 ;
  assign y3606 = ~n17862 ;
  assign y3607 = ~n17863 ;
  assign y3608 = ~n17866 ;
  assign y3609 = ~n17868 ;
  assign y3610 = n17872 ;
  assign y3611 = n17876 ;
  assign y3612 = ~n17881 ;
  assign y3613 = ~n17882 ;
  assign y3614 = n17884 ;
  assign y3615 = n17887 ;
  assign y3616 = ~n17891 ;
  assign y3617 = n17892 ;
  assign y3618 = ~1'b0 ;
  assign y3619 = n17897 ;
  assign y3620 = ~n17901 ;
  assign y3621 = ~n17903 ;
  assign y3622 = ~n17907 ;
  assign y3623 = ~n17909 ;
  assign y3624 = n17913 ;
  assign y3625 = n17918 ;
  assign y3626 = ~n17919 ;
  assign y3627 = ~n17921 ;
  assign y3628 = ~n17922 ;
  assign y3629 = n17924 ;
  assign y3630 = n17926 ;
  assign y3631 = n17930 ;
  assign y3632 = n17932 ;
  assign y3633 = ~n17935 ;
  assign y3634 = n17937 ;
  assign y3635 = n17939 ;
  assign y3636 = ~n17946 ;
  assign y3637 = n17949 ;
  assign y3638 = n17952 ;
  assign y3639 = ~n17959 ;
  assign y3640 = ~n17964 ;
  assign y3641 = ~n17970 ;
  assign y3642 = n17972 ;
  assign y3643 = ~n17974 ;
  assign y3644 = n17978 ;
  assign y3645 = ~n17979 ;
  assign y3646 = ~n17980 ;
  assign y3647 = ~n17982 ;
  assign y3648 = n17987 ;
  assign y3649 = n17993 ;
  assign y3650 = n18004 ;
  assign y3651 = n18007 ;
  assign y3652 = n18009 ;
  assign y3653 = ~n18010 ;
  assign y3654 = n18019 ;
  assign y3655 = n18022 ;
  assign y3656 = ~n18024 ;
  assign y3657 = n18028 ;
  assign y3658 = n18029 ;
  assign y3659 = ~1'b0 ;
  assign y3660 = n18030 ;
  assign y3661 = ~n18035 ;
  assign y3662 = n18038 ;
  assign y3663 = ~n18042 ;
  assign y3664 = n18043 ;
  assign y3665 = n18047 ;
  assign y3666 = n18051 ;
  assign y3667 = ~n18052 ;
  assign y3668 = n18055 ;
  assign y3669 = ~n18057 ;
  assign y3670 = ~n18058 ;
  assign y3671 = n18059 ;
  assign y3672 = n10578 ;
  assign y3673 = n18064 ;
  assign y3674 = n18067 ;
  assign y3675 = ~n18068 ;
  assign y3676 = ~1'b0 ;
  assign y3677 = ~1'b0 ;
  assign y3678 = n18069 ;
  assign y3679 = ~n18072 ;
  assign y3680 = ~n18075 ;
  assign y3681 = ~n18076 ;
  assign y3682 = n18079 ;
  assign y3683 = ~n18080 ;
  assign y3684 = ~n18082 ;
  assign y3685 = n18083 ;
  assign y3686 = ~n18085 ;
  assign y3687 = ~n18088 ;
  assign y3688 = n18089 ;
  assign y3689 = n18094 ;
  assign y3690 = n18102 ;
  assign y3691 = n18106 ;
  assign y3692 = n18110 ;
  assign y3693 = ~n18111 ;
  assign y3694 = ~n18112 ;
  assign y3695 = ~n18128 ;
  assign y3696 = n18129 ;
  assign y3697 = ~n18135 ;
  assign y3698 = n18137 ;
  assign y3699 = n18141 ;
  assign y3700 = ~n18142 ;
  assign y3701 = n18143 ;
  assign y3702 = ~n18144 ;
  assign y3703 = n18159 ;
  assign y3704 = n18162 ;
  assign y3705 = ~n18163 ;
  assign y3706 = ~n18173 ;
  assign y3707 = ~n18174 ;
  assign y3708 = n18175 ;
  assign y3709 = n18179 ;
  assign y3710 = n18181 ;
  assign y3711 = ~1'b0 ;
  assign y3712 = n18183 ;
  assign y3713 = n18186 ;
  assign y3714 = ~n18188 ;
  assign y3715 = n18192 ;
  assign y3716 = ~n18195 ;
  assign y3717 = n18196 ;
  assign y3718 = ~n18200 ;
  assign y3719 = n18202 ;
  assign y3720 = ~n18208 ;
  assign y3721 = ~n18214 ;
  assign y3722 = ~n18216 ;
  assign y3723 = ~1'b0 ;
  assign y3724 = n18217 ;
  assign y3725 = ~1'b0 ;
  assign y3726 = n18223 ;
  assign y3727 = ~n18229 ;
  assign y3728 = ~n18231 ;
  assign y3729 = ~n18233 ;
  assign y3730 = ~n18241 ;
  assign y3731 = ~n18247 ;
  assign y3732 = ~n18255 ;
  assign y3733 = n18261 ;
  assign y3734 = ~n18263 ;
  assign y3735 = ~n18266 ;
  assign y3736 = ~n18271 ;
  assign y3737 = n18272 ;
  assign y3738 = n18275 ;
  assign y3739 = n18278 ;
  assign y3740 = n18279 ;
  assign y3741 = n18281 ;
  assign y3742 = ~n18283 ;
  assign y3743 = n18285 ;
  assign y3744 = n18290 ;
  assign y3745 = n18298 ;
  assign y3746 = ~n18307 ;
  assign y3747 = n18313 ;
  assign y3748 = n18324 ;
  assign y3749 = n18328 ;
  assign y3750 = ~n18330 ;
  assign y3751 = ~n18331 ;
  assign y3752 = n18333 ;
  assign y3753 = ~n18334 ;
  assign y3754 = n18337 ;
  assign y3755 = ~n18341 ;
  assign y3756 = ~n18343 ;
  assign y3757 = n18346 ;
  assign y3758 = n18348 ;
  assign y3759 = n18353 ;
  assign y3760 = ~n18354 ;
  assign y3761 = ~n18359 ;
  assign y3762 = ~1'b0 ;
  assign y3763 = n18360 ;
  assign y3764 = n18362 ;
  assign y3765 = n18363 ;
  assign y3766 = ~n18364 ;
  assign y3767 = ~n18370 ;
  assign y3768 = ~n18371 ;
  assign y3769 = ~n18374 ;
  assign y3770 = ~n18377 ;
  assign y3771 = n18381 ;
  assign y3772 = ~n18387 ;
  assign y3773 = n18389 ;
  assign y3774 = n18399 ;
  assign y3775 = ~n18402 ;
  assign y3776 = ~1'b0 ;
  assign y3777 = ~n18408 ;
  assign y3778 = ~n18409 ;
  assign y3779 = n18422 ;
  assign y3780 = ~n18425 ;
  assign y3781 = ~n18433 ;
  assign y3782 = ~n18434 ;
  assign y3783 = ~n18435 ;
  assign y3784 = n18440 ;
  assign y3785 = ~n18442 ;
  assign y3786 = n18444 ;
  assign y3787 = ~1'b0 ;
  assign y3788 = ~1'b0 ;
  assign y3789 = ~n18446 ;
  assign y3790 = n18449 ;
  assign y3791 = ~n18452 ;
  assign y3792 = ~n18463 ;
  assign y3793 = n18464 ;
  assign y3794 = n18472 ;
  assign y3795 = n18474 ;
  assign y3796 = n18477 ;
  assign y3797 = n18485 ;
  assign y3798 = n18489 ;
  assign y3799 = ~n18494 ;
  assign y3800 = ~1'b0 ;
  assign y3801 = ~n18498 ;
  assign y3802 = n18502 ;
  assign y3803 = n18509 ;
  assign y3804 = n18510 ;
  assign y3805 = n18513 ;
  assign y3806 = ~n18516 ;
  assign y3807 = ~n18520 ;
  assign y3808 = ~n18521 ;
  assign y3809 = ~n18527 ;
  assign y3810 = ~n18529 ;
  assign y3811 = n18534 ;
  assign y3812 = ~n18536 ;
  assign y3813 = ~n18545 ;
  assign y3814 = n18547 ;
  assign y3815 = n18549 ;
  assign y3816 = ~n18550 ;
  assign y3817 = ~n18551 ;
  assign y3818 = ~n18555 ;
  assign y3819 = n18561 ;
  assign y3820 = n18564 ;
  assign y3821 = n18574 ;
  assign y3822 = ~n18586 ;
  assign y3823 = ~n18587 ;
  assign y3824 = ~n18590 ;
  assign y3825 = ~n18591 ;
  assign y3826 = n18594 ;
  assign y3827 = n18596 ;
  assign y3828 = ~n18601 ;
  assign y3829 = n18603 ;
  assign y3830 = n18605 ;
  assign y3831 = ~n18607 ;
  assign y3832 = ~n18610 ;
  assign y3833 = n18615 ;
  assign y3834 = ~n18618 ;
  assign y3835 = ~n18626 ;
  assign y3836 = ~n18628 ;
  assign y3837 = ~n18629 ;
  assign y3838 = n18634 ;
  assign y3839 = ~n18635 ;
  assign y3840 = ~n18637 ;
  assign y3841 = ~n18639 ;
  assign y3842 = ~n18641 ;
  assign y3843 = ~n18643 ;
  assign y3844 = ~n18648 ;
  assign y3845 = n18651 ;
  assign y3846 = ~n18653 ;
  assign y3847 = ~n18658 ;
  assign y3848 = ~n18664 ;
  assign y3849 = ~n18675 ;
  assign y3850 = n18681 ;
  assign y3851 = n18687 ;
  assign y3852 = n18688 ;
  assign y3853 = n18697 ;
  assign y3854 = ~n18700 ;
  assign y3855 = ~1'b0 ;
  assign y3856 = n18703 ;
  assign y3857 = ~n18704 ;
  assign y3858 = ~n18705 ;
  assign y3859 = ~n18707 ;
  assign y3860 = n10055 ;
  assign y3861 = ~n18709 ;
  assign y3862 = ~n18710 ;
  assign y3863 = n18724 ;
  assign y3864 = ~n18727 ;
  assign y3865 = ~n18732 ;
  assign y3866 = ~n18733 ;
  assign y3867 = n18738 ;
  assign y3868 = ~n18742 ;
  assign y3869 = ~n18743 ;
  assign y3870 = n18746 ;
  assign y3871 = n18751 ;
  assign y3872 = n18755 ;
  assign y3873 = n18759 ;
  assign y3874 = n18765 ;
  assign y3875 = n18767 ;
  assign y3876 = n18769 ;
  assign y3877 = ~1'b0 ;
  assign y3878 = n18770 ;
  assign y3879 = n18771 ;
  assign y3880 = n18772 ;
  assign y3881 = n18780 ;
  assign y3882 = n18783 ;
  assign y3883 = ~n18785 ;
  assign y3884 = n18788 ;
  assign y3885 = ~n18795 ;
  assign y3886 = ~n18797 ;
  assign y3887 = n18800 ;
  assign y3888 = ~n18803 ;
  assign y3889 = n18804 ;
  assign y3890 = ~n18806 ;
  assign y3891 = ~n18809 ;
  assign y3892 = n18810 ;
  assign y3893 = ~n18811 ;
  assign y3894 = ~n18814 ;
  assign y3895 = n18817 ;
  assign y3896 = n18820 ;
  assign y3897 = ~n18821 ;
  assign y3898 = ~n18823 ;
  assign y3899 = n18827 ;
  assign y3900 = n18828 ;
  assign y3901 = n18829 ;
  assign y3902 = ~n18831 ;
  assign y3903 = n18832 ;
  assign y3904 = n18833 ;
  assign y3905 = n18834 ;
  assign y3906 = n18837 ;
  assign y3907 = ~n18839 ;
  assign y3908 = n18840 ;
  assign y3909 = ~n18843 ;
  assign y3910 = n18846 ;
  assign y3911 = n18847 ;
  assign y3912 = n18848 ;
  assign y3913 = n18849 ;
  assign y3914 = n18851 ;
  assign y3915 = ~1'b0 ;
  assign y3916 = n18853 ;
  assign y3917 = ~n18856 ;
  assign y3918 = ~n18858 ;
  assign y3919 = n18861 ;
  assign y3920 = ~n18862 ;
  assign y3921 = ~n18864 ;
  assign y3922 = n18865 ;
  assign y3923 = n18866 ;
  assign y3924 = ~n18869 ;
  assign y3925 = ~n18872 ;
  assign y3926 = n18875 ;
  assign y3927 = ~n18879 ;
  assign y3928 = n18888 ;
  assign y3929 = n18892 ;
  assign y3930 = ~n18893 ;
  assign y3931 = n18896 ;
  assign y3932 = ~n18899 ;
  assign y3933 = ~n18903 ;
  assign y3934 = n18905 ;
  assign y3935 = n18908 ;
  assign y3936 = ~n18915 ;
  assign y3937 = ~n18920 ;
  assign y3938 = ~1'b0 ;
  assign y3939 = ~n18929 ;
  assign y3940 = n18930 ;
  assign y3941 = ~n18932 ;
  assign y3942 = ~n18941 ;
  assign y3943 = n18944 ;
  assign y3944 = ~n18945 ;
  assign y3945 = ~n18946 ;
  assign y3946 = ~n18950 ;
  assign y3947 = ~n18952 ;
  assign y3948 = ~n18955 ;
  assign y3949 = ~n18956 ;
  assign y3950 = ~n18962 ;
  assign y3951 = ~n18965 ;
  assign y3952 = n18969 ;
  assign y3953 = n18974 ;
  assign y3954 = n18978 ;
  assign y3955 = n18987 ;
  assign y3956 = ~n18988 ;
  assign y3957 = ~n18991 ;
  assign y3958 = n18992 ;
  assign y3959 = ~n18993 ;
  assign y3960 = n18995 ;
  assign y3961 = ~n18997 ;
  assign y3962 = ~n18998 ;
  assign y3963 = ~n19001 ;
  assign y3964 = ~n19003 ;
  assign y3965 = n19006 ;
  assign y3966 = n19008 ;
  assign y3967 = ~n19010 ;
  assign y3968 = ~n19011 ;
  assign y3969 = ~n19015 ;
  assign y3970 = ~n19018 ;
  assign y3971 = n19022 ;
  assign y3972 = n19023 ;
  assign y3973 = ~n19028 ;
  assign y3974 = n19029 ;
  assign y3975 = n19030 ;
  assign y3976 = n19031 ;
  assign y3977 = ~n19035 ;
  assign y3978 = ~n19039 ;
  assign y3979 = ~n19042 ;
  assign y3980 = ~n19044 ;
  assign y3981 = n19045 ;
  assign y3982 = ~n19046 ;
  assign y3983 = ~n19048 ;
  assign y3984 = n19049 ;
  assign y3985 = ~n19050 ;
  assign y3986 = n19051 ;
  assign y3987 = ~n19054 ;
  assign y3988 = ~n19061 ;
  assign y3989 = n19065 ;
  assign y3990 = n19066 ;
  assign y3991 = ~n19067 ;
  assign y3992 = n19069 ;
  assign y3993 = n19072 ;
  assign y3994 = ~n19078 ;
  assign y3995 = ~n19079 ;
  assign y3996 = ~n19081 ;
  assign y3997 = ~1'b0 ;
  assign y3998 = ~n19084 ;
  assign y3999 = n19088 ;
  assign y4000 = n19097 ;
  assign y4001 = n19098 ;
  assign y4002 = ~n19099 ;
  assign y4003 = n19100 ;
  assign y4004 = ~n19101 ;
  assign y4005 = n19107 ;
  assign y4006 = n19108 ;
  assign y4007 = n19112 ;
  assign y4008 = n19122 ;
  assign y4009 = ~n19125 ;
  assign y4010 = ~n19128 ;
  assign y4011 = ~n19129 ;
  assign y4012 = ~n19130 ;
  assign y4013 = ~n19132 ;
  assign y4014 = n19134 ;
  assign y4015 = n19136 ;
  assign y4016 = n19145 ;
  assign y4017 = ~n19146 ;
  assign y4018 = n19147 ;
  assign y4019 = ~n19148 ;
  assign y4020 = ~n19151 ;
  assign y4021 = n19157 ;
  assign y4022 = ~n19167 ;
  assign y4023 = n19172 ;
  assign y4024 = ~n19173 ;
  assign y4025 = ~n19179 ;
  assign y4026 = ~n19181 ;
  assign y4027 = ~n19188 ;
  assign y4028 = n19190 ;
  assign y4029 = n19191 ;
  assign y4030 = ~n19192 ;
  assign y4031 = ~n19194 ;
  assign y4032 = n19200 ;
  assign y4033 = n19203 ;
  assign y4034 = n19205 ;
  assign y4035 = n19207 ;
  assign y4036 = n19209 ;
  assign y4037 = n19211 ;
  assign y4038 = ~n19214 ;
  assign y4039 = ~n19218 ;
  assign y4040 = n19222 ;
  assign y4041 = ~n19227 ;
  assign y4042 = n19229 ;
  assign y4043 = ~n19234 ;
  assign y4044 = n19238 ;
  assign y4045 = ~1'b0 ;
  assign y4046 = n19240 ;
  assign y4047 = n19242 ;
  assign y4048 = n19243 ;
  assign y4049 = n19248 ;
  assign y4050 = ~n19252 ;
  assign y4051 = n19254 ;
  assign y4052 = ~1'b0 ;
  assign y4053 = ~n19255 ;
  assign y4054 = ~n19256 ;
  assign y4055 = n19258 ;
  assign y4056 = ~n19263 ;
  assign y4057 = ~n19264 ;
  assign y4058 = ~n19278 ;
  assign y4059 = ~n19279 ;
  assign y4060 = n19280 ;
  assign y4061 = ~n19285 ;
  assign y4062 = ~n19291 ;
  assign y4063 = n19292 ;
  assign y4064 = ~n19298 ;
  assign y4065 = ~n19302 ;
  assign y4066 = n19307 ;
  assign y4067 = n19309 ;
  assign y4068 = ~n19312 ;
  assign y4069 = n19317 ;
  assign y4070 = n19327 ;
  assign y4071 = ~n19332 ;
  assign y4072 = n19335 ;
  assign y4073 = n19341 ;
  assign y4074 = ~n19342 ;
  assign y4075 = ~1'b0 ;
  assign y4076 = n19344 ;
  assign y4077 = n19347 ;
  assign y4078 = ~n19355 ;
  assign y4079 = n19373 ;
  assign y4080 = ~n19377 ;
  assign y4081 = ~1'b0 ;
  assign y4082 = ~1'b0 ;
  assign y4083 = ~n19378 ;
  assign y4084 = n19380 ;
  assign y4085 = n19382 ;
  assign y4086 = ~1'b0 ;
  assign y4087 = ~n19383 ;
  assign y4088 = n19387 ;
  assign y4089 = n19389 ;
  assign y4090 = n19390 ;
  assign y4091 = n19392 ;
  assign y4092 = ~1'b0 ;
  assign y4093 = n19397 ;
  assign y4094 = ~n19400 ;
  assign y4095 = ~n19401 ;
  assign y4096 = n19402 ;
  assign y4097 = ~1'b0 ;
  assign y4098 = ~n19404 ;
  assign y4099 = n19408 ;
  assign y4100 = ~n19412 ;
  assign y4101 = ~n19415 ;
  assign y4102 = ~n19427 ;
  assign y4103 = n19432 ;
  assign y4104 = n19437 ;
  assign y4105 = n19438 ;
  assign y4106 = ~n19439 ;
  assign y4107 = ~n19448 ;
  assign y4108 = n19453 ;
  assign y4109 = ~n19456 ;
  assign y4110 = ~n19458 ;
  assign y4111 = n19463 ;
  assign y4112 = ~n19466 ;
  assign y4113 = ~n19471 ;
  assign y4114 = n19478 ;
  assign y4115 = n19479 ;
  assign y4116 = ~n19484 ;
  assign y4117 = ~1'b0 ;
  assign y4118 = n19486 ;
  assign y4119 = n19487 ;
  assign y4120 = n19490 ;
  assign y4121 = ~1'b0 ;
  assign y4122 = n19494 ;
  assign y4123 = n19496 ;
  assign y4124 = ~n19499 ;
  assign y4125 = n19503 ;
  assign y4126 = ~n19516 ;
  assign y4127 = n19518 ;
  assign y4128 = ~1'b0 ;
  assign y4129 = ~n19521 ;
  assign y4130 = n19525 ;
  assign y4131 = ~n19528 ;
  assign y4132 = ~n19529 ;
  assign y4133 = ~n19535 ;
  assign y4134 = n19536 ;
  assign y4135 = n19538 ;
  assign y4136 = ~n19539 ;
  assign y4137 = n19543 ;
  assign y4138 = n19547 ;
  assign y4139 = ~1'b0 ;
  assign y4140 = n19552 ;
  assign y4141 = n19553 ;
  assign y4142 = n19556 ;
  assign y4143 = ~n19558 ;
  assign y4144 = ~n19560 ;
  assign y4145 = ~1'b0 ;
  assign y4146 = ~n19564 ;
  assign y4147 = n19570 ;
  assign y4148 = ~n19573 ;
  assign y4149 = n19574 ;
  assign y4150 = ~n19578 ;
  assign y4151 = ~n19583 ;
  assign y4152 = n19589 ;
  assign y4153 = n19591 ;
  assign y4154 = n19592 ;
  assign y4155 = n19595 ;
  assign y4156 = ~n19596 ;
  assign y4157 = ~n19600 ;
  assign y4158 = ~n19602 ;
  assign y4159 = n19604 ;
  assign y4160 = n19605 ;
  assign y4161 = ~n19609 ;
  assign y4162 = n19612 ;
  assign y4163 = n19614 ;
  assign y4164 = ~n19618 ;
  assign y4165 = ~n19619 ;
  assign y4166 = ~n19622 ;
  assign y4167 = n19625 ;
  assign y4168 = n19627 ;
  assign y4169 = n19633 ;
  assign y4170 = ~n19635 ;
  assign y4171 = ~n19639 ;
  assign y4172 = ~n19642 ;
  assign y4173 = n19644 ;
  assign y4174 = n19647 ;
  assign y4175 = ~n19649 ;
  assign y4176 = ~1'b0 ;
  assign y4177 = n19650 ;
  assign y4178 = n19652 ;
  assign y4179 = ~n19654 ;
  assign y4180 = ~1'b0 ;
  assign y4181 = ~n19657 ;
  assign y4182 = n19661 ;
  assign y4183 = ~n19663 ;
  assign y4184 = ~n19669 ;
  assign y4185 = n19676 ;
  assign y4186 = n19677 ;
  assign y4187 = ~n19680 ;
  assign y4188 = n19682 ;
  assign y4189 = ~n19691 ;
  assign y4190 = n19694 ;
  assign y4191 = ~n19696 ;
  assign y4192 = ~n19697 ;
  assign y4193 = n19700 ;
  assign y4194 = ~n19703 ;
  assign y4195 = ~n19704 ;
  assign y4196 = ~n19705 ;
  assign y4197 = n19706 ;
  assign y4198 = ~n19707 ;
  assign y4199 = ~n19711 ;
  assign y4200 = n19717 ;
  assign y4201 = ~1'b0 ;
  assign y4202 = n19718 ;
  assign y4203 = ~n19720 ;
  assign y4204 = n19724 ;
  assign y4205 = ~n19730 ;
  assign y4206 = n19736 ;
  assign y4207 = ~n19738 ;
  assign y4208 = ~n19739 ;
  assign y4209 = ~n19748 ;
  assign y4210 = n19751 ;
  assign y4211 = ~n19756 ;
  assign y4212 = n19763 ;
  assign y4213 = ~n19767 ;
  assign y4214 = ~n19768 ;
  assign y4215 = ~n19771 ;
  assign y4216 = ~n19778 ;
  assign y4217 = n19779 ;
  assign y4218 = n19789 ;
  assign y4219 = ~n19797 ;
  assign y4220 = n19804 ;
  assign y4221 = ~n19808 ;
  assign y4222 = ~n19811 ;
  assign y4223 = n19813 ;
  assign y4224 = ~n19817 ;
  assign y4225 = n19821 ;
  assign y4226 = n19822 ;
  assign y4227 = n19824 ;
  assign y4228 = ~1'b0 ;
  assign y4229 = ~n19827 ;
  assign y4230 = ~n19828 ;
  assign y4231 = ~n19831 ;
  assign y4232 = n4970 ;
  assign y4233 = n19834 ;
  assign y4234 = n19840 ;
  assign y4235 = ~n19841 ;
  assign y4236 = n19842 ;
  assign y4237 = ~n19845 ;
  assign y4238 = ~n19846 ;
  assign y4239 = n19848 ;
  assign y4240 = n19849 ;
  assign y4241 = n19852 ;
  assign y4242 = ~n19857 ;
  assign y4243 = n19858 ;
  assign y4244 = ~n19860 ;
  assign y4245 = ~n19861 ;
  assign y4246 = n19862 ;
  assign y4247 = ~n19864 ;
  assign y4248 = ~n19866 ;
  assign y4249 = n19867 ;
  assign y4250 = ~n19871 ;
  assign y4251 = ~n19872 ;
  assign y4252 = n19877 ;
  assign y4253 = ~n19880 ;
  assign y4254 = n19881 ;
  assign y4255 = n19883 ;
  assign y4256 = n19892 ;
  assign y4257 = ~n19897 ;
  assign y4258 = n19898 ;
  assign y4259 = n19901 ;
  assign y4260 = n19904 ;
  assign y4261 = n19905 ;
  assign y4262 = ~n19907 ;
  assign y4263 = n19910 ;
  assign y4264 = n19916 ;
  assign y4265 = ~1'b0 ;
  assign y4266 = ~n19918 ;
  assign y4267 = n19927 ;
  assign y4268 = ~n19930 ;
  assign y4269 = ~n19932 ;
  assign y4270 = n19933 ;
  assign y4271 = ~n19941 ;
  assign y4272 = ~n19942 ;
  assign y4273 = ~n19943 ;
  assign y4274 = n19949 ;
  assign y4275 = ~1'b0 ;
  assign y4276 = ~1'b0 ;
  assign y4277 = ~n19950 ;
  assign y4278 = ~n19953 ;
  assign y4279 = ~n19954 ;
  assign y4280 = ~n19957 ;
  assign y4281 = ~n19961 ;
  assign y4282 = n19962 ;
  assign y4283 = ~n19970 ;
  assign y4284 = ~n19971 ;
  assign y4285 = n19972 ;
  assign y4286 = ~n19974 ;
  assign y4287 = ~n19976 ;
  assign y4288 = ~n19977 ;
  assign y4289 = n19979 ;
  assign y4290 = ~n19981 ;
  assign y4291 = ~n19982 ;
  assign y4292 = n4678 ;
  assign y4293 = ~n19983 ;
  assign y4294 = n19984 ;
  assign y4295 = ~n19988 ;
  assign y4296 = ~n19995 ;
  assign y4297 = n19998 ;
  assign y4298 = ~n19999 ;
  assign y4299 = ~n20000 ;
  assign y4300 = ~n20006 ;
  assign y4301 = n20008 ;
  assign y4302 = n20012 ;
  assign y4303 = ~n20014 ;
  assign y4304 = ~n20017 ;
  assign y4305 = ~n20024 ;
  assign y4306 = ~n20029 ;
  assign y4307 = n20031 ;
  assign y4308 = n20035 ;
  assign y4309 = n20037 ;
  assign y4310 = ~n20046 ;
  assign y4311 = n20050 ;
  assign y4312 = ~n20052 ;
  assign y4313 = ~n20055 ;
  assign y4314 = ~n20056 ;
  assign y4315 = ~n20060 ;
  assign y4316 = ~n20063 ;
  assign y4317 = n20065 ;
  assign y4318 = n20070 ;
  assign y4319 = ~n20071 ;
  assign y4320 = ~1'b0 ;
  assign y4321 = n20073 ;
  assign y4322 = ~n20074 ;
  assign y4323 = n12687 ;
  assign y4324 = n20076 ;
  assign y4325 = ~n20080 ;
  assign y4326 = ~n20083 ;
  assign y4327 = n20087 ;
  assign y4328 = ~n20090 ;
  assign y4329 = n20092 ;
  assign y4330 = ~n20093 ;
  assign y4331 = ~n20094 ;
  assign y4332 = ~n20097 ;
  assign y4333 = n20099 ;
  assign y4334 = ~n20100 ;
  assign y4335 = n20109 ;
  assign y4336 = ~n20110 ;
  assign y4337 = ~n20111 ;
  assign y4338 = ~n20116 ;
  assign y4339 = ~1'b0 ;
  assign y4340 = ~n20118 ;
  assign y4341 = n20121 ;
  assign y4342 = n20122 ;
  assign y4343 = ~n20123 ;
  assign y4344 = n20126 ;
  assign y4345 = n20128 ;
  assign y4346 = ~n20129 ;
  assign y4347 = ~n20133 ;
  assign y4348 = n20134 ;
  assign y4349 = ~n20140 ;
  assign y4350 = ~n20141 ;
  assign y4351 = ~n20142 ;
  assign y4352 = n20143 ;
  assign y4353 = ~n20144 ;
  assign y4354 = ~n20149 ;
  assign y4355 = n20154 ;
  assign y4356 = ~n20155 ;
  assign y4357 = n20161 ;
  assign y4358 = n20165 ;
  assign y4359 = n20170 ;
  assign y4360 = n20172 ;
  assign y4361 = n20173 ;
  assign y4362 = ~n20174 ;
  assign y4363 = ~n20175 ;
  assign y4364 = ~n20180 ;
  assign y4365 = ~n20182 ;
  assign y4366 = n20184 ;
  assign y4367 = n20186 ;
  assign y4368 = ~n20193 ;
  assign y4369 = n20195 ;
  assign y4370 = n20199 ;
  assign y4371 = n20202 ;
  assign y4372 = ~n20204 ;
  assign y4373 = n20211 ;
  assign y4374 = ~n20215 ;
  assign y4375 = ~n20221 ;
  assign y4376 = n20222 ;
  assign y4377 = ~n20223 ;
  assign y4378 = n20228 ;
  assign y4379 = ~n20237 ;
  assign y4380 = n20241 ;
  assign y4381 = ~n20242 ;
  assign y4382 = ~n20243 ;
  assign y4383 = ~n20247 ;
  assign y4384 = ~n20249 ;
  assign y4385 = n20257 ;
  assign y4386 = n20259 ;
  assign y4387 = n20263 ;
  assign y4388 = ~n20264 ;
  assign y4389 = ~n20266 ;
  assign y4390 = n20267 ;
  assign y4391 = n20270 ;
  assign y4392 = n20271 ;
  assign y4393 = ~n20278 ;
  assign y4394 = n20280 ;
  assign y4395 = ~n20282 ;
  assign y4396 = ~n20286 ;
  assign y4397 = n20287 ;
  assign y4398 = n20290 ;
  assign y4399 = ~1'b0 ;
  assign y4400 = ~n20297 ;
  assign y4401 = ~n20299 ;
  assign y4402 = ~n20303 ;
  assign y4403 = ~n20309 ;
  assign y4404 = ~n20311 ;
  assign y4405 = n20314 ;
  assign y4406 = ~n20318 ;
  assign y4407 = ~n20320 ;
  assign y4408 = ~1'b0 ;
  assign y4409 = ~n20321 ;
  assign y4410 = ~n20323 ;
  assign y4411 = n20324 ;
  assign y4412 = ~n20325 ;
  assign y4413 = n20329 ;
  assign y4414 = ~n20331 ;
  assign y4415 = ~n20332 ;
  assign y4416 = n20335 ;
  assign y4417 = n20338 ;
  assign y4418 = n20339 ;
  assign y4419 = n20341 ;
  assign y4420 = n20349 ;
  assign y4421 = ~n20351 ;
  assign y4422 = n20356 ;
  assign y4423 = ~n20360 ;
  assign y4424 = ~n20361 ;
  assign y4425 = ~n20364 ;
  assign y4426 = ~n20366 ;
  assign y4427 = ~n20368 ;
  assign y4428 = n20369 ;
  assign y4429 = ~n20370 ;
  assign y4430 = n20371 ;
  assign y4431 = n20374 ;
  assign y4432 = ~n20375 ;
  assign y4433 = ~n20377 ;
  assign y4434 = ~n20387 ;
  assign y4435 = ~n20394 ;
  assign y4436 = n20399 ;
  assign y4437 = n20403 ;
  assign y4438 = ~n20404 ;
  assign y4439 = n20407 ;
  assign y4440 = n20408 ;
  assign y4441 = n20411 ;
  assign y4442 = n20416 ;
  assign y4443 = ~n20420 ;
  assign y4444 = n20427 ;
  assign y4445 = n20429 ;
  assign y4446 = n20430 ;
  assign y4447 = ~n20434 ;
  assign y4448 = n20437 ;
  assign y4449 = ~n20440 ;
  assign y4450 = n20445 ;
  assign y4451 = ~n20446 ;
  assign y4452 = ~n20448 ;
  assign y4453 = ~1'b0 ;
  assign y4454 = ~n20450 ;
  assign y4455 = ~n20454 ;
  assign y4456 = n20459 ;
  assign y4457 = ~n20461 ;
  assign y4458 = ~n20464 ;
  assign y4459 = ~n20471 ;
  assign y4460 = ~n20472 ;
  assign y4461 = n20473 ;
  assign y4462 = ~n20479 ;
  assign y4463 = ~n20480 ;
  assign y4464 = n20481 ;
  assign y4465 = ~n20487 ;
  assign y4466 = ~n20488 ;
  assign y4467 = n20493 ;
  assign y4468 = ~n20500 ;
  assign y4469 = ~n20502 ;
  assign y4470 = ~n20505 ;
  assign y4471 = ~1'b0 ;
  assign y4472 = ~n20506 ;
  assign y4473 = ~n20507 ;
  assign y4474 = ~n20509 ;
  assign y4475 = n20510 ;
  assign y4476 = ~1'b0 ;
  assign y4477 = ~n20511 ;
  assign y4478 = n20519 ;
  assign y4479 = n20521 ;
  assign y4480 = ~n20527 ;
  assign y4481 = n20530 ;
  assign y4482 = n20533 ;
  assign y4483 = n20537 ;
  assign y4484 = n20539 ;
  assign y4485 = ~n20545 ;
  assign y4486 = ~n20546 ;
  assign y4487 = n20549 ;
  assign y4488 = ~n20550 ;
  assign y4489 = n20551 ;
  assign y4490 = ~n20555 ;
  assign y4491 = ~n20557 ;
  assign y4492 = ~1'b0 ;
  assign y4493 = n20562 ;
  assign y4494 = ~n20567 ;
  assign y4495 = ~n20569 ;
  assign y4496 = n20572 ;
  assign y4497 = ~n20574 ;
  assign y4498 = ~1'b0 ;
  assign y4499 = ~n20580 ;
  assign y4500 = ~n20586 ;
  assign y4501 = ~n20589 ;
  assign y4502 = n20590 ;
  assign y4503 = ~n20593 ;
  assign y4504 = n20594 ;
  assign y4505 = ~n20596 ;
  assign y4506 = n20607 ;
  assign y4507 = ~n20610 ;
  assign y4508 = n20613 ;
  assign y4509 = n20617 ;
  assign y4510 = n20619 ;
  assign y4511 = ~n20624 ;
  assign y4512 = ~n20625 ;
  assign y4513 = n20626 ;
  assign y4514 = n20628 ;
  assign y4515 = ~n20630 ;
  assign y4516 = n20633 ;
  assign y4517 = n20634 ;
  assign y4518 = n20637 ;
  assign y4519 = n20641 ;
  assign y4520 = ~n20644 ;
  assign y4521 = ~n20653 ;
  assign y4522 = n20658 ;
  assign y4523 = ~n20661 ;
  assign y4524 = ~n20666 ;
  assign y4525 = ~n20669 ;
  assign y4526 = ~n20671 ;
  assign y4527 = n20673 ;
  assign y4528 = n20677 ;
  assign y4529 = n20679 ;
  assign y4530 = n20682 ;
  assign y4531 = ~n20684 ;
  assign y4532 = ~n20685 ;
  assign y4533 = ~n20686 ;
  assign y4534 = ~n20695 ;
  assign y4535 = n20696 ;
  assign y4536 = ~1'b0 ;
  assign y4537 = n20698 ;
  assign y4538 = ~n20704 ;
  assign y4539 = n20710 ;
  assign y4540 = n20717 ;
  assign y4541 = n20721 ;
  assign y4542 = n20731 ;
  assign y4543 = n20734 ;
  assign y4544 = n20736 ;
  assign y4545 = ~n20740 ;
  assign y4546 = ~n20742 ;
  assign y4547 = ~n20745 ;
  assign y4548 = n20747 ;
  assign y4549 = n20753 ;
  assign y4550 = ~n20756 ;
  assign y4551 = n20757 ;
  assign y4552 = ~n20759 ;
  assign y4553 = n20763 ;
  assign y4554 = n20766 ;
  assign y4555 = ~n20769 ;
  assign y4556 = ~n20771 ;
  assign y4557 = ~1'b0 ;
  assign y4558 = ~n20772 ;
  assign y4559 = ~n20773 ;
  assign y4560 = n20775 ;
  assign y4561 = ~n20777 ;
  assign y4562 = n20779 ;
  assign y4563 = n20784 ;
  assign y4564 = ~1'b0 ;
  assign y4565 = n20786 ;
  assign y4566 = ~n20788 ;
  assign y4567 = ~n20790 ;
  assign y4568 = ~n20791 ;
  assign y4569 = n20793 ;
  assign y4570 = ~n20796 ;
  assign y4571 = ~n20801 ;
  assign y4572 = n20803 ;
  assign y4573 = n20810 ;
  assign y4574 = n20811 ;
  assign y4575 = ~n20813 ;
  assign y4576 = ~n20815 ;
  assign y4577 = ~n20818 ;
  assign y4578 = ~n20822 ;
  assign y4579 = ~n20824 ;
  assign y4580 = ~1'b0 ;
  assign y4581 = n20826 ;
  assign y4582 = ~n20827 ;
  assign y4583 = ~n20830 ;
  assign y4584 = n20831 ;
  assign y4585 = ~1'b0 ;
  assign y4586 = ~n20832 ;
  assign y4587 = n20835 ;
  assign y4588 = n20836 ;
  assign y4589 = ~n20840 ;
  assign y4590 = n20843 ;
  assign y4591 = ~n20845 ;
  assign y4592 = ~n20847 ;
  assign y4593 = ~n20850 ;
  assign y4594 = ~n20852 ;
  assign y4595 = ~n20854 ;
  assign y4596 = n20856 ;
  assign y4597 = ~n20860 ;
  assign y4598 = ~n20866 ;
  assign y4599 = ~n20867 ;
  assign y4600 = n20870 ;
  assign y4601 = ~n20874 ;
  assign y4602 = n20875 ;
  assign y4603 = n20883 ;
  assign y4604 = ~1'b0 ;
  assign y4605 = ~n20891 ;
  assign y4606 = n20892 ;
  assign y4607 = n20893 ;
  assign y4608 = ~n20895 ;
  assign y4609 = ~n20898 ;
  assign y4610 = ~n20899 ;
  assign y4611 = ~n20900 ;
  assign y4612 = n20903 ;
  assign y4613 = ~n20904 ;
  assign y4614 = ~1'b0 ;
  assign y4615 = ~n20905 ;
  assign y4616 = ~n20906 ;
  assign y4617 = ~n20907 ;
  assign y4618 = ~n20915 ;
  assign y4619 = n20921 ;
  assign y4620 = ~1'b0 ;
  assign y4621 = ~n20922 ;
  assign y4622 = n20925 ;
  assign y4623 = ~n20928 ;
  assign y4624 = ~n20933 ;
  assign y4625 = n20934 ;
  assign y4626 = ~n20937 ;
  assign y4627 = n20938 ;
  assign y4628 = n20940 ;
  assign y4629 = n20943 ;
  assign y4630 = ~1'b0 ;
  assign y4631 = n20944 ;
  assign y4632 = n20949 ;
  assign y4633 = ~n20954 ;
  assign y4634 = ~n20959 ;
  assign y4635 = ~n20961 ;
  assign y4636 = ~n20965 ;
  assign y4637 = ~n20966 ;
  assign y4638 = ~1'b0 ;
  assign y4639 = n20968 ;
  assign y4640 = n20972 ;
  assign y4641 = n20973 ;
  assign y4642 = n20974 ;
  assign y4643 = n20975 ;
  assign y4644 = n20976 ;
  assign y4645 = ~n20977 ;
  assign y4646 = n20978 ;
  assign y4647 = ~n20980 ;
  assign y4648 = ~n20985 ;
  assign y4649 = n20992 ;
  assign y4650 = ~n20993 ;
  assign y4651 = ~n20994 ;
  assign y4652 = ~n20995 ;
  assign y4653 = n20996 ;
  assign y4654 = n21001 ;
  assign y4655 = n21003 ;
  assign y4656 = ~n21005 ;
  assign y4657 = ~n21010 ;
  assign y4658 = ~n21012 ;
  assign y4659 = ~n21014 ;
  assign y4660 = n21020 ;
  assign y4661 = n21026 ;
  assign y4662 = n21027 ;
  assign y4663 = ~n21028 ;
  assign y4664 = ~n21030 ;
  assign y4665 = ~n21031 ;
  assign y4666 = ~n21033 ;
  assign y4667 = ~n21040 ;
  assign y4668 = n21042 ;
  assign y4669 = n21044 ;
  assign y4670 = n21047 ;
  assign y4671 = n21053 ;
  assign y4672 = ~n21056 ;
  assign y4673 = n21058 ;
  assign y4674 = ~n21060 ;
  assign y4675 = ~n21064 ;
  assign y4676 = n21069 ;
  assign y4677 = ~n21079 ;
  assign y4678 = ~n21084 ;
  assign y4679 = ~n21086 ;
  assign y4680 = n21090 ;
  assign y4681 = ~1'b0 ;
  assign y4682 = ~1'b0 ;
  assign y4683 = ~n21093 ;
  assign y4684 = n21094 ;
  assign y4685 = ~n21097 ;
  assign y4686 = ~n21099 ;
  assign y4687 = n21100 ;
  assign y4688 = ~n21101 ;
  assign y4689 = n21103 ;
  assign y4690 = ~1'b0 ;
  assign y4691 = ~n21104 ;
  assign y4692 = ~n21105 ;
  assign y4693 = ~n21107 ;
  assign y4694 = ~n21113 ;
  assign y4695 = ~n21114 ;
  assign y4696 = ~n21118 ;
  assign y4697 = n21121 ;
  assign y4698 = n21122 ;
  assign y4699 = ~n21125 ;
  assign y4700 = n21129 ;
  assign y4701 = ~n21132 ;
  assign y4702 = ~n21133 ;
  assign y4703 = n21134 ;
  assign y4704 = n21135 ;
  assign y4705 = ~n21136 ;
  assign y4706 = ~n21137 ;
  assign y4707 = n21138 ;
  assign y4708 = ~n21139 ;
  assign y4709 = n21140 ;
  assign y4710 = n21142 ;
  assign y4711 = ~1'b0 ;
  assign y4712 = n21144 ;
  assign y4713 = n21145 ;
  assign y4714 = ~n21150 ;
  assign y4715 = n21151 ;
  assign y4716 = n21153 ;
  assign y4717 = n21155 ;
  assign y4718 = ~n21159 ;
  assign y4719 = ~n21160 ;
  assign y4720 = ~n21166 ;
  assign y4721 = ~n21169 ;
  assign y4722 = n21174 ;
  assign y4723 = ~n21176 ;
  assign y4724 = ~n21178 ;
  assign y4725 = ~n21180 ;
  assign y4726 = ~n21181 ;
  assign y4727 = n21187 ;
  assign y4728 = ~n21189 ;
  assign y4729 = ~n21192 ;
  assign y4730 = ~n21195 ;
  assign y4731 = n21198 ;
  assign y4732 = ~n21203 ;
  assign y4733 = ~n21212 ;
  assign y4734 = n21217 ;
  assign y4735 = n21220 ;
  assign y4736 = n21223 ;
  assign y4737 = n21226 ;
  assign y4738 = n21230 ;
  assign y4739 = ~n21233 ;
  assign y4740 = ~n21234 ;
  assign y4741 = n21236 ;
  assign y4742 = n21238 ;
  assign y4743 = ~n21240 ;
  assign y4744 = ~n21242 ;
  assign y4745 = ~1'b0 ;
  assign y4746 = ~n21243 ;
  assign y4747 = ~n21247 ;
  assign y4748 = ~n21250 ;
  assign y4749 = ~n21266 ;
  assign y4750 = ~n21267 ;
  assign y4751 = ~n21275 ;
  assign y4752 = ~n21277 ;
  assign y4753 = n21278 ;
  assign y4754 = n21281 ;
  assign y4755 = ~n21283 ;
  assign y4756 = ~n21285 ;
  assign y4757 = ~n21286 ;
  assign y4758 = ~n21290 ;
  assign y4759 = ~1'b0 ;
  assign y4760 = n21293 ;
  assign y4761 = ~n21294 ;
  assign y4762 = n21295 ;
  assign y4763 = ~n21300 ;
  assign y4764 = n21301 ;
  assign y4765 = ~n21302 ;
  assign y4766 = n21305 ;
  assign y4767 = ~n21308 ;
  assign y4768 = n21311 ;
  assign y4769 = n21318 ;
  assign y4770 = ~n21321 ;
  assign y4771 = ~n21325 ;
  assign y4772 = n21329 ;
  assign y4773 = n21331 ;
  assign y4774 = ~n21335 ;
  assign y4775 = n21336 ;
  assign y4776 = ~n21344 ;
  assign y4777 = ~n21350 ;
  assign y4778 = ~n21353 ;
  assign y4779 = ~n21357 ;
  assign y4780 = ~n21359 ;
  assign y4781 = n21365 ;
  assign y4782 = ~n21366 ;
  assign y4783 = ~n21370 ;
  assign y4784 = ~n21375 ;
  assign y4785 = ~n21377 ;
  assign y4786 = ~n21379 ;
  assign y4787 = n21383 ;
  assign y4788 = ~n21385 ;
  assign y4789 = ~n21394 ;
  assign y4790 = n21397 ;
  assign y4791 = ~n21399 ;
  assign y4792 = n21402 ;
  assign y4793 = ~n21410 ;
  assign y4794 = n21412 ;
  assign y4795 = ~n21413 ;
  assign y4796 = ~1'b0 ;
  assign y4797 = n21416 ;
  assign y4798 = n21418 ;
  assign y4799 = ~n21419 ;
  assign y4800 = n21421 ;
  assign y4801 = n21427 ;
  assign y4802 = ~n21429 ;
  assign y4803 = ~n21433 ;
  assign y4804 = ~n21439 ;
  assign y4805 = ~n21441 ;
  assign y4806 = n21443 ;
  assign y4807 = ~n21444 ;
  assign y4808 = n21448 ;
  assign y4809 = ~n21449 ;
  assign y4810 = n21453 ;
  assign y4811 = n21459 ;
  assign y4812 = ~n21463 ;
  assign y4813 = n21465 ;
  assign y4814 = n21466 ;
  assign y4815 = ~n21467 ;
  assign y4816 = n21469 ;
  assign y4817 = ~1'b0 ;
  assign y4818 = n21471 ;
  assign y4819 = n21485 ;
  assign y4820 = ~n21488 ;
  assign y4821 = ~n21490 ;
  assign y4822 = ~1'b0 ;
  assign y4823 = ~n21495 ;
  assign y4824 = ~n21496 ;
  assign y4825 = ~n21498 ;
  assign y4826 = n21504 ;
  assign y4827 = n21510 ;
  assign y4828 = ~n21511 ;
  assign y4829 = ~n21515 ;
  assign y4830 = ~1'b0 ;
  assign y4831 = ~n21520 ;
  assign y4832 = ~n21521 ;
  assign y4833 = ~n21523 ;
  assign y4834 = n21528 ;
  assign y4835 = ~n21529 ;
  assign y4836 = n21531 ;
  assign y4837 = n21537 ;
  assign y4838 = ~n21542 ;
  assign y4839 = n21547 ;
  assign y4840 = n21551 ;
  assign y4841 = n21559 ;
  assign y4842 = ~n21562 ;
  assign y4843 = n21564 ;
  assign y4844 = n21566 ;
  assign y4845 = n21568 ;
  assign y4846 = ~n21569 ;
  assign y4847 = n21572 ;
  assign y4848 = n21579 ;
  assign y4849 = n21583 ;
  assign y4850 = ~1'b0 ;
  assign y4851 = ~n21584 ;
  assign y4852 = ~n21591 ;
  assign y4853 = n21593 ;
  assign y4854 = n21595 ;
  assign y4855 = n21599 ;
  assign y4856 = ~1'b0 ;
  assign y4857 = n21603 ;
  assign y4858 = n21604 ;
  assign y4859 = n21605 ;
  assign y4860 = ~n21608 ;
  assign y4861 = n21610 ;
  assign y4862 = n21612 ;
  assign y4863 = ~n21613 ;
  assign y4864 = n21616 ;
  assign y4865 = ~n21618 ;
  assign y4866 = ~n21619 ;
  assign y4867 = ~n21620 ;
  assign y4868 = n21623 ;
  assign y4869 = ~n21624 ;
  assign y4870 = ~n21626 ;
  assign y4871 = n21627 ;
  assign y4872 = n21628 ;
  assign y4873 = n21632 ;
  assign y4874 = n21633 ;
  assign y4875 = ~n21635 ;
  assign y4876 = n21637 ;
  assign y4877 = n21639 ;
  assign y4878 = n21642 ;
  assign y4879 = ~n21643 ;
  assign y4880 = n21644 ;
  assign y4881 = n21645 ;
  assign y4882 = n21647 ;
  assign y4883 = n21651 ;
  assign y4884 = ~n21654 ;
  assign y4885 = n21657 ;
  assign y4886 = n21660 ;
  assign y4887 = ~n21666 ;
  assign y4888 = n21667 ;
  assign y4889 = ~n21669 ;
  assign y4890 = ~1'b0 ;
  assign y4891 = n21670 ;
  assign y4892 = ~n21672 ;
  assign y4893 = n21675 ;
  assign y4894 = n21676 ;
  assign y4895 = ~n21678 ;
  assign y4896 = ~n21681 ;
  assign y4897 = ~n21683 ;
  assign y4898 = n21684 ;
  assign y4899 = n21685 ;
  assign y4900 = ~n21687 ;
  assign y4901 = n21688 ;
  assign y4902 = n21690 ;
  assign y4903 = n21691 ;
  assign y4904 = ~n21692 ;
  assign y4905 = ~n21694 ;
  assign y4906 = n21697 ;
  assign y4907 = ~n21700 ;
  assign y4908 = ~n21706 ;
  assign y4909 = ~n21709 ;
  assign y4910 = ~n21713 ;
  assign y4911 = ~n21714 ;
  assign y4912 = n21718 ;
  assign y4913 = ~n21723 ;
  assign y4914 = n21725 ;
  assign y4915 = n21729 ;
  assign y4916 = ~n21732 ;
  assign y4917 = ~n21734 ;
  assign y4918 = ~n21737 ;
  assign y4919 = n21741 ;
  assign y4920 = ~1'b0 ;
  assign y4921 = ~1'b0 ;
  assign y4922 = n21745 ;
  assign y4923 = ~n21747 ;
  assign y4924 = ~n21750 ;
  assign y4925 = ~1'b0 ;
  assign y4926 = ~n21751 ;
  assign y4927 = n21755 ;
  assign y4928 = n21757 ;
  assign y4929 = ~n21767 ;
  assign y4930 = n21773 ;
  assign y4931 = ~n21777 ;
  assign y4932 = ~n21778 ;
  assign y4933 = ~n21779 ;
  assign y4934 = n21783 ;
  assign y4935 = n21794 ;
  assign y4936 = ~1'b0 ;
  assign y4937 = n21796 ;
  assign y4938 = n21799 ;
  assign y4939 = n21800 ;
  assign y4940 = ~n21801 ;
  assign y4941 = ~n21808 ;
  assign y4942 = n21811 ;
  assign y4943 = ~n21814 ;
  assign y4944 = n21815 ;
  assign y4945 = n21818 ;
  assign y4946 = n21822 ;
  assign y4947 = n21823 ;
  assign y4948 = ~n21824 ;
  assign y4949 = n21826 ;
  assign y4950 = n21829 ;
  assign y4951 = n21834 ;
  assign y4952 = ~n21839 ;
  assign y4953 = ~n21842 ;
  assign y4954 = ~n21847 ;
  assign y4955 = ~n21852 ;
  assign y4956 = ~n21857 ;
  assign y4957 = ~n21858 ;
  assign y4958 = n21859 ;
  assign y4959 = n21860 ;
  assign y4960 = n21865 ;
  assign y4961 = ~1'b0 ;
  assign y4962 = ~n21866 ;
  assign y4963 = n21867 ;
  assign y4964 = n21868 ;
  assign y4965 = ~n21869 ;
  assign y4966 = n21872 ;
  assign y4967 = ~n21873 ;
  assign y4968 = n21874 ;
  assign y4969 = ~1'b0 ;
  assign y4970 = ~n21876 ;
  assign y4971 = ~n21879 ;
  assign y4972 = n21880 ;
  assign y4973 = n155 ;
  assign y4974 = ~n21883 ;
  assign y4975 = n21885 ;
  assign y4976 = n21887 ;
  assign y4977 = ~n21890 ;
  assign y4978 = ~n21892 ;
  assign y4979 = ~n21896 ;
  assign y4980 = ~n21902 ;
  assign y4981 = ~n21905 ;
  assign y4982 = ~n21906 ;
  assign y4983 = ~n21913 ;
  assign y4984 = n21918 ;
  assign y4985 = n21920 ;
  assign y4986 = ~n21921 ;
  assign y4987 = ~n21930 ;
  assign y4988 = n21931 ;
  assign y4989 = n21932 ;
  assign y4990 = ~n21936 ;
  assign y4991 = n21938 ;
  assign y4992 = n21941 ;
  assign y4993 = ~n21942 ;
  assign y4994 = n21943 ;
  assign y4995 = n21946 ;
  assign y4996 = ~n21953 ;
  assign y4997 = n21962 ;
  assign y4998 = n21967 ;
  assign y4999 = ~n21971 ;
  assign y5000 = ~n21972 ;
  assign y5001 = ~n21975 ;
  assign y5002 = ~n21981 ;
  assign y5003 = ~n21983 ;
  assign y5004 = ~n21989 ;
  assign y5005 = ~n21990 ;
  assign y5006 = ~n21993 ;
  assign y5007 = n21994 ;
  assign y5008 = n21995 ;
  assign y5009 = n21996 ;
  assign y5010 = ~n21997 ;
  assign y5011 = n21999 ;
  assign y5012 = ~n22000 ;
  assign y5013 = ~1'b0 ;
  assign y5014 = n22007 ;
  assign y5015 = ~n22008 ;
  assign y5016 = ~n22012 ;
  assign y5017 = n22015 ;
  assign y5018 = ~1'b0 ;
  assign y5019 = ~n22019 ;
  assign y5020 = n22020 ;
  assign y5021 = ~n22021 ;
  assign y5022 = n22025 ;
  assign y5023 = ~n22027 ;
  assign y5024 = ~n22028 ;
  assign y5025 = n22029 ;
  assign y5026 = ~1'b0 ;
  assign y5027 = ~n22034 ;
  assign y5028 = n22036 ;
  assign y5029 = n22038 ;
  assign y5030 = n22039 ;
  assign y5031 = n14243 ;
  assign y5032 = ~n22044 ;
  assign y5033 = ~n22045 ;
  assign y5034 = n22051 ;
  assign y5035 = ~n22055 ;
  assign y5036 = n22056 ;
  assign y5037 = n22057 ;
  assign y5038 = n22073 ;
  assign y5039 = ~n22075 ;
  assign y5040 = n22076 ;
  assign y5041 = ~n22077 ;
  assign y5042 = n22079 ;
  assign y5043 = n22080 ;
  assign y5044 = n22084 ;
  assign y5045 = ~n22090 ;
  assign y5046 = ~n22091 ;
  assign y5047 = ~n22092 ;
  assign y5048 = n22095 ;
  assign y5049 = ~n22097 ;
  assign y5050 = ~n22098 ;
  assign y5051 = ~1'b0 ;
  assign y5052 = ~n22102 ;
  assign y5053 = n22111 ;
  assign y5054 = ~n22112 ;
  assign y5055 = ~n22114 ;
  assign y5056 = ~n22119 ;
  assign y5057 = ~n22120 ;
  assign y5058 = n22122 ;
  assign y5059 = ~1'b0 ;
  assign y5060 = ~n22125 ;
  assign y5061 = ~n22127 ;
  assign y5062 = n22129 ;
  assign y5063 = ~n22132 ;
  assign y5064 = ~1'b0 ;
  assign y5065 = n22133 ;
  assign y5066 = ~n22134 ;
  assign y5067 = ~n22135 ;
  assign y5068 = ~n22142 ;
  assign y5069 = ~n22149 ;
  assign y5070 = n22153 ;
  assign y5071 = ~n22161 ;
  assign y5072 = n22163 ;
  assign y5073 = n22166 ;
  assign y5074 = ~n22168 ;
  assign y5075 = n22172 ;
  assign y5076 = ~n22173 ;
  assign y5077 = n22175 ;
  assign y5078 = n22186 ;
  assign y5079 = ~1'b0 ;
  assign y5080 = n22187 ;
  assign y5081 = ~n22191 ;
  assign y5082 = n22198 ;
  assign y5083 = n22199 ;
  assign y5084 = ~n22200 ;
  assign y5085 = n22202 ;
  assign y5086 = n22204 ;
  assign y5087 = ~n22205 ;
  assign y5088 = ~n22209 ;
  assign y5089 = ~n22212 ;
  assign y5090 = ~n22223 ;
  assign y5091 = ~n22225 ;
  assign y5092 = ~n22229 ;
  assign y5093 = ~n22230 ;
  assign y5094 = n22231 ;
  assign y5095 = ~n22234 ;
  assign y5096 = ~n22235 ;
  assign y5097 = n22237 ;
  assign y5098 = n22242 ;
  assign y5099 = ~n22243 ;
  assign y5100 = n22245 ;
  assign y5101 = n22246 ;
  assign y5102 = n22247 ;
  assign y5103 = n22252 ;
  assign y5104 = n22254 ;
  assign y5105 = n22255 ;
  assign y5106 = ~n22257 ;
  assign y5107 = ~n22260 ;
  assign y5108 = ~n22264 ;
  assign y5109 = ~n22266 ;
  assign y5110 = ~n22273 ;
  assign y5111 = n22275 ;
  assign y5112 = ~n22281 ;
  assign y5113 = n22284 ;
  assign y5114 = ~1'b0 ;
  assign y5115 = n22286 ;
  assign y5116 = ~n22288 ;
  assign y5117 = n22291 ;
  assign y5118 = ~n22292 ;
  assign y5119 = n22294 ;
  assign y5120 = ~n22295 ;
  assign y5121 = n22298 ;
  assign y5122 = n22299 ;
  assign y5123 = n22301 ;
  assign y5124 = ~n22302 ;
  assign y5125 = ~n22303 ;
  assign y5126 = n22304 ;
  assign y5127 = ~n22306 ;
  assign y5128 = ~1'b0 ;
  assign y5129 = ~n22307 ;
  assign y5130 = n22309 ;
  assign y5131 = ~n22310 ;
  assign y5132 = ~n22313 ;
  assign y5133 = ~n22314 ;
  assign y5134 = ~n22317 ;
  assign y5135 = ~n22318 ;
  assign y5136 = ~n22321 ;
  assign y5137 = ~n22323 ;
  assign y5138 = n22325 ;
  assign y5139 = n22326 ;
  assign y5140 = n22327 ;
  assign y5141 = n22328 ;
  assign y5142 = ~n22331 ;
  assign y5143 = ~n22333 ;
  assign y5144 = n22336 ;
  assign y5145 = n22337 ;
  assign y5146 = n22339 ;
  assign y5147 = ~n22341 ;
  assign y5148 = ~n22351 ;
  assign y5149 = ~n22356 ;
  assign y5150 = n22357 ;
  assign y5151 = ~n22363 ;
  assign y5152 = ~n22367 ;
  assign y5153 = n22372 ;
  assign y5154 = ~1'b0 ;
  assign y5155 = ~n22374 ;
  assign y5156 = n22380 ;
  assign y5157 = ~n22387 ;
  assign y5158 = n22388 ;
  assign y5159 = n22389 ;
  assign y5160 = n22390 ;
  assign y5161 = n22392 ;
  assign y5162 = ~1'b0 ;
  assign y5163 = ~n22393 ;
  assign y5164 = n22396 ;
  assign y5165 = n22404 ;
  assign y5166 = ~n22406 ;
  assign y5167 = ~n22407 ;
  assign y5168 = n22411 ;
  assign y5169 = ~n22412 ;
  assign y5170 = n22416 ;
  assign y5171 = n22417 ;
  assign y5172 = n22419 ;
  assign y5173 = ~n22425 ;
  assign y5174 = ~n22429 ;
  assign y5175 = ~n22433 ;
  assign y5176 = n22435 ;
  assign y5177 = ~n22440 ;
  assign y5178 = ~n22442 ;
  assign y5179 = n22445 ;
  assign y5180 = ~n22449 ;
  assign y5181 = ~n22450 ;
  assign y5182 = ~n22462 ;
  assign y5183 = n22465 ;
  assign y5184 = ~n22468 ;
  assign y5185 = ~n22469 ;
  assign y5186 = ~1'b0 ;
  assign y5187 = n22475 ;
  assign y5188 = n22476 ;
  assign y5189 = ~n22481 ;
  assign y5190 = n22482 ;
  assign y5191 = n22483 ;
  assign y5192 = n22485 ;
  assign y5193 = ~n22487 ;
  assign y5194 = ~1'b0 ;
  assign y5195 = n22488 ;
  assign y5196 = ~n22490 ;
  assign y5197 = n22492 ;
  assign y5198 = ~n22494 ;
  assign y5199 = ~n22495 ;
  assign y5200 = ~n22498 ;
  assign y5201 = n22499 ;
  assign y5202 = n22501 ;
  assign y5203 = ~n22503 ;
  assign y5204 = ~n22505 ;
  assign y5205 = ~n22506 ;
  assign y5206 = n22510 ;
  assign y5207 = ~n22513 ;
  assign y5208 = n22514 ;
  assign y5209 = n22515 ;
  assign y5210 = ~n22519 ;
  assign y5211 = n22522 ;
  assign y5212 = n22525 ;
  assign y5213 = ~n22531 ;
  assign y5214 = ~n22532 ;
  assign y5215 = n22537 ;
  assign y5216 = ~n22540 ;
  assign y5217 = n22542 ;
  assign y5218 = n22543 ;
  assign y5219 = ~n22544 ;
  assign y5220 = ~n22549 ;
  assign y5221 = n22551 ;
  assign y5222 = n22553 ;
  assign y5223 = ~n22554 ;
  assign y5224 = n22559 ;
  assign y5225 = n22563 ;
  assign y5226 = ~n22566 ;
  assign y5227 = n22574 ;
  assign y5228 = n22579 ;
  assign y5229 = n22584 ;
  assign y5230 = ~n22587 ;
  assign y5231 = ~n22588 ;
  assign y5232 = ~n22593 ;
  assign y5233 = ~n22595 ;
  assign y5234 = n22601 ;
  assign y5235 = ~n22606 ;
  assign y5236 = ~1'b0 ;
  assign y5237 = n22607 ;
  assign y5238 = n22614 ;
  assign y5239 = n22615 ;
  assign y5240 = n22618 ;
  assign y5241 = n22628 ;
  assign y5242 = n22630 ;
  assign y5243 = n22634 ;
  assign y5244 = ~n22637 ;
  assign y5245 = ~n22638 ;
  assign y5246 = ~n22639 ;
  assign y5247 = n22647 ;
  assign y5248 = n22648 ;
  assign y5249 = ~n22651 ;
  assign y5250 = n22655 ;
  assign y5251 = n22656 ;
  assign y5252 = ~n22660 ;
  assign y5253 = ~n22662 ;
  assign y5254 = n22665 ;
  assign y5255 = n22671 ;
  assign y5256 = n22672 ;
  assign y5257 = n22674 ;
  assign y5258 = n22678 ;
  assign y5259 = n22684 ;
  assign y5260 = n22687 ;
  assign y5261 = ~n22692 ;
  assign y5262 = n22695 ;
  assign y5263 = n22700 ;
  assign y5264 = n22702 ;
  assign y5265 = n22705 ;
  assign y5266 = ~n22709 ;
  assign y5267 = n22712 ;
  assign y5268 = ~n22714 ;
  assign y5269 = ~n22716 ;
  assign y5270 = ~n22717 ;
  assign y5271 = n22722 ;
  assign y5272 = ~n22727 ;
  assign y5273 = n22734 ;
  assign y5274 = ~n22739 ;
  assign y5275 = n22742 ;
  assign y5276 = ~n22743 ;
  assign y5277 = n22745 ;
  assign y5278 = n22746 ;
  assign y5279 = ~n22749 ;
  assign y5280 = ~n22751 ;
  assign y5281 = ~n22753 ;
  assign y5282 = n22754 ;
  assign y5283 = n22763 ;
  assign y5284 = ~n22765 ;
  assign y5285 = ~n22767 ;
  assign y5286 = ~n22770 ;
  assign y5287 = ~1'b0 ;
  assign y5288 = ~n22771 ;
  assign y5289 = n22776 ;
  assign y5290 = ~n22778 ;
  assign y5291 = ~n22779 ;
  assign y5292 = ~1'b0 ;
  assign y5293 = ~n22784 ;
  assign y5294 = ~n22787 ;
  assign y5295 = ~n22792 ;
  assign y5296 = ~n22793 ;
  assign y5297 = n22795 ;
  assign y5298 = ~n22797 ;
  assign y5299 = ~n22800 ;
  assign y5300 = ~n22802 ;
  assign y5301 = ~n22810 ;
  assign y5302 = ~1'b0 ;
  assign y5303 = n22814 ;
  assign y5304 = ~n22817 ;
  assign y5305 = n22821 ;
  assign y5306 = ~1'b0 ;
  assign y5307 = ~1'b0 ;
  assign y5308 = ~n22828 ;
  assign y5309 = n22830 ;
  assign y5310 = n22832 ;
  assign y5311 = ~n22838 ;
  assign y5312 = ~n22842 ;
  assign y5313 = n22846 ;
  assign y5314 = ~n22852 ;
  assign y5315 = n22855 ;
  assign y5316 = ~n22856 ;
  assign y5317 = n22857 ;
  assign y5318 = ~n22860 ;
  assign y5319 = ~n22865 ;
  assign y5320 = ~n22866 ;
  assign y5321 = ~n22870 ;
  assign y5322 = ~n22874 ;
  assign y5323 = ~1'b0 ;
  assign y5324 = n22876 ;
  assign y5325 = ~n22877 ;
  assign y5326 = ~n22878 ;
  assign y5327 = ~n22879 ;
  assign y5328 = ~n22882 ;
  assign y5329 = n22883 ;
  assign y5330 = ~n22896 ;
  assign y5331 = ~n22898 ;
  assign y5332 = ~n22901 ;
  assign y5333 = n22904 ;
  assign y5334 = ~n22908 ;
  assign y5335 = n22910 ;
  assign y5336 = ~n22913 ;
  assign y5337 = ~n22916 ;
  assign y5338 = ~n22919 ;
  assign y5339 = n22920 ;
  assign y5340 = n22923 ;
  assign y5341 = n22926 ;
  assign y5342 = n22927 ;
  assign y5343 = ~n22930 ;
  assign y5344 = ~n22935 ;
  assign y5345 = n22936 ;
  assign y5346 = ~n22937 ;
  assign y5347 = ~n22938 ;
  assign y5348 = n22940 ;
  assign y5349 = n22942 ;
  assign y5350 = n22946 ;
  assign y5351 = n22948 ;
  assign y5352 = n22949 ;
  assign y5353 = n22950 ;
  assign y5354 = n22953 ;
  assign y5355 = ~n22961 ;
  assign y5356 = ~n22966 ;
  assign y5357 = n22969 ;
  assign y5358 = n22970 ;
  assign y5359 = n22972 ;
  assign y5360 = n22974 ;
  assign y5361 = n22975 ;
  assign y5362 = ~n22976 ;
  assign y5363 = ~n22977 ;
  assign y5364 = ~n22978 ;
  assign y5365 = ~n22980 ;
  assign y5366 = n22984 ;
  assign y5367 = n22985 ;
  assign y5368 = ~n22986 ;
  assign y5369 = ~n22989 ;
  assign y5370 = n22990 ;
  assign y5371 = ~n22992 ;
  assign y5372 = ~n23000 ;
  assign y5373 = ~n23001 ;
  assign y5374 = ~n23006 ;
  assign y5375 = ~n23009 ;
  assign y5376 = ~n23014 ;
  assign y5377 = n23016 ;
  assign y5378 = ~n23017 ;
  assign y5379 = ~n23018 ;
  assign y5380 = ~n23019 ;
  assign y5381 = ~n23021 ;
  assign y5382 = n23027 ;
  assign y5383 = n23031 ;
  assign y5384 = ~n23032 ;
  assign y5385 = ~n23042 ;
  assign y5386 = ~n23044 ;
  assign y5387 = ~n23049 ;
  assign y5388 = ~n23050 ;
  assign y5389 = ~n23051 ;
  assign y5390 = ~1'b0 ;
  assign y5391 = ~n23052 ;
  assign y5392 = ~n23053 ;
  assign y5393 = n23058 ;
  assign y5394 = ~n23061 ;
  assign y5395 = ~n23062 ;
  assign y5396 = ~n23067 ;
  assign y5397 = n23068 ;
  assign y5398 = ~n23073 ;
  assign y5399 = n23080 ;
  assign y5400 = n23086 ;
  assign y5401 = ~n23088 ;
  assign y5402 = ~n23092 ;
  assign y5403 = ~n23093 ;
  assign y5404 = ~n23096 ;
  assign y5405 = n23098 ;
  assign y5406 = ~n23099 ;
  assign y5407 = ~n23102 ;
  assign y5408 = ~n23103 ;
  assign y5409 = n23107 ;
  assign y5410 = n23115 ;
  assign y5411 = ~n23116 ;
  assign y5412 = ~n23122 ;
  assign y5413 = n23124 ;
  assign y5414 = n23125 ;
  assign y5415 = n23126 ;
  assign y5416 = n23127 ;
  assign y5417 = n23132 ;
  assign y5418 = ~n23133 ;
  assign y5419 = n23135 ;
  assign y5420 = n23136 ;
  assign y5421 = ~n23138 ;
  assign y5422 = n23139 ;
  assign y5423 = n23140 ;
  assign y5424 = ~n23146 ;
  assign y5425 = n23148 ;
  assign y5426 = n23151 ;
  assign y5427 = ~n23155 ;
  assign y5428 = ~n23156 ;
  assign y5429 = ~n23157 ;
  assign y5430 = ~n23159 ;
  assign y5431 = ~n23162 ;
  assign y5432 = ~n23163 ;
  assign y5433 = ~n23167 ;
  assign y5434 = ~1'b0 ;
  assign y5435 = n23168 ;
  assign y5436 = n23170 ;
  assign y5437 = ~n23173 ;
  assign y5438 = n23177 ;
  assign y5439 = n23178 ;
  assign y5440 = ~n23179 ;
  assign y5441 = ~n23180 ;
  assign y5442 = n23181 ;
  assign y5443 = ~n23183 ;
  assign y5444 = ~n23186 ;
  assign y5445 = n23191 ;
  assign y5446 = ~n23194 ;
  assign y5447 = n23196 ;
  assign y5448 = ~n23199 ;
  assign y5449 = ~n23206 ;
  assign y5450 = n23208 ;
  assign y5451 = n23211 ;
  assign y5452 = ~n23215 ;
  assign y5453 = n23216 ;
  assign y5454 = ~n23219 ;
  assign y5455 = n23221 ;
  assign y5456 = ~1'b0 ;
  assign y5457 = ~n23224 ;
  assign y5458 = n23225 ;
  assign y5459 = ~n23231 ;
  assign y5460 = ~n23232 ;
  assign y5461 = n23234 ;
  assign y5462 = n23236 ;
  assign y5463 = ~n23237 ;
  assign y5464 = ~n23238 ;
  assign y5465 = ~n23239 ;
  assign y5466 = n23242 ;
  assign y5467 = ~n23243 ;
  assign y5468 = n23244 ;
  assign y5469 = n23246 ;
  assign y5470 = n23250 ;
  assign y5471 = ~n23252 ;
  assign y5472 = n23254 ;
  assign y5473 = n23258 ;
  assign y5474 = ~n23265 ;
  assign y5475 = ~n23266 ;
  assign y5476 = ~n23267 ;
  assign y5477 = n23271 ;
  assign y5478 = ~n23272 ;
  assign y5479 = n23276 ;
  assign y5480 = n23279 ;
  assign y5481 = ~n23284 ;
  assign y5482 = ~n23285 ;
  assign y5483 = ~1'b0 ;
  assign y5484 = n23295 ;
  assign y5485 = n23297 ;
  assign y5486 = n23303 ;
  assign y5487 = ~n23307 ;
  assign y5488 = n23309 ;
  assign y5489 = ~n23313 ;
  assign y5490 = ~n23314 ;
  assign y5491 = n23315 ;
  assign y5492 = ~n23317 ;
  assign y5493 = n23319 ;
  assign y5494 = n23320 ;
  assign y5495 = n23321 ;
  assign y5496 = n23323 ;
  assign y5497 = ~n23325 ;
  assign y5498 = ~n23329 ;
  assign y5499 = ~1'b0 ;
  assign y5500 = ~n23333 ;
  assign y5501 = ~n23337 ;
  assign y5502 = n23345 ;
  assign y5503 = ~n23347 ;
  assign y5504 = ~n23350 ;
  assign y5505 = n23354 ;
  assign y5506 = n23355 ;
  assign y5507 = ~n23360 ;
  assign y5508 = ~n23363 ;
  assign y5509 = n23365 ;
  assign y5510 = ~n23370 ;
  assign y5511 = n23371 ;
  assign y5512 = ~n23374 ;
  assign y5513 = n23377 ;
  assign y5514 = n23379 ;
  assign y5515 = ~n23381 ;
  assign y5516 = n23383 ;
  assign y5517 = ~n23385 ;
  assign y5518 = n23387 ;
  assign y5519 = n23388 ;
  assign y5520 = n23391 ;
  assign y5521 = n23393 ;
  assign y5522 = ~n23396 ;
  assign y5523 = ~n23398 ;
  assign y5524 = ~n23400 ;
  assign y5525 = ~n23403 ;
  assign y5526 = ~n23405 ;
  assign y5527 = n23409 ;
  assign y5528 = ~n23410 ;
  assign y5529 = ~n23412 ;
  assign y5530 = ~n23414 ;
  assign y5531 = n23417 ;
  assign y5532 = n23418 ;
  assign y5533 = ~n23420 ;
  assign y5534 = ~n23427 ;
  assign y5535 = n23429 ;
  assign y5536 = n23435 ;
  assign y5537 = ~n23438 ;
  assign y5538 = ~n23441 ;
  assign y5539 = ~1'b0 ;
  assign y5540 = n23442 ;
  assign y5541 = ~n23445 ;
  assign y5542 = n23447 ;
  assign y5543 = ~n23453 ;
  assign y5544 = n23454 ;
  assign y5545 = n23459 ;
  assign y5546 = n23461 ;
  assign y5547 = n23463 ;
  assign y5548 = ~n23465 ;
  assign y5549 = n23470 ;
  assign y5550 = ~n23477 ;
  assign y5551 = ~n23480 ;
  assign y5552 = n23483 ;
  assign y5553 = n23485 ;
  assign y5554 = n23487 ;
  assign y5555 = ~n23488 ;
  assign y5556 = n23492 ;
  assign y5557 = n23493 ;
  assign y5558 = n23494 ;
  assign y5559 = n23495 ;
  assign y5560 = ~n23496 ;
  assign y5561 = n23498 ;
  assign y5562 = ~n23503 ;
  assign y5563 = ~n23505 ;
  assign y5564 = n23508 ;
  assign y5565 = ~n23509 ;
  assign y5566 = n23510 ;
  assign y5567 = n23516 ;
  assign y5568 = n23518 ;
  assign y5569 = ~n23523 ;
  assign y5570 = n23524 ;
  assign y5571 = ~n23525 ;
  assign y5572 = n23530 ;
  assign y5573 = n23536 ;
  assign y5574 = n23540 ;
  assign y5575 = ~n23542 ;
  assign y5576 = ~1'b0 ;
  assign y5577 = ~n23544 ;
  assign y5578 = ~n23546 ;
  assign y5579 = ~n23548 ;
  assign y5580 = n23551 ;
  assign y5581 = ~1'b0 ;
  assign y5582 = ~n23552 ;
  assign y5583 = n23556 ;
  assign y5584 = n23559 ;
  assign y5585 = n23566 ;
  assign y5586 = ~n23574 ;
  assign y5587 = ~n23575 ;
  assign y5588 = ~n23578 ;
  assign y5589 = ~n23582 ;
  assign y5590 = n23583 ;
  assign y5591 = n23588 ;
  assign y5592 = n23590 ;
  assign y5593 = n23591 ;
  assign y5594 = ~n23595 ;
  assign y5595 = ~n23601 ;
  assign y5596 = ~n23602 ;
  assign y5597 = ~n23606 ;
  assign y5598 = n23607 ;
  assign y5599 = n23614 ;
  assign y5600 = ~n23616 ;
  assign y5601 = ~1'b0 ;
  assign y5602 = n23619 ;
  assign y5603 = ~n23623 ;
  assign y5604 = n23629 ;
  assign y5605 = ~n23631 ;
  assign y5606 = n23636 ;
  assign y5607 = n23637 ;
  assign y5608 = ~n23639 ;
  assign y5609 = n23640 ;
  assign y5610 = n23644 ;
  assign y5611 = ~n23647 ;
  assign y5612 = n23649 ;
  assign y5613 = ~n23650 ;
  assign y5614 = n23652 ;
  assign y5615 = ~n23655 ;
  assign y5616 = ~n23661 ;
  assign y5617 = ~n23664 ;
  assign y5618 = ~n23666 ;
  assign y5619 = n23671 ;
  assign y5620 = ~n23673 ;
  assign y5621 = n23674 ;
  assign y5622 = ~n23676 ;
  assign y5623 = ~n23678 ;
  assign y5624 = n23679 ;
  assign y5625 = ~n9195 ;
  assign y5626 = ~n23680 ;
  assign y5627 = ~n23683 ;
  assign y5628 = n23685 ;
  assign y5629 = ~n23688 ;
  assign y5630 = ~n23690 ;
  assign y5631 = ~n23692 ;
  assign y5632 = n23694 ;
  assign y5633 = n23695 ;
  assign y5634 = n23699 ;
  assign y5635 = ~n23700 ;
  assign y5636 = n23702 ;
  assign y5637 = ~n23705 ;
  assign y5638 = ~n23707 ;
  assign y5639 = ~n23719 ;
  assign y5640 = ~n23720 ;
  assign y5641 = n23721 ;
  assign y5642 = ~n23722 ;
  assign y5643 = ~n23723 ;
  assign y5644 = ~n23725 ;
  assign y5645 = n23726 ;
  assign y5646 = ~n23733 ;
  assign y5647 = ~n23735 ;
  assign y5648 = n23739 ;
  assign y5649 = n23742 ;
  assign y5650 = ~n23744 ;
  assign y5651 = n23749 ;
  assign y5652 = ~n23751 ;
  assign y5653 = ~n23753 ;
  assign y5654 = ~n23757 ;
  assign y5655 = ~n23758 ;
  assign y5656 = n23760 ;
  assign y5657 = n23761 ;
  assign y5658 = n23765 ;
  assign y5659 = ~1'b0 ;
  assign y5660 = n23768 ;
  assign y5661 = ~n23771 ;
  assign y5662 = ~n23774 ;
  assign y5663 = n23775 ;
  assign y5664 = n23777 ;
  assign y5665 = ~n23778 ;
  assign y5666 = n23779 ;
  assign y5667 = n23782 ;
  assign y5668 = n16263 ;
  assign y5669 = ~n23783 ;
  assign y5670 = ~n23784 ;
  assign y5671 = ~n23786 ;
  assign y5672 = ~n23788 ;
  assign y5673 = ~n23790 ;
  assign y5674 = ~n23792 ;
  assign y5675 = ~n23798 ;
  assign y5676 = ~n23802 ;
  assign y5677 = ~n23807 ;
  assign y5678 = ~n23812 ;
  assign y5679 = n23815 ;
  assign y5680 = ~n23818 ;
  assign y5681 = ~n23819 ;
  assign y5682 = ~1'b0 ;
  assign y5683 = ~n23820 ;
  assign y5684 = ~n23826 ;
  assign y5685 = ~n23827 ;
  assign y5686 = n23829 ;
  assign y5687 = ~n23832 ;
  assign y5688 = ~1'b0 ;
  assign y5689 = ~n23835 ;
  assign y5690 = ~n23836 ;
  assign y5691 = ~n23837 ;
  assign y5692 = n23838 ;
  assign y5693 = ~n23841 ;
  assign y5694 = ~1'b0 ;
  assign y5695 = ~n23844 ;
  assign y5696 = ~n23845 ;
  assign y5697 = ~n23851 ;
  assign y5698 = ~n23855 ;
  assign y5699 = ~n23857 ;
  assign y5700 = n23858 ;
  assign y5701 = ~n23863 ;
  assign y5702 = ~1'b0 ;
  assign y5703 = n23864 ;
  assign y5704 = ~n23865 ;
  assign y5705 = ~n23866 ;
  assign y5706 = ~n23871 ;
  assign y5707 = ~n23872 ;
  assign y5708 = ~n23873 ;
  assign y5709 = ~1'b0 ;
  assign y5710 = ~1'b0 ;
  assign y5711 = n23875 ;
  assign y5712 = ~n23877 ;
  assign y5713 = ~n23879 ;
  assign y5714 = ~n23880 ;
  assign y5715 = n23881 ;
  assign y5716 = n23886 ;
  assign y5717 = n23888 ;
  assign y5718 = ~n23891 ;
  assign y5719 = ~n23892 ;
  assign y5720 = n23894 ;
  assign y5721 = ~n23896 ;
  assign y5722 = n23905 ;
  assign y5723 = ~1'b0 ;
  assign y5724 = ~n23906 ;
  assign y5725 = n23913 ;
  assign y5726 = n23917 ;
  assign y5727 = n23919 ;
  assign y5728 = ~n23920 ;
  assign y5729 = n23921 ;
  assign y5730 = n23926 ;
  assign y5731 = ~n23928 ;
  assign y5732 = n23940 ;
  assign y5733 = n23941 ;
  assign y5734 = n23943 ;
  assign y5735 = n23950 ;
  assign y5736 = n23956 ;
  assign y5737 = ~n23957 ;
  assign y5738 = ~1'b0 ;
  assign y5739 = ~n23960 ;
  assign y5740 = ~n23968 ;
  assign y5741 = n23970 ;
  assign y5742 = n23974 ;
  assign y5743 = ~n23976 ;
  assign y5744 = ~n23978 ;
  assign y5745 = n23982 ;
  assign y5746 = n23986 ;
  assign y5747 = n23988 ;
  assign y5748 = n23995 ;
  assign y5749 = n24003 ;
  assign y5750 = ~n24004 ;
  assign y5751 = n24006 ;
  assign y5752 = n24009 ;
  assign y5753 = ~1'b0 ;
  assign y5754 = ~1'b0 ;
  assign y5755 = ~n24010 ;
  assign y5756 = n24012 ;
  assign y5757 = n24015 ;
  assign y5758 = ~n24016 ;
  assign y5759 = n24018 ;
  assign y5760 = ~n24020 ;
  assign y5761 = ~n24023 ;
  assign y5762 = n24024 ;
  assign y5763 = ~n24027 ;
  assign y5764 = ~n24028 ;
  assign y5765 = ~n24032 ;
  assign y5766 = n24033 ;
  assign y5767 = ~n24044 ;
  assign y5768 = ~1'b0 ;
  assign y5769 = n24046 ;
  assign y5770 = ~n24047 ;
  assign y5771 = ~n24048 ;
  assign y5772 = n24051 ;
  assign y5773 = ~n24053 ;
  assign y5774 = n24057 ;
  assign y5775 = ~n24064 ;
  assign y5776 = ~n24066 ;
  assign y5777 = ~n24067 ;
  assign y5778 = n24073 ;
  assign y5779 = ~n24074 ;
  assign y5780 = n24075 ;
  assign y5781 = n24076 ;
  assign y5782 = ~n24077 ;
  assign y5783 = n24078 ;
  assign y5784 = n24079 ;
  assign y5785 = ~1'b0 ;
  assign y5786 = n24081 ;
  assign y5787 = n24082 ;
  assign y5788 = ~n24083 ;
  assign y5789 = n24087 ;
  assign y5790 = n24089 ;
  assign y5791 = ~n24093 ;
  assign y5792 = ~n24094 ;
  assign y5793 = ~n24097 ;
  assign y5794 = n24098 ;
  assign y5795 = ~n24102 ;
  assign y5796 = n24104 ;
  assign y5797 = ~n24105 ;
  assign y5798 = n24107 ;
  assign y5799 = n24111 ;
  assign y5800 = ~n24112 ;
  assign y5801 = ~n24115 ;
  assign y5802 = ~n24120 ;
  assign y5803 = ~n24121 ;
  assign y5804 = n24124 ;
  assign y5805 = n24126 ;
  assign y5806 = n24135 ;
  assign y5807 = n24137 ;
  assign y5808 = n24138 ;
  assign y5809 = n24140 ;
  assign y5810 = ~n24142 ;
  assign y5811 = ~n24143 ;
  assign y5812 = n24147 ;
  assign y5813 = n24149 ;
  assign y5814 = ~n24151 ;
  assign y5815 = ~n24157 ;
  assign y5816 = ~n24160 ;
  assign y5817 = n24162 ;
  assign y5818 = ~n24165 ;
  assign y5819 = n24167 ;
  assign y5820 = ~n24172 ;
  assign y5821 = ~n24174 ;
  assign y5822 = ~n24175 ;
  assign y5823 = n24176 ;
  assign y5824 = n24180 ;
  assign y5825 = ~n24189 ;
  assign y5826 = ~n24192 ;
  assign y5827 = n24200 ;
  assign y5828 = ~n24202 ;
  assign y5829 = n24204 ;
  assign y5830 = ~n24205 ;
  assign y5831 = ~n24208 ;
  assign y5832 = n24213 ;
  assign y5833 = ~n24220 ;
  assign y5834 = n24223 ;
  assign y5835 = ~n24226 ;
  assign y5836 = n24229 ;
  assign y5837 = n24232 ;
  assign y5838 = n24237 ;
  assign y5839 = n24242 ;
  assign y5840 = n24243 ;
  assign y5841 = ~n24244 ;
  assign y5842 = ~n24248 ;
  assign y5843 = ~n24253 ;
  assign y5844 = n24256 ;
  assign y5845 = ~n24258 ;
  assign y5846 = ~1'b0 ;
  assign y5847 = ~n24259 ;
  assign y5848 = n24260 ;
  assign y5849 = n24263 ;
  assign y5850 = n24264 ;
  assign y5851 = n24266 ;
  assign y5852 = ~n24268 ;
  assign y5853 = ~n24269 ;
  assign y5854 = ~n24271 ;
  assign y5855 = n24275 ;
  assign y5856 = n24279 ;
  assign y5857 = n24280 ;
  assign y5858 = n24281 ;
  assign y5859 = n24284 ;
  assign y5860 = n24286 ;
  assign y5861 = ~n24288 ;
  assign y5862 = ~n24292 ;
  assign y5863 = n24294 ;
  assign y5864 = ~n24295 ;
  assign y5865 = ~n24305 ;
  assign y5866 = n24307 ;
  assign y5867 = ~n24310 ;
  assign y5868 = ~n24311 ;
  assign y5869 = ~n24316 ;
  assign y5870 = ~n24318 ;
  assign y5871 = ~n24319 ;
  assign y5872 = n24320 ;
  assign y5873 = ~n24321 ;
  assign y5874 = n24322 ;
  assign y5875 = n24331 ;
  assign y5876 = ~1'b0 ;
  assign y5877 = ~n24335 ;
  assign y5878 = ~n24338 ;
  assign y5879 = ~n24340 ;
  assign y5880 = n24343 ;
  assign y5881 = ~n24346 ;
  assign y5882 = ~n24350 ;
  assign y5883 = n24351 ;
  assign y5884 = ~n24355 ;
  assign y5885 = n24357 ;
  assign y5886 = ~n24361 ;
  assign y5887 = ~n24363 ;
  assign y5888 = ~n24364 ;
  assign y5889 = n24370 ;
  assign y5890 = n24373 ;
  assign y5891 = ~n24376 ;
  assign y5892 = ~n24381 ;
  assign y5893 = ~n24384 ;
  assign y5894 = n24385 ;
  assign y5895 = n24388 ;
  assign y5896 = ~n24389 ;
  assign y5897 = ~n24394 ;
  assign y5898 = ~n24397 ;
  assign y5899 = n24398 ;
  assign y5900 = n24401 ;
  assign y5901 = ~n24402 ;
  assign y5902 = ~n24403 ;
  assign y5903 = ~n24405 ;
  assign y5904 = ~n24406 ;
  assign y5905 = n24407 ;
  assign y5906 = ~n24409 ;
  assign y5907 = n24415 ;
  assign y5908 = ~n24417 ;
  assign y5909 = ~n24418 ;
  assign y5910 = ~n24421 ;
  assign y5911 = ~n24422 ;
  assign y5912 = ~n24427 ;
  assign y5913 = n24428 ;
  assign y5914 = ~n24429 ;
  assign y5915 = n24432 ;
  assign y5916 = n24434 ;
  assign y5917 = ~n24437 ;
  assign y5918 = ~n24438 ;
  assign y5919 = ~n24442 ;
  assign y5920 = n24443 ;
  assign y5921 = ~n24446 ;
  assign y5922 = ~n24448 ;
  assign y5923 = n24451 ;
  assign y5924 = ~n24452 ;
  assign y5925 = n24462 ;
  assign y5926 = ~n24463 ;
  assign y5927 = n24467 ;
  assign y5928 = n24468 ;
  assign y5929 = n24471 ;
  assign y5930 = ~n24476 ;
  assign y5931 = ~1'b0 ;
  assign y5932 = n24477 ;
  assign y5933 = n24479 ;
  assign y5934 = n24485 ;
  assign y5935 = n24489 ;
  assign y5936 = ~n24492 ;
  assign y5937 = ~n24496 ;
  assign y5938 = n24499 ;
  assign y5939 = ~n24500 ;
  assign y5940 = n24502 ;
  assign y5941 = ~1'b0 ;
  assign y5942 = n24503 ;
  assign y5943 = n24507 ;
  assign y5944 = ~n24509 ;
  assign y5945 = ~n24511 ;
  assign y5946 = n24512 ;
  assign y5947 = ~n24515 ;
  assign y5948 = n24517 ;
  assign y5949 = ~n24520 ;
  assign y5950 = n24521 ;
  assign y5951 = ~n24527 ;
  assign y5952 = ~n24532 ;
  assign y5953 = ~n24533 ;
  assign y5954 = n24539 ;
  assign y5955 = n24540 ;
  assign y5956 = ~n24541 ;
  assign y5957 = ~n24542 ;
  assign y5958 = n24546 ;
  assign y5959 = ~n24548 ;
  assign y5960 = n24550 ;
  assign y5961 = ~n24551 ;
  assign y5962 = n24552 ;
  assign y5963 = ~n24553 ;
  assign y5964 = n24554 ;
  assign y5965 = ~n24556 ;
  assign y5966 = ~n24559 ;
  assign y5967 = n24564 ;
  assign y5968 = ~n24566 ;
  assign y5969 = n24567 ;
  assign y5970 = n24570 ;
  assign y5971 = ~n24572 ;
  assign y5972 = n24573 ;
  assign y5973 = n24577 ;
  assign y5974 = n24581 ;
  assign y5975 = ~n24583 ;
  assign y5976 = ~n24590 ;
  assign y5977 = n24591 ;
  assign y5978 = ~n24595 ;
  assign y5979 = ~n24597 ;
  assign y5980 = n24600 ;
  assign y5981 = n24605 ;
  assign y5982 = n24609 ;
  assign y5983 = ~n24610 ;
  assign y5984 = ~n24613 ;
  assign y5985 = ~n24619 ;
  assign y5986 = n24622 ;
  assign y5987 = ~n24624 ;
  assign y5988 = ~n24629 ;
  assign y5989 = ~n24630 ;
  assign y5990 = ~1'b0 ;
  assign y5991 = n24632 ;
  assign y5992 = ~n24636 ;
  assign y5993 = n24638 ;
  assign y5994 = n24640 ;
  assign y5995 = n24643 ;
  assign y5996 = ~n24649 ;
  assign y5997 = ~1'b0 ;
  assign y5998 = ~n9990 ;
  assign y5999 = n24655 ;
  assign y6000 = n24656 ;
  assign y6001 = ~n24659 ;
  assign y6002 = n24660 ;
  assign y6003 = ~n24662 ;
  assign y6004 = ~n24664 ;
  assign y6005 = ~n24665 ;
  assign y6006 = ~n24667 ;
  assign y6007 = n24670 ;
  assign y6008 = n24675 ;
  assign y6009 = n24681 ;
  assign y6010 = n24683 ;
  assign y6011 = n24685 ;
  assign y6012 = ~n24690 ;
  assign y6013 = n24695 ;
  assign y6014 = ~n24696 ;
  assign y6015 = ~n24702 ;
  assign y6016 = n24705 ;
  assign y6017 = ~n24709 ;
  assign y6018 = n24711 ;
  assign y6019 = ~n24713 ;
  assign y6020 = ~n24716 ;
  assign y6021 = ~n24724 ;
  assign y6022 = ~n24728 ;
  assign y6023 = ~n24730 ;
  assign y6024 = n24732 ;
  assign y6025 = n24735 ;
  assign y6026 = ~n24737 ;
  assign y6027 = n24741 ;
  assign y6028 = ~n24747 ;
  assign y6029 = n24749 ;
  assign y6030 = ~n24750 ;
  assign y6031 = ~n24753 ;
  assign y6032 = n24754 ;
  assign y6033 = n24758 ;
  assign y6034 = n24762 ;
  assign y6035 = n24764 ;
  assign y6036 = ~1'b0 ;
  assign y6037 = n24766 ;
  assign y6038 = n24767 ;
  assign y6039 = n24768 ;
  assign y6040 = n24769 ;
  assign y6041 = n24772 ;
  assign y6042 = ~n24777 ;
  assign y6043 = n24778 ;
  assign y6044 = n24780 ;
  assign y6045 = n24782 ;
  assign y6046 = ~n24785 ;
  assign y6047 = n24786 ;
  assign y6048 = ~n24791 ;
  assign y6049 = ~n24792 ;
  assign y6050 = n24800 ;
  assign y6051 = n24804 ;
  assign y6052 = ~n24808 ;
  assign y6053 = ~n24811 ;
  assign y6054 = n24814 ;
  assign y6055 = n24816 ;
  assign y6056 = n24817 ;
  assign y6057 = ~n24818 ;
  assign y6058 = n24821 ;
  assign y6059 = ~n24822 ;
  assign y6060 = ~n24827 ;
  assign y6061 = n24830 ;
  assign y6062 = n24835 ;
  assign y6063 = n24839 ;
  assign y6064 = n24840 ;
  assign y6065 = ~n24841 ;
  assign y6066 = n24847 ;
  assign y6067 = n24848 ;
  assign y6068 = ~n24850 ;
  assign y6069 = ~n24851 ;
  assign y6070 = ~n24852 ;
  assign y6071 = n24857 ;
  assign y6072 = ~n24859 ;
  assign y6073 = n24862 ;
  assign y6074 = ~n24868 ;
  assign y6075 = ~n24869 ;
  assign y6076 = ~n24871 ;
  assign y6077 = n24873 ;
  assign y6078 = ~n24877 ;
  assign y6079 = n24878 ;
  assign y6080 = n24881 ;
  assign y6081 = ~n24882 ;
  assign y6082 = ~n24885 ;
  assign y6083 = n24892 ;
  assign y6084 = n24898 ;
  assign y6085 = ~n24903 ;
  assign y6086 = ~n24907 ;
  assign y6087 = n24912 ;
  assign y6088 = n24915 ;
  assign y6089 = n24919 ;
  assign y6090 = ~n24920 ;
  assign y6091 = ~n24924 ;
  assign y6092 = ~n24927 ;
  assign y6093 = n24929 ;
  assign y6094 = ~n24930 ;
  assign y6095 = ~n24931 ;
  assign y6096 = n24935 ;
  assign y6097 = ~n24936 ;
  assign y6098 = n24938 ;
  assign y6099 = ~1'b0 ;
  assign y6100 = n24940 ;
  assign y6101 = ~n24942 ;
  assign y6102 = n24944 ;
  assign y6103 = ~n24945 ;
  assign y6104 = n24947 ;
  assign y6105 = ~n24948 ;
  assign y6106 = n24952 ;
  assign y6107 = n24955 ;
  assign y6108 = ~n24966 ;
  assign y6109 = ~n24968 ;
  assign y6110 = ~n24970 ;
  assign y6111 = n24971 ;
  assign y6112 = n24973 ;
  assign y6113 = ~n24974 ;
  assign y6114 = ~n24978 ;
  assign y6115 = n24979 ;
  assign y6116 = n24980 ;
  assign y6117 = ~1'b0 ;
  assign y6118 = n24983 ;
  assign y6119 = ~n24985 ;
  assign y6120 = ~n24988 ;
  assign y6121 = ~n24989 ;
  assign y6122 = ~n24990 ;
  assign y6123 = n24996 ;
  assign y6124 = ~n24997 ;
  assign y6125 = ~n24998 ;
  assign y6126 = ~n25000 ;
  assign y6127 = ~1'b0 ;
  assign y6128 = ~n25002 ;
  assign y6129 = n25004 ;
  assign y6130 = ~n25006 ;
  assign y6131 = ~n25009 ;
  assign y6132 = ~n25010 ;
  assign y6133 = n25014 ;
  assign y6134 = ~n25015 ;
  assign y6135 = n25020 ;
  assign y6136 = n25022 ;
  assign y6137 = ~n25023 ;
  assign y6138 = n25024 ;
  assign y6139 = n25033 ;
  assign y6140 = ~n25036 ;
  assign y6141 = ~n25038 ;
  assign y6142 = n25042 ;
  assign y6143 = ~n25044 ;
  assign y6144 = ~n25047 ;
  assign y6145 = ~1'b0 ;
  assign y6146 = ~n25051 ;
  assign y6147 = ~n25052 ;
  assign y6148 = n25056 ;
  assign y6149 = n25057 ;
  assign y6150 = n25062 ;
  assign y6151 = n25063 ;
  assign y6152 = n25066 ;
  assign y6153 = n25070 ;
  assign y6154 = ~n25072 ;
  assign y6155 = ~1'b0 ;
  assign y6156 = n25073 ;
  assign y6157 = ~n25074 ;
  assign y6158 = ~n25078 ;
  assign y6159 = ~n25080 ;
  assign y6160 = n25081 ;
  assign y6161 = n25083 ;
  assign y6162 = ~1'b0 ;
  assign y6163 = n25085 ;
  assign y6164 = ~n25088 ;
  assign y6165 = n25092 ;
  assign y6166 = n25097 ;
  assign y6167 = ~n25098 ;
  assign y6168 = n25100 ;
  assign y6169 = ~n25103 ;
  assign y6170 = n25105 ;
  assign y6171 = ~n25108 ;
  assign y6172 = ~n25111 ;
  assign y6173 = n25113 ;
  assign y6174 = ~n25114 ;
  assign y6175 = n25116 ;
  assign y6176 = ~n25117 ;
  assign y6177 = ~n25118 ;
  assign y6178 = n25120 ;
  assign y6179 = ~n25123 ;
  assign y6180 = n25126 ;
  assign y6181 = ~1'b0 ;
  assign y6182 = n25127 ;
  assign y6183 = n25128 ;
  assign y6184 = n25129 ;
  assign y6185 = ~n2176 ;
  assign y6186 = ~n25130 ;
  assign y6187 = ~n25132 ;
  assign y6188 = n25140 ;
  assign y6189 = n25142 ;
  assign y6190 = ~n25143 ;
  assign y6191 = n25144 ;
  assign y6192 = ~n25146 ;
  assign y6193 = ~n25147 ;
  assign y6194 = ~n25150 ;
  assign y6195 = ~1'b0 ;
  assign y6196 = ~n25160 ;
  assign y6197 = ~n25166 ;
  assign y6198 = n25167 ;
  assign y6199 = ~n25168 ;
  assign y6200 = ~n25172 ;
  assign y6201 = n25174 ;
  assign y6202 = n25175 ;
  assign y6203 = n25176 ;
  assign y6204 = ~n25178 ;
  assign y6205 = n25179 ;
  assign y6206 = ~n25180 ;
  assign y6207 = ~n25184 ;
  assign y6208 = n25188 ;
  assign y6209 = n25193 ;
  assign y6210 = n25194 ;
  assign y6211 = ~n25195 ;
  assign y6212 = n25196 ;
  assign y6213 = ~n25201 ;
  assign y6214 = n25204 ;
  assign y6215 = ~n25206 ;
  assign y6216 = ~n25207 ;
  assign y6217 = n25209 ;
  assign y6218 = ~n25214 ;
  assign y6219 = n25218 ;
  assign y6220 = n25219 ;
  assign y6221 = n25220 ;
  assign y6222 = ~1'b0 ;
  assign y6223 = ~1'b0 ;
  assign y6224 = n25231 ;
  assign y6225 = n25235 ;
  assign y6226 = n25237 ;
  assign y6227 = ~n25238 ;
  assign y6228 = ~n25242 ;
  assign y6229 = n25247 ;
  assign y6230 = n25250 ;
  assign y6231 = ~1'b0 ;
  assign y6232 = n25253 ;
  assign y6233 = ~n25258 ;
  assign y6234 = n25260 ;
  assign y6235 = ~n25262 ;
  assign y6236 = n25264 ;
  assign y6237 = n25267 ;
  assign y6238 = n25269 ;
  assign y6239 = n25270 ;
  assign y6240 = n25272 ;
  assign y6241 = ~n25279 ;
  assign y6242 = ~n25280 ;
  assign y6243 = n25281 ;
  assign y6244 = n25282 ;
  assign y6245 = ~1'b0 ;
  assign y6246 = n25285 ;
  assign y6247 = n25293 ;
  assign y6248 = n25298 ;
  assign y6249 = ~n25299 ;
  assign y6250 = n25301 ;
  assign y6251 = n25303 ;
  assign y6252 = ~n25308 ;
  assign y6253 = ~1'b0 ;
  assign y6254 = n25309 ;
  assign y6255 = ~n25310 ;
  assign y6256 = ~n25311 ;
  assign y6257 = n25312 ;
  assign y6258 = ~n25314 ;
  assign y6259 = ~n25323 ;
  assign y6260 = ~1'b0 ;
  assign y6261 = n25324 ;
  assign y6262 = ~n25325 ;
  assign y6263 = n25326 ;
  assign y6264 = ~n25329 ;
  assign y6265 = ~n25335 ;
  assign y6266 = ~n25337 ;
  assign y6267 = n25338 ;
  assign y6268 = n25340 ;
  assign y6269 = ~n25343 ;
  assign y6270 = ~n25345 ;
  assign y6271 = ~n25347 ;
  assign y6272 = n25348 ;
  assign y6273 = ~n25351 ;
  assign y6274 = ~n25357 ;
  assign y6275 = ~1'b0 ;
  assign y6276 = n25360 ;
  assign y6277 = ~n25361 ;
  assign y6278 = n25368 ;
  assign y6279 = ~n25373 ;
  assign y6280 = n25374 ;
  assign y6281 = n25377 ;
  assign y6282 = ~n25378 ;
  assign y6283 = ~n25380 ;
  assign y6284 = ~n25386 ;
  assign y6285 = n25389 ;
  assign y6286 = n25392 ;
  assign y6287 = ~1'b0 ;
  assign y6288 = ~n25395 ;
  assign y6289 = n25404 ;
  assign y6290 = n25406 ;
  assign y6291 = n25411 ;
  assign y6292 = ~n25413 ;
  assign y6293 = ~n25416 ;
  assign y6294 = n25419 ;
  assign y6295 = ~n25422 ;
  assign y6296 = n25430 ;
  assign y6297 = ~n25431 ;
  assign y6298 = ~n25432 ;
  assign y6299 = ~n25433 ;
  assign y6300 = ~n25436 ;
  assign y6301 = ~n25440 ;
  assign y6302 = ~1'b0 ;
  assign y6303 = ~n25441 ;
  assign y6304 = n25446 ;
  assign y6305 = ~n25447 ;
  assign y6306 = n624 ;
  assign y6307 = n25450 ;
  assign y6308 = ~n25453 ;
  assign y6309 = n25454 ;
  assign y6310 = n25457 ;
  assign y6311 = ~n25458 ;
  assign y6312 = n25459 ;
  assign y6313 = n25461 ;
  assign y6314 = ~n25465 ;
  assign y6315 = n25467 ;
  assign y6316 = ~n25473 ;
  assign y6317 = n25479 ;
  assign y6318 = n25482 ;
  assign y6319 = ~n25483 ;
  assign y6320 = ~n25484 ;
  assign y6321 = ~n25485 ;
  assign y6322 = ~n25487 ;
  assign y6323 = n25488 ;
  assign y6324 = ~n25495 ;
  assign y6325 = ~n25500 ;
  assign y6326 = ~1'b0 ;
  assign y6327 = ~1'b0 ;
  assign y6328 = n25501 ;
  assign y6329 = ~n25503 ;
  assign y6330 = ~n25512 ;
  assign y6331 = ~n25515 ;
  assign y6332 = ~n25517 ;
  assign y6333 = n25521 ;
  assign y6334 = n25523 ;
  assign y6335 = ~n25526 ;
  assign y6336 = ~n25530 ;
  assign y6337 = n25531 ;
  assign y6338 = ~1'b0 ;
  assign y6339 = n25534 ;
  assign y6340 = n25537 ;
  assign y6341 = n25541 ;
  assign y6342 = n25545 ;
  assign y6343 = n25548 ;
  assign y6344 = ~n25549 ;
  assign y6345 = ~n25550 ;
  assign y6346 = n25551 ;
  assign y6347 = n25555 ;
  assign y6348 = n25559 ;
  assign y6349 = n25560 ;
  assign y6350 = n25561 ;
  assign y6351 = n25562 ;
  assign y6352 = ~n25570 ;
  assign y6353 = n25574 ;
  assign y6354 = n25577 ;
  assign y6355 = ~1'b0 ;
  assign y6356 = n25578 ;
  assign y6357 = n25584 ;
  assign y6358 = n25587 ;
  assign y6359 = ~n25588 ;
  assign y6360 = ~n25594 ;
  assign y6361 = n25597 ;
  assign y6362 = ~n25599 ;
  assign y6363 = ~1'b0 ;
  assign y6364 = n25602 ;
  assign y6365 = ~n25606 ;
  assign y6366 = ~n25608 ;
  assign y6367 = ~n25609 ;
  assign y6368 = ~n25617 ;
  assign y6369 = ~n25618 ;
  assign y6370 = ~n25619 ;
  assign y6371 = n25622 ;
  assign y6372 = n25624 ;
  assign y6373 = n25626 ;
  assign y6374 = n25629 ;
  assign y6375 = ~n25631 ;
  assign y6376 = ~n25632 ;
  assign y6377 = n25635 ;
  assign y6378 = ~n25636 ;
  assign y6379 = ~n25637 ;
  assign y6380 = ~n25639 ;
  assign y6381 = ~n25641 ;
  assign y6382 = ~n25643 ;
  assign y6383 = ~n25645 ;
  assign y6384 = ~n25647 ;
  assign y6385 = ~n25652 ;
  assign y6386 = ~n25653 ;
  assign y6387 = n25658 ;
  assign y6388 = n25659 ;
  assign y6389 = n25663 ;
  assign y6390 = n25666 ;
  assign y6391 = ~n25670 ;
  assign y6392 = n25673 ;
  assign y6393 = ~n25677 ;
  assign y6394 = n25678 ;
  assign y6395 = ~n25679 ;
  assign y6396 = ~n25681 ;
  assign y6397 = n25685 ;
  assign y6398 = ~n25687 ;
  assign y6399 = ~n25689 ;
  assign y6400 = ~n25692 ;
  assign y6401 = n25693 ;
  assign y6402 = n25694 ;
  assign y6403 = n25696 ;
  assign y6404 = ~n25698 ;
  assign y6405 = n25700 ;
  assign y6406 = ~n25702 ;
  assign y6407 = ~n25704 ;
  assign y6408 = ~n25706 ;
  assign y6409 = ~n25707 ;
  assign y6410 = n25716 ;
  assign y6411 = ~n25717 ;
  assign y6412 = ~n25722 ;
  assign y6413 = ~n25725 ;
  assign y6414 = ~n25726 ;
  assign y6415 = n25728 ;
  assign y6416 = ~n25729 ;
  assign y6417 = ~n25732 ;
  assign y6418 = ~1'b0 ;
  assign y6419 = n25737 ;
  assign y6420 = n25740 ;
  assign y6421 = n25742 ;
  assign y6422 = n25745 ;
  assign y6423 = ~n25748 ;
  assign y6424 = n25749 ;
  assign y6425 = n25751 ;
  assign y6426 = n25755 ;
  assign y6427 = n25756 ;
  assign y6428 = ~n25759 ;
  assign y6429 = n25761 ;
  assign y6430 = n25763 ;
  assign y6431 = n25768 ;
  assign y6432 = ~n25771 ;
  assign y6433 = n25778 ;
  assign y6434 = ~n25783 ;
  assign y6435 = n25786 ;
  assign y6436 = ~n25788 ;
  assign y6437 = ~n25790 ;
  assign y6438 = ~n25791 ;
  assign y6439 = ~n25794 ;
  assign y6440 = ~n25798 ;
  assign y6441 = n25803 ;
  assign y6442 = ~n25808 ;
  assign y6443 = n25809 ;
  assign y6444 = n25816 ;
  assign y6445 = ~n25818 ;
  assign y6446 = n25821 ;
  assign y6447 = ~n25822 ;
  assign y6448 = n25823 ;
  assign y6449 = ~n25827 ;
  assign y6450 = ~n15552 ;
  assign y6451 = ~n25829 ;
  assign y6452 = ~n25830 ;
  assign y6453 = n25831 ;
  assign y6454 = ~n25836 ;
  assign y6455 = ~n25837 ;
  assign y6456 = ~n25841 ;
  assign y6457 = ~n25842 ;
  assign y6458 = n25843 ;
  assign y6459 = n25850 ;
  assign y6460 = ~n25851 ;
  assign y6461 = ~n25853 ;
  assign y6462 = ~n25854 ;
  assign y6463 = n25859 ;
  assign y6464 = n25862 ;
  assign y6465 = n25866 ;
  assign y6466 = n25870 ;
  assign y6467 = n25878 ;
  assign y6468 = ~n25880 ;
  assign y6469 = n25882 ;
  assign y6470 = ~n25884 ;
  assign y6471 = n25886 ;
  assign y6472 = ~n25890 ;
  assign y6473 = n25893 ;
  assign y6474 = ~n25894 ;
  assign y6475 = ~n25895 ;
  assign y6476 = n25899 ;
  assign y6477 = ~n25901 ;
  assign y6478 = n25902 ;
  assign y6479 = ~n25903 ;
  assign y6480 = n25904 ;
  assign y6481 = n25907 ;
  assign y6482 = n25912 ;
  assign y6483 = ~n25916 ;
  assign y6484 = n25919 ;
  assign y6485 = ~n25925 ;
  assign y6486 = ~n25930 ;
  assign y6487 = ~n25931 ;
  assign y6488 = ~n25932 ;
  assign y6489 = n25935 ;
  assign y6490 = ~n25936 ;
  assign y6491 = ~n25940 ;
  assign y6492 = ~n25941 ;
  assign y6493 = ~n25942 ;
  assign y6494 = n25944 ;
  assign y6495 = ~n25946 ;
  assign y6496 = ~n25951 ;
  assign y6497 = ~n25952 ;
  assign y6498 = n25953 ;
  assign y6499 = ~n25957 ;
  assign y6500 = ~n25962 ;
  assign y6501 = ~n25967 ;
  assign y6502 = ~n25970 ;
  assign y6503 = ~n25974 ;
  assign y6504 = ~n25975 ;
  assign y6505 = n25976 ;
  assign y6506 = ~n25977 ;
  assign y6507 = ~n25980 ;
  assign y6508 = ~n25983 ;
  assign y6509 = ~n25986 ;
  assign y6510 = ~n25988 ;
  assign y6511 = ~n25992 ;
  assign y6512 = n25995 ;
  assign y6513 = ~n25999 ;
  assign y6514 = n26000 ;
  assign y6515 = ~n26002 ;
  assign y6516 = n26005 ;
  assign y6517 = ~1'b0 ;
  assign y6518 = ~n26006 ;
  assign y6519 = n26009 ;
  assign y6520 = n26010 ;
  assign y6521 = n26012 ;
  assign y6522 = n26029 ;
  assign y6523 = n26032 ;
  assign y6524 = n26036 ;
  assign y6525 = n26040 ;
  assign y6526 = ~n26041 ;
  assign y6527 = n26042 ;
  assign y6528 = ~1'b0 ;
  assign y6529 = ~1'b0 ;
  assign y6530 = ~n26045 ;
  assign y6531 = n26050 ;
  assign y6532 = ~n26051 ;
  assign y6533 = n26053 ;
  assign y6534 = ~n26054 ;
  assign y6535 = ~n26056 ;
  assign y6536 = ~n26060 ;
  assign y6537 = ~n26061 ;
  assign y6538 = ~n26063 ;
  assign y6539 = ~1'b0 ;
  assign y6540 = ~n26066 ;
  assign y6541 = n26067 ;
  assign y6542 = ~n26068 ;
  assign y6543 = ~n26072 ;
  assign y6544 = n26073 ;
  assign y6545 = n26075 ;
  assign y6546 = ~n26079 ;
  assign y6547 = ~n26083 ;
  assign y6548 = n26085 ;
  assign y6549 = ~1'b0 ;
  assign y6550 = ~n26087 ;
  assign y6551 = n26095 ;
  assign y6552 = n26097 ;
  assign y6553 = ~n26100 ;
  assign y6554 = n26101 ;
  assign y6555 = n26108 ;
  assign y6556 = n26109 ;
  assign y6557 = ~n26114 ;
  assign y6558 = n26118 ;
  assign y6559 = n26119 ;
  assign y6560 = n26120 ;
  assign y6561 = n26121 ;
  assign y6562 = n26122 ;
  assign y6563 = n26124 ;
  assign y6564 = ~n26125 ;
  assign y6565 = n26131 ;
  assign y6566 = n26132 ;
  assign y6567 = n26133 ;
  assign y6568 = ~n26134 ;
  assign y6569 = n26137 ;
  assign y6570 = n26140 ;
  assign y6571 = ~n26141 ;
  assign y6572 = ~n26143 ;
  assign y6573 = ~1'b0 ;
  assign y6574 = n26145 ;
  assign y6575 = ~n26148 ;
  assign y6576 = n26149 ;
  assign y6577 = ~n26151 ;
  assign y6578 = n26152 ;
  assign y6579 = ~n26155 ;
  assign y6580 = ~n26157 ;
  assign y6581 = n26159 ;
  assign y6582 = ~n26160 ;
  assign y6583 = n26161 ;
  assign y6584 = ~n26165 ;
  assign y6585 = n26168 ;
  assign y6586 = n26169 ;
  assign y6587 = ~n26172 ;
  assign y6588 = n26178 ;
  assign y6589 = ~n26179 ;
  assign y6590 = ~n26181 ;
  assign y6591 = n26184 ;
  assign y6592 = ~n26186 ;
  assign y6593 = ~1'b0 ;
  assign y6594 = n26187 ;
  assign y6595 = ~n26189 ;
  assign y6596 = ~n26192 ;
  assign y6597 = n26196 ;
  assign y6598 = n26197 ;
  assign y6599 = ~n26201 ;
  assign y6600 = n26208 ;
  assign y6601 = n26210 ;
  assign y6602 = ~n26212 ;
  assign y6603 = ~n26218 ;
  assign y6604 = ~n26219 ;
  assign y6605 = n26221 ;
  assign y6606 = n26224 ;
  assign y6607 = n26225 ;
  assign y6608 = ~n26231 ;
  assign y6609 = ~n26233 ;
  assign y6610 = n26237 ;
  assign y6611 = ~n26242 ;
  assign y6612 = ~n26245 ;
  assign y6613 = n26248 ;
  assign y6614 = n26249 ;
  assign y6615 = n26251 ;
  assign y6616 = n26253 ;
  assign y6617 = n26256 ;
  assign y6618 = n26258 ;
  assign y6619 = n26260 ;
  assign y6620 = ~n26263 ;
  assign y6621 = ~n26267 ;
  assign y6622 = n26268 ;
  assign y6623 = ~n26271 ;
  assign y6624 = n26274 ;
  assign y6625 = n26278 ;
  assign y6626 = n26281 ;
  assign y6627 = ~n26282 ;
  assign y6628 = n26286 ;
  assign y6629 = ~1'b0 ;
  assign y6630 = n26295 ;
  assign y6631 = n26299 ;
  assign y6632 = ~1'b0 ;
  assign y6633 = n26301 ;
  assign y6634 = ~n26303 ;
  assign y6635 = ~n26306 ;
  assign y6636 = ~n26310 ;
  assign y6637 = ~1'b0 ;
  assign y6638 = ~n26313 ;
  assign y6639 = ~n26315 ;
  assign y6640 = ~n26316 ;
  assign y6641 = n26318 ;
  assign y6642 = n26323 ;
  assign y6643 = n26327 ;
  assign y6644 = n26331 ;
  assign y6645 = n26332 ;
  assign y6646 = ~n26334 ;
  assign y6647 = 1'b0 ;
  assign y6648 = ~n26338 ;
  assign y6649 = ~n26344 ;
  assign y6650 = ~n26346 ;
  assign y6651 = ~n26347 ;
  assign y6652 = ~n26350 ;
  assign y6653 = ~n26356 ;
  assign y6654 = ~n26359 ;
  assign y6655 = n26362 ;
  assign y6656 = ~n26364 ;
  assign y6657 = n26365 ;
  assign y6658 = n26368 ;
  assign y6659 = n26372 ;
  assign y6660 = ~n26373 ;
  assign y6661 = n26375 ;
  assign y6662 = ~n26378 ;
  assign y6663 = ~n26382 ;
  assign y6664 = n26385 ;
  assign y6665 = ~n26388 ;
  assign y6666 = ~n26392 ;
  assign y6667 = n26401 ;
  assign y6668 = ~n26402 ;
  assign y6669 = ~n26403 ;
  assign y6670 = n26408 ;
  assign y6671 = n26412 ;
  assign y6672 = ~n26414 ;
  assign y6673 = ~n26415 ;
  assign y6674 = ~n26416 ;
  assign y6675 = ~n26419 ;
  assign y6676 = ~n26425 ;
  assign y6677 = ~n26426 ;
  assign y6678 = ~n26429 ;
  assign y6679 = ~1'b0 ;
  assign y6680 = n26431 ;
  assign y6681 = ~n26432 ;
  assign y6682 = n26433 ;
  assign y6683 = ~n26437 ;
  assign y6684 = n26442 ;
  assign y6685 = ~n26444 ;
  assign y6686 = ~n26448 ;
  assign y6687 = ~n26450 ;
  assign y6688 = ~n26454 ;
  assign y6689 = ~1'b0 ;
  assign y6690 = ~n26457 ;
  assign y6691 = n26458 ;
  assign y6692 = ~n26460 ;
  assign y6693 = n26462 ;
  assign y6694 = ~n26464 ;
  assign y6695 = ~n26465 ;
  assign y6696 = n26466 ;
  assign y6697 = n26468 ;
  assign y6698 = ~n26469 ;
  assign y6699 = ~n26470 ;
  assign y6700 = n26471 ;
  assign y6701 = n26478 ;
  assign y6702 = ~n26479 ;
  assign y6703 = n26480 ;
  assign y6704 = ~n26483 ;
  assign y6705 = n26486 ;
  assign y6706 = ~n26487 ;
  assign y6707 = n26493 ;
  assign y6708 = ~n26494 ;
  assign y6709 = n26496 ;
  assign y6710 = n26497 ;
  assign y6711 = n26498 ;
  assign y6712 = n26500 ;
  assign y6713 = ~n26502 ;
  assign y6714 = ~n26507 ;
  assign y6715 = ~n26511 ;
  assign y6716 = n26518 ;
  assign y6717 = n26520 ;
  assign y6718 = ~n26523 ;
  assign y6719 = n26525 ;
  assign y6720 = ~1'b0 ;
  assign y6721 = ~n26527 ;
  assign y6722 = n26535 ;
  assign y6723 = ~n26538 ;
  assign y6724 = ~n26539 ;
  assign y6725 = n26543 ;
  assign y6726 = ~n26544 ;
  assign y6727 = ~n26546 ;
  assign y6728 = n26549 ;
  assign y6729 = n26550 ;
  assign y6730 = n26551 ;
  assign y6731 = ~n26552 ;
  assign y6732 = n26553 ;
  assign y6733 = n26556 ;
  assign y6734 = n26564 ;
  assign y6735 = ~n26565 ;
  assign y6736 = ~1'b0 ;
  assign y6737 = n26569 ;
  assign y6738 = n26571 ;
  assign y6739 = ~n26573 ;
  assign y6740 = n26574 ;
  assign y6741 = ~n26576 ;
  assign y6742 = ~n26579 ;
  assign y6743 = n26586 ;
  assign y6744 = n26589 ;
  assign y6745 = n15082 ;
  assign y6746 = ~1'b0 ;
  assign y6747 = ~n26593 ;
  assign y6748 = ~n26596 ;
  assign y6749 = ~n26597 ;
  assign y6750 = ~n26599 ;
  assign y6751 = n26600 ;
  assign y6752 = ~n26601 ;
  assign y6753 = ~n26612 ;
  assign y6754 = ~1'b0 ;
  assign y6755 = ~n26618 ;
  assign y6756 = n26626 ;
  assign y6757 = n26627 ;
  assign y6758 = n26629 ;
  assign y6759 = ~n26636 ;
  assign y6760 = ~n5168 ;
  assign y6761 = n26638 ;
  assign y6762 = ~n26642 ;
  assign y6763 = ~n26643 ;
  assign y6764 = n26645 ;
  assign y6765 = ~n26648 ;
  assign y6766 = ~n26650 ;
  assign y6767 = n26651 ;
  assign y6768 = ~n26657 ;
  assign y6769 = n26658 ;
  assign y6770 = ~n26660 ;
  assign y6771 = ~n26661 ;
  assign y6772 = n26665 ;
  assign y6773 = n26666 ;
  assign y6774 = n26667 ;
  assign y6775 = ~n26675 ;
  assign y6776 = ~n26678 ;
  assign y6777 = n26681 ;
  assign y6778 = n26683 ;
  assign y6779 = ~1'b0 ;
  assign y6780 = ~n26684 ;
  assign y6781 = ~n26685 ;
  assign y6782 = n26686 ;
  assign y6783 = n26687 ;
  assign y6784 = n26691 ;
  assign y6785 = n26696 ;
  assign y6786 = n26697 ;
  assign y6787 = n26699 ;
  assign y6788 = ~n26700 ;
  assign y6789 = n26702 ;
  assign y6790 = n26704 ;
  assign y6791 = ~n26705 ;
  assign y6792 = ~n26706 ;
  assign y6793 = n26708 ;
  assign y6794 = ~n26710 ;
  assign y6795 = ~n10291 ;
  assign y6796 = n26712 ;
  assign y6797 = n26716 ;
  assign y6798 = ~n26718 ;
  assign y6799 = ~n26721 ;
  assign y6800 = n26722 ;
  assign y6801 = ~n26724 ;
  assign y6802 = ~n26725 ;
  assign y6803 = ~n26727 ;
  assign y6804 = ~n26729 ;
  assign y6805 = n26730 ;
  assign y6806 = n26735 ;
  assign y6807 = n26739 ;
  assign y6808 = ~n26742 ;
  assign y6809 = n26744 ;
  assign y6810 = ~n26748 ;
  assign y6811 = ~n26750 ;
  assign y6812 = n26752 ;
  assign y6813 = n26754 ;
  assign y6814 = ~n26757 ;
  assign y6815 = n26758 ;
  assign y6816 = ~n26761 ;
  assign y6817 = n26764 ;
  assign y6818 = ~n26769 ;
  assign y6819 = n26775 ;
  assign y6820 = ~n26778 ;
  assign y6821 = ~1'b0 ;
  assign y6822 = ~n26779 ;
  assign y6823 = ~n26782 ;
  assign y6824 = ~n26786 ;
  assign y6825 = ~n26787 ;
  assign y6826 = n26789 ;
  assign y6827 = n26794 ;
  assign y6828 = ~n26798 ;
  assign y6829 = n26800 ;
  assign y6830 = ~n26802 ;
  assign y6831 = ~n26803 ;
  assign y6832 = n26805 ;
  assign y6833 = ~n26808 ;
  assign y6834 = n26815 ;
  assign y6835 = ~n26816 ;
  assign y6836 = n26818 ;
  assign y6837 = ~1'b0 ;
  assign y6838 = ~1'b0 ;
  assign y6839 = n26819 ;
  assign y6840 = ~n26825 ;
  assign y6841 = n26828 ;
  assign y6842 = n26829 ;
  assign y6843 = ~n26831 ;
  assign y6844 = ~n26834 ;
  assign y6845 = ~n26835 ;
  assign y6846 = ~n26836 ;
  assign y6847 = ~n26839 ;
  assign y6848 = ~n26841 ;
  assign y6849 = ~n26842 ;
  assign y6850 = n26846 ;
  assign y6851 = n26852 ;
  assign y6852 = ~n26854 ;
  assign y6853 = n26858 ;
  assign y6854 = ~n26860 ;
  assign y6855 = ~n26864 ;
  assign y6856 = ~n26866 ;
  assign y6857 = n26869 ;
  assign y6858 = ~n26870 ;
  assign y6859 = n26874 ;
  assign y6860 = n26875 ;
  assign y6861 = ~n26876 ;
  assign y6862 = ~n26878 ;
  assign y6863 = n26881 ;
  assign y6864 = ~n26884 ;
  assign y6865 = n26886 ;
  assign y6866 = ~n26888 ;
  assign y6867 = n26889 ;
  assign y6868 = n26890 ;
  assign y6869 = ~n26892 ;
  assign y6870 = n26893 ;
  assign y6871 = ~n26894 ;
  assign y6872 = n26895 ;
  assign y6873 = ~n26902 ;
  assign y6874 = n26904 ;
  assign y6875 = ~n26908 ;
  assign y6876 = ~1'b0 ;
  assign y6877 = ~n26910 ;
  assign y6878 = ~n26911 ;
  assign y6879 = n26913 ;
  assign y6880 = n26915 ;
  assign y6881 = ~n26917 ;
  assign y6882 = n26919 ;
  assign y6883 = n26920 ;
  assign y6884 = ~n26924 ;
  assign y6885 = ~n26926 ;
  assign y6886 = n26927 ;
  assign y6887 = ~1'b0 ;
  assign y6888 = n26930 ;
  assign y6889 = n26933 ;
  assign y6890 = n26934 ;
  assign y6891 = ~n26935 ;
  assign y6892 = n26936 ;
  assign y6893 = n26939 ;
  assign y6894 = ~n26947 ;
  assign y6895 = n26952 ;
  assign y6896 = ~n26954 ;
  assign y6897 = ~n26957 ;
  assign y6898 = n26960 ;
  assign y6899 = ~n26962 ;
  assign y6900 = n26964 ;
  assign y6901 = ~n26968 ;
  assign y6902 = ~n26970 ;
  assign y6903 = ~n26975 ;
  assign y6904 = n26981 ;
  assign y6905 = n26984 ;
  assign y6906 = n26986 ;
  assign y6907 = n26989 ;
  assign y6908 = ~n26993 ;
  assign y6909 = n27000 ;
  assign y6910 = ~n27004 ;
  assign y6911 = ~n27008 ;
  assign y6912 = ~n27012 ;
  assign y6913 = ~n27014 ;
  assign y6914 = ~n27018 ;
  assign y6915 = ~n27022 ;
  assign y6916 = ~n27024 ;
  assign y6917 = ~n27029 ;
  assign y6918 = n8823 ;
  assign y6919 = ~n27031 ;
  assign y6920 = n27034 ;
  assign y6921 = n27035 ;
  assign y6922 = n27037 ;
  assign y6923 = ~n27038 ;
  assign y6924 = n27046 ;
  assign y6925 = n27048 ;
  assign y6926 = ~n27049 ;
  assign y6927 = n27051 ;
  assign y6928 = n27059 ;
  assign y6929 = n27060 ;
  assign y6930 = n27061 ;
  assign y6931 = ~n27063 ;
  assign y6932 = n27064 ;
  assign y6933 = n27066 ;
  assign y6934 = ~1'b0 ;
  assign y6935 = ~n27069 ;
  assign y6936 = n27070 ;
  assign y6937 = ~n27073 ;
  assign y6938 = n27074 ;
  assign y6939 = ~n27078 ;
  assign y6940 = ~n27079 ;
  assign y6941 = n27081 ;
  assign y6942 = ~n27082 ;
  assign y6943 = ~1'b0 ;
  assign y6944 = n27084 ;
  assign y6945 = n27088 ;
  assign y6946 = n27090 ;
  assign y6947 = ~n27091 ;
  assign y6948 = ~n27092 ;
  assign y6949 = n27094 ;
  assign y6950 = ~n27096 ;
  assign y6951 = ~n27097 ;
  assign y6952 = n27100 ;
  assign y6953 = ~n27104 ;
  assign y6954 = n27105 ;
  assign y6955 = n27107 ;
  assign y6956 = n27108 ;
  assign y6957 = ~n27109 ;
  assign y6958 = n27110 ;
  assign y6959 = n27111 ;
  assign y6960 = ~n27114 ;
  assign y6961 = ~1'b0 ;
  assign y6962 = n27116 ;
  assign y6963 = ~n27118 ;
  assign y6964 = n27119 ;
  assign y6965 = ~n27120 ;
  assign y6966 = ~n27123 ;
  assign y6967 = ~n27125 ;
  assign y6968 = ~n27127 ;
  assign y6969 = ~n27132 ;
  assign y6970 = n27133 ;
  assign y6971 = n27136 ;
  assign y6972 = n27137 ;
  assign y6973 = ~n27138 ;
  assign y6974 = ~n27140 ;
  assign y6975 = n27141 ;
  assign y6976 = ~n27142 ;
  assign y6977 = n27143 ;
  assign y6978 = ~n27151 ;
  assign y6979 = n27155 ;
  assign y6980 = n27157 ;
  assign y6981 = ~n27160 ;
  assign y6982 = n27162 ;
  assign y6983 = ~n27165 ;
  assign y6984 = ~n27170 ;
  assign y6985 = n27177 ;
  assign y6986 = ~n27178 ;
  assign y6987 = n27182 ;
  assign y6988 = n27185 ;
  assign y6989 = ~n27186 ;
  assign y6990 = ~n27189 ;
  assign y6991 = ~n27190 ;
  assign y6992 = ~1'b0 ;
  assign y6993 = ~n27191 ;
  assign y6994 = ~n27192 ;
  assign y6995 = n27193 ;
  assign y6996 = ~n27195 ;
  assign y6997 = ~n27196 ;
  assign y6998 = ~n27198 ;
  assign y6999 = ~n27200 ;
  assign y7000 = ~1'b0 ;
  assign y7001 = ~n27202 ;
  assign y7002 = ~n27206 ;
  assign y7003 = n27207 ;
  assign y7004 = ~n27208 ;
  assign y7005 = ~n27209 ;
  assign y7006 = n27210 ;
  assign y7007 = n27212 ;
  assign y7008 = n27216 ;
  assign y7009 = ~n27219 ;
  assign y7010 = ~n27221 ;
  assign y7011 = ~n27222 ;
  assign y7012 = ~n27223 ;
  assign y7013 = ~n27225 ;
  assign y7014 = n27226 ;
  assign y7015 = n27229 ;
  assign y7016 = ~n27232 ;
  assign y7017 = n27234 ;
  assign y7018 = ~n27236 ;
  assign y7019 = ~n27238 ;
  assign y7020 = ~n27240 ;
  assign y7021 = n27241 ;
  assign y7022 = ~n27249 ;
  assign y7023 = ~n27251 ;
  assign y7024 = ~n27252 ;
  assign y7025 = ~n27253 ;
  assign y7026 = ~n27255 ;
  assign y7027 = n27256 ;
  assign y7028 = ~1'b0 ;
  assign y7029 = ~1'b0 ;
  assign y7030 = n27257 ;
  assign y7031 = ~n27258 ;
  assign y7032 = n27260 ;
  assign y7033 = ~n27261 ;
  assign y7034 = ~n27263 ;
  assign y7035 = n27265 ;
  assign y7036 = ~n27273 ;
  assign y7037 = n27274 ;
  assign y7038 = ~1'b0 ;
  assign y7039 = ~n27277 ;
  assign y7040 = ~n27283 ;
  assign y7041 = ~n27286 ;
  assign y7042 = ~n27287 ;
  assign y7043 = ~n27288 ;
  assign y7044 = ~n27289 ;
  assign y7045 = ~n27293 ;
  assign y7046 = n27299 ;
  assign y7047 = n27301 ;
  assign y7048 = n27302 ;
  assign y7049 = n27306 ;
  assign y7050 = ~n27309 ;
  assign y7051 = n27311 ;
  assign y7052 = ~n27313 ;
  assign y7053 = n27316 ;
  assign y7054 = n27318 ;
  assign y7055 = ~n27323 ;
  assign y7056 = ~1'b0 ;
  assign y7057 = n27325 ;
  assign y7058 = n27326 ;
  assign y7059 = n27328 ;
  assign y7060 = n27333 ;
  assign y7061 = ~n27335 ;
  assign y7062 = ~n27340 ;
  assign y7063 = n27343 ;
  assign y7064 = n27348 ;
  assign y7065 = n27350 ;
  assign y7066 = n27352 ;
  assign y7067 = n27353 ;
  assign y7068 = n27362 ;
  assign y7069 = n27364 ;
  assign y7070 = ~n27365 ;
  assign y7071 = ~n27367 ;
  assign y7072 = n27368 ;
  assign y7073 = n27370 ;
  assign y7074 = n27371 ;
  assign y7075 = ~n27373 ;
  assign y7076 = ~n27376 ;
  assign y7077 = n27378 ;
  assign y7078 = ~n27382 ;
  assign y7079 = ~n27385 ;
  assign y7080 = n27387 ;
  assign y7081 = n27389 ;
  assign y7082 = n27393 ;
  assign y7083 = ~n27395 ;
  assign y7084 = n27397 ;
  assign y7085 = ~n27400 ;
  assign y7086 = ~n27401 ;
  assign y7087 = n27406 ;
  assign y7088 = n27407 ;
  assign y7089 = ~n27408 ;
  assign y7090 = ~n27409 ;
  assign y7091 = n27411 ;
  assign y7092 = ~n27413 ;
  assign y7093 = n27414 ;
  assign y7094 = ~n27417 ;
  assign y7095 = n27423 ;
  assign y7096 = ~n27428 ;
  assign y7097 = ~n27429 ;
  assign y7098 = ~n27431 ;
  assign y7099 = ~n9791 ;
  assign y7100 = ~n27432 ;
  assign y7101 = n27434 ;
  assign y7102 = ~1'b0 ;
  assign y7103 = ~n27436 ;
  assign y7104 = n27437 ;
  assign y7105 = n27443 ;
  assign y7106 = n27444 ;
  assign y7107 = ~n27445 ;
  assign y7108 = ~n27447 ;
  assign y7109 = n27452 ;
  assign y7110 = ~1'b0 ;
  assign y7111 = ~n27454 ;
  assign y7112 = ~n27455 ;
  assign y7113 = ~n27459 ;
  assign y7114 = ~n27460 ;
  assign y7115 = ~n27461 ;
  assign y7116 = n27466 ;
  assign y7117 = ~n27468 ;
  assign y7118 = n27478 ;
  assign y7119 = ~1'b0 ;
  assign y7120 = n27480 ;
  assign y7121 = ~n27489 ;
  assign y7122 = n27492 ;
  assign y7123 = ~n27493 ;
  assign y7124 = n27496 ;
  assign y7125 = n27497 ;
  assign y7126 = ~n27499 ;
  assign y7127 = ~1'b0 ;
  assign y7128 = ~1'b0 ;
  assign y7129 = ~n27502 ;
  assign y7130 = ~n27503 ;
  assign y7131 = ~n27507 ;
  assign y7132 = ~n27511 ;
  assign y7133 = n27516 ;
  assign y7134 = ~n27519 ;
  assign y7135 = ~n27521 ;
  assign y7136 = ~n27523 ;
  assign y7137 = n27524 ;
  assign y7138 = n27527 ;
  assign y7139 = ~n27535 ;
  assign y7140 = ~n27537 ;
  assign y7141 = n27541 ;
  assign y7142 = ~n27542 ;
  assign y7143 = ~n27544 ;
  assign y7144 = ~n27548 ;
  assign y7145 = n27550 ;
  assign y7146 = n27553 ;
  assign y7147 = ~n27554 ;
  assign y7148 = n27555 ;
  assign y7149 = ~n27562 ;
  assign y7150 = n27564 ;
  assign y7151 = n27566 ;
  assign y7152 = n27571 ;
  assign y7153 = n27573 ;
  assign y7154 = ~n27578 ;
  assign y7155 = n27583 ;
  assign y7156 = n27584 ;
  assign y7157 = ~n27586 ;
  assign y7158 = n27590 ;
  assign y7159 = n27591 ;
  assign y7160 = n27592 ;
  assign y7161 = n27596 ;
  assign y7162 = ~n27599 ;
  assign y7163 = n27600 ;
  assign y7164 = n27604 ;
  assign y7165 = ~n27607 ;
  assign y7166 = ~n27610 ;
  assign y7167 = ~n27612 ;
  assign y7168 = ~n27613 ;
  assign y7169 = ~n27618 ;
  assign y7170 = ~n27626 ;
  assign y7171 = ~n8472 ;
  assign y7172 = ~n27628 ;
  assign y7173 = n27630 ;
  assign y7174 = n27632 ;
  assign y7175 = ~1'b0 ;
  assign y7176 = ~n27635 ;
  assign y7177 = n27636 ;
  assign y7178 = n27637 ;
  assign y7179 = n27640 ;
  assign y7180 = n27644 ;
  assign y7181 = ~n27645 ;
  assign y7182 = ~n27646 ;
  assign y7183 = ~1'b0 ;
  assign y7184 = ~n27652 ;
  assign y7185 = ~n27656 ;
  assign y7186 = n27657 ;
  assign y7187 = n27658 ;
  assign y7188 = n27661 ;
  assign y7189 = n27665 ;
  assign y7190 = ~1'b0 ;
  assign y7191 = ~1'b0 ;
  assign y7192 = n27667 ;
  assign y7193 = n27672 ;
  assign y7194 = ~n27674 ;
  assign y7195 = n27676 ;
  assign y7196 = n27680 ;
  assign y7197 = ~n27682 ;
  assign y7198 = n27685 ;
  assign y7199 = ~n27686 ;
  assign y7200 = ~1'b0 ;
  assign y7201 = n27688 ;
  assign y7202 = ~n27691 ;
  assign y7203 = n27697 ;
  assign y7204 = ~n27701 ;
  assign y7205 = ~n27704 ;
  assign y7206 = ~n27705 ;
  assign y7207 = n27706 ;
  assign y7208 = ~1'b0 ;
  assign y7209 = ~n27712 ;
  assign y7210 = n27715 ;
  assign y7211 = n27716 ;
  assign y7212 = ~n27717 ;
  assign y7213 = n27718 ;
  assign y7214 = n27719 ;
  assign y7215 = n27720 ;
  assign y7216 = ~n27724 ;
  assign y7217 = ~n27726 ;
  assign y7218 = ~n27728 ;
  assign y7219 = ~n27732 ;
  assign y7220 = n27734 ;
  assign y7221 = n27736 ;
  assign y7222 = n27737 ;
  assign y7223 = ~n27741 ;
  assign y7224 = n27746 ;
  assign y7225 = ~n27748 ;
  assign y7226 = ~n27753 ;
  assign y7227 = ~1'b0 ;
  assign y7228 = n27754 ;
  assign y7229 = ~n27756 ;
  assign y7230 = ~n27758 ;
  assign y7231 = n27761 ;
  assign y7232 = ~n27764 ;
  assign y7233 = n27766 ;
  assign y7234 = ~1'b0 ;
  assign y7235 = ~n27772 ;
  assign y7236 = n27773 ;
  assign y7237 = ~n27774 ;
  assign y7238 = ~n27775 ;
  assign y7239 = ~n27776 ;
  assign y7240 = n27777 ;
  assign y7241 = n27779 ;
  assign y7242 = ~n27780 ;
  assign y7243 = ~n27782 ;
  assign y7244 = n27783 ;
  assign y7245 = n27787 ;
  assign y7246 = ~n27790 ;
  assign y7247 = ~1'b0 ;
  assign y7248 = n27791 ;
  assign y7249 = ~n27795 ;
  assign y7250 = ~n27796 ;
  assign y7251 = ~n27802 ;
  assign y7252 = n27803 ;
  assign y7253 = ~n27804 ;
  assign y7254 = ~n27806 ;
  assign y7255 = ~n27808 ;
  assign y7256 = n27811 ;
  assign y7257 = n27813 ;
  assign y7258 = n27815 ;
  assign y7259 = n27817 ;
  assign y7260 = ~n27820 ;
  assign y7261 = n27824 ;
  assign y7262 = n27825 ;
  assign y7263 = ~n27827 ;
  assign y7264 = ~n27831 ;
  assign y7265 = ~n27834 ;
  assign y7266 = ~n27836 ;
  assign y7267 = n27837 ;
  assign y7268 = ~n27843 ;
  assign y7269 = ~n27844 ;
  assign y7270 = ~n27845 ;
  assign y7271 = n27847 ;
  assign y7272 = n27853 ;
  assign y7273 = ~n27856 ;
  assign y7274 = n27857 ;
  assign y7275 = n27860 ;
  assign y7276 = ~n27868 ;
  assign y7277 = n27875 ;
  assign y7278 = n27876 ;
  assign y7279 = n27879 ;
  assign y7280 = n27880 ;
  assign y7281 = n27881 ;
  assign y7282 = ~n27883 ;
  assign y7283 = ~n27886 ;
  assign y7284 = n27887 ;
  assign y7285 = n27890 ;
  assign y7286 = n27896 ;
  assign y7287 = ~n27899 ;
  assign y7288 = n27900 ;
  assign y7289 = ~n27902 ;
  assign y7290 = ~n27906 ;
  assign y7291 = ~n27916 ;
  assign y7292 = n27918 ;
  assign y7293 = ~n27919 ;
  assign y7294 = n27920 ;
  assign y7295 = n27921 ;
  assign y7296 = ~n27924 ;
  assign y7297 = n27925 ;
  assign y7298 = n27927 ;
  assign y7299 = ~n27929 ;
  assign y7300 = ~n27930 ;
  assign y7301 = n27931 ;
  assign y7302 = n27935 ;
  assign y7303 = n27936 ;
  assign y7304 = n27938 ;
  assign y7305 = n27943 ;
  assign y7306 = ~n27945 ;
  assign y7307 = n27946 ;
  assign y7308 = ~n27950 ;
  assign y7309 = ~n27956 ;
  assign y7310 = n27957 ;
  assign y7311 = n27958 ;
  assign y7312 = n27959 ;
  assign y7313 = n27963 ;
  assign y7314 = n27965 ;
  assign y7315 = ~n27967 ;
  assign y7316 = ~n27971 ;
  assign y7317 = ~1'b0 ;
  assign y7318 = n27974 ;
  assign y7319 = n27975 ;
  assign y7320 = ~n27977 ;
  assign y7321 = ~n27980 ;
  assign y7322 = ~n27981 ;
  assign y7323 = ~n27986 ;
  assign y7324 = ~n27987 ;
  assign y7325 = ~n27988 ;
  assign y7326 = ~1'b0 ;
  assign y7327 = ~n27990 ;
  assign y7328 = n27991 ;
  assign y7329 = n27992 ;
  assign y7330 = n27993 ;
  assign y7331 = n27994 ;
  assign y7332 = n27995 ;
  assign y7333 = n27996 ;
  assign y7334 = ~n28001 ;
  assign y7335 = ~n28003 ;
  assign y7336 = ~n28006 ;
  assign y7337 = n28008 ;
  assign y7338 = ~n28009 ;
  assign y7339 = n28011 ;
  assign y7340 = n28012 ;
  assign y7341 = ~n28013 ;
  assign y7342 = ~n28014 ;
  assign y7343 = n28015 ;
  assign y7344 = n28020 ;
  assign y7345 = ~n28028 ;
  assign y7346 = ~n28030 ;
  assign y7347 = ~n28034 ;
  assign y7348 = ~n28035 ;
  assign y7349 = n28036 ;
  assign y7350 = ~n28037 ;
  assign y7351 = ~n28039 ;
  assign y7352 = ~n28040 ;
  assign y7353 = ~n28043 ;
  assign y7354 = n28054 ;
  assign y7355 = ~n28055 ;
  assign y7356 = n28058 ;
  assign y7357 = ~n28060 ;
  assign y7358 = n28064 ;
  assign y7359 = n28065 ;
  assign y7360 = ~n28071 ;
  assign y7361 = n28073 ;
  assign y7362 = n28077 ;
  assign y7363 = ~n28078 ;
  assign y7364 = ~n28080 ;
  assign y7365 = ~n28085 ;
  assign y7366 = ~1'b0 ;
  assign y7367 = ~1'b0 ;
  assign y7368 = ~n28086 ;
  assign y7369 = n28087 ;
  assign y7370 = ~n28089 ;
  assign y7371 = ~n28090 ;
  assign y7372 = n28093 ;
  assign y7373 = ~n28097 ;
  assign y7374 = ~n28098 ;
  assign y7375 = n28101 ;
  assign y7376 = ~n28103 ;
  assign y7377 = ~n28105 ;
  assign y7378 = n28108 ;
  assign y7379 = ~n28109 ;
  assign y7380 = n28110 ;
  assign y7381 = n28112 ;
  assign y7382 = ~n28113 ;
  assign y7383 = n28119 ;
  assign y7384 = n28120 ;
  assign y7385 = ~n28124 ;
  assign y7386 = ~n28126 ;
  assign y7387 = ~n28129 ;
  assign y7388 = ~n28133 ;
  assign y7389 = n28138 ;
  assign y7390 = n28139 ;
  assign y7391 = ~n28142 ;
  assign y7392 = n28143 ;
  assign y7393 = ~n28144 ;
  assign y7394 = ~n28146 ;
  assign y7395 = ~1'b0 ;
  assign y7396 = ~1'b0 ;
  assign y7397 = ~n28147 ;
  assign y7398 = ~n28148 ;
  assign y7399 = ~n28149 ;
  assign y7400 = n28153 ;
  assign y7401 = n28155 ;
  assign y7402 = n28156 ;
  assign y7403 = n28160 ;
  assign y7404 = n28161 ;
  assign y7405 = n28166 ;
  assign y7406 = ~n28169 ;
  assign y7407 = ~n28171 ;
  assign y7408 = n28172 ;
  assign y7409 = ~n28178 ;
  assign y7410 = ~n28179 ;
  assign y7411 = ~n28181 ;
  assign y7412 = n28182 ;
  assign y7413 = ~n28186 ;
  assign y7414 = n28188 ;
  assign y7415 = n28200 ;
  assign y7416 = n28203 ;
  assign y7417 = n28204 ;
  assign y7418 = n28208 ;
  assign y7419 = ~n28210 ;
  assign y7420 = ~n28211 ;
  assign y7421 = ~n28212 ;
  assign y7422 = n28218 ;
  assign y7423 = n28221 ;
  assign y7424 = n28223 ;
  assign y7425 = ~n28226 ;
  assign y7426 = ~n28231 ;
  assign y7427 = n28234 ;
  assign y7428 = n28236 ;
  assign y7429 = ~n28237 ;
  assign y7430 = n28242 ;
  assign y7431 = ~n28246 ;
  assign y7432 = ~1'b0 ;
  assign y7433 = ~1'b0 ;
  assign y7434 = n28249 ;
  assign y7435 = ~n28252 ;
  assign y7436 = ~n28258 ;
  assign y7437 = ~n28259 ;
  assign y7438 = ~n28260 ;
  assign y7439 = n28262 ;
  assign y7440 = ~n28267 ;
  assign y7441 = ~n28268 ;
  assign y7442 = ~n28270 ;
  assign y7443 = ~1'b0 ;
  assign y7444 = ~n28274 ;
  assign y7445 = n28277 ;
  assign y7446 = ~n28283 ;
  assign y7447 = n28285 ;
  assign y7448 = n28291 ;
  assign y7449 = ~n28294 ;
  assign y7450 = n28296 ;
  assign y7451 = ~n28297 ;
  assign y7452 = ~n28298 ;
  assign y7453 = ~1'b0 ;
  assign y7454 = n28299 ;
  assign y7455 = ~n28300 ;
  assign y7456 = ~n28307 ;
  assign y7457 = ~n28309 ;
  assign y7458 = ~1'b0 ;
  assign y7459 = ~n28310 ;
  assign y7460 = n28311 ;
  assign y7461 = n28313 ;
  assign y7462 = n28316 ;
  assign y7463 = n28317 ;
  assign y7464 = n28321 ;
  assign y7465 = n28324 ;
  assign y7466 = n28327 ;
  assign y7467 = n28328 ;
  assign y7468 = n28330 ;
  assign y7469 = ~n28332 ;
  assign y7470 = n28333 ;
  assign y7471 = ~1'b0 ;
  assign y7472 = n28337 ;
  assign y7473 = n28338 ;
  assign y7474 = n28339 ;
  assign y7475 = n28340 ;
  assign y7476 = n28344 ;
  assign y7477 = n28348 ;
  assign y7478 = ~n28350 ;
  assign y7479 = ~n28355 ;
  assign y7480 = n28356 ;
  assign y7481 = n28361 ;
  assign y7482 = ~n28364 ;
  assign y7483 = ~n28370 ;
  assign y7484 = n28372 ;
  assign y7485 = ~n28375 ;
  assign y7486 = ~n28382 ;
  assign y7487 = n28383 ;
  assign y7488 = n28384 ;
  assign y7489 = ~1'b0 ;
  assign y7490 = ~n28386 ;
  assign y7491 = n28387 ;
  assign y7492 = ~n28388 ;
  assign y7493 = ~n28389 ;
  assign y7494 = n28392 ;
  assign y7495 = ~n28394 ;
  assign y7496 = ~1'b0 ;
  assign y7497 = n28395 ;
  assign y7498 = ~n28398 ;
  assign y7499 = n28400 ;
  assign y7500 = ~n28402 ;
  assign y7501 = ~n28403 ;
  assign y7502 = ~n28408 ;
  assign y7503 = n28410 ;
  assign y7504 = ~n28412 ;
  assign y7505 = ~1'b0 ;
  assign y7506 = ~n28414 ;
  assign y7507 = n28420 ;
  assign y7508 = n28422 ;
  assign y7509 = ~n28423 ;
  assign y7510 = ~n28424 ;
  assign y7511 = ~n28431 ;
  assign y7512 = n28433 ;
  assign y7513 = n28434 ;
  assign y7514 = ~1'b0 ;
  assign y7515 = ~1'b0 ;
  assign y7516 = ~n28438 ;
  assign y7517 = n28440 ;
  assign y7518 = ~n28441 ;
  assign y7519 = n28444 ;
  assign y7520 = n28445 ;
  assign y7521 = n28446 ;
  assign y7522 = n28451 ;
  assign y7523 = ~1'b0 ;
  assign y7524 = ~n28453 ;
  assign y7525 = n28456 ;
  assign y7526 = n28458 ;
  assign y7527 = ~n28459 ;
  assign y7528 = ~n28463 ;
  assign y7529 = n28467 ;
  assign y7530 = n28468 ;
  assign y7531 = ~n28472 ;
  assign y7532 = ~1'b0 ;
  assign y7533 = n28474 ;
  assign y7534 = ~n28487 ;
  assign y7535 = ~n28489 ;
  assign y7536 = n28493 ;
  assign y7537 = n28494 ;
  assign y7538 = ~n28496 ;
  assign y7539 = ~n28497 ;
  assign y7540 = n28500 ;
  assign y7541 = n28503 ;
  assign y7542 = ~1'b0 ;
  assign y7543 = n28505 ;
  assign y7544 = n28507 ;
  assign y7545 = ~n28509 ;
  assign y7546 = n28510 ;
  assign y7547 = n28514 ;
  assign y7548 = n28518 ;
  assign y7549 = n28522 ;
  assign y7550 = ~n28523 ;
  assign y7551 = ~n28524 ;
  assign y7552 = ~n28526 ;
  assign y7553 = ~n28529 ;
  assign y7554 = n28531 ;
  assign y7555 = n28535 ;
  assign y7556 = n28536 ;
  assign y7557 = ~n28540 ;
  assign y7558 = ~n28542 ;
  assign y7559 = ~n28544 ;
  assign y7560 = ~n28551 ;
  assign y7561 = n28554 ;
  assign y7562 = ~1'b0 ;
  assign y7563 = ~1'b0 ;
  assign y7564 = ~n28555 ;
  assign y7565 = ~n28557 ;
  assign y7566 = n28559 ;
  assign y7567 = ~n28560 ;
  assign y7568 = ~n28561 ;
  assign y7569 = ~n28562 ;
  assign y7570 = n28563 ;
  assign y7571 = ~n28567 ;
  assign y7572 = ~1'b0 ;
  assign y7573 = ~n28570 ;
  assign y7574 = ~n28571 ;
  assign y7575 = n28574 ;
  assign y7576 = n28577 ;
  assign y7577 = ~n28582 ;
  assign y7578 = n28583 ;
  assign y7579 = ~n28589 ;
  assign y7580 = n28594 ;
  assign y7581 = ~n28595 ;
  assign y7582 = ~n28597 ;
  assign y7583 = n28602 ;
  assign y7584 = n28610 ;
  assign y7585 = n28611 ;
  assign y7586 = n28612 ;
  assign y7587 = ~n28618 ;
  assign y7588 = ~n28619 ;
  assign y7589 = n28620 ;
  assign y7590 = n28621 ;
  assign y7591 = n28622 ;
  assign y7592 = ~1'b0 ;
  assign y7593 = n28625 ;
  assign y7594 = ~n28626 ;
  assign y7595 = ~n28633 ;
  assign y7596 = ~n28636 ;
  assign y7597 = ~n28641 ;
  assign y7598 = ~n28642 ;
  assign y7599 = n28644 ;
  assign y7600 = n28646 ;
  assign y7601 = ~n28647 ;
  assign y7602 = ~n28648 ;
  assign y7603 = ~n28649 ;
  assign y7604 = ~n28650 ;
  assign y7605 = ~n28651 ;
  assign y7606 = n28655 ;
  assign y7607 = ~n28665 ;
  assign y7608 = n28666 ;
  assign y7609 = n28670 ;
  assign y7610 = ~n28671 ;
  assign y7611 = ~n28672 ;
  assign y7612 = ~n28673 ;
  assign y7613 = ~n28677 ;
  assign y7614 = ~n28680 ;
  assign y7615 = ~n28682 ;
  assign y7616 = ~n28684 ;
  assign y7617 = ~n28685 ;
  assign y7618 = n28686 ;
  assign y7619 = ~n28690 ;
  assign y7620 = n28691 ;
  assign y7621 = ~n28694 ;
  assign y7622 = ~n28697 ;
  assign y7623 = ~n28701 ;
  assign y7624 = ~n28704 ;
  assign y7625 = ~1'b0 ;
  assign y7626 = n28705 ;
  assign y7627 = ~n28706 ;
  assign y7628 = n28708 ;
  assign y7629 = n28709 ;
  assign y7630 = n28710 ;
  assign y7631 = n28711 ;
  assign y7632 = ~n28712 ;
  assign y7633 = n28713 ;
  assign y7634 = n28714 ;
  assign y7635 = n28718 ;
  assign y7636 = n28720 ;
  assign y7637 = ~n28726 ;
  assign y7638 = ~n28729 ;
  assign y7639 = n28731 ;
  assign y7640 = ~n28735 ;
  assign y7641 = ~n28736 ;
  assign y7642 = ~n28737 ;
  assign y7643 = ~n28738 ;
  assign y7644 = ~n28739 ;
  assign y7645 = ~n28741 ;
  assign y7646 = ~1'b0 ;
  assign y7647 = ~1'b0 ;
  assign y7648 = ~n28750 ;
  assign y7649 = ~n28752 ;
  assign y7650 = ~n28756 ;
  assign y7651 = n28757 ;
  assign y7652 = n28759 ;
  assign y7653 = ~n28760 ;
  assign y7654 = n28762 ;
  assign y7655 = n28763 ;
  assign y7656 = n28765 ;
  assign y7657 = ~n28766 ;
  assign y7658 = ~n28769 ;
  assign y7659 = ~n28770 ;
  assign y7660 = n28773 ;
  assign y7661 = n28776 ;
  assign y7662 = n28779 ;
  assign y7663 = ~n28782 ;
  assign y7664 = ~n28785 ;
  assign y7665 = ~n28789 ;
  assign y7666 = n28794 ;
  assign y7667 = n28796 ;
  assign y7668 = n28797 ;
  assign y7669 = ~n28801 ;
  assign y7670 = n28805 ;
  assign y7671 = ~n28808 ;
  assign y7672 = n28812 ;
  assign y7673 = ~n28813 ;
  assign y7674 = n28814 ;
  assign y7675 = ~n28821 ;
  assign y7676 = ~n28824 ;
  assign y7677 = ~n28825 ;
  assign y7678 = ~n28829 ;
  assign y7679 = n28831 ;
  assign y7680 = n28835 ;
  assign y7681 = ~n28836 ;
  assign y7682 = n28837 ;
  assign y7683 = n28838 ;
  assign y7684 = n28839 ;
  assign y7685 = n28840 ;
  assign y7686 = ~n28842 ;
  assign y7687 = n28845 ;
  assign y7688 = ~1'b0 ;
  assign y7689 = n28847 ;
  assign y7690 = ~n28848 ;
  assign y7691 = n28851 ;
  assign y7692 = ~n28854 ;
  assign y7693 = ~n28855 ;
  assign y7694 = n28856 ;
  assign y7695 = n28863 ;
  assign y7696 = n28864 ;
  assign y7697 = ~n28870 ;
  assign y7698 = ~n28880 ;
  assign y7699 = ~n28881 ;
  assign y7700 = ~n28882 ;
  assign y7701 = ~n28884 ;
  assign y7702 = n28889 ;
  assign y7703 = n28891 ;
  assign y7704 = ~n28894 ;
  assign y7705 = ~n28896 ;
  assign y7706 = ~n28897 ;
  assign y7707 = n28899 ;
  assign y7708 = n28904 ;
  assign y7709 = ~n28905 ;
  assign y7710 = ~n28906 ;
  assign y7711 = n28909 ;
  assign y7712 = ~n28911 ;
  assign y7713 = n28916 ;
  assign y7714 = n28917 ;
  assign y7715 = n28918 ;
  assign y7716 = ~n28919 ;
  assign y7717 = n28922 ;
  assign y7718 = ~n28927 ;
  assign y7719 = ~n28931 ;
  assign y7720 = n28933 ;
  assign y7721 = ~n28936 ;
  assign y7722 = n28938 ;
  assign y7723 = ~n28941 ;
  assign y7724 = n28942 ;
  assign y7725 = ~n28943 ;
  assign y7726 = n28948 ;
  assign y7727 = ~n28949 ;
  assign y7728 = ~n28951 ;
  assign y7729 = ~n28956 ;
  assign y7730 = ~n28960 ;
  assign y7731 = ~n28972 ;
  assign y7732 = n28973 ;
  assign y7733 = ~n28977 ;
  assign y7734 = ~n28978 ;
  assign y7735 = ~n28979 ;
  assign y7736 = n28981 ;
  assign y7737 = ~1'b0 ;
  assign y7738 = ~n28983 ;
  assign y7739 = n28986 ;
  assign y7740 = n28987 ;
  assign y7741 = ~n28989 ;
  assign y7742 = ~n28991 ;
  assign y7743 = n28995 ;
  assign y7744 = n28997 ;
  assign y7745 = n29001 ;
  assign y7746 = ~n29002 ;
  assign y7747 = n29003 ;
  assign y7748 = n29004 ;
  assign y7749 = n29005 ;
  assign y7750 = n29006 ;
  assign y7751 = ~n29007 ;
  assign y7752 = n29009 ;
  assign y7753 = n29013 ;
  assign y7754 = n29014 ;
  assign y7755 = ~n29015 ;
  assign y7756 = ~n29018 ;
  assign y7757 = n29019 ;
  assign y7758 = ~n29028 ;
  assign y7759 = n29030 ;
  assign y7760 = ~n29032 ;
  assign y7761 = n29033 ;
  assign y7762 = ~n29039 ;
  assign y7763 = ~n29041 ;
  assign y7764 = ~n29042 ;
  assign y7765 = ~n29043 ;
  assign y7766 = ~n29044 ;
  assign y7767 = n29045 ;
  assign y7768 = ~n29046 ;
  assign y7769 = n29048 ;
  assign y7770 = n29051 ;
  assign y7771 = n29054 ;
  assign y7772 = n29056 ;
  assign y7773 = n29058 ;
  assign y7774 = ~n29060 ;
  assign y7775 = ~n29061 ;
  assign y7776 = ~n29063 ;
  assign y7777 = ~n29068 ;
  assign y7778 = n29073 ;
  assign y7779 = n29076 ;
  assign y7780 = n29077 ;
  assign y7781 = ~n29080 ;
  assign y7782 = n29082 ;
  assign y7783 = n29087 ;
  assign y7784 = ~n29088 ;
  assign y7785 = n29089 ;
  assign y7786 = ~n29091 ;
  assign y7787 = ~n29092 ;
  assign y7788 = ~n29093 ;
  assign y7789 = ~1'b0 ;
  assign y7790 = ~1'b0 ;
  assign y7791 = ~n29097 ;
  assign y7792 = ~n29100 ;
  assign y7793 = ~n29101 ;
  assign y7794 = n29102 ;
  assign y7795 = ~n29103 ;
  assign y7796 = ~n29109 ;
  assign y7797 = ~n29112 ;
  assign y7798 = n29118 ;
  assign y7799 = n29120 ;
  assign y7800 = ~n29127 ;
  assign y7801 = ~n29130 ;
  assign y7802 = n29131 ;
  assign y7803 = n29134 ;
  assign y7804 = n29135 ;
  assign y7805 = n29136 ;
  assign y7806 = ~n29138 ;
  assign y7807 = n29140 ;
  assign y7808 = n29141 ;
  assign y7809 = n29142 ;
  assign y7810 = n29144 ;
  assign y7811 = ~1'b0 ;
  assign y7812 = n29145 ;
  assign y7813 = ~n29146 ;
  assign y7814 = n29149 ;
  assign y7815 = n29151 ;
  assign y7816 = ~n29156 ;
  assign y7817 = ~n29158 ;
  assign y7818 = ~n29162 ;
  assign y7819 = ~n29163 ;
  assign y7820 = ~n29166 ;
  assign y7821 = n29168 ;
  assign y7822 = n29169 ;
  assign y7823 = n29171 ;
  assign y7824 = ~n29177 ;
  assign y7825 = n29180 ;
  assign y7826 = n29181 ;
  assign y7827 = ~n29182 ;
  assign y7828 = ~n29184 ;
  assign y7829 = n29187 ;
  assign y7830 = n29198 ;
  assign y7831 = ~1'b0 ;
  assign y7832 = n29199 ;
  assign y7833 = n29204 ;
  assign y7834 = n29209 ;
  assign y7835 = n29212 ;
  assign y7836 = n29214 ;
  assign y7837 = n29215 ;
  assign y7838 = n29219 ;
  assign y7839 = n29220 ;
  assign y7840 = n29222 ;
  assign y7841 = n29224 ;
  assign y7842 = ~n29228 ;
  assign y7843 = n29230 ;
  assign y7844 = ~n29232 ;
  assign y7845 = n29235 ;
  assign y7846 = ~n29236 ;
  assign y7847 = ~n29237 ;
  assign y7848 = n29247 ;
  assign y7849 = ~n29248 ;
  assign y7850 = ~n29251 ;
  assign y7851 = n29257 ;
  assign y7852 = ~n29263 ;
  assign y7853 = ~n29265 ;
  assign y7854 = ~n29267 ;
  assign y7855 = ~n29269 ;
  assign y7856 = n29273 ;
  assign y7857 = ~n29274 ;
  assign y7858 = ~n29278 ;
  assign y7859 = ~1'b0 ;
  assign y7860 = ~n29279 ;
  assign y7861 = ~n29291 ;
  assign y7862 = ~n29293 ;
  assign y7863 = n29298 ;
  assign y7864 = n29303 ;
  assign y7865 = ~n29304 ;
  assign y7866 = ~n29308 ;
  assign y7867 = ~n29310 ;
  assign y7868 = n29314 ;
  assign y7869 = ~1'b0 ;
  assign y7870 = ~n29316 ;
  assign y7871 = n29317 ;
  assign y7872 = ~n29319 ;
  assign y7873 = n29321 ;
  assign y7874 = n29322 ;
  assign y7875 = n29326 ;
  assign y7876 = n29328 ;
  assign y7877 = n29329 ;
  assign y7878 = ~n29333 ;
  assign y7879 = n29335 ;
  assign y7880 = ~1'b0 ;
  assign y7881 = ~n29336 ;
  assign y7882 = n29337 ;
  assign y7883 = n29339 ;
  assign y7884 = n29341 ;
  assign y7885 = n29345 ;
  assign y7886 = n29347 ;
  assign y7887 = ~n29350 ;
  assign y7888 = n29356 ;
  assign y7889 = n29358 ;
  assign y7890 = n29360 ;
  assign y7891 = ~n29362 ;
  assign y7892 = n29363 ;
  assign y7893 = ~n29365 ;
  assign y7894 = n29376 ;
  assign y7895 = ~n29382 ;
  assign y7896 = n29383 ;
  assign y7897 = ~n29386 ;
  assign y7898 = n29388 ;
  assign y7899 = ~n29392 ;
  assign y7900 = n29396 ;
  assign y7901 = n29398 ;
  assign y7902 = ~n29399 ;
  assign y7903 = ~n29401 ;
  assign y7904 = n29403 ;
  assign y7905 = n29405 ;
  assign y7906 = ~n29409 ;
  assign y7907 = n29411 ;
  assign y7908 = ~n29413 ;
  assign y7909 = ~n29415 ;
  assign y7910 = n29418 ;
  assign y7911 = n29422 ;
  assign y7912 = ~n29425 ;
  assign y7913 = n29428 ;
  assign y7914 = ~n29436 ;
  assign y7915 = n29443 ;
  assign y7916 = ~n29445 ;
  assign y7917 = n29447 ;
  assign y7918 = ~n29448 ;
  assign y7919 = ~n29451 ;
  assign y7920 = n29454 ;
  assign y7921 = n29456 ;
  assign y7922 = n26633 ;
  assign y7923 = n29457 ;
  assign y7924 = n29461 ;
  assign y7925 = ~n29463 ;
  assign y7926 = n29465 ;
  assign y7927 = ~n29468 ;
  assign y7928 = n29469 ;
  assign y7929 = ~n29471 ;
  assign y7930 = ~1'b0 ;
  assign y7931 = n29472 ;
  assign y7932 = ~n29475 ;
  assign y7933 = n29477 ;
  assign y7934 = n29478 ;
  assign y7935 = n29479 ;
  assign y7936 = n29483 ;
  assign y7937 = n29486 ;
  assign y7938 = n29488 ;
  assign y7939 = ~n29491 ;
  assign y7940 = n29493 ;
  assign y7941 = n29495 ;
  assign y7942 = ~n29496 ;
  assign y7943 = ~n29499 ;
  assign y7944 = n29500 ;
  assign y7945 = n29503 ;
  assign y7946 = n29504 ;
  assign y7947 = ~n29506 ;
  assign y7948 = ~n29510 ;
  assign y7949 = n29512 ;
  assign y7950 = ~1'b0 ;
  assign y7951 = n29514 ;
  assign y7952 = n29520 ;
  assign y7953 = n29521 ;
  assign y7954 = n29524 ;
  assign y7955 = n29526 ;
  assign y7956 = ~n29529 ;
  assign y7957 = n29530 ;
  assign y7958 = n29533 ;
  assign y7959 = n29536 ;
  assign y7960 = n29542 ;
  assign y7961 = n29545 ;
  assign y7962 = ~1'b0 ;
  assign y7963 = n29546 ;
  assign y7964 = ~n29550 ;
  assign y7965 = ~n29551 ;
  assign y7966 = ~n29552 ;
  assign y7967 = n29553 ;
  assign y7968 = n29554 ;
  assign y7969 = n29555 ;
  assign y7970 = n29556 ;
  assign y7971 = n29557 ;
  assign y7972 = n29560 ;
  assign y7973 = n29563 ;
  assign y7974 = n29565 ;
  assign y7975 = ~n29568 ;
  assign y7976 = ~n29570 ;
  assign y7977 = n29571 ;
  assign y7978 = n29575 ;
  assign y7979 = n29576 ;
  assign y7980 = n29578 ;
  assign y7981 = ~n29581 ;
  assign y7982 = ~n29583 ;
  assign y7983 = ~1'b0 ;
  assign y7984 = ~n29586 ;
  assign y7985 = ~n29587 ;
  assign y7986 = n29589 ;
  assign y7987 = n29596 ;
  assign y7988 = ~n29598 ;
  assign y7989 = ~n29601 ;
  assign y7990 = ~1'b0 ;
  assign y7991 = ~1'b0 ;
  assign y7992 = ~n29603 ;
  assign y7993 = ~n29606 ;
  assign y7994 = n29612 ;
  assign y7995 = n29614 ;
  assign y7996 = n29615 ;
  assign y7997 = n29623 ;
  assign y7998 = n29629 ;
  assign y7999 = n29631 ;
  assign y8000 = n29632 ;
  assign y8001 = n29637 ;
  assign y8002 = n29639 ;
  assign y8003 = ~n29646 ;
  assign y8004 = n29648 ;
  assign y8005 = n29655 ;
  assign y8006 = ~n29658 ;
  assign y8007 = ~n29660 ;
  assign y8008 = n29661 ;
  assign y8009 = n29664 ;
  assign y8010 = n29665 ;
  assign y8011 = ~n29669 ;
  assign y8012 = ~n29675 ;
  assign y8013 = ~n29682 ;
  assign y8014 = ~n29685 ;
  assign y8015 = ~n29686 ;
  assign y8016 = n29687 ;
  assign y8017 = ~n29688 ;
  assign y8018 = n29689 ;
  assign y8019 = ~n29691 ;
  assign y8020 = n29693 ;
  assign y8021 = ~1'b0 ;
  assign y8022 = ~n29695 ;
  assign y8023 = n29697 ;
  assign y8024 = ~n29698 ;
  assign y8025 = n29703 ;
  assign y8026 = ~n29705 ;
  assign y8027 = n29709 ;
  assign y8028 = n29711 ;
  assign y8029 = ~n29713 ;
  assign y8030 = ~n29715 ;
  assign y8031 = n29716 ;
  assign y8032 = n29723 ;
  assign y8033 = ~n29724 ;
  assign y8034 = n29726 ;
  assign y8035 = ~n29730 ;
  assign y8036 = n29733 ;
  assign y8037 = ~n29734 ;
  assign y8038 = n29741 ;
  assign y8039 = n29745 ;
  assign y8040 = ~1'b0 ;
  assign y8041 = ~n29747 ;
  assign y8042 = ~n29748 ;
  assign y8043 = n29749 ;
  assign y8044 = ~n29750 ;
  assign y8045 = n29753 ;
  assign y8046 = ~n29756 ;
  assign y8047 = n29758 ;
  assign y8048 = ~n29760 ;
  assign y8049 = ~n29770 ;
  assign y8050 = ~1'b0 ;
  assign y8051 = ~n29772 ;
  assign y8052 = n29773 ;
  assign y8053 = n29774 ;
  assign y8054 = n29775 ;
  assign y8055 = n29778 ;
  assign y8056 = n29779 ;
  assign y8057 = n29780 ;
  assign y8058 = n29781 ;
  assign y8059 = n29785 ;
  assign y8060 = ~n29789 ;
  assign y8061 = n29792 ;
  assign y8062 = ~n29795 ;
  assign y8063 = ~n29796 ;
  assign y8064 = n29797 ;
  assign y8065 = ~n29802 ;
  assign y8066 = ~n29803 ;
  assign y8067 = ~n29806 ;
  assign y8068 = ~n29807 ;
  assign y8069 = ~n29809 ;
  assign y8070 = ~1'b0 ;
  assign y8071 = n29811 ;
  assign y8072 = n29814 ;
  assign y8073 = ~n29815 ;
  assign y8074 = n29816 ;
  assign y8075 = n29817 ;
  assign y8076 = n29818 ;
  assign y8077 = n29820 ;
  assign y8078 = ~n29822 ;
  assign y8079 = n29825 ;
  assign y8080 = n29826 ;
  assign y8081 = ~n29827 ;
  assign y8082 = n29834 ;
  assign y8083 = n29835 ;
  assign y8084 = n29842 ;
  assign y8085 = n29844 ;
  assign y8086 = n29845 ;
  assign y8087 = n29847 ;
  assign y8088 = n29850 ;
  assign y8089 = ~n29854 ;
  assign y8090 = n29859 ;
  assign y8091 = n29860 ;
  assign y8092 = ~n29862 ;
  assign y8093 = n29867 ;
  assign y8094 = ~n29868 ;
  assign y8095 = ~n29870 ;
  assign y8096 = n29873 ;
  assign y8097 = ~1'b0 ;
  assign y8098 = n29877 ;
  assign y8099 = n29880 ;
  assign y8100 = ~n29882 ;
  assign y8101 = ~n29885 ;
  assign y8102 = n29886 ;
  assign y8103 = ~n29887 ;
  assign y8104 = ~n29888 ;
  assign y8105 = n29890 ;
  assign y8106 = n29893 ;
  assign y8107 = n29895 ;
  assign y8108 = n29898 ;
  assign y8109 = ~n29899 ;
  assign y8110 = n29901 ;
  assign y8111 = n29903 ;
  assign y8112 = ~n29904 ;
  assign y8113 = ~n29906 ;
  assign y8114 = ~n29912 ;
  assign y8115 = ~n29913 ;
  assign y8116 = n29918 ;
  assign y8117 = n29919 ;
  assign y8118 = ~1'b0 ;
  assign y8119 = ~n29926 ;
  assign y8120 = ~n29928 ;
  assign y8121 = n29931 ;
  assign y8122 = ~n29935 ;
  assign y8123 = ~n29940 ;
  assign y8124 = n29941 ;
  assign y8125 = ~n29942 ;
  assign y8126 = n29944 ;
  assign y8127 = n29948 ;
  assign y8128 = n29952 ;
  assign y8129 = ~n29953 ;
  assign y8130 = ~n29956 ;
  assign y8131 = ~n29957 ;
  assign y8132 = ~n29958 ;
  assign y8133 = n29959 ;
  assign y8134 = n29960 ;
  assign y8135 = ~n29962 ;
  assign y8136 = n29965 ;
  assign y8137 = ~n29969 ;
  assign y8138 = ~1'b0 ;
  assign y8139 = ~n29974 ;
  assign y8140 = n29975 ;
  assign y8141 = n29978 ;
  assign y8142 = ~n29981 ;
  assign y8143 = n29986 ;
  assign y8144 = ~n29993 ;
  assign y8145 = ~n29997 ;
  assign y8146 = n30000 ;
  assign y8147 = ~n30003 ;
  assign y8148 = ~1'b0 ;
  assign y8149 = ~1'b0 ;
  assign y8150 = ~n30005 ;
  assign y8151 = ~n30006 ;
  assign y8152 = n30009 ;
  assign y8153 = n30013 ;
  assign y8154 = ~n30017 ;
  assign y8155 = n30023 ;
  assign y8156 = n30024 ;
  assign y8157 = n30032 ;
  assign y8158 = n30037 ;
  assign y8159 = n30039 ;
  assign y8160 = ~n30041 ;
  assign y8161 = n30048 ;
  assign y8162 = ~n30049 ;
  assign y8163 = ~n30050 ;
  assign y8164 = ~n30051 ;
  assign y8165 = n30053 ;
  assign y8166 = ~n30057 ;
  assign y8167 = n30058 ;
  assign y8168 = ~n30060 ;
  assign y8169 = ~1'b0 ;
  assign y8170 = ~n30061 ;
  assign y8171 = ~n30062 ;
  assign y8172 = ~n30063 ;
  assign y8173 = ~n30068 ;
  assign y8174 = n30070 ;
  assign y8175 = n30071 ;
  assign y8176 = n30072 ;
  assign y8177 = n30076 ;
  assign y8178 = n30078 ;
  assign y8179 = ~1'b0 ;
  assign y8180 = ~n30079 ;
  assign y8181 = ~n30082 ;
  assign y8182 = ~n30087 ;
  assign y8183 = ~n30088 ;
  assign y8184 = ~n30089 ;
  assign y8185 = n30091 ;
  assign y8186 = n30092 ;
  assign y8187 = ~n30093 ;
  assign y8188 = n30094 ;
  assign y8189 = ~1'b0 ;
  assign y8190 = ~n30098 ;
  assign y8191 = ~n30099 ;
  assign y8192 = ~n30100 ;
  assign y8193 = n30102 ;
  assign y8194 = n30103 ;
  assign y8195 = n30108 ;
  assign y8196 = ~n30109 ;
  assign y8197 = ~n30113 ;
  assign y8198 = ~n30114 ;
  assign y8199 = ~n30115 ;
  assign y8200 = ~1'b0 ;
  assign y8201 = n30116 ;
  assign y8202 = ~n30117 ;
  assign y8203 = n30120 ;
  assign y8204 = ~n30122 ;
  assign y8205 = n30123 ;
  assign y8206 = n30125 ;
  assign y8207 = ~n30128 ;
  assign y8208 = n30130 ;
  assign y8209 = ~n30131 ;
  assign y8210 = n30137 ;
  assign y8211 = ~n30139 ;
  assign y8212 = ~n30140 ;
  assign y8213 = ~n30141 ;
  assign y8214 = ~n30142 ;
  assign y8215 = ~n30144 ;
  assign y8216 = n30147 ;
  assign y8217 = n30151 ;
  assign y8218 = ~n30154 ;
  assign y8219 = n30156 ;
  assign y8220 = ~n30160 ;
  assign y8221 = ~n30162 ;
  assign y8222 = ~n30164 ;
  assign y8223 = ~n30165 ;
  assign y8224 = n30166 ;
  assign y8225 = ~n30168 ;
  assign y8226 = ~n30170 ;
  assign y8227 = ~n30173 ;
  assign y8228 = n30175 ;
  assign y8229 = n30180 ;
  assign y8230 = ~n30181 ;
  assign y8231 = ~n30182 ;
  assign y8232 = ~n30185 ;
  assign y8233 = ~1'b0 ;
  assign y8234 = ~n30188 ;
  assign y8235 = ~n30190 ;
  assign y8236 = n30193 ;
  assign y8237 = ~n30199 ;
  assign y8238 = n30201 ;
  assign y8239 = ~n30204 ;
  assign y8240 = ~n30213 ;
  assign y8241 = n30214 ;
  assign y8242 = ~1'b0 ;
  assign y8243 = n30215 ;
  assign y8244 = n30216 ;
  assign y8245 = n30218 ;
  assign y8246 = n30223 ;
  assign y8247 = ~n30227 ;
  assign y8248 = n30231 ;
  assign y8249 = ~n30233 ;
  assign y8250 = ~n30236 ;
  assign y8251 = n30237 ;
  assign y8252 = ~n30239 ;
  assign y8253 = ~n30241 ;
  assign y8254 = ~n30242 ;
  assign y8255 = ~n30245 ;
  assign y8256 = n30246 ;
  assign y8257 = ~n30248 ;
  assign y8258 = n30250 ;
  assign y8259 = ~n30251 ;
  assign y8260 = n30252 ;
  assign y8261 = ~n30254 ;
  assign y8262 = n30256 ;
  assign y8263 = ~1'b0 ;
  assign y8264 = ~n30261 ;
  assign y8265 = n30266 ;
  assign y8266 = ~n30267 ;
  assign y8267 = n30268 ;
  assign y8268 = ~n30270 ;
  assign y8269 = ~n30271 ;
  assign y8270 = n30272 ;
  assign y8271 = n30274 ;
  assign y8272 = ~n30276 ;
  assign y8273 = n30280 ;
  assign y8274 = ~n30285 ;
  assign y8275 = ~n30286 ;
  assign y8276 = n30288 ;
  assign y8277 = n30291 ;
  assign y8278 = n30294 ;
  assign y8279 = n30295 ;
  assign y8280 = ~n30297 ;
  assign y8281 = ~n30301 ;
  assign y8282 = n30303 ;
  assign y8283 = n30309 ;
  assign y8284 = ~n30310 ;
  assign y8285 = ~n30311 ;
  assign y8286 = n30312 ;
  assign y8287 = n30313 ;
  assign y8288 = ~n30316 ;
  assign y8289 = n30317 ;
  assign y8290 = n30318 ;
  assign y8291 = n30320 ;
  assign y8292 = n30330 ;
  assign y8293 = n30332 ;
  assign y8294 = ~n30334 ;
  assign y8295 = ~n30338 ;
  assign y8296 = ~n30339 ;
  assign y8297 = ~n30341 ;
  assign y8298 = ~n30342 ;
  assign y8299 = ~n30343 ;
  assign y8300 = n30346 ;
  assign y8301 = ~n30349 ;
  assign y8302 = ~n30350 ;
  assign y8303 = n30358 ;
  assign y8304 = ~n30363 ;
  assign y8305 = n30365 ;
  assign y8306 = n30366 ;
  assign y8307 = n30369 ;
  assign y8308 = ~n30370 ;
  assign y8309 = n30373 ;
  assign y8310 = ~n30374 ;
  assign y8311 = ~n30375 ;
  assign y8312 = n30377 ;
  assign y8313 = n30382 ;
  assign y8314 = ~1'b0 ;
  assign y8315 = ~1'b0 ;
  assign y8316 = n30387 ;
  assign y8317 = n30388 ;
  assign y8318 = n30395 ;
  assign y8319 = n30396 ;
  assign y8320 = ~n30399 ;
  assign y8321 = ~n30405 ;
  assign y8322 = n30407 ;
  assign y8323 = n30408 ;
  assign y8324 = ~n30409 ;
  assign y8325 = ~n30412 ;
  assign y8326 = ~1'b0 ;
  assign y8327 = ~n30413 ;
  assign y8328 = n30414 ;
  assign y8329 = n30415 ;
  assign y8330 = ~n30416 ;
  assign y8331 = ~n30417 ;
  assign y8332 = ~n30422 ;
  assign y8333 = ~n30423 ;
  assign y8334 = n30424 ;
  assign y8335 = ~1'b0 ;
  assign y8336 = n30426 ;
  assign y8337 = ~n30427 ;
  assign y8338 = ~n30429 ;
  assign y8339 = n30430 ;
  assign y8340 = n30431 ;
  assign y8341 = ~n30433 ;
  assign y8342 = n30434 ;
  assign y8343 = ~n30437 ;
  assign y8344 = n30439 ;
  assign y8345 = ~n30442 ;
  assign y8346 = ~n30445 ;
  assign y8347 = n30448 ;
  assign y8348 = ~n30450 ;
  assign y8349 = n30451 ;
  assign y8350 = ~n30452 ;
  assign y8351 = ~n30453 ;
  assign y8352 = n30455 ;
  assign y8353 = ~n30457 ;
  assign y8354 = ~n30459 ;
  assign y8355 = ~n30460 ;
  assign y8356 = n30463 ;
  assign y8357 = ~1'b0 ;
  assign y8358 = ~n30465 ;
  assign y8359 = n30469 ;
  assign y8360 = n30470 ;
  assign y8361 = ~n30472 ;
  assign y8362 = ~n30479 ;
  assign y8363 = ~n30480 ;
  assign y8364 = ~n30481 ;
  assign y8365 = n30483 ;
  assign y8366 = ~n30484 ;
  assign y8367 = ~n30487 ;
  assign y8368 = ~n30493 ;
  assign y8369 = n30494 ;
  assign y8370 = n30496 ;
  assign y8371 = ~n30500 ;
  assign y8372 = ~n30501 ;
  assign y8373 = ~n30503 ;
  assign y8374 = n30504 ;
  assign y8375 = n30505 ;
  assign y8376 = ~n30506 ;
  assign y8377 = ~n30507 ;
  assign y8378 = ~n30515 ;
  assign y8379 = n30517 ;
  assign y8380 = ~n30518 ;
  assign y8381 = n30519 ;
  assign y8382 = n30520 ;
  assign y8383 = n30521 ;
  assign y8384 = ~n30522 ;
  assign y8385 = n30526 ;
  assign y8386 = ~n30529 ;
  assign y8387 = ~n30530 ;
  assign y8388 = n30531 ;
  assign y8389 = ~n30534 ;
  assign y8390 = n30536 ;
  assign y8391 = n30538 ;
  assign y8392 = ~n30541 ;
  assign y8393 = ~n30542 ;
  assign y8394 = n30543 ;
  assign y8395 = n30546 ;
  assign y8396 = n30547 ;
  assign y8397 = ~n30549 ;
  assign y8398 = ~n30553 ;
  assign y8399 = ~n30554 ;
  assign y8400 = n30556 ;
  assign y8401 = n30558 ;
  assign y8402 = n30563 ;
  assign y8403 = ~n30566 ;
  assign y8404 = n30568 ;
  assign y8405 = n30570 ;
  assign y8406 = n30571 ;
  assign y8407 = n30575 ;
  assign y8408 = n30576 ;
  assign y8409 = ~n30577 ;
  assign y8410 = ~n30578 ;
  assign y8411 = ~1'b0 ;
  assign y8412 = ~n30580 ;
  assign y8413 = ~n30581 ;
  assign y8414 = n30582 ;
  assign y8415 = ~n30584 ;
  assign y8416 = n30585 ;
  assign y8417 = n30589 ;
  assign y8418 = n30591 ;
  assign y8419 = ~n30592 ;
  assign y8420 = ~n30593 ;
  assign y8421 = n30595 ;
  assign y8422 = n30596 ;
  assign y8423 = n30598 ;
  assign y8424 = n30601 ;
  assign y8425 = n30602 ;
  assign y8426 = n30603 ;
  assign y8427 = n30605 ;
  assign y8428 = ~n30606 ;
  assign y8429 = n30608 ;
  assign y8430 = ~n30610 ;
  assign y8431 = n30611 ;
  assign y8432 = ~n30613 ;
  assign y8433 = n30617 ;
  assign y8434 = n30619 ;
  assign y8435 = n30623 ;
  assign y8436 = ~n30624 ;
  assign y8437 = n30625 ;
  assign y8438 = ~n30627 ;
  assign y8439 = n30630 ;
  assign y8440 = n30634 ;
  assign y8441 = ~n30644 ;
  assign y8442 = ~1'b0 ;
  assign y8443 = ~1'b0 ;
  assign y8444 = ~n30645 ;
  assign y8445 = ~n30647 ;
  assign y8446 = n30648 ;
  assign y8447 = ~n30649 ;
  assign y8448 = ~n30654 ;
  assign y8449 = ~n30656 ;
  assign y8450 = n30657 ;
  assign y8451 = n30659 ;
  assign y8452 = ~n30660 ;
  assign y8453 = n30662 ;
  assign y8454 = ~1'b0 ;
  assign y8455 = ~n30663 ;
  assign y8456 = ~n30665 ;
  assign y8457 = n30666 ;
  assign y8458 = n30669 ;
  assign y8459 = ~n30672 ;
  assign y8460 = ~n30675 ;
  assign y8461 = ~n30679 ;
  assign y8462 = ~n30682 ;
  assign y8463 = ~1'b0 ;
  assign y8464 = n30686 ;
  assign y8465 = ~n30687 ;
  assign y8466 = n30692 ;
  assign y8467 = n30697 ;
  assign y8468 = ~n30700 ;
  assign y8469 = ~n30701 ;
  assign y8470 = ~n30710 ;
  assign y8471 = n30715 ;
  assign y8472 = n30718 ;
  assign y8473 = ~n30720 ;
  assign y8474 = ~n30722 ;
  assign y8475 = n30724 ;
  assign y8476 = ~n30728 ;
  assign y8477 = ~n30729 ;
  assign y8478 = n30730 ;
  assign y8479 = n30731 ;
  assign y8480 = ~n30734 ;
  assign y8481 = ~n30736 ;
  assign y8482 = n30739 ;
  assign y8483 = n30741 ;
  assign y8484 = n30743 ;
  assign y8485 = ~n30746 ;
  assign y8486 = ~n30751 ;
  assign y8487 = ~n30753 ;
  assign y8488 = n30755 ;
  assign y8489 = n30764 ;
  assign y8490 = n30767 ;
  assign y8491 = ~n30770 ;
  assign y8492 = ~n30771 ;
  assign y8493 = ~n30773 ;
  assign y8494 = n30779 ;
  assign y8495 = ~1'b0 ;
  assign y8496 = n30781 ;
  assign y8497 = n30785 ;
  assign y8498 = n30786 ;
  assign y8499 = n30790 ;
  assign y8500 = ~n30794 ;
  assign y8501 = n30795 ;
  assign y8502 = n30796 ;
  assign y8503 = ~n30797 ;
  assign y8504 = ~n30799 ;
  assign y8505 = n30801 ;
  assign y8506 = n30803 ;
  assign y8507 = n30804 ;
  assign y8508 = ~n30806 ;
  assign y8509 = ~n30807 ;
  assign y8510 = n30808 ;
  assign y8511 = n30813 ;
  assign y8512 = ~n30816 ;
  assign y8513 = n30817 ;
  assign y8514 = ~n30818 ;
  assign y8515 = ~n30819 ;
  assign y8516 = n30824 ;
  assign y8517 = n30828 ;
  assign y8518 = ~n30836 ;
  assign y8519 = n30837 ;
  assign y8520 = n30842 ;
  assign y8521 = ~n30843 ;
  assign y8522 = ~n30846 ;
  assign y8523 = n30848 ;
  assign y8524 = n30854 ;
  assign y8525 = ~n30857 ;
  assign y8526 = n30859 ;
  assign y8527 = n30861 ;
  assign y8528 = ~n30864 ;
  assign y8529 = ~n30865 ;
  assign y8530 = ~n30867 ;
  assign y8531 = n30868 ;
  assign y8532 = ~n30869 ;
  assign y8533 = ~n30872 ;
  assign y8534 = ~n30874 ;
  assign y8535 = n30879 ;
  assign y8536 = n30883 ;
  assign y8537 = n30885 ;
  assign y8538 = ~n30886 ;
  assign y8539 = ~n30890 ;
  assign y8540 = ~n30893 ;
  assign y8541 = ~n30895 ;
  assign y8542 = ~n30897 ;
  assign y8543 = n30898 ;
  assign y8544 = n30900 ;
  assign y8545 = n30904 ;
  assign y8546 = ~n30905 ;
  assign y8547 = ~n30909 ;
  assign y8548 = ~1'b0 ;
  assign y8549 = n30911 ;
  assign y8550 = ~n30913 ;
  assign y8551 = n30915 ;
  assign y8552 = n30916 ;
  assign y8553 = ~n30917 ;
  assign y8554 = ~n30918 ;
  assign y8555 = ~n30919 ;
  assign y8556 = ~n30920 ;
  assign y8557 = ~n30921 ;
  assign y8558 = n30923 ;
  assign y8559 = n30925 ;
  assign y8560 = n30926 ;
  assign y8561 = ~n30929 ;
  assign y8562 = ~n30931 ;
  assign y8563 = ~n30932 ;
  assign y8564 = n30934 ;
  assign y8565 = n30937 ;
  assign y8566 = n30939 ;
  assign y8567 = n30942 ;
  assign y8568 = ~n30944 ;
  assign y8569 = n30946 ;
  assign y8570 = n30950 ;
  assign y8571 = n30951 ;
  assign y8572 = ~n30953 ;
  assign y8573 = ~n30954 ;
  assign y8574 = n30956 ;
  assign y8575 = ~n30957 ;
  assign y8576 = n30958 ;
  assign y8577 = ~n30959 ;
  assign y8578 = n30961 ;
  assign y8579 = ~n30962 ;
  assign y8580 = n30964 ;
  assign y8581 = ~1'b0 ;
  assign y8582 = n30968 ;
  assign y8583 = ~n30970 ;
  assign y8584 = n30971 ;
  assign y8585 = n30976 ;
  assign y8586 = n30977 ;
  assign y8587 = ~n30979 ;
  assign y8588 = ~n30982 ;
  assign y8589 = ~n30984 ;
  assign y8590 = n30985 ;
  assign y8591 = ~1'b0 ;
  assign y8592 = ~n30987 ;
  assign y8593 = n30993 ;
  assign y8594 = n30995 ;
  assign y8595 = ~n30998 ;
  assign y8596 = n31001 ;
  assign y8597 = n31004 ;
  assign y8598 = ~n31007 ;
  assign y8599 = n31009 ;
  assign y8600 = ~n31013 ;
  assign y8601 = ~n31014 ;
  assign y8602 = n31019 ;
  assign y8603 = ~1'b0 ;
  assign y8604 = ~n31020 ;
  assign y8605 = ~n31021 ;
  assign y8606 = ~n31022 ;
  assign y8607 = n31023 ;
  assign y8608 = n31024 ;
  assign y8609 = ~n31030 ;
  assign y8610 = ~n31031 ;
  assign y8611 = n31032 ;
  assign y8612 = ~n31037 ;
  assign y8613 = n31043 ;
  assign y8614 = ~n31045 ;
  assign y8615 = n31048 ;
  assign y8616 = n31049 ;
  assign y8617 = ~n31050 ;
  assign y8618 = n31052 ;
  assign y8619 = n31055 ;
  assign y8620 = n31057 ;
  assign y8621 = ~n31062 ;
  assign y8622 = ~n31064 ;
  assign y8623 = n31067 ;
  assign y8624 = ~n31069 ;
  assign y8625 = n31074 ;
  assign y8626 = n31077 ;
  assign y8627 = ~n31080 ;
  assign y8628 = n31083 ;
  assign y8629 = n31084 ;
  assign y8630 = ~n31087 ;
  assign y8631 = ~n31088 ;
  assign y8632 = n31091 ;
  assign y8633 = ~n31096 ;
  assign y8634 = ~1'b0 ;
  assign y8635 = ~n31098 ;
  assign y8636 = n31101 ;
  assign y8637 = ~n31102 ;
  assign y8638 = n31103 ;
  assign y8639 = n31107 ;
  assign y8640 = ~n31108 ;
  assign y8641 = n31109 ;
  assign y8642 = ~n31115 ;
  assign y8643 = ~1'b0 ;
  assign y8644 = ~1'b0 ;
  assign y8645 = ~n31116 ;
  assign y8646 = n31118 ;
  assign y8647 = ~n31120 ;
  assign y8648 = n31121 ;
  assign y8649 = ~n31122 ;
  assign y8650 = n31125 ;
  assign y8651 = ~n31126 ;
  assign y8652 = ~n31129 ;
  assign y8653 = ~n31131 ;
  assign y8654 = ~n31133 ;
  assign y8655 = n31136 ;
  assign y8656 = ~n31139 ;
  assign y8657 = ~n31143 ;
  assign y8658 = ~n31148 ;
  assign y8659 = ~n31150 ;
  assign y8660 = ~n31151 ;
  assign y8661 = ~n31152 ;
  assign y8662 = n31153 ;
  assign y8663 = n31155 ;
  assign y8664 = n31157 ;
  assign y8665 = ~n31159 ;
  assign y8666 = ~1'b0 ;
  assign y8667 = n31162 ;
  assign y8668 = ~n31169 ;
  assign y8669 = n31170 ;
  assign y8670 = n31179 ;
  assign y8671 = ~n31185 ;
  assign y8672 = n31186 ;
  assign y8673 = ~n31188 ;
  assign y8674 = ~n31196 ;
  assign y8675 = ~n31197 ;
  assign y8676 = n31200 ;
  assign y8677 = n31202 ;
  assign y8678 = ~n31203 ;
  assign y8679 = ~n31206 ;
  assign y8680 = n31208 ;
  assign y8681 = ~n31209 ;
  assign y8682 = ~n31212 ;
  assign y8683 = ~n31214 ;
  assign y8684 = n31217 ;
  assign y8685 = n31223 ;
  assign y8686 = n31224 ;
  assign y8687 = ~n31226 ;
  assign y8688 = n31228 ;
  assign y8689 = n31229 ;
  assign y8690 = ~n31230 ;
  assign y8691 = n31233 ;
  assign y8692 = ~n31238 ;
  assign y8693 = ~n31239 ;
  assign y8694 = ~n31241 ;
  assign y8695 = ~n31245 ;
  assign y8696 = n31250 ;
  assign y8697 = ~n31251 ;
  assign y8698 = ~1'b0 ;
  assign y8699 = ~n31256 ;
  assign y8700 = ~n31257 ;
  assign y8701 = n31259 ;
  assign y8702 = n31261 ;
  assign y8703 = n31264 ;
  assign y8704 = n31265 ;
  assign y8705 = ~n31270 ;
  assign y8706 = n31271 ;
  assign y8707 = ~n31274 ;
  assign y8708 = n31276 ;
  assign y8709 = ~1'b0 ;
  assign y8710 = n31277 ;
  assign y8711 = ~n31278 ;
  assign y8712 = n31279 ;
  assign y8713 = ~n31281 ;
  assign y8714 = n31282 ;
  assign y8715 = n31285 ;
  assign y8716 = ~n31289 ;
  assign y8717 = ~n31290 ;
  assign y8718 = ~n31293 ;
  assign y8719 = ~1'b0 ;
  assign y8720 = ~1'b0 ;
  assign y8721 = ~n31297 ;
  assign y8722 = n31300 ;
  assign y8723 = ~n31301 ;
  assign y8724 = n31302 ;
  assign y8725 = ~n31303 ;
  assign y8726 = ~n31308 ;
  assign y8727 = ~n31310 ;
  assign y8728 = n31311 ;
  assign y8729 = ~n31313 ;
  assign y8730 = ~1'b0 ;
  assign y8731 = n31316 ;
  assign y8732 = ~n31318 ;
  assign y8733 = ~n31326 ;
  assign y8734 = ~n31328 ;
  assign y8735 = n31333 ;
  assign y8736 = ~n31339 ;
  assign y8737 = ~n31341 ;
  assign y8738 = n31343 ;
  assign y8739 = n31345 ;
  assign y8740 = n31346 ;
  assign y8741 = ~1'b0 ;
  assign y8742 = n31348 ;
  assign y8743 = n31350 ;
  assign y8744 = n31353 ;
  assign y8745 = n31354 ;
  assign y8746 = n31355 ;
  assign y8747 = n31357 ;
  assign y8748 = n31359 ;
  assign y8749 = n31362 ;
  assign y8750 = n31363 ;
  assign y8751 = n31368 ;
  assign y8752 = ~1'b0 ;
  assign y8753 = ~n31370 ;
  assign y8754 = ~n31373 ;
  assign y8755 = n31375 ;
  assign y8756 = n31377 ;
  assign y8757 = n31379 ;
  assign y8758 = n31381 ;
  assign y8759 = ~n31382 ;
  assign y8760 = ~n31387 ;
  assign y8761 = ~n31388 ;
  assign y8762 = n31390 ;
  assign y8763 = n31392 ;
  assign y8764 = n31394 ;
  assign y8765 = ~n31396 ;
  assign y8766 = ~n31397 ;
  assign y8767 = ~n31403 ;
  assign y8768 = n31404 ;
  assign y8769 = ~n31405 ;
  assign y8770 = ~n31412 ;
  assign y8771 = ~n31413 ;
  assign y8772 = ~n31417 ;
  assign y8773 = ~n31422 ;
  assign y8774 = n31426 ;
  assign y8775 = ~n31427 ;
  assign y8776 = n31435 ;
  assign y8777 = ~n31436 ;
  assign y8778 = n31437 ;
  assign y8779 = n31440 ;
  assign y8780 = n31441 ;
  assign y8781 = ~n31442 ;
  assign y8782 = n31443 ;
  assign y8783 = ~n31450 ;
  assign y8784 = ~1'b0 ;
  assign y8785 = ~n31452 ;
  assign y8786 = n31458 ;
  assign y8787 = n31459 ;
  assign y8788 = n31461 ;
  assign y8789 = n31462 ;
  assign y8790 = n31466 ;
  assign y8791 = ~n31469 ;
  assign y8792 = ~n31470 ;
  assign y8793 = ~n31473 ;
  assign y8794 = n31474 ;
  assign y8795 = ~n31478 ;
  assign y8796 = ~1'b0 ;
  assign y8797 = n31479 ;
  assign y8798 = ~n31480 ;
  assign y8799 = ~n31481 ;
  assign y8800 = ~n31484 ;
  assign y8801 = ~n31487 ;
  assign y8802 = n31488 ;
  assign y8803 = n31494 ;
  assign y8804 = ~n31495 ;
  assign y8805 = ~n31496 ;
  assign y8806 = ~n31498 ;
  assign y8807 = n31501 ;
  assign y8808 = n31503 ;
  assign y8809 = ~n31508 ;
  assign y8810 = n31509 ;
  assign y8811 = ~n31512 ;
  assign y8812 = ~n31516 ;
  assign y8813 = n31517 ;
  assign y8814 = n31519 ;
  assign y8815 = ~n31523 ;
  assign y8816 = ~n31526 ;
  assign y8817 = n31528 ;
  assign y8818 = n31530 ;
  assign y8819 = ~n31531 ;
  assign y8820 = ~n31532 ;
  assign y8821 = ~n31533 ;
  assign y8822 = ~n31538 ;
  assign y8823 = n31547 ;
  assign y8824 = ~n31549 ;
  assign y8825 = ~n31550 ;
  assign y8826 = n31551 ;
  assign y8827 = ~n31552 ;
  assign y8828 = ~n31555 ;
  assign y8829 = ~1'b0 ;
  assign y8830 = ~n31556 ;
  assign y8831 = ~n31558 ;
  assign y8832 = ~n31559 ;
  assign y8833 = n31560 ;
  assign y8834 = n31562 ;
  assign y8835 = n31564 ;
  assign y8836 = n31565 ;
  assign y8837 = n31568 ;
  assign y8838 = ~n31570 ;
  assign y8839 = ~n31572 ;
  assign y8840 = ~1'b0 ;
  assign y8841 = n31573 ;
  assign y8842 = ~n31575 ;
  assign y8843 = ~n31576 ;
  assign y8844 = ~n31577 ;
  assign y8845 = n31579 ;
  assign y8846 = n31580 ;
  assign y8847 = n31581 ;
  assign y8848 = ~n31582 ;
  assign y8849 = n31583 ;
  assign y8850 = n31585 ;
  assign y8851 = ~1'b0 ;
  assign y8852 = ~n31586 ;
  assign y8853 = ~n31589 ;
  assign y8854 = n31591 ;
  assign y8855 = ~n31592 ;
  assign y8856 = ~n31595 ;
  assign y8857 = ~n31596 ;
  assign y8858 = ~n31598 ;
  assign y8859 = ~n31599 ;
  assign y8860 = n31604 ;
  assign y8861 = ~n31608 ;
  assign y8862 = n31610 ;
  assign y8863 = ~n31611 ;
  assign y8864 = ~n31613 ;
  assign y8865 = ~n31615 ;
  assign y8866 = n31617 ;
  assign y8867 = n31620 ;
  assign y8868 = n31624 ;
  assign y8869 = ~n31626 ;
  assign y8870 = ~n31627 ;
  assign y8871 = ~n31629 ;
  assign y8872 = ~1'b0 ;
  assign y8873 = ~n31631 ;
  assign y8874 = ~n31632 ;
  assign y8875 = n31633 ;
  assign y8876 = ~n31635 ;
  assign y8877 = ~n31636 ;
  assign y8878 = n31637 ;
  assign y8879 = ~n31639 ;
  assign y8880 = n31641 ;
  assign y8881 = n31643 ;
  assign y8882 = n31646 ;
  assign y8883 = ~n31649 ;
  assign y8884 = ~1'b0 ;
  assign y8885 = n31658 ;
  assign y8886 = n31659 ;
  assign y8887 = ~n31660 ;
  assign y8888 = n31661 ;
  assign y8889 = n25224 ;
  assign y8890 = ~n31662 ;
  assign y8891 = n31666 ;
  assign y8892 = ~n31667 ;
  assign y8893 = n31669 ;
  assign y8894 = ~n31671 ;
  assign y8895 = ~1'b0 ;
  assign y8896 = n31673 ;
  assign y8897 = n31675 ;
  assign y8898 = ~n31680 ;
  assign y8899 = n31682 ;
  assign y8900 = n31684 ;
  assign y8901 = n31686 ;
  assign y8902 = ~n31687 ;
  assign y8903 = ~n31688 ;
  assign y8904 = ~n31690 ;
  assign y8905 = ~1'b0 ;
  assign y8906 = ~n31692 ;
  assign y8907 = ~n31693 ;
  assign y8908 = n31694 ;
  assign y8909 = n31695 ;
  assign y8910 = ~n31696 ;
  assign y8911 = ~n31697 ;
  assign y8912 = n31701 ;
  assign y8913 = ~n31702 ;
  assign y8914 = ~n31703 ;
  assign y8915 = n31704 ;
  assign y8916 = ~1'b0 ;
  assign y8917 = n31706 ;
  assign y8918 = n31711 ;
  assign y8919 = ~n31712 ;
  assign y8920 = ~n31719 ;
  assign y8921 = n31721 ;
  assign y8922 = ~n31724 ;
  assign y8923 = ~n31729 ;
  assign y8924 = ~n31731 ;
  assign y8925 = ~n31732 ;
  assign y8926 = ~n31738 ;
  assign y8927 = ~1'b0 ;
  assign y8928 = ~1'b0 ;
endmodule
